
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (NOP, ADDS, LLS, LRS, ADD, SUB, ANDR, ORR, XORR, SNE, SLE, SGE, 
   BEQZ, BNEZ, SUBI, ANDI, ORI, XORI, SLLI, SRLI, SNEI, SLEI, SGEI, LW, SW, 
   SUBU, SUBUI, ADDU, ADDUI, SRA1, SEQ, SLT, SGT, SLTU, SGTU, SGEU, LHI, JR, 
   JALR, SRAI, SEQI, SLTI, SGTI, LB, LBU, LHU, SB, SLTUI, SGTUI, SGEUI);
attribute ENUM_ENCODING of aluOp : type is 
   "000000 000001 000010 000011 000100 000101 000110 000111 001000 001001 001010 001011 001100 001101 001110 001111 010000 010001 010010 010011 010100 010101 010110 010111 011000 011001 011010 011011 011100 011101 011110 011111 100000 100001 100010 100011 100100 100101 100110 100111 101000 101001 101010 101011 101100 101101 101110 101111 110000 110001";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 6 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 6 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "000000" => return NOP;
         when "000001" => return ADDS;
         when "000010" => return LLS;
         when "000011" => return LRS;
         when "000100" => return ADD;
         when "000101" => return SUB;
         when "000110" => return ANDR;
         when "000111" => return ORR;
         when "001000" => return XORR;
         when "001001" => return SNE;
         when "001010" => return SLE;
         when "001011" => return SGE;
         when "001100" => return BEQZ;
         when "001101" => return BNEZ;
         when "001110" => return SUBI;
         when "001111" => return ANDI;
         when "010000" => return ORI;
         when "010001" => return XORI;
         when "010010" => return SLLI;
         when "010011" => return SRLI;
         when "010100" => return SNEI;
         when "010101" => return SLEI;
         when "010110" => return SGEI;
         when "010111" => return LW;
         when "011000" => return SW;
         when "011001" => return SUBU;
         when "011010" => return SUBUI;
         when "011011" => return ADDU;
         when "011100" => return ADDUI;
         when "011101" => return SRA1;
         when "011110" => return SEQ;
         when "011111" => return SLT;
         when "100000" => return SGT;
         when "100001" => return SLTU;
         when "100010" => return SGTU;
         when "100011" => return SGEU;
         when "100100" => return LHI;
         when "100101" => return JR;
         when "100110" => return JALR;
         when "100111" => return SRAI;
         when "101000" => return SEQI;
         when "101001" => return SLTI;
         when "101010" => return SGTI;
         when "101011" => return LB;
         when "101100" => return LBU;
         when "101101" => return LHU;
         when "101110" => return SB;
         when "101111" => return SLTUI;
         when "110000" => return SGTUI;
         when "110001" => return SGEUI;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "000000";
         when ADDS => return "000001";
         when LLS => return "000010";
         when LRS => return "000011";
         when ADD => return "000100";
         when SUB => return "000101";
         when ANDR => return "000110";
         when ORR => return "000111";
         when XORR => return "001000";
         when SNE => return "001001";
         when SLE => return "001010";
         when SGE => return "001011";
         when BEQZ => return "001100";
         when BNEZ => return "001101";
         when SUBI => return "001110";
         when ANDI => return "001111";
         when ORI => return "010000";
         when XORI => return "010001";
         when SLLI => return "010010";
         when SRLI => return "010011";
         when SNEI => return "010100";
         when SLEI => return "010101";
         when SGEI => return "010110";
         when LW => return "010111";
         when SW => return "011000";
         when SUBU => return "011001";
         when SUBUI => return "011010";
         when ADDU => return "011011";
         when ADDUI => return "011100";
         when SRA1 => return "011101";
         when SEQ => return "011110";
         when SLT => return "011111";
         when SGT => return "100000";
         when SLTU => return "100001";
         when SGTU => return "100010";
         when SGEU => return "100011";
         when LHI => return "100100";
         when JR => return "100101";
         when JALR => return "100110";
         when SRAI => return "100111";
         when SEQI => return "101000";
         when SLTI => return "101001";
         when SGTI => return "101010";
         when LB => return "101011";
         when LBU => return "101100";
         when LHU => return "101101";
         when SB => return "101110";
         when SLTUI => return "101111";
         when SGTUI => return "110000";
         when SGEUI => return "110001";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "000000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_rbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_rbsh_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rbsh_0 is

   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal MR_int_1_31_port, MR_int_1_30_port, MR_int_1_29_port, 
      MR_int_1_28_port, MR_int_1_27_port, MR_int_1_26_port, MR_int_1_25_port, 
      MR_int_1_24_port, MR_int_1_23_port, MR_int_1_22_port, MR_int_1_21_port, 
      MR_int_1_20_port, MR_int_1_19_port, MR_int_1_18_port, MR_int_1_17_port, 
      MR_int_1_16_port, MR_int_1_15_port, MR_int_1_14_port, MR_int_1_13_port, 
      MR_int_1_12_port, MR_int_1_11_port, MR_int_1_10_port, MR_int_1_9_port, 
      MR_int_1_8_port, MR_int_1_7_port, MR_int_1_6_port, MR_int_1_5_port, 
      MR_int_1_4_port, MR_int_1_3_port, MR_int_1_2_port, MR_int_1_1_port, 
      MR_int_1_0_port, MR_int_2_31_port, MR_int_2_30_port, MR_int_2_29_port, 
      MR_int_2_28_port, MR_int_2_27_port, MR_int_2_26_port, MR_int_2_25_port, 
      MR_int_2_24_port, MR_int_2_23_port, MR_int_2_22_port, MR_int_2_21_port, 
      MR_int_2_20_port, MR_int_2_19_port, MR_int_2_18_port, MR_int_2_17_port, 
      MR_int_2_16_port, MR_int_2_15_port, MR_int_2_14_port, MR_int_2_13_port, 
      MR_int_2_12_port, MR_int_2_11_port, MR_int_2_10_port, MR_int_2_9_port, 
      MR_int_2_8_port, MR_int_2_7_port, MR_int_2_6_port, MR_int_2_5_port, 
      MR_int_2_4_port, MR_int_2_3_port, MR_int_2_2_port, MR_int_2_1_port, 
      MR_int_2_0_port, MR_int_3_31_port, MR_int_3_30_port, MR_int_3_29_port, 
      MR_int_3_28_port, MR_int_3_27_port, MR_int_3_26_port, MR_int_3_25_port, 
      MR_int_3_24_port, MR_int_3_23_port, MR_int_3_22_port, MR_int_3_21_port, 
      MR_int_3_20_port, MR_int_3_19_port, MR_int_3_18_port, MR_int_3_17_port, 
      MR_int_3_16_port, MR_int_3_15_port, MR_int_3_14_port, MR_int_3_13_port, 
      MR_int_3_12_port, MR_int_3_11_port, MR_int_3_10_port, MR_int_3_9_port, 
      MR_int_3_8_port, MR_int_3_7_port, MR_int_3_6_port, MR_int_3_5_port, 
      MR_int_3_4_port, MR_int_3_3_port, MR_int_3_2_port, MR_int_3_1_port, 
      MR_int_3_0_port, MR_int_4_31_port, MR_int_4_30_port, MR_int_4_29_port, 
      MR_int_4_28_port, MR_int_4_27_port, MR_int_4_26_port, MR_int_4_25_port, 
      MR_int_4_24_port, MR_int_4_23_port, MR_int_4_22_port, MR_int_4_21_port, 
      MR_int_4_20_port, MR_int_4_19_port, MR_int_4_18_port, MR_int_4_17_port, 
      MR_int_4_16_port, MR_int_4_15_port, MR_int_4_14_port, MR_int_4_13_port, 
      MR_int_4_12_port, MR_int_4_11_port, MR_int_4_10_port, MR_int_4_9_port, 
      MR_int_4_8_port, MR_int_4_7_port, MR_int_4_6_port, MR_int_4_5_port, 
      MR_int_4_4_port, MR_int_4_3_port, MR_int_4_2_port, MR_int_4_1_port, 
      MR_int_4_0_port, n1, n2, n3 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => MR_int_4_31_port, B => MR_int_4_15_port, S 
                           => n3, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => MR_int_4_30_port, B => MR_int_4_14_port, S 
                           => n3, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => MR_int_4_29_port, B => MR_int_4_13_port, S 
                           => n3, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => MR_int_4_28_port, B => MR_int_4_12_port, S 
                           => n3, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => MR_int_4_27_port, B => MR_int_4_11_port, S 
                           => n3, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => MR_int_4_26_port, B => MR_int_4_10_port, S 
                           => n3, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => MR_int_4_25_port, B => MR_int_4_9_port, S 
                           => n3, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => MR_int_4_24_port, B => MR_int_4_8_port, S 
                           => n3, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => MR_int_4_23_port, B => MR_int_4_7_port, S 
                           => n2, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => MR_int_4_22_port, B => MR_int_4_6_port, S 
                           => n2, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => MR_int_4_21_port, B => MR_int_4_5_port, S 
                           => n2, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => MR_int_4_20_port, B => MR_int_4_4_port, S 
                           => n2, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => MR_int_4_19_port, B => MR_int_4_3_port, S 
                           => n2, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => MR_int_4_18_port, B => MR_int_4_2_port, S 
                           => n2, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => MR_int_4_17_port, B => MR_int_4_1_port, S 
                           => n2, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => MR_int_4_16_port, B => MR_int_4_0_port, S 
                           => n2, Z => B(16));
   M1_4_15 : MUX2_X1 port map( A => MR_int_4_15_port, B => MR_int_4_31_port, S 
                           => n2, Z => B(15));
   M1_4_14 : MUX2_X1 port map( A => MR_int_4_14_port, B => MR_int_4_30_port, S 
                           => n2, Z => B(14));
   M1_4_13 : MUX2_X1 port map( A => MR_int_4_13_port, B => MR_int_4_29_port, S 
                           => n2, Z => B(13));
   M1_4_12 : MUX2_X1 port map( A => MR_int_4_12_port, B => MR_int_4_28_port, S 
                           => n2, Z => B(12));
   M1_4_11 : MUX2_X1 port map( A => MR_int_4_11_port, B => MR_int_4_27_port, S 
                           => n1, Z => B(11));
   M1_4_10 : MUX2_X1 port map( A => MR_int_4_10_port, B => MR_int_4_26_port, S 
                           => n1, Z => B(10));
   M1_4_9 : MUX2_X1 port map( A => MR_int_4_9_port, B => MR_int_4_25_port, S =>
                           n1, Z => B(9));
   M1_4_8 : MUX2_X1 port map( A => MR_int_4_8_port, B => MR_int_4_24_port, S =>
                           n1, Z => B(8));
   M1_4_7 : MUX2_X1 port map( A => MR_int_4_7_port, B => MR_int_4_23_port, S =>
                           n1, Z => B(7));
   M1_4_6 : MUX2_X1 port map( A => MR_int_4_6_port, B => MR_int_4_22_port, S =>
                           n1, Z => B(6));
   M1_4_5 : MUX2_X1 port map( A => MR_int_4_5_port, B => MR_int_4_21_port, S =>
                           n1, Z => B(5));
   M1_4_4 : MUX2_X1 port map( A => MR_int_4_4_port, B => MR_int_4_20_port, S =>
                           n1, Z => B(4));
   M1_4_3 : MUX2_X1 port map( A => MR_int_4_3_port, B => MR_int_4_19_port, S =>
                           n1, Z => B(3));
   M1_4_2 : MUX2_X1 port map( A => MR_int_4_2_port, B => MR_int_4_18_port, S =>
                           n1, Z => B(2));
   M1_4_1 : MUX2_X1 port map( A => MR_int_4_1_port, B => MR_int_4_17_port, S =>
                           n1, Z => B(1));
   M1_4_0 : MUX2_X1 port map( A => MR_int_4_0_port, B => MR_int_4_16_port, S =>
                           n1, Z => B(0));
   M1_3_31_0 : MUX2_X1 port map( A => MR_int_3_31_port, B => MR_int_3_7_port, S
                           => SH(3), Z => MR_int_4_31_port);
   M1_3_30_0 : MUX2_X1 port map( A => MR_int_3_30_port, B => MR_int_3_6_port, S
                           => SH(3), Z => MR_int_4_30_port);
   M1_3_29_0 : MUX2_X1 port map( A => MR_int_3_29_port, B => MR_int_3_5_port, S
                           => SH(3), Z => MR_int_4_29_port);
   M1_3_28_0 : MUX2_X1 port map( A => MR_int_3_28_port, B => MR_int_3_4_port, S
                           => SH(3), Z => MR_int_4_28_port);
   M1_3_27_0 : MUX2_X1 port map( A => MR_int_3_27_port, B => MR_int_3_3_port, S
                           => SH(3), Z => MR_int_4_27_port);
   M1_3_26_0 : MUX2_X1 port map( A => MR_int_3_26_port, B => MR_int_3_2_port, S
                           => SH(3), Z => MR_int_4_26_port);
   M1_3_25_0 : MUX2_X1 port map( A => MR_int_3_25_port, B => MR_int_3_1_port, S
                           => SH(3), Z => MR_int_4_25_port);
   M1_3_24_0 : MUX2_X1 port map( A => MR_int_3_24_port, B => MR_int_3_0_port, S
                           => SH(3), Z => MR_int_4_24_port);
   M1_3_23_0 : MUX2_X1 port map( A => MR_int_3_23_port, B => MR_int_3_31_port, 
                           S => SH(3), Z => MR_int_4_23_port);
   M1_3_22_0 : MUX2_X1 port map( A => MR_int_3_22_port, B => MR_int_3_30_port, 
                           S => SH(3), Z => MR_int_4_22_port);
   M1_3_21_0 : MUX2_X1 port map( A => MR_int_3_21_port, B => MR_int_3_29_port, 
                           S => SH(3), Z => MR_int_4_21_port);
   M1_3_20_0 : MUX2_X1 port map( A => MR_int_3_20_port, B => MR_int_3_28_port, 
                           S => SH(3), Z => MR_int_4_20_port);
   M1_3_19_0 : MUX2_X1 port map( A => MR_int_3_19_port, B => MR_int_3_27_port, 
                           S => SH(3), Z => MR_int_4_19_port);
   M1_3_18_0 : MUX2_X1 port map( A => MR_int_3_18_port, B => MR_int_3_26_port, 
                           S => SH(3), Z => MR_int_4_18_port);
   M1_3_17_0 : MUX2_X1 port map( A => MR_int_3_17_port, B => MR_int_3_25_port, 
                           S => SH(3), Z => MR_int_4_17_port);
   M1_3_16_0 : MUX2_X1 port map( A => MR_int_3_16_port, B => MR_int_3_24_port, 
                           S => SH(3), Z => MR_int_4_16_port);
   M1_3_15_0 : MUX2_X1 port map( A => MR_int_3_15_port, B => MR_int_3_23_port, 
                           S => SH(3), Z => MR_int_4_15_port);
   M1_3_14_0 : MUX2_X1 port map( A => MR_int_3_14_port, B => MR_int_3_22_port, 
                           S => SH(3), Z => MR_int_4_14_port);
   M1_3_13_0 : MUX2_X1 port map( A => MR_int_3_13_port, B => MR_int_3_21_port, 
                           S => SH(3), Z => MR_int_4_13_port);
   M1_3_12_0 : MUX2_X1 port map( A => MR_int_3_12_port, B => MR_int_3_20_port, 
                           S => SH(3), Z => MR_int_4_12_port);
   M1_3_11_0 : MUX2_X1 port map( A => MR_int_3_11_port, B => MR_int_3_19_port, 
                           S => SH(3), Z => MR_int_4_11_port);
   M1_3_10_0 : MUX2_X1 port map( A => MR_int_3_10_port, B => MR_int_3_18_port, 
                           S => SH(3), Z => MR_int_4_10_port);
   M1_3_9_0 : MUX2_X1 port map( A => MR_int_3_9_port, B => MR_int_3_17_port, S 
                           => SH(3), Z => MR_int_4_9_port);
   M1_3_8_0 : MUX2_X1 port map( A => MR_int_3_8_port, B => MR_int_3_16_port, S 
                           => SH(3), Z => MR_int_4_8_port);
   M1_3_7 : MUX2_X1 port map( A => MR_int_3_7_port, B => MR_int_3_15_port, S =>
                           SH(3), Z => MR_int_4_7_port);
   M1_3_6 : MUX2_X1 port map( A => MR_int_3_6_port, B => MR_int_3_14_port, S =>
                           SH(3), Z => MR_int_4_6_port);
   M1_3_5 : MUX2_X1 port map( A => MR_int_3_5_port, B => MR_int_3_13_port, S =>
                           SH(3), Z => MR_int_4_5_port);
   M1_3_4 : MUX2_X1 port map( A => MR_int_3_4_port, B => MR_int_3_12_port, S =>
                           SH(3), Z => MR_int_4_4_port);
   M1_3_3 : MUX2_X1 port map( A => MR_int_3_3_port, B => MR_int_3_11_port, S =>
                           SH(3), Z => MR_int_4_3_port);
   M1_3_2 : MUX2_X1 port map( A => MR_int_3_2_port, B => MR_int_3_10_port, S =>
                           SH(3), Z => MR_int_4_2_port);
   M1_3_1 : MUX2_X1 port map( A => MR_int_3_1_port, B => MR_int_3_9_port, S => 
                           SH(3), Z => MR_int_4_1_port);
   M1_3_0 : MUX2_X1 port map( A => MR_int_3_0_port, B => MR_int_3_8_port, S => 
                           SH(3), Z => MR_int_4_0_port);
   M1_2_31_0 : MUX2_X1 port map( A => MR_int_2_31_port, B => MR_int_2_3_port, S
                           => SH(2), Z => MR_int_3_31_port);
   M1_2_30_0 : MUX2_X1 port map( A => MR_int_2_30_port, B => MR_int_2_2_port, S
                           => SH(2), Z => MR_int_3_30_port);
   M1_2_29_0 : MUX2_X1 port map( A => MR_int_2_29_port, B => MR_int_2_1_port, S
                           => SH(2), Z => MR_int_3_29_port);
   M1_2_28_0 : MUX2_X1 port map( A => MR_int_2_28_port, B => MR_int_2_0_port, S
                           => SH(2), Z => MR_int_3_28_port);
   M1_2_27_0 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, 
                           S => SH(2), Z => MR_int_3_27_port);
   M1_2_26_0 : MUX2_X1 port map( A => MR_int_2_26_port, B => MR_int_2_30_port, 
                           S => SH(2), Z => MR_int_3_26_port);
   M1_2_25_0 : MUX2_X1 port map( A => MR_int_2_25_port, B => MR_int_2_29_port, 
                           S => SH(2), Z => MR_int_3_25_port);
   M1_2_24_0 : MUX2_X1 port map( A => MR_int_2_24_port, B => MR_int_2_28_port, 
                           S => SH(2), Z => MR_int_3_24_port);
   M1_2_23_0 : MUX2_X1 port map( A => MR_int_2_23_port, B => MR_int_2_27_port, 
                           S => SH(2), Z => MR_int_3_23_port);
   M1_2_22_0 : MUX2_X1 port map( A => MR_int_2_22_port, B => MR_int_2_26_port, 
                           S => SH(2), Z => MR_int_3_22_port);
   M1_2_21_0 : MUX2_X1 port map( A => MR_int_2_21_port, B => MR_int_2_25_port, 
                           S => SH(2), Z => MR_int_3_21_port);
   M1_2_20_0 : MUX2_X1 port map( A => MR_int_2_20_port, B => MR_int_2_24_port, 
                           S => SH(2), Z => MR_int_3_20_port);
   M1_2_19_0 : MUX2_X1 port map( A => MR_int_2_19_port, B => MR_int_2_23_port, 
                           S => SH(2), Z => MR_int_3_19_port);
   M1_2_18_0 : MUX2_X1 port map( A => MR_int_2_18_port, B => MR_int_2_22_port, 
                           S => SH(2), Z => MR_int_3_18_port);
   M1_2_17_0 : MUX2_X1 port map( A => MR_int_2_17_port, B => MR_int_2_21_port, 
                           S => SH(2), Z => MR_int_3_17_port);
   M1_2_16_0 : MUX2_X1 port map( A => MR_int_2_16_port, B => MR_int_2_20_port, 
                           S => SH(2), Z => MR_int_3_16_port);
   M1_2_15_0 : MUX2_X1 port map( A => MR_int_2_15_port, B => MR_int_2_19_port, 
                           S => SH(2), Z => MR_int_3_15_port);
   M1_2_14_0 : MUX2_X1 port map( A => MR_int_2_14_port, B => MR_int_2_18_port, 
                           S => SH(2), Z => MR_int_3_14_port);
   M1_2_13_0 : MUX2_X1 port map( A => MR_int_2_13_port, B => MR_int_2_17_port, 
                           S => SH(2), Z => MR_int_3_13_port);
   M1_2_12_0 : MUX2_X1 port map( A => MR_int_2_12_port, B => MR_int_2_16_port, 
                           S => SH(2), Z => MR_int_3_12_port);
   M1_2_11_0 : MUX2_X1 port map( A => MR_int_2_11_port, B => MR_int_2_15_port, 
                           S => SH(2), Z => MR_int_3_11_port);
   M1_2_10_0 : MUX2_X1 port map( A => MR_int_2_10_port, B => MR_int_2_14_port, 
                           S => SH(2), Z => MR_int_3_10_port);
   M1_2_9_0 : MUX2_X1 port map( A => MR_int_2_9_port, B => MR_int_2_13_port, S 
                           => SH(2), Z => MR_int_3_9_port);
   M1_2_8_0 : MUX2_X1 port map( A => MR_int_2_8_port, B => MR_int_2_12_port, S 
                           => SH(2), Z => MR_int_3_8_port);
   M1_2_7_0 : MUX2_X1 port map( A => MR_int_2_7_port, B => MR_int_2_11_port, S 
                           => SH(2), Z => MR_int_3_7_port);
   M1_2_6_0 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_10_port, S 
                           => SH(2), Z => MR_int_3_6_port);
   M1_2_5_0 : MUX2_X1 port map( A => MR_int_2_5_port, B => MR_int_2_9_port, S 
                           => SH(2), Z => MR_int_3_5_port);
   M1_2_4_0 : MUX2_X1 port map( A => MR_int_2_4_port, B => MR_int_2_8_port, S 
                           => SH(2), Z => MR_int_3_4_port);
   M1_2_3 : MUX2_X1 port map( A => MR_int_2_3_port, B => MR_int_2_7_port, S => 
                           SH(2), Z => MR_int_3_3_port);
   M1_2_2 : MUX2_X1 port map( A => MR_int_2_2_port, B => MR_int_2_6_port, S => 
                           SH(2), Z => MR_int_3_2_port);
   M1_2_1 : MUX2_X1 port map( A => MR_int_2_1_port, B => MR_int_2_5_port, S => 
                           SH(2), Z => MR_int_3_1_port);
   M1_2_0 : MUX2_X1 port map( A => MR_int_2_0_port, B => MR_int_2_4_port, S => 
                           SH(2), Z => MR_int_3_0_port);
   M1_1_31_0 : MUX2_X1 port map( A => MR_int_1_31_port, B => MR_int_1_1_port, S
                           => SH(1), Z => MR_int_2_31_port);
   M1_1_30_0 : MUX2_X1 port map( A => MR_int_1_30_port, B => MR_int_1_0_port, S
                           => SH(1), Z => MR_int_2_30_port);
   M1_1_29_0 : MUX2_X1 port map( A => MR_int_1_29_port, B => MR_int_1_31_port, 
                           S => SH(1), Z => MR_int_2_29_port);
   M1_1_28_0 : MUX2_X1 port map( A => MR_int_1_28_port, B => MR_int_1_30_port, 
                           S => SH(1), Z => MR_int_2_28_port);
   M1_1_27_0 : MUX2_X1 port map( A => MR_int_1_27_port, B => MR_int_1_29_port, 
                           S => SH(1), Z => MR_int_2_27_port);
   M1_1_26_0 : MUX2_X1 port map( A => MR_int_1_26_port, B => MR_int_1_28_port, 
                           S => SH(1), Z => MR_int_2_26_port);
   M1_1_25_0 : MUX2_X1 port map( A => MR_int_1_25_port, B => MR_int_1_27_port, 
                           S => SH(1), Z => MR_int_2_25_port);
   M1_1_24_0 : MUX2_X1 port map( A => MR_int_1_24_port, B => MR_int_1_26_port, 
                           S => SH(1), Z => MR_int_2_24_port);
   M1_1_23_0 : MUX2_X1 port map( A => MR_int_1_23_port, B => MR_int_1_25_port, 
                           S => SH(1), Z => MR_int_2_23_port);
   M1_1_22_0 : MUX2_X1 port map( A => MR_int_1_22_port, B => MR_int_1_24_port, 
                           S => SH(1), Z => MR_int_2_22_port);
   M1_1_21_0 : MUX2_X1 port map( A => MR_int_1_21_port, B => MR_int_1_23_port, 
                           S => SH(1), Z => MR_int_2_21_port);
   M1_1_20_0 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_22_port, 
                           S => SH(1), Z => MR_int_2_20_port);
   M1_1_19_0 : MUX2_X1 port map( A => MR_int_1_19_port, B => MR_int_1_21_port, 
                           S => SH(1), Z => MR_int_2_19_port);
   M1_1_18_0 : MUX2_X1 port map( A => MR_int_1_18_port, B => MR_int_1_20_port, 
                           S => SH(1), Z => MR_int_2_18_port);
   M1_1_17_0 : MUX2_X1 port map( A => MR_int_1_17_port, B => MR_int_1_19_port, 
                           S => SH(1), Z => MR_int_2_17_port);
   M1_1_16_0 : MUX2_X1 port map( A => MR_int_1_16_port, B => MR_int_1_18_port, 
                           S => SH(1), Z => MR_int_2_16_port);
   M1_1_15_0 : MUX2_X1 port map( A => MR_int_1_15_port, B => MR_int_1_17_port, 
                           S => SH(1), Z => MR_int_2_15_port);
   M1_1_14_0 : MUX2_X1 port map( A => MR_int_1_14_port, B => MR_int_1_16_port, 
                           S => SH(1), Z => MR_int_2_14_port);
   M1_1_13_0 : MUX2_X1 port map( A => MR_int_1_13_port, B => MR_int_1_15_port, 
                           S => SH(1), Z => MR_int_2_13_port);
   M1_1_12_0 : MUX2_X1 port map( A => MR_int_1_12_port, B => MR_int_1_14_port, 
                           S => SH(1), Z => MR_int_2_12_port);
   M1_1_11_0 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_13_port, 
                           S => SH(1), Z => MR_int_2_11_port);
   M1_1_10_0 : MUX2_X1 port map( A => MR_int_1_10_port, B => MR_int_1_12_port, 
                           S => SH(1), Z => MR_int_2_10_port);
   M1_1_9_0 : MUX2_X1 port map( A => MR_int_1_9_port, B => MR_int_1_11_port, S 
                           => SH(1), Z => MR_int_2_9_port);
   M1_1_8_0 : MUX2_X1 port map( A => MR_int_1_8_port, B => MR_int_1_10_port, S 
                           => SH(1), Z => MR_int_2_8_port);
   M1_1_7_0 : MUX2_X1 port map( A => MR_int_1_7_port, B => MR_int_1_9_port, S 
                           => SH(1), Z => MR_int_2_7_port);
   M1_1_6_0 : MUX2_X1 port map( A => MR_int_1_6_port, B => MR_int_1_8_port, S 
                           => SH(1), Z => MR_int_2_6_port);
   M1_1_5_0 : MUX2_X1 port map( A => MR_int_1_5_port, B => MR_int_1_7_port, S 
                           => SH(1), Z => MR_int_2_5_port);
   M1_1_4_0 : MUX2_X1 port map( A => MR_int_1_4_port, B => MR_int_1_6_port, S 
                           => SH(1), Z => MR_int_2_4_port);
   M1_1_3_0 : MUX2_X1 port map( A => MR_int_1_3_port, B => MR_int_1_5_port, S 
                           => SH(1), Z => MR_int_2_3_port);
   M1_1_2_0 : MUX2_X1 port map( A => MR_int_1_2_port, B => MR_int_1_4_port, S 
                           => SH(1), Z => MR_int_2_2_port);
   M1_1_1 : MUX2_X1 port map( A => MR_int_1_1_port, B => MR_int_1_3_port, S => 
                           SH(1), Z => MR_int_2_1_port);
   M1_1_0 : MUX2_X1 port map( A => MR_int_1_0_port, B => MR_int_1_2_port, S => 
                           SH(1), Z => MR_int_2_0_port);
   M1_0_31_0 : MUX2_X1 port map( A => A(31), B => A(0), S => SH(0), Z => 
                           MR_int_1_31_port);
   M1_0_30_0 : MUX2_X1 port map( A => A(30), B => A(31), S => SH(0), Z => 
                           MR_int_1_30_port);
   M1_0_29_0 : MUX2_X1 port map( A => A(29), B => A(30), S => SH(0), Z => 
                           MR_int_1_29_port);
   M1_0_28_0 : MUX2_X1 port map( A => A(28), B => A(29), S => SH(0), Z => 
                           MR_int_1_28_port);
   M1_0_27_0 : MUX2_X1 port map( A => A(27), B => A(28), S => SH(0), Z => 
                           MR_int_1_27_port);
   M1_0_26_0 : MUX2_X1 port map( A => A(26), B => A(27), S => SH(0), Z => 
                           MR_int_1_26_port);
   M1_0_25_0 : MUX2_X1 port map( A => A(25), B => A(26), S => SH(0), Z => 
                           MR_int_1_25_port);
   M1_0_24_0 : MUX2_X1 port map( A => A(24), B => A(25), S => SH(0), Z => 
                           MR_int_1_24_port);
   M1_0_23_0 : MUX2_X1 port map( A => A(23), B => A(24), S => SH(0), Z => 
                           MR_int_1_23_port);
   M1_0_22_0 : MUX2_X1 port map( A => A(22), B => A(23), S => SH(0), Z => 
                           MR_int_1_22_port);
   M1_0_21_0 : MUX2_X1 port map( A => A(21), B => A(22), S => SH(0), Z => 
                           MR_int_1_21_port);
   M1_0_20_0 : MUX2_X1 port map( A => A(20), B => A(21), S => SH(0), Z => 
                           MR_int_1_20_port);
   M1_0_19_0 : MUX2_X1 port map( A => A(19), B => A(20), S => SH(0), Z => 
                           MR_int_1_19_port);
   M1_0_18_0 : MUX2_X1 port map( A => A(18), B => A(19), S => SH(0), Z => 
                           MR_int_1_18_port);
   M1_0_17_0 : MUX2_X1 port map( A => A(17), B => A(18), S => SH(0), Z => 
                           MR_int_1_17_port);
   M1_0_16_0 : MUX2_X1 port map( A => A(16), B => A(17), S => SH(0), Z => 
                           MR_int_1_16_port);
   M1_0_15_0 : MUX2_X1 port map( A => A(15), B => A(16), S => SH(0), Z => 
                           MR_int_1_15_port);
   M1_0_14_0 : MUX2_X1 port map( A => A(14), B => A(15), S => SH(0), Z => 
                           MR_int_1_14_port);
   M1_0_13_0 : MUX2_X1 port map( A => A(13), B => A(14), S => SH(0), Z => 
                           MR_int_1_13_port);
   M1_0_12_0 : MUX2_X1 port map( A => A(12), B => A(13), S => SH(0), Z => 
                           MR_int_1_12_port);
   M1_0_11_0 : MUX2_X1 port map( A => A(11), B => A(12), S => SH(0), Z => 
                           MR_int_1_11_port);
   M1_0_10_0 : MUX2_X1 port map( A => A(10), B => A(11), S => SH(0), Z => 
                           MR_int_1_10_port);
   M1_0_9_0 : MUX2_X1 port map( A => A(9), B => A(10), S => SH(0), Z => 
                           MR_int_1_9_port);
   M1_0_8_0 : MUX2_X1 port map( A => A(8), B => A(9), S => SH(0), Z => 
                           MR_int_1_8_port);
   M1_0_7_0 : MUX2_X1 port map( A => A(7), B => A(8), S => SH(0), Z => 
                           MR_int_1_7_port);
   M1_0_6_0 : MUX2_X1 port map( A => A(6), B => A(7), S => SH(0), Z => 
                           MR_int_1_6_port);
   M1_0_5_0 : MUX2_X1 port map( A => A(5), B => A(6), S => SH(0), Z => 
                           MR_int_1_5_port);
   M1_0_4_0 : MUX2_X1 port map( A => A(4), B => A(5), S => SH(0), Z => 
                           MR_int_1_4_port);
   M1_0_3_0 : MUX2_X1 port map( A => A(3), B => A(4), S => SH(0), Z => 
                           MR_int_1_3_port);
   M1_0_2_0 : MUX2_X1 port map( A => A(2), B => A(3), S => SH(0), Z => 
                           MR_int_1_2_port);
   M1_0_1_0 : MUX2_X1 port map( A => A(1), B => A(2), S => SH(0), Z => 
                           MR_int_1_1_port);
   M1_0_0 : MUX2_X1 port map( A => A(0), B => A(1), S => SH(0), Z => 
                           MR_int_1_0_port);
   U2 : CLKBUF_X3 port map( A => SH(4), Z => n1);
   U3 : CLKBUF_X3 port map( A => SH(4), Z => n2);
   U4 : CLKBUF_X3 port map( A => SH(4), Z => n3);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_lbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_lbsh_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_lbsh_0 is

   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n1, n2, n3 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n3, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n3, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n3, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n3, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n3, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n3, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n3, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n3, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n2, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n2, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n2, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n2, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n2, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n2, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n2, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n2, Z => B(16));
   M0_4_15 : MUX2_X1 port map( A => ML_int_4_15_port, B => ML_int_4_31_port, S 
                           => n2, Z => B(15));
   M0_4_14 : MUX2_X1 port map( A => ML_int_4_14_port, B => ML_int_4_30_port, S 
                           => n2, Z => B(14));
   M0_4_13 : MUX2_X1 port map( A => ML_int_4_13_port, B => ML_int_4_29_port, S 
                           => n2, Z => B(13));
   M0_4_12 : MUX2_X1 port map( A => ML_int_4_12_port, B => ML_int_4_28_port, S 
                           => n2, Z => B(12));
   M0_4_11 : MUX2_X1 port map( A => ML_int_4_11_port, B => ML_int_4_27_port, S 
                           => n1, Z => B(11));
   M0_4_10 : MUX2_X1 port map( A => ML_int_4_10_port, B => ML_int_4_26_port, S 
                           => n1, Z => B(10));
   M0_4_9 : MUX2_X1 port map( A => ML_int_4_9_port, B => ML_int_4_25_port, S =>
                           n1, Z => B(9));
   M0_4_8 : MUX2_X1 port map( A => ML_int_4_8_port, B => ML_int_4_24_port, S =>
                           n1, Z => B(8));
   M0_4_7 : MUX2_X1 port map( A => ML_int_4_7_port, B => ML_int_4_23_port, S =>
                           n1, Z => B(7));
   M0_4_6 : MUX2_X1 port map( A => ML_int_4_6_port, B => ML_int_4_22_port, S =>
                           n1, Z => B(6));
   M0_4_5 : MUX2_X1 port map( A => ML_int_4_5_port, B => ML_int_4_21_port, S =>
                           n1, Z => B(5));
   M0_4_4 : MUX2_X1 port map( A => ML_int_4_4_port, B => ML_int_4_20_port, S =>
                           n1, Z => B(4));
   M0_4_3 : MUX2_X1 port map( A => ML_int_4_3_port, B => ML_int_4_19_port, S =>
                           n1, Z => B(3));
   M0_4_2 : MUX2_X1 port map( A => ML_int_4_2_port, B => ML_int_4_18_port, S =>
                           n1, Z => B(2));
   M0_4_1 : MUX2_X1 port map( A => ML_int_4_1_port, B => ML_int_4_17_port, S =>
                           n1, Z => B(1));
   M0_4_0 : MUX2_X1 port map( A => ML_int_4_0_port, B => ML_int_4_16_port, S =>
                           n1, Z => B(0));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => SH(3), Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => SH(3), Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => SH(3), Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => SH(3), Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => SH(3), Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => SH(3), Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => SH(3), Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => SH(3), Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => SH(3), Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => SH(3), Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => SH(3), Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => SH(3), Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => SH(3), Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => SH(3), Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => SH(3), Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => SH(3), Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => SH(3), Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => SH(3), Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => SH(3), Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => SH(3), Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           SH(3), Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           SH(3), Z => ML_int_4_8_port);
   M0_3_7 : MUX2_X1 port map( A => ML_int_3_7_port, B => ML_int_3_31_port, S =>
                           SH(3), Z => ML_int_4_7_port);
   M0_3_6 : MUX2_X1 port map( A => ML_int_3_6_port, B => ML_int_3_30_port, S =>
                           SH(3), Z => ML_int_4_6_port);
   M0_3_5 : MUX2_X1 port map( A => ML_int_3_5_port, B => ML_int_3_29_port, S =>
                           SH(3), Z => ML_int_4_5_port);
   M0_3_4 : MUX2_X1 port map( A => ML_int_3_4_port, B => ML_int_3_28_port, S =>
                           SH(3), Z => ML_int_4_4_port);
   M0_3_3 : MUX2_X1 port map( A => ML_int_3_3_port, B => ML_int_3_27_port, S =>
                           SH(3), Z => ML_int_4_3_port);
   M0_3_2 : MUX2_X1 port map( A => ML_int_3_2_port, B => ML_int_3_26_port, S =>
                           SH(3), Z => ML_int_4_2_port);
   M0_3_1 : MUX2_X1 port map( A => ML_int_3_1_port, B => ML_int_3_25_port, S =>
                           SH(3), Z => ML_int_4_1_port);
   M0_3_0 : MUX2_X1 port map( A => ML_int_3_0_port, B => ML_int_3_24_port, S =>
                           SH(3), Z => ML_int_4_0_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => SH(2), Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => SH(2), Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => SH(2), Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => SH(2), Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => SH(2), Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => SH(2), Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => SH(2), Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => SH(2), Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => SH(2), Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => SH(2), Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => SH(2), Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => SH(2), Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => SH(2), Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => SH(2), Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => SH(2), Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => SH(2), Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => SH(2), Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => SH(2), Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           SH(2), Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           SH(2), Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           SH(2), Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           SH(2), Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           SH(2), Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           SH(2), Z => ML_int_3_4_port);
   M0_2_3 : MUX2_X1 port map( A => ML_int_2_3_port, B => ML_int_2_31_port, S =>
                           SH(2), Z => ML_int_3_3_port);
   M0_2_2 : MUX2_X1 port map( A => ML_int_2_2_port, B => ML_int_2_30_port, S =>
                           SH(2), Z => ML_int_3_2_port);
   M0_2_1 : MUX2_X1 port map( A => ML_int_2_1_port, B => ML_int_2_29_port, S =>
                           SH(2), Z => ML_int_3_1_port);
   M0_2_0 : MUX2_X1 port map( A => ML_int_2_0_port, B => ML_int_2_28_port, S =>
                           SH(2), Z => ML_int_3_0_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => SH(1), Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => SH(1), Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => SH(1), Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => SH(1), Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => SH(1), Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => SH(1), Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => SH(1), Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => SH(1), Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => SH(1), Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => SH(1), Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           SH(1), Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           SH(1), Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           SH(1), Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           SH(1), Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           SH(1), Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           SH(1), Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           SH(1), Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           SH(1), Z => ML_int_2_2_port);
   M0_1_1 : MUX2_X1 port map( A => ML_int_1_1_port, B => ML_int_1_31_port, S =>
                           SH(1), Z => ML_int_2_1_port);
   M0_1_0 : MUX2_X1 port map( A => ML_int_1_0_port, B => ML_int_1_30_port, S =>
                           SH(1), Z => ML_int_2_0_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => SH(0), Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => SH(0), Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => SH(0), Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => SH(0), Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => SH(0), Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => SH(0), Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => SH(0), Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => SH(0), Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => SH(0), Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => SH(0), Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => SH(0), Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => SH(0), Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => SH(0), Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => SH(0), Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => SH(0), Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => SH(0), Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => SH(0), Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => SH(0), Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => SH(0), Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => SH(0), Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => SH(0), Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => SH(0), Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => SH(0), Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => SH(0), Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => SH(0), Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => SH(0), Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => SH(0), Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => SH(0), Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => SH(0), Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => SH(0), Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => SH(0), Z => 
                           ML_int_1_1_port);
   M0_0_0 : MUX2_X1 port map( A => A(0), B => A(31), S => SH(0), Z => 
                           ML_int_1_0_port);
   U2 : CLKBUF_X3 port map( A => SH(4), Z => n1);
   U3 : CLKBUF_X3 port map( A => SH(4), Z => n2);
   U4 : CLKBUF_X3 port map( A => SH(4), Z => n3);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sra_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sra_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172 : std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U2 : NOR2_X2 port map( A1 => n131, A2 => SH(0), ZN => n52);
   U3 : AOI221_X4 port map( B1 => n52, B2 => A(6), C1 => n53, C2 => A(7), A => 
                           n171, ZN => n35);
   U4 : AOI221_X4 port map( B1 => n52, B2 => A(14), C1 => n53, C2 => A(15), A 
                           => n162, ZN => n135);
   U5 : AOI221_X4 port map( B1 => n52, B2 => A(10), C1 => n53, C2 => A(11), A 
                           => n158, ZN => n13);
   U6 : AOI221_X4 port map( B1 => n52, B2 => A(12), C1 => n53, C2 => A(13), A 
                           => n155, ZN => n64);
   U7 : AOI221_X4 port map( B1 => n52, B2 => A(16), C1 => n53, C2 => A(17), A 
                           => n152, ZN => n116);
   U8 : NOR2_X2 port map( A1 => n172, A2 => n131, ZN => n53);
   U9 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n75);
   U10 : INV_X1 port map( A => SH(4), ZN => n1);
   U11 : INV_X1 port map( A => SH(4), ZN => n2);
   U12 : OAI221_X1 port map( B1 => n3, B2 => n4, C1 => n5, C2 => n1, A => n6, 
                           ZN => B_9_port);
   U13 : AOI222_X1 port map( A1 => n7, A2 => n8, B1 => n9, B2 => n10, C1 => n11
                           , C2 => n12, ZN => n6);
   U14 : OAI221_X1 port map( B1 => n13, B2 => n4, C1 => n14, C2 => n1, A => n15
                           , ZN => B_8_port);
   U15 : AOI222_X1 port map( A1 => n7, A2 => n16, B1 => n9, B2 => n17, C1 => 
                           n11, C2 => n18, ZN => n15);
   U16 : OAI221_X1 port map( B1 => n19, B2 => n4, C1 => n20, C2 => n1, A => n21
                           , ZN => B_7_port);
   U17 : AOI222_X1 port map( A1 => n7, A2 => n22, B1 => n9, B2 => n23, C1 => 
                           n11, C2 => n24, ZN => n21);
   U18 : OAI221_X1 port map( B1 => n25, B2 => n4, C1 => n26, C2 => n1, A => n27
                           , ZN => B_6_port);
   U19 : AOI222_X1 port map( A1 => n7, A2 => n28, B1 => n9, B2 => n29, C1 => 
                           n11, C2 => n30, ZN => n27);
   U20 : OAI221_X1 port map( B1 => n31, B2 => n4, C1 => n32, C2 => n1, A => n33
                           , ZN => B_5_port);
   U21 : AOI222_X1 port map( A1 => n7, A2 => n34, B1 => n9, B2 => n8, C1 => n11
                           , C2 => n10, ZN => n33);
   U22 : OAI221_X1 port map( B1 => n35, B2 => n4, C1 => n36, C2 => n1, A => n37
                           , ZN => B_4_port);
   U23 : AOI222_X1 port map( A1 => n7, A2 => n38, B1 => n9, B2 => n16, C1 => 
                           n11, C2 => n17, ZN => n37);
   U24 : OAI221_X1 port map( B1 => n19, B2 => n39, C1 => n40, C2 => n1, A => 
                           n41, ZN => B_3_port);
   U25 : AOI222_X1 port map( A1 => n11, A2 => n23, B1 => n42, B2 => n43, C1 => 
                           n9, C2 => n22, ZN => n41);
   U26 : INV_X1 port map( A => n44, ZN => n22);
   U27 : OAI221_X1 port map( B1 => n45, B2 => n46, C1 => n47, C2 => n48, A => 
                           n49, ZN => n43);
   U28 : AOI22_X1 port map( A1 => A(4), A2 => n50, B1 => A(3), B2 => n51, ZN =>
                           n49);
   U29 : AOI221_X1 port map( B1 => n52, B2 => A(9), C1 => n53, C2 => A(10), A 
                           => n54, ZN => n19);
   U30 : OAI22_X1 port map( A1 => n55, A2 => n56, B1 => n57, B2 => n58, ZN => 
                           n54);
   U31 : OAI21_X1 port map( B1 => SH(4), B2 => n59, A => n60, ZN => B_30_port);
   U32 : OAI221_X1 port map( B1 => n25, B2 => n39, C1 => n61, C2 => n1, A => 
                           n62, ZN => B_2_port);
   U33 : AOI222_X1 port map( A1 => n11, A2 => n29, B1 => n42, B2 => n63, C1 => 
                           n9, C2 => n28, ZN => n62);
   U34 : INV_X1 port map( A => n64, ZN => n28);
   U35 : OAI221_X1 port map( B1 => n45, B2 => n65, C1 => n47, C2 => n46, A => 
                           n66, ZN => n63);
   U36 : AOI22_X1 port map( A1 => A(3), A2 => n50, B1 => A(2), B2 => n51, ZN =>
                           n66);
   U37 : AOI221_X1 port map( B1 => n52, B2 => A(8), C1 => n53, C2 => A(9), A =>
                           n67, ZN => n25);
   U38 : OAI22_X1 port map( A1 => n57, A2 => n56, B1 => n48, B2 => n58, ZN => 
                           n67);
   U39 : INV_X1 port map( A => A(7), ZN => n57);
   U40 : OAI21_X1 port map( B1 => SH(4), B2 => n68, A => n60, ZN => B_29_port);
   U41 : OAI21_X1 port map( B1 => SH(4), B2 => n69, A => n60, ZN => B_28_port);
   U42 : OAI21_X1 port map( B1 => SH(4), B2 => n70, A => n60, ZN => B_27_port);
   U43 : OAI21_X1 port map( B1 => SH(4), B2 => n71, A => n60, ZN => B_26_port);
   U44 : OAI21_X1 port map( B1 => SH(4), B2 => n5, A => n60, ZN => B_25_port);
   U45 : AOI221_X1 port map( B1 => n72, B2 => n73, C1 => n74, C2 => n75, A => 
                           n76, ZN => n5);
   U46 : OAI21_X1 port map( B1 => SH(4), B2 => n14, A => n60, ZN => B_24_port);
   U47 : AOI221_X1 port map( B1 => n77, B2 => n73, C1 => n78, C2 => n75, A => 
                           n76, ZN => n14);
   U48 : OAI21_X1 port map( B1 => SH(4), B2 => n20, A => n60, ZN => B_23_port);
   U49 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n80, C2 => n75, A => 
                           n76, ZN => n20);
   U50 : OAI21_X1 port map( B1 => SH(4), B2 => n26, A => n60, ZN => B_22_port);
   U51 : AOI221_X1 port map( B1 => n81, B2 => n73, C1 => n82, C2 => n75, A => 
                           n83, ZN => n26);
   U52 : INV_X1 port map( A => n84, ZN => n83);
   U53 : AOI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n84);
   U54 : OAI21_X1 port map( B1 => SH(4), B2 => n32, A => n60, ZN => B_21_port);
   U55 : AOI221_X1 port map( B1 => n74, B2 => n73, C1 => n12, C2 => n75, A => 
                           n88, ZN => n32);
   U56 : INV_X1 port map( A => n89, ZN => n88);
   U57 : AOI21_X1 port map( B1 => n85, B2 => n72, A => n87, ZN => n89);
   U58 : OAI21_X1 port map( B1 => SH(4), B2 => n36, A => n60, ZN => B_20_port);
   U59 : AOI221_X1 port map( B1 => n78, B2 => n73, C1 => n18, C2 => n75, A => 
                           n90, ZN => n36);
   U60 : INV_X1 port map( A => n91, ZN => n90);
   U61 : AOI21_X1 port map( B1 => n85, B2 => n77, A => n87, ZN => n91);
   U62 : OAI221_X1 port map( B1 => n31, B2 => n39, C1 => n92, C2 => n1, A => 
                           n93, ZN => B_1_port);
   U63 : AOI222_X1 port map( A1 => n11, A2 => n8, B1 => n42, B2 => n94, C1 => 
                           n9, C2 => n34, ZN => n93);
   U64 : INV_X1 port map( A => n3, ZN => n34);
   U65 : AOI221_X1 port map( B1 => n52, B2 => A(11), C1 => n53, C2 => A(12), A 
                           => n95, ZN => n3);
   U66 : OAI22_X1 port map( A1 => n96, A2 => n56, B1 => n97, B2 => n58, ZN => 
                           n95);
   U67 : OAI221_X1 port map( B1 => n45, B2 => n98, C1 => n47, C2 => n65, A => 
                           n99, ZN => n94);
   U68 : AOI22_X1 port map( A1 => A(2), A2 => n50, B1 => A(1), B2 => n51, ZN =>
                           n99);
   U69 : INV_X1 port map( A => n100, ZN => n8);
   U70 : AOI221_X1 port map( B1 => n52, B2 => A(7), C1 => n53, C2 => A(8), A =>
                           n101, ZN => n31);
   U71 : OAI22_X1 port map( A1 => n48, A2 => n56, B1 => n46, B2 => n58, ZN => 
                           n101);
   U72 : INV_X1 port map( A => A(6), ZN => n48);
   U73 : OAI21_X1 port map( B1 => SH(4), B2 => n40, A => n60, ZN => B_19_port);
   U74 : AOI221_X1 port map( B1 => n80, B2 => n73, C1 => n24, C2 => n75, A => 
                           n102, ZN => n40);
   U75 : INV_X1 port map( A => n103, ZN => n102);
   U76 : AOI21_X1 port map( B1 => n85, B2 => n79, A => n87, ZN => n103);
   U77 : NOR2_X1 port map( A1 => n104, A2 => n105, ZN => n87);
   U78 : OAI21_X1 port map( B1 => SH(4), B2 => n61, A => n60, ZN => B_18_port);
   U79 : AOI221_X1 port map( B1 => n86, B2 => n106, C1 => n81, C2 => n85, A => 
                           n107, ZN => n61);
   U80 : INV_X1 port map( A => n108, ZN => n107);
   U81 : AOI22_X1 port map( A1 => n73, A2 => n82, B1 => n75, B2 => n30, ZN => 
                           n108);
   U82 : OAI21_X1 port map( B1 => SH(4), B2 => n92, A => n60, ZN => B_17_port);
   U83 : AOI221_X1 port map( B1 => n12, B2 => n73, C1 => n10, C2 => n75, A => 
                           n109, ZN => n92);
   U84 : INV_X1 port map( A => n110, ZN => n109);
   U85 : AOI22_X1 port map( A1 => n106, A2 => n72, B1 => n85, B2 => n74, ZN => 
                           n110);
   U86 : OAI21_X1 port map( B1 => SH(4), B2 => n111, A => n60, ZN => B_16_port)
                           ;
   U87 : OAI221_X1 port map( B1 => n112, B2 => n39, C1 => n113, C2 => n4, A => 
                           n114, ZN => B_15_port);
   U88 : AOI221_X1 port map( B1 => n11, B2 => n79, C1 => n9, C2 => n80, A => 
                           n115, ZN => n114);
   U89 : INV_X1 port map( A => n60, ZN => n115);
   U90 : NAND2_X1 port map( A1 => SH(4), A2 => A(31), ZN => n60);
   U91 : INV_X1 port map( A => n23, ZN => n113);
   U92 : INV_X1 port map( A => n24, ZN => n112);
   U93 : OAI221_X1 port map( B1 => n116, B2 => n4, C1 => n59, C2 => n1, A => 
                           n117, ZN => B_14_port);
   U94 : AOI222_X1 port map( A1 => n7, A2 => n30, B1 => n9, B2 => n82, C1 => 
                           n11, C2 => n81, ZN => n117);
   U95 : AOI21_X1 port map( B1 => n86, B2 => n75, A => n118, ZN => n59);
   U96 : OAI221_X1 port map( B1 => n100, B2 => n4, C1 => n68, C2 => n2, A => 
                           n119, ZN => B_13_port);
   U97 : AOI222_X1 port map( A1 => n7, A2 => n10, B1 => n9, B2 => n12, C1 => 
                           n11, C2 => n74, ZN => n119);
   U98 : OAI221_X1 port map( B1 => n45, B2 => n120, C1 => n47, C2 => n121, A =>
                           n122, ZN => n74);
   U99 : AOI22_X1 port map( A1 => A(26), A2 => n50, B1 => A(25), B2 => n51, ZN 
                           => n122);
   U100 : OAI221_X1 port map( B1 => n45, B2 => n123, C1 => n47, C2 => n124, A 
                           => n125, ZN => n12);
   U101 : AOI22_X1 port map( A1 => A(22), A2 => n50, B1 => A(21), B2 => n51, ZN
                           => n125);
   U102 : INV_X1 port map( A => A(23), ZN => n123);
   U103 : OAI221_X1 port map( B1 => n45, B2 => n126, C1 => n47, C2 => n127, A 
                           => n128, ZN => n10);
   U104 : AOI22_X1 port map( A1 => A(18), A2 => n50, B1 => A(17), B2 => n51, ZN
                           => n128);
   U105 : AOI21_X1 port map( B1 => n72, B2 => n75, A => n118, ZN => n68);
   U106 : OAI222_X1 port map( A1 => n58, A2 => n129, B1 => n56, B2 => n130, C1 
                           => n131, C2 => n132, ZN => n72);
   U107 : AOI221_X1 port map( B1 => n52, B2 => A(15), C1 => n53, C2 => A(16), A
                           => n133, ZN => n100);
   U108 : INV_X1 port map( A => n134, ZN => n133);
   U109 : AOI22_X1 port map( A1 => A(14), A2 => n50, B1 => A(13), B2 => n51, ZN
                           => n134);
   U110 : OAI221_X1 port map( B1 => n135, B2 => n4, C1 => n69, C2 => n2, A => 
                           n136, ZN => B_12_port);
   U111 : AOI222_X1 port map( A1 => n7, A2 => n17, B1 => n9, B2 => n18, C1 => 
                           n11, C2 => n78, ZN => n136);
   U112 : AOI21_X1 port map( B1 => n77, B2 => n75, A => n118, ZN => n69);
   U113 : OAI221_X1 port map( B1 => n44, B2 => n4, C1 => n70, C2 => n2, A => 
                           n137, ZN => B_11_port);
   U114 : AOI222_X1 port map( A1 => n7, A2 => n23, B1 => n9, B2 => n24, C1 => 
                           n11, C2 => n80, ZN => n137);
   U115 : OAI221_X1 port map( B1 => n45, B2 => n138, C1 => n47, C2 => n139, A 
                           => n140, ZN => n80);
   U116 : AOI22_X1 port map( A1 => A(24), A2 => n50, B1 => A(23), B2 => n51, ZN
                           => n140);
   U117 : OAI221_X1 port map( B1 => n127, B2 => n56, C1 => n126, C2 => n58, A 
                           => n141, ZN => n24);
   U118 : AOI22_X1 port map( A1 => A(21), A2 => n52, B1 => A(22), B2 => n53, ZN
                           => n141);
   U119 : OAI221_X1 port map( B1 => n45, B2 => n142, C1 => n47, C2 => n143, A 
                           => n144, ZN => n23);
   U120 : AOI22_X1 port map( A1 => A(16), A2 => n50, B1 => A(15), B2 => n51, ZN
                           => n144);
   U121 : INV_X1 port map( A => A(17), ZN => n142);
   U122 : AOI21_X1 port map( B1 => n79, B2 => n75, A => n118, ZN => n70);
   U123 : OAI21_X1 port map( B1 => n105, B2 => n132, A => n104, ZN => n118);
   U124 : OAI221_X1 port map( B1 => n45, B2 => n129, C1 => n47, C2 => n130, A 
                           => n145, ZN => n79);
   U125 : AOI22_X1 port map( A1 => A(28), A2 => n50, B1 => A(27), B2 => n51, ZN
                           => n145);
   U126 : AOI221_X1 port map( B1 => n52, B2 => A(13), C1 => n53, C2 => A(14), A
                           => n146, ZN => n44);
   U127 : OAI22_X1 port map( A1 => n147, A2 => n56, B1 => n148, B2 => n58, ZN 
                           => n146);
   U128 : INV_X1 port map( A => A(12), ZN => n147);
   U129 : OAI221_X1 port map( B1 => n64, B2 => n4, C1 => n71, C2 => n2, A => 
                           n149, ZN => B_10_port);
   U130 : AOI222_X1 port map( A1 => n7, A2 => n29, B1 => n9, B2 => n30, C1 => 
                           n11, C2 => n82, ZN => n149);
   U131 : OAI221_X1 port map( B1 => n45, B2 => n124, C1 => n47, C2 => n138, A 
                           => n150, ZN => n82);
   U132 : AOI22_X1 port map( A1 => A(23), A2 => n50, B1 => A(22), B2 => n51, ZN
                           => n150);
   U133 : INV_X1 port map( A => A(25), ZN => n138);
   U134 : INV_X1 port map( A => A(24), ZN => n124);
   U135 : OAI221_X1 port map( B1 => n126, B2 => n56, C1 => n143, C2 => n58, A 
                           => n151, ZN => n30);
   U136 : AOI22_X1 port map( A1 => A(20), A2 => n52, B1 => A(21), B2 => n53, ZN
                           => n151);
   U137 : INV_X1 port map( A => n116, ZN => n29);
   U138 : INV_X1 port map( A => n153, ZN => n152);
   U139 : AOI22_X1 port map( A1 => A(15), A2 => n50, B1 => A(14), B2 => n51, ZN
                           => n153);
   U140 : INV_X1 port map( A => n39, ZN => n7);
   U141 : AOI221_X1 port map( B1 => n86, B2 => n73, C1 => n81, C2 => n75, A => 
                           n76, ZN => n71);
   U142 : INV_X1 port map( A => n104, ZN => n76);
   U143 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n104);
   U144 : OAI221_X1 port map( B1 => n45, B2 => n121, C1 => n47, C2 => n129, A 
                           => n154, ZN => n81);
   U145 : AOI22_X1 port map( A1 => A(27), A2 => n50, B1 => A(26), B2 => n51, ZN
                           => n154);
   U146 : INV_X1 port map( A => A(29), ZN => n129);
   U147 : INV_X1 port map( A => A(28), ZN => n121);
   U148 : MUX2_X1 port map( A => A(30), B => A(31), S => n58, Z => n86);
   U149 : OAI22_X1 port map( A1 => n148, A2 => n56, B1 => n96, B2 => n58, ZN =>
                           n155);
   U150 : INV_X1 port map( A => A(10), ZN => n96);
   U151 : INV_X1 port map( A => A(11), ZN => n148);
   U152 : OAI221_X1 port map( B1 => n35, B2 => n39, C1 => n111, C2 => n2, A => 
                           n156, ZN => B_0_port);
   U153 : AOI222_X1 port map( A1 => n11, A2 => n16, B1 => n42, B2 => n157, C1 
                           => n9, C2 => n38, ZN => n156);
   U154 : INV_X1 port map( A => n13, ZN => n38);
   U155 : OAI22_X1 port map( A1 => n97, A2 => n56, B1 => n55, B2 => n58, ZN => 
                           n158);
   U156 : INV_X1 port map( A => A(8), ZN => n55);
   U157 : INV_X1 port map( A => A(9), ZN => n97);
   U158 : AND2_X1 port map( A1 => n159, A2 => n105, ZN => n9);
   U159 : OAI221_X1 port map( B1 => n45, B2 => n160, C1 => n47, C2 => n98, A =>
                           n161, ZN => n157);
   U160 : AOI22_X1 port map( A1 => A(1), A2 => n50, B1 => A(0), B2 => n51, ZN 
                           => n161);
   U161 : INV_X1 port map( A => A(3), ZN => n98);
   U162 : INV_X1 port map( A => A(2), ZN => n160);
   U163 : INV_X1 port map( A => n4, ZN => n42);
   U164 : NAND2_X1 port map( A1 => n75, A2 => n1, ZN => n4);
   U165 : INV_X1 port map( A => n135, ZN => n16);
   U166 : INV_X1 port map( A => n163, ZN => n162);
   U167 : AOI22_X1 port map( A1 => A(13), A2 => n50, B1 => A(12), B2 => n51, ZN
                           => n163);
   U168 : AND2_X1 port map( A1 => SH(2), A2 => n159, ZN => n11);
   U169 : AND2_X1 port map( A1 => SH(3), A2 => n2, ZN => n159);
   U170 : AOI221_X1 port map( B1 => n18, B2 => n73, C1 => n17, C2 => n75, A => 
                           n164, ZN => n111);
   U171 : INV_X1 port map( A => n165, ZN => n164);
   U172 : AOI22_X1 port map( A1 => n106, A2 => n77, B1 => n85, B2 => n78, ZN =>
                           n165);
   U173 : OAI221_X1 port map( B1 => n45, B2 => n139, C1 => n47, C2 => n120, A 
                           => n166, ZN => n78);
   U174 : AOI22_X1 port map( A1 => A(25), A2 => n50, B1 => A(24), B2 => n51, ZN
                           => n166);
   U175 : INV_X1 port map( A => A(27), ZN => n120);
   U176 : INV_X1 port map( A => A(26), ZN => n139);
   U177 : AND2_X1 port map( A1 => SH(3), A2 => n105, ZN => n85);
   U178 : OAI221_X1 port map( B1 => n45, B2 => n130, C1 => n47, C2 => n132, A 
                           => n167, ZN => n77);
   U179 : AOI22_X1 port map( A1 => A(29), A2 => n50, B1 => A(28), B2 => n51, ZN
                           => n167);
   U180 : INV_X1 port map( A => A(31), ZN => n132);
   U181 : INV_X1 port map( A => A(30), ZN => n130);
   U182 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n106);
   U183 : OAI221_X1 port map( B1 => n45, B2 => n143, C1 => n126, C2 => n47, A 
                           => n168, ZN => n17);
   U184 : AOI22_X1 port map( A1 => A(17), A2 => n50, B1 => A(16), B2 => n51, ZN
                           => n168);
   U185 : INV_X1 port map( A => n58, ZN => n51);
   U186 : INV_X1 port map( A => n56, ZN => n50);
   U187 : INV_X1 port map( A => n53, ZN => n47);
   U188 : INV_X1 port map( A => A(19), ZN => n126);
   U189 : INV_X1 port map( A => A(18), ZN => n143);
   U190 : INV_X1 port map( A => n52, ZN => n45);
   U191 : OAI221_X1 port map( B1 => n56, B2 => n169, C1 => n127, C2 => n58, A 
                           => n170, ZN => n18);
   U192 : AOI22_X1 port map( A1 => A(22), A2 => n52, B1 => A(23), B2 => n53, ZN
                           => n170);
   U193 : INV_X1 port map( A => A(20), ZN => n127);
   U194 : INV_X1 port map( A => A(21), ZN => n169);
   U195 : NAND2_X1 port map( A1 => n73, A2 => n1, ZN => n39);
   U196 : NOR2_X1 port map( A1 => n105, A2 => SH(3), ZN => n73);
   U197 : INV_X1 port map( A => SH(2), ZN => n105);
   U198 : OAI22_X1 port map( A1 => n46, A2 => n56, B1 => n65, B2 => n58, ZN => 
                           n171);
   U199 : NAND2_X1 port map( A1 => n172, A2 => n131, ZN => n58);
   U200 : INV_X1 port map( A => A(4), ZN => n65);
   U201 : NAND2_X1 port map( A1 => SH(0), A2 => n131, ZN => n56);
   U202 : INV_X1 port map( A => A(5), ZN => n46);
   U203 : INV_X1 port map( A => SH(0), ZN => n172);
   U204 : INV_X1 port map( A => SH(1), ZN => n131);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW_rash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rash_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163 : std_logic;

begin
   
   U3 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n51);
   U4 : NOR2_X2 port map( A1 => n163, A2 => SH(1), ZN => n50);
   U5 : INV_X1 port map( A => SH(4), ZN => n1);
   U6 : INV_X1 port map( A => SH(4), ZN => n2);
   U7 : OAI221_X1 port map( B1 => n3, B2 => n4, C1 => n5, C2 => n1, A => n6, ZN
                           => B(9));
   U8 : AOI222_X1 port map( A1 => n7, A2 => n8, B1 => n9, B2 => n10, C1 => n11,
                           C2 => n12, ZN => n6);
   U9 : OAI221_X1 port map( B1 => n13, B2 => n4, C1 => n14, C2 => n1, A => n15,
                           ZN => B(8));
   U10 : AOI222_X1 port map( A1 => n7, A2 => n16, B1 => n9, B2 => n17, C1 => 
                           n11, C2 => n18, ZN => n15);
   U11 : OAI221_X1 port map( B1 => n19, B2 => n4, C1 => n20, C2 => n1, A => n21
                           , ZN => B(7));
   U12 : AOI222_X1 port map( A1 => n7, A2 => n22, B1 => n9, B2 => n23, C1 => 
                           n11, C2 => n24, ZN => n21);
   U13 : OAI221_X1 port map( B1 => n25, B2 => n4, C1 => n26, C2 => n1, A => n27
                           , ZN => B(6));
   U14 : AOI222_X1 port map( A1 => n7, A2 => n28, B1 => n9, B2 => n29, C1 => 
                           n11, C2 => n30, ZN => n27);
   U15 : OAI221_X1 port map( B1 => n31, B2 => n4, C1 => n32, C2 => n1, A => n33
                           , ZN => B(5));
   U16 : AOI222_X1 port map( A1 => n7, A2 => n34, B1 => n9, B2 => n8, C1 => n11
                           , C2 => n10, ZN => n33);
   U17 : OAI221_X1 port map( B1 => n35, B2 => n4, C1 => n36, C2 => n1, A => n37
                           , ZN => B(4));
   U18 : AOI222_X1 port map( A1 => n7, A2 => n38, B1 => n9, B2 => n16, C1 => 
                           n11, C2 => n17, ZN => n37);
   U19 : OAI221_X1 port map( B1 => n19, B2 => n39, C1 => n40, C2 => n1, A => 
                           n41, ZN => B(3));
   U20 : AOI222_X1 port map( A1 => n11, A2 => n23, B1 => n42, B2 => n43, C1 => 
                           n9, C2 => n22, ZN => n41);
   U21 : INV_X1 port map( A => n44, ZN => n22);
   U22 : OAI221_X1 port map( B1 => n45, B2 => n46, C1 => n47, C2 => n48, A => 
                           n49, ZN => n43);
   U23 : AOI22_X1 port map( A1 => A(4), A2 => n50, B1 => A(3), B2 => n51, ZN =>
                           n49);
   U24 : AOI221_X1 port map( B1 => n52, B2 => A(10), C1 => n53, C2 => A(9), A 
                           => n54, ZN => n19);
   U25 : OAI22_X1 port map( A1 => n55, A2 => n56, B1 => n57, B2 => n58, ZN => 
                           n54);
   U26 : AND2_X1 port map( A1 => n42, A2 => n59, ZN => B(31));
   U27 : AND2_X1 port map( A1 => n60, A2 => n42, ZN => B(30));
   U28 : OAI221_X1 port map( B1 => n25, B2 => n39, C1 => n61, C2 => n2, A => 
                           n62, ZN => B(2));
   U29 : AOI222_X1 port map( A1 => n11, A2 => n29, B1 => n42, B2 => n63, C1 => 
                           n9, C2 => n28, ZN => n62);
   U30 : INV_X1 port map( A => n64, ZN => n28);
   U31 : OAI221_X1 port map( B1 => n45, B2 => n48, C1 => n47, C2 => n65, A => 
                           n66, ZN => n63);
   U32 : AOI22_X1 port map( A1 => A(3), A2 => n50, B1 => A(2), B2 => n51, ZN =>
                           n66);
   U33 : AOI221_X1 port map( B1 => n52, B2 => A(9), C1 => n53, C2 => A(8), A =>
                           n67, ZN => n25);
   U34 : OAI22_X1 port map( A1 => n57, A2 => n56, B1 => n46, B2 => n58, ZN => 
                           n67);
   U35 : INV_X1 port map( A => A(7), ZN => n57);
   U36 : AND2_X1 port map( A1 => n68, A2 => n42, ZN => B(29));
   U37 : AND2_X1 port map( A1 => n69, A2 => n42, ZN => B(28));
   U38 : NOR3_X1 port map( A1 => n70, A2 => SH(4), A3 => SH(3), ZN => B(27));
   U39 : NOR2_X1 port map( A1 => SH(4), A2 => n71, ZN => B(26));
   U40 : NOR2_X1 port map( A1 => SH(4), A2 => n5, ZN => B(25));
   U41 : AOI22_X1 port map( A1 => n72, A2 => n73, B1 => n68, B2 => n74, ZN => 
                           n5);
   U42 : NOR2_X1 port map( A1 => SH(4), A2 => n14, ZN => B(24));
   U43 : AOI22_X1 port map( A1 => n75, A2 => n73, B1 => n69, B2 => n74, ZN => 
                           n14);
   U44 : NOR2_X1 port map( A1 => SH(4), A2 => n20, ZN => B(23));
   U45 : AOI222_X1 port map( A1 => n76, A2 => n74, B1 => n59, B2 => n77, C1 => 
                           n78, C2 => n73, ZN => n20);
   U46 : NOR2_X1 port map( A1 => SH(4), A2 => n26, ZN => B(22));
   U47 : AOI222_X1 port map( A1 => n79, A2 => n74, B1 => n60, B2 => n77, C1 => 
                           n80, C2 => n73, ZN => n26);
   U48 : NOR2_X1 port map( A1 => SH(4), A2 => n32, ZN => B(21));
   U49 : AOI222_X1 port map( A1 => n72, A2 => n74, B1 => n68, B2 => n77, C1 => 
                           n12, C2 => n73, ZN => n32);
   U50 : NOR2_X1 port map( A1 => SH(4), A2 => n36, ZN => B(20));
   U51 : AOI222_X1 port map( A1 => n75, A2 => n74, B1 => n69, B2 => n77, C1 => 
                           n18, C2 => n73, ZN => n36);
   U52 : OAI221_X1 port map( B1 => n31, B2 => n39, C1 => n81, C2 => n2, A => 
                           n82, ZN => B(1));
   U53 : AOI222_X1 port map( A1 => n11, A2 => n8, B1 => n42, B2 => n83, C1 => 
                           n9, C2 => n34, ZN => n82);
   U54 : INV_X1 port map( A => n3, ZN => n34);
   U55 : AOI221_X1 port map( B1 => n52, B2 => A(12), C1 => n53, C2 => A(11), A 
                           => n84, ZN => n3);
   U56 : OAI22_X1 port map( A1 => n85, A2 => n56, B1 => n86, B2 => n58, ZN => 
                           n84);
   U57 : OAI221_X1 port map( B1 => n45, B2 => n65, C1 => n47, C2 => n87, A => 
                           n88, ZN => n83);
   U58 : AOI22_X1 port map( A1 => A(2), A2 => n50, B1 => A(1), B2 => n51, ZN =>
                           n88);
   U59 : AOI221_X1 port map( B1 => n52, B2 => A(8), C1 => n53, C2 => A(7), A =>
                           n89, ZN => n31);
   U60 : OAI22_X1 port map( A1 => n46, A2 => n56, B1 => n48, B2 => n58, ZN => 
                           n89);
   U61 : INV_X1 port map( A => A(6), ZN => n46);
   U62 : NOR2_X1 port map( A1 => SH(4), A2 => n40, ZN => B(19));
   U63 : AOI222_X1 port map( A1 => n24, A2 => n73, B1 => n78, B2 => n74, C1 => 
                           n90, C2 => SH(3), ZN => n40);
   U64 : NOR2_X1 port map( A1 => SH(4), A2 => n61, ZN => B(18));
   U65 : AOI221_X1 port map( B1 => n80, B2 => n74, C1 => n30, C2 => n73, A => 
                           n91, ZN => n61);
   U66 : INV_X1 port map( A => n92, ZN => n91);
   U67 : AOI22_X1 port map( A1 => n93, A2 => n60, B1 => n77, B2 => n79, ZN => 
                           n92);
   U68 : NOR2_X1 port map( A1 => SH(4), A2 => n81, ZN => B(17));
   U69 : AOI221_X1 port map( B1 => n12, B2 => n74, C1 => n10, C2 => n73, A => 
                           n94, ZN => n81);
   U70 : INV_X1 port map( A => n95, ZN => n94);
   U71 : AOI22_X1 port map( A1 => n93, A2 => n68, B1 => n77, B2 => n72, ZN => 
                           n95);
   U72 : NOR2_X1 port map( A1 => SH(4), A2 => n96, ZN => B(16));
   U73 : OAI221_X1 port map( B1 => n97, B2 => n39, C1 => n98, C2 => n4, A => 
                           n99, ZN => B(15));
   U74 : AOI222_X1 port map( A1 => n11, A2 => n76, B1 => n100, B2 => n59, C1 =>
                           n9, C2 => n78, ZN => n99);
   U75 : INV_X1 port map( A => n24, ZN => n97);
   U76 : OAI221_X1 port map( B1 => n101, B2 => n39, C1 => n102, C2 => n4, A => 
                           n103, ZN => B(14));
   U77 : AOI222_X1 port map( A1 => n11, A2 => n79, B1 => n100, B2 => n60, C1 =>
                           n9, C2 => n80, ZN => n103);
   U78 : INV_X1 port map( A => n29, ZN => n102);
   U79 : INV_X1 port map( A => n30, ZN => n101);
   U80 : OAI221_X1 port map( B1 => n104, B2 => n39, C1 => n105, C2 => n4, A => 
                           n106, ZN => B(13));
   U81 : AOI222_X1 port map( A1 => n11, A2 => n72, B1 => n100, B2 => n68, C1 =>
                           n9, C2 => n12, ZN => n106);
   U82 : OAI221_X1 port map( B1 => n45, B2 => n107, C1 => n47, C2 => n108, A =>
                           n109, ZN => n12);
   U83 : AOI22_X1 port map( A1 => A(22), A2 => n50, B1 => A(21), B2 => n51, ZN 
                           => n109);
   U84 : INV_X1 port map( A => A(23), ZN => n108);
   U85 : OAI222_X1 port map( A1 => n56, A2 => n110, B1 => n47, B2 => n111, C1 
                           => n58, C2 => n112, ZN => n68);
   U86 : OAI221_X1 port map( B1 => n45, B2 => n113, C1 => n47, C2 => n114, A =>
                           n115, ZN => n72);
   U87 : AOI22_X1 port map( A1 => A(26), A2 => n50, B1 => A(25), B2 => n51, ZN 
                           => n115);
   U88 : INV_X1 port map( A => n8, ZN => n105);
   U89 : OAI221_X1 port map( B1 => n45, B2 => n116, C1 => n47, C2 => n117, A =>
                           n118, ZN => n8);
   U90 : AOI22_X1 port map( A1 => A(14), A2 => n50, B1 => A(13), B2 => n51, ZN 
                           => n118);
   U91 : INV_X1 port map( A => n10, ZN => n104);
   U92 : OAI221_X1 port map( B1 => n45, B2 => n119, C1 => n47, C2 => n120, A =>
                           n121, ZN => n10);
   U93 : AOI22_X1 port map( A1 => A(18), A2 => n50, B1 => A(17), B2 => n51, ZN 
                           => n121);
   U94 : INV_X1 port map( A => n122, ZN => B(12));
   U95 : AOI221_X1 port map( B1 => n17, B2 => n7, C1 => n16, C2 => n42, A => 
                           n123, ZN => n122);
   U96 : INV_X1 port map( A => n124, ZN => n123);
   U97 : AOI222_X1 port map( A1 => n11, A2 => n75, B1 => n100, B2 => n69, C1 =>
                           n9, C2 => n18, ZN => n124);
   U98 : NOR2_X1 port map( A1 => n1, A2 => n125, ZN => n100);
   U99 : OAI221_X1 port map( B1 => n98, B2 => n39, C1 => n44, C2 => n4, A => 
                           n126, ZN => B(11));
   U100 : AOI221_X1 port map( B1 => n11, B2 => n78, C1 => n9, C2 => n24, A => 
                           n127, ZN => n126);
   U101 : NOR3_X1 port map( A1 => n1, A2 => SH(3), A3 => n70, ZN => n127);
   U102 : INV_X1 port map( A => n90, ZN => n70);
   U103 : MUX2_X1 port map( A => n76, B => n59, S => SH(2), Z => n90);
   U104 : NOR2_X1 port map( A1 => n111, A2 => n58, ZN => n59);
   U105 : OAI221_X1 port map( B1 => n45, B2 => n110, C1 => n47, C2 => n112, A 
                           => n128, ZN => n76);
   U106 : AOI22_X1 port map( A1 => A(28), A2 => n50, B1 => A(27), B2 => n51, ZN
                           => n128);
   U107 : OAI221_X1 port map( B1 => n119, B2 => n56, C1 => n120, C2 => n58, A 
                           => n129, ZN => n24);
   U108 : AOI22_X1 port map( A1 => A(22), A2 => n52, B1 => A(21), B2 => n53, ZN
                           => n129);
   U109 : OAI221_X1 port map( B1 => n45, B2 => n130, C1 => n47, C2 => n131, A 
                           => n132, ZN => n78);
   U110 : AOI22_X1 port map( A1 => A(24), A2 => n50, B1 => A(23), B2 => n51, ZN
                           => n132);
   U111 : AOI221_X1 port map( B1 => n52, B2 => A(14), C1 => n53, C2 => A(13), A
                           => n133, ZN => n44);
   U112 : OAI22_X1 port map( A1 => n134, A2 => n56, B1 => n135, B2 => n58, ZN 
                           => n133);
   U113 : INV_X1 port map( A => A(12), ZN => n134);
   U114 : INV_X1 port map( A => n23, ZN => n98);
   U115 : OAI221_X1 port map( B1 => n45, B2 => n136, C1 => n47, C2 => n137, A 
                           => n138, ZN => n23);
   U116 : AOI22_X1 port map( A1 => A(16), A2 => n50, B1 => A(15), B2 => n51, ZN
                           => n138);
   U117 : OAI221_X1 port map( B1 => n64, B2 => n4, C1 => n71, C2 => n2, A => 
                           n139, ZN => B(10));
   U118 : AOI222_X1 port map( A1 => n7, A2 => n29, B1 => n9, B2 => n30, C1 => 
                           n11, C2 => n80, ZN => n139);
   U119 : OAI221_X1 port map( B1 => n45, B2 => n131, C1 => n47, C2 => n107, A 
                           => n140, ZN => n80);
   U120 : AOI22_X1 port map( A1 => A(23), A2 => n50, B1 => A(22), B2 => n51, ZN
                           => n140);
   U121 : INV_X1 port map( A => A(24), ZN => n107);
   U122 : INV_X1 port map( A => A(25), ZN => n131);
   U123 : OAI221_X1 port map( B1 => n45, B2 => n141, C1 => n119, C2 => n47, A 
                           => n142, ZN => n30);
   U124 : AOI22_X1 port map( A1 => n50, A2 => A(19), B1 => n51, B2 => A(18), ZN
                           => n142);
   U125 : OAI221_X1 port map( B1 => n45, B2 => n137, C1 => n47, C2 => n116, A 
                           => n143, ZN => n29);
   U126 : AOI22_X1 port map( A1 => A(15), A2 => n50, B1 => A(14), B2 => n51, ZN
                           => n143);
   U127 : INV_X1 port map( A => A(16), ZN => n116);
   U128 : INV_X1 port map( A => A(17), ZN => n137);
   U129 : INV_X1 port map( A => n39, ZN => n7);
   U130 : AOI22_X1 port map( A1 => n79, A2 => n73, B1 => n60, B2 => n74, ZN => 
                           n71);
   U131 : OAI22_X1 port map( A1 => n58, A2 => n110, B1 => n56, B2 => n111, ZN 
                           => n60);
   U132 : OAI221_X1 port map( B1 => n45, B2 => n112, C1 => n47, C2 => n113, A 
                           => n144, ZN => n79);
   U133 : AOI22_X1 port map( A1 => A(27), A2 => n50, B1 => A(26), B2 => n51, ZN
                           => n144);
   U134 : INV_X1 port map( A => A(28), ZN => n113);
   U135 : INV_X1 port map( A => A(29), ZN => n112);
   U136 : AOI221_X1 port map( B1 => n52, B2 => A(13), C1 => n53, C2 => A(12), A
                           => n145, ZN => n64);
   U137 : OAI22_X1 port map( A1 => n135, A2 => n56, B1 => n85, B2 => n58, ZN =>
                           n145);
   U138 : INV_X1 port map( A => A(10), ZN => n85);
   U139 : INV_X1 port map( A => A(11), ZN => n135);
   U140 : OAI221_X1 port map( B1 => n35, B2 => n39, C1 => n96, C2 => n1, A => 
                           n146, ZN => B(0));
   U141 : AOI222_X1 port map( A1 => n11, A2 => n16, B1 => n42, B2 => n147, C1 
                           => n9, C2 => n38, ZN => n146);
   U142 : INV_X1 port map( A => n13, ZN => n38);
   U143 : AOI221_X1 port map( B1 => n52, B2 => A(11), C1 => n53, C2 => A(10), A
                           => n148, ZN => n13);
   U144 : OAI22_X1 port map( A1 => n86, A2 => n56, B1 => n55, B2 => n58, ZN => 
                           n148);
   U145 : INV_X1 port map( A => A(8), ZN => n55);
   U146 : INV_X1 port map( A => A(9), ZN => n86);
   U147 : AND2_X1 port map( A1 => n149, A2 => n150, ZN => n9);
   U148 : OAI221_X1 port map( B1 => n45, B2 => n87, C1 => n47, C2 => n151, A =>
                           n152, ZN => n147);
   U149 : AOI22_X1 port map( A1 => A(1), A2 => n50, B1 => A(0), B2 => n51, ZN 
                           => n152);
   U150 : INV_X1 port map( A => A(2), ZN => n151);
   U151 : INV_X1 port map( A => A(3), ZN => n87);
   U152 : INV_X1 port map( A => n4, ZN => n42);
   U153 : NAND2_X1 port map( A1 => n73, A2 => n1, ZN => n4);
   U154 : OAI221_X1 port map( B1 => n45, B2 => n117, C1 => n47, C2 => n153, A 
                           => n154, ZN => n16);
   U155 : AOI22_X1 port map( A1 => A(13), A2 => n50, B1 => A(12), B2 => n51, ZN
                           => n154);
   U156 : INV_X1 port map( A => A(14), ZN => n153);
   U157 : INV_X1 port map( A => A(15), ZN => n117);
   U158 : AND2_X1 port map( A1 => SH(2), A2 => n149, ZN => n11);
   U159 : NOR2_X1 port map( A1 => n155, A2 => SH(4), ZN => n149);
   U160 : AOI221_X1 port map( B1 => n18, B2 => n74, C1 => n17, C2 => n73, A => 
                           n156, ZN => n96);
   U161 : INV_X1 port map( A => n157, ZN => n156);
   U162 : AOI22_X1 port map( A1 => n93, A2 => n69, B1 => n77, B2 => n75, ZN => 
                           n157);
   U163 : OAI221_X1 port map( B1 => n45, B2 => n114, C1 => n47, C2 => n130, A 
                           => n158, ZN => n75);
   U164 : AOI22_X1 port map( A1 => A(25), A2 => n50, B1 => A(24), B2 => n51, ZN
                           => n158);
   U165 : INV_X1 port map( A => A(26), ZN => n130);
   U166 : INV_X1 port map( A => A(27), ZN => n114);
   U167 : NOR2_X1 port map( A1 => n155, A2 => SH(2), ZN => n77);
   U168 : OAI221_X1 port map( B1 => n45, B2 => n111, C1 => n47, C2 => n110, A 
                           => n159, ZN => n69);
   U169 : AOI22_X1 port map( A1 => A(29), A2 => n50, B1 => A(28), B2 => n51, ZN
                           => n159);
   U170 : INV_X1 port map( A => A(30), ZN => n110);
   U171 : INV_X1 port map( A => A(31), ZN => n111);
   U172 : NOR2_X1 port map( A1 => n150, A2 => n155, ZN => n93);
   U173 : INV_X1 port map( A => n125, ZN => n73);
   U174 : NAND2_X1 port map( A1 => n150, A2 => n155, ZN => n125);
   U175 : INV_X1 port map( A => SH(3), ZN => n155);
   U176 : OAI221_X1 port map( B1 => n45, B2 => n120, C1 => n47, C2 => n136, A 
                           => n160, ZN => n17);
   U177 : AOI22_X1 port map( A1 => A(17), A2 => n50, B1 => A(16), B2 => n51, ZN
                           => n160);
   U178 : INV_X1 port map( A => A(18), ZN => n136);
   U179 : INV_X1 port map( A => A(19), ZN => n120);
   U180 : OAI221_X1 port map( B1 => n56, B2 => n141, C1 => n119, C2 => n58, A 
                           => n161, ZN => n18);
   U181 : AOI22_X1 port map( A1 => A(23), A2 => n52, B1 => A(22), B2 => n53, ZN
                           => n161);
   U182 : INV_X1 port map( A => A(20), ZN => n119);
   U183 : INV_X1 port map( A => A(21), ZN => n141);
   U184 : NAND2_X1 port map( A1 => n74, A2 => n1, ZN => n39);
   U185 : NOR2_X1 port map( A1 => n150, A2 => SH(3), ZN => n74);
   U186 : INV_X1 port map( A => SH(2), ZN => n150);
   U187 : AOI221_X1 port map( B1 => n52, B2 => A(7), C1 => n53, C2 => A(6), A 
                           => n162, ZN => n35);
   U188 : OAI22_X1 port map( A1 => n48, A2 => n56, B1 => n65, B2 => n58, ZN => 
                           n162);
   U189 : INV_X1 port map( A => n51, ZN => n58);
   U190 : INV_X1 port map( A => A(4), ZN => n65);
   U191 : INV_X1 port map( A => n50, ZN => n56);
   U192 : INV_X1 port map( A => A(5), ZN => n48);
   U193 : INV_X1 port map( A => n47, ZN => n53);
   U194 : NAND2_X1 port map( A1 => SH(1), A2 => n163, ZN => n47);
   U195 : INV_X1 port map( A => SH(0), ZN => n163);
   U196 : INV_X1 port map( A => n45, ZN => n52);
   U197 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n45);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_sla_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sla_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sla_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178 : std_logic;

begin
   B <= ( B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, A(0) );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n76);
   U3 : NAND2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n27);
   U4 : OAI221_X4 port map( B1 => n25, B2 => n169, C1 => n27, C2 => n152, A => 
                           n176, ZN => n102);
   U5 : OAI221_X4 port map( B1 => n25, B2 => n164, C1 => n27, C2 => n171, A => 
                           n172, ZN => n97);
   U6 : OAI221_X4 port map( B1 => n25, B2 => n162, C1 => n27, C2 => n169, A => 
                           n170, ZN => n95);
   U7 : OAI221_X4 port map( B1 => n25, B2 => n153, C1 => n27, C2 => n164, A => 
                           n165, ZN => n88);
   U8 : OAI221_X4 port map( B1 => n25, B2 => n150, C1 => n27, C2 => n162, A => 
                           n163, ZN => n86);
   U9 : NAND2_X2 port map( A1 => SH(1), A2 => n178, ZN => n25);
   U10 : INV_X1 port map( A => n31, ZN => n1);
   U11 : INV_X2 port map( A => n1, ZN => n2);
   U12 : INV_X1 port map( A => n30, ZN => n3);
   U13 : INV_X2 port map( A => n3, ZN => n4);
   U14 : INV_X1 port map( A => SH(4), ZN => n5);
   U15 : INV_X1 port map( A => SH(4), ZN => n6);
   U16 : OAI21_X1 port map( B1 => SH(4), B2 => n7, A => n8, ZN => B_9_port);
   U17 : OAI21_X1 port map( B1 => SH(4), B2 => n9, A => n8, ZN => B_8_port);
   U18 : OAI21_X1 port map( B1 => SH(4), B2 => n10, A => n8, ZN => B_7_port);
   U19 : OAI21_X1 port map( B1 => SH(4), B2 => n11, A => n8, ZN => B_6_port);
   U20 : OAI21_X1 port map( B1 => SH(4), B2 => n12, A => n8, ZN => B_5_port);
   U21 : OAI21_X1 port map( B1 => SH(4), B2 => n13, A => n8, ZN => B_4_port);
   U22 : OAI21_X1 port map( B1 => SH(4), B2 => n14, A => n8, ZN => B_3_port);
   U23 : OAI221_X1 port map( B1 => n15, B2 => n16, C1 => n17, C2 => n5, A => 
                           n18, ZN => B_31_port);
   U24 : AOI222_X1 port map( A1 => n19, A2 => n20, B1 => n21, B2 => n22, C1 => 
                           n23, C2 => n24, ZN => n18);
   U25 : OAI221_X1 port map( B1 => n25, B2 => n26, C1 => n27, C2 => n28, A => 
                           n29, ZN => n22);
   U26 : AOI22_X1 port map( A1 => A(30), A2 => n4, B1 => A(31), B2 => n2, ZN =>
                           n29);
   U27 : INV_X1 port map( A => A(29), ZN => n26);
   U28 : OAI221_X1 port map( B1 => n32, B2 => n16, C1 => n33, C2 => n5, A => 
                           n34, ZN => B_30_port);
   U29 : AOI222_X1 port map( A1 => n19, A2 => n35, B1 => n21, B2 => n36, C1 => 
                           n23, C2 => n37, ZN => n34);
   U30 : OAI221_X1 port map( B1 => n25, B2 => n28, C1 => n27, C2 => n38, A => 
                           n39, ZN => n36);
   U31 : AOI22_X1 port map( A1 => A(29), A2 => n4, B1 => A(30), B2 => n2, ZN =>
                           n39);
   U32 : INV_X1 port map( A => A(28), ZN => n28);
   U33 : OAI21_X1 port map( B1 => SH(4), B2 => n40, A => n8, ZN => B_2_port);
   U34 : OAI221_X1 port map( B1 => n41, B2 => n16, C1 => n42, C2 => n5, A => 
                           n43, ZN => B_29_port);
   U35 : AOI222_X1 port map( A1 => n19, A2 => n44, B1 => n21, B2 => n45, C1 => 
                           n23, C2 => n46, ZN => n43);
   U36 : OAI221_X1 port map( B1 => n25, B2 => n38, C1 => n27, C2 => n47, A => 
                           n48, ZN => n45);
   U37 : AOI22_X1 port map( A1 => A(28), A2 => n4, B1 => A(29), B2 => n2, ZN =>
                           n48);
   U38 : INV_X1 port map( A => A(27), ZN => n38);
   U39 : OAI221_X1 port map( B1 => n49, B2 => n16, C1 => n50, C2 => n5, A => 
                           n51, ZN => B_28_port);
   U40 : AOI222_X1 port map( A1 => n19, A2 => n52, B1 => n21, B2 => n53, C1 => 
                           n23, C2 => n54, ZN => n51);
   U41 : OAI221_X1 port map( B1 => n25, B2 => n47, C1 => n27, C2 => n55, A => 
                           n56, ZN => n53);
   U42 : AOI22_X1 port map( A1 => A(27), A2 => n4, B1 => A(28), B2 => n2, ZN =>
                           n56);
   U43 : INV_X1 port map( A => A(26), ZN => n47);
   U44 : INV_X1 port map( A => n57, ZN => n21);
   U45 : OAI221_X1 port map( B1 => n15, B2 => n57, C1 => n58, C2 => n5, A => 
                           n59, ZN => B_27_port);
   U46 : AOI222_X1 port map( A1 => n60, A2 => n24, B1 => n23, B2 => n20, C1 => 
                           n19, C2 => n61, ZN => n59);
   U47 : INV_X1 port map( A => n62, ZN => n15);
   U48 : OAI221_X1 port map( B1 => n25, B2 => n55, C1 => n27, C2 => n63, A => 
                           n64, ZN => n62);
   U49 : AOI22_X1 port map( A1 => A(26), A2 => n4, B1 => A(27), B2 => n2, ZN =>
                           n64);
   U50 : INV_X1 port map( A => A(25), ZN => n55);
   U51 : OAI221_X1 port map( B1 => n32, B2 => n57, C1 => n65, C2 => n5, A => 
                           n66, ZN => B_26_port);
   U52 : AOI222_X1 port map( A1 => n60, A2 => n37, B1 => n23, B2 => n35, C1 => 
                           n19, C2 => n67, ZN => n66);
   U53 : INV_X1 port map( A => n68, ZN => n32);
   U54 : OAI221_X1 port map( B1 => n25, B2 => n63, C1 => n27, C2 => n69, A => 
                           n70, ZN => n68);
   U55 : AOI22_X1 port map( A1 => A(25), A2 => n4, B1 => A(26), B2 => n2, ZN =>
                           n70);
   U56 : INV_X1 port map( A => A(24), ZN => n63);
   U57 : OAI221_X1 port map( B1 => n41, B2 => n57, C1 => n7, C2 => n5, A => n71
                           , ZN => B_25_port);
   U58 : AOI222_X1 port map( A1 => n60, A2 => n46, B1 => n23, B2 => n44, C1 => 
                           n19, C2 => n72, ZN => n71);
   U59 : AOI221_X1 port map( B1 => n73, B2 => n74, C1 => n75, C2 => n76, A => 
                           n77, ZN => n7);
   U60 : INV_X1 port map( A => n78, ZN => n77);
   U61 : AOI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => n78);
   U62 : INV_X1 port map( A => n82, ZN => n41);
   U63 : OAI221_X1 port map( B1 => n25, B2 => n69, C1 => n27, C2 => n83, A => 
                           n84, ZN => n82);
   U64 : AOI22_X1 port map( A1 => A(24), A2 => n4, B1 => A(25), B2 => n2, ZN =>
                           n84);
   U65 : INV_X1 port map( A => A(23), ZN => n69);
   U66 : OAI221_X1 port map( B1 => n49, B2 => n57, C1 => n9, C2 => n5, A => n85
                           , ZN => B_24_port);
   U67 : AOI222_X1 port map( A1 => n60, A2 => n54, B1 => n23, B2 => n52, C1 => 
                           n19, C2 => n86, ZN => n85);
   U68 : AOI221_X1 port map( B1 => n87, B2 => n74, C1 => n88, C2 => n76, A => 
                           n89, ZN => n9);
   U69 : INV_X1 port map( A => n90, ZN => n49);
   U70 : OAI221_X1 port map( B1 => n25, B2 => n83, C1 => n27, C2 => n91, A => 
                           n92, ZN => n90);
   U71 : AOI22_X1 port map( A1 => A(23), A2 => n4, B1 => A(24), B2 => n2, ZN =>
                           n92);
   U72 : INV_X1 port map( A => A(22), ZN => n83);
   U73 : OAI221_X1 port map( B1 => n93, B2 => n57, C1 => n10, C2 => n5, A => 
                           n94, ZN => B_23_port);
   U74 : AOI222_X1 port map( A1 => n60, A2 => n20, B1 => n23, B2 => n61, C1 => 
                           n19, C2 => n95, ZN => n94);
   U75 : AOI221_X1 port map( B1 => n96, B2 => n74, C1 => n97, C2 => n76, A => 
                           n89, ZN => n10);
   U76 : INV_X1 port map( A => n24, ZN => n93);
   U77 : OAI221_X1 port map( B1 => n25, B2 => n91, C1 => n27, C2 => n98, A => 
                           n99, ZN => n24);
   U78 : AOI22_X1 port map( A1 => A(22), A2 => n4, B1 => A(23), B2 => n2, ZN =>
                           n99);
   U79 : INV_X1 port map( A => A(21), ZN => n91);
   U80 : OAI221_X1 port map( B1 => n100, B2 => n57, C1 => n11, C2 => n5, A => 
                           n101, ZN => B_22_port);
   U81 : AOI222_X1 port map( A1 => n60, A2 => n35, B1 => n23, B2 => n67, C1 => 
                           n19, C2 => n102, ZN => n101);
   U82 : AOI221_X1 port map( B1 => n103, B2 => n74, C1 => n104, C2 => n76, A =>
                           n89, ZN => n11);
   U83 : INV_X1 port map( A => n37, ZN => n100);
   U84 : OAI221_X1 port map( B1 => n25, B2 => n98, C1 => n27, C2 => n105, A => 
                           n106, ZN => n37);
   U85 : AOI22_X1 port map( A1 => A(21), A2 => n4, B1 => A(22), B2 => n2, ZN =>
                           n106);
   U86 : INV_X1 port map( A => A(20), ZN => n98);
   U87 : OAI221_X1 port map( B1 => n107, B2 => n57, C1 => n12, C2 => n6, A => 
                           n108, ZN => B_21_port);
   U88 : AOI222_X1 port map( A1 => n60, A2 => n44, B1 => n23, B2 => n72, C1 => 
                           n19, C2 => n75, ZN => n108);
   U89 : AOI221_X1 port map( B1 => n80, B2 => n74, C1 => n73, C2 => n76, A => 
                           n89, ZN => n12);
   U90 : INV_X1 port map( A => n109, ZN => n89);
   U91 : INV_X1 port map( A => n46, ZN => n107);
   U92 : OAI221_X1 port map( B1 => n25, B2 => n105, C1 => n27, C2 => n110, A =>
                           n111, ZN => n46);
   U93 : AOI22_X1 port map( A1 => A(20), A2 => n4, B1 => A(21), B2 => n2, ZN =>
                           n111);
   U94 : INV_X1 port map( A => A(19), ZN => n105);
   U95 : OAI221_X1 port map( B1 => n112, B2 => n57, C1 => n13, C2 => n6, A => 
                           n113, ZN => B_20_port);
   U96 : AOI222_X1 port map( A1 => n60, A2 => n52, B1 => n23, B2 => n86, C1 => 
                           n19, C2 => n88, ZN => n113);
   U97 : AOI21_X1 port map( B1 => n87, B2 => n76, A => n114, ZN => n13);
   U98 : INV_X1 port map( A => n54, ZN => n112);
   U99 : OAI221_X1 port map( B1 => n25, B2 => n110, C1 => n27, C2 => n115, A =>
                           n116, ZN => n54);
   U100 : AOI22_X1 port map( A1 => A(19), A2 => n4, B1 => A(20), B2 => n2, ZN 
                           => n116);
   U101 : INV_X1 port map( A => A(18), ZN => n110);
   U102 : OAI21_X1 port map( B1 => SH(4), B2 => n117, A => n8, ZN => B_1_port);
   U103 : OAI221_X1 port map( B1 => n118, B2 => n57, C1 => n14, C2 => n6, A => 
                           n119, ZN => B_19_port);
   U104 : AOI222_X1 port map( A1 => n60, A2 => n61, B1 => n23, B2 => n95, C1 =>
                           n19, C2 => n97, ZN => n119);
   U105 : AOI21_X1 port map( B1 => n96, B2 => n76, A => n114, ZN => n14);
   U106 : INV_X1 port map( A => n20, ZN => n118);
   U107 : OAI221_X1 port map( B1 => n25, B2 => n115, C1 => n27, C2 => n120, A 
                           => n121, ZN => n20);
   U108 : AOI22_X1 port map( A1 => A(18), A2 => n4, B1 => A(19), B2 => n2, ZN 
                           => n121);
   U109 : INV_X1 port map( A => A(17), ZN => n115);
   U110 : OAI221_X1 port map( B1 => n122, B2 => n57, C1 => n40, C2 => n6, A => 
                           n123, ZN => B_18_port);
   U111 : AOI222_X1 port map( A1 => n60, A2 => n67, B1 => n23, B2 => n102, C1 
                           => n19, C2 => n104, ZN => n123);
   U112 : AOI21_X1 port map( B1 => n103, B2 => n76, A => n114, ZN => n40);
   U113 : INV_X1 port map( A => n35, ZN => n122);
   U114 : OAI221_X1 port map( B1 => n25, B2 => n120, C1 => n27, C2 => n124, A 
                           => n125, ZN => n35);
   U115 : AOI22_X1 port map( A1 => A(17), A2 => n4, B1 => A(18), B2 => n2, ZN 
                           => n125);
   U116 : INV_X1 port map( A => A(16), ZN => n120);
   U117 : OAI221_X1 port map( B1 => n126, B2 => n57, C1 => n117, C2 => n6, A =>
                           n127, ZN => B_17_port);
   U118 : AOI222_X1 port map( A1 => n60, A2 => n72, B1 => n23, B2 => n75, C1 =>
                           n19, C2 => n73, ZN => n127);
   U119 : INV_X1 port map( A => n16, ZN => n60);
   U120 : AOI21_X1 port map( B1 => n80, B2 => n76, A => n114, ZN => n117);
   U121 : OAI21_X1 port map( B1 => n128, B2 => n129, A => n109, ZN => n114);
   U122 : INV_X1 port map( A => n44, ZN => n126);
   U123 : OAI221_X1 port map( B1 => n25, B2 => n124, C1 => n27, C2 => n130, A 
                           => n131, ZN => n44);
   U124 : AOI22_X1 port map( A1 => A(16), A2 => n4, B1 => A(17), B2 => n2, ZN 
                           => n131);
   U125 : INV_X1 port map( A => A(15), ZN => n124);
   U126 : OAI221_X1 port map( B1 => n132, B2 => n16, C1 => n133, C2 => n57, A 
                           => n134, ZN => B_16_port);
   U127 : AOI221_X1 port map( B1 => n19, B2 => n87, C1 => n23, C2 => n88, A => 
                           n135, ZN => n134);
   U128 : INV_X1 port map( A => n8, ZN => n135);
   U129 : AND2_X1 port map( A1 => n136, A2 => n129, ZN => n23);
   U130 : AND2_X1 port map( A1 => n136, A2 => SH(2), ZN => n19);
   U131 : AND2_X1 port map( A1 => SH(3), A2 => n6, ZN => n136);
   U132 : NAND2_X1 port map( A1 => n76, A2 => n5, ZN => n57);
   U133 : INV_X1 port map( A => n52, ZN => n133);
   U134 : OAI221_X1 port map( B1 => n25, B2 => n130, C1 => n27, C2 => n137, A 
                           => n138, ZN => n52);
   U135 : AOI22_X1 port map( A1 => A(15), A2 => n4, B1 => A(16), B2 => n2, ZN 
                           => n138);
   U136 : INV_X1 port map( A => A(14), ZN => n130);
   U137 : NAND2_X1 port map( A1 => n74, A2 => n5, ZN => n16);
   U138 : INV_X1 port map( A => n86, ZN => n132);
   U139 : OAI21_X1 port map( B1 => SH(4), B2 => n17, A => n8, ZN => B_15_port);
   U140 : AOI221_X1 port map( B1 => n95, B2 => n74, C1 => n61, C2 => n76, A => 
                           n139, ZN => n17);
   U141 : INV_X1 port map( A => n140, ZN => n139);
   U142 : AOI22_X1 port map( A1 => n141, A2 => n96, B1 => n79, B2 => n97, ZN =>
                           n140);
   U143 : OAI221_X1 port map( B1 => n25, B2 => n137, C1 => n27, C2 => n142, A 
                           => n143, ZN => n61);
   U144 : AOI22_X1 port map( A1 => A(14), A2 => n4, B1 => A(15), B2 => n2, ZN 
                           => n143);
   U145 : INV_X1 port map( A => A(13), ZN => n137);
   U146 : OAI21_X1 port map( B1 => SH(4), B2 => n33, A => n8, ZN => B_14_port);
   U147 : AOI221_X1 port map( B1 => n102, B2 => n74, C1 => n67, C2 => n76, A =>
                           n144, ZN => n33);
   U148 : INV_X1 port map( A => n145, ZN => n144);
   U149 : AOI22_X1 port map( A1 => n141, A2 => n103, B1 => n79, B2 => n104, ZN 
                           => n145);
   U150 : OAI221_X1 port map( B1 => n25, B2 => n142, C1 => n27, C2 => n146, A 
                           => n147, ZN => n67);
   U151 : AOI22_X1 port map( A1 => A(13), A2 => n4, B1 => A(14), B2 => n2, ZN 
                           => n147);
   U152 : INV_X1 port map( A => A(12), ZN => n142);
   U153 : OAI21_X1 port map( B1 => SH(4), B2 => n42, A => n8, ZN => B_13_port);
   U154 : AOI221_X1 port map( B1 => n80, B2 => n141, C1 => n73, C2 => n79, A =>
                           n148, ZN => n42);
   U155 : INV_X1 port map( A => n149, ZN => n148);
   U156 : AOI22_X1 port map( A1 => n74, A2 => n75, B1 => n76, B2 => n72, ZN => 
                           n149);
   U157 : OAI221_X1 port map( B1 => n25, B2 => n146, C1 => n27, C2 => n150, A 
                           => n151, ZN => n72);
   U158 : AOI22_X1 port map( A1 => A(12), A2 => n4, B1 => A(13), B2 => n2, ZN 
                           => n151);
   U159 : INV_X1 port map( A => A(11), ZN => n146);
   U160 : OAI221_X1 port map( B1 => n25, B2 => n152, C1 => n27, C2 => n153, A 
                           => n154, ZN => n75);
   U161 : AOI22_X1 port map( A1 => A(8), A2 => n4, B1 => A(9), B2 => n2, ZN => 
                           n154);
   U162 : OAI221_X1 port map( B1 => n25, B2 => n155, C1 => n27, C2 => n156, A 
                           => n157, ZN => n73);
   U163 : AOI22_X1 port map( A1 => A(4), A2 => n4, B1 => A(5), B2 => n2, ZN => 
                           n157);
   U164 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n141);
   U165 : MUX2_X1 port map( A => A(0), B => A(1), S => n2, Z => n80);
   U166 : OAI21_X1 port map( B1 => SH(4), B2 => n50, A => n8, ZN => B_12_port);
   U167 : AOI221_X1 port map( B1 => n88, B2 => n74, C1 => n86, C2 => n76, A => 
                           n158, ZN => n50);
   U168 : INV_X1 port map( A => n159, ZN => n158);
   U169 : AOI21_X1 port map( B1 => n79, B2 => n87, A => n81, ZN => n159);
   U170 : OAI221_X1 port map( B1 => n25, B2 => n156, C1 => n160, C2 => n27, A 
                           => n161, ZN => n87);
   U171 : AOI22_X1 port map( A1 => n4, A2 => A(3), B1 => A(4), B2 => n2, ZN => 
                           n161);
   U172 : INV_X1 port map( A => A(2), ZN => n156);
   U173 : AOI22_X1 port map( A1 => A(11), A2 => n4, B1 => A(12), B2 => n2, ZN 
                           => n163);
   U174 : INV_X1 port map( A => A(10), ZN => n150);
   U175 : AOI22_X1 port map( A1 => A(7), A2 => n4, B1 => A(8), B2 => n2, ZN => 
                           n165);
   U176 : INV_X1 port map( A => A(6), ZN => n153);
   U177 : OAI21_X1 port map( B1 => SH(4), B2 => n58, A => n8, ZN => B_11_port);
   U178 : AOI221_X1 port map( B1 => n97, B2 => n74, C1 => n95, C2 => n76, A => 
                           n166, ZN => n58);
   U179 : INV_X1 port map( A => n167, ZN => n166);
   U180 : AOI21_X1 port map( B1 => n79, B2 => n96, A => n81, ZN => n167);
   U181 : OAI221_X1 port map( B1 => n160, B2 => n25, C1 => n128, C2 => n27, A 
                           => n168, ZN => n96);
   U182 : AOI22_X1 port map( A1 => n4, A2 => A(2), B1 => A(3), B2 => n2, ZN => 
                           n168);
   U183 : INV_X1 port map( A => A(0), ZN => n128);
   U184 : INV_X1 port map( A => A(1), ZN => n160);
   U185 : AOI22_X1 port map( A1 => A(10), A2 => n4, B1 => A(11), B2 => n2, ZN 
                           => n170);
   U186 : INV_X1 port map( A => A(9), ZN => n162);
   U187 : AOI22_X1 port map( A1 => A(6), A2 => n4, B1 => A(7), B2 => n2, ZN => 
                           n172);
   U188 : INV_X1 port map( A => A(5), ZN => n164);
   U189 : OAI21_X1 port map( B1 => SH(4), B2 => n65, A => n8, ZN => B_10_port);
   U190 : NAND2_X1 port map( A1 => SH(4), A2 => A(0), ZN => n8);
   U191 : AOI221_X1 port map( B1 => n104, B2 => n74, C1 => n102, C2 => n76, A 
                           => n173, ZN => n65);
   U192 : INV_X1 port map( A => n174, ZN => n173);
   U193 : AOI21_X1 port map( B1 => n79, B2 => n103, A => n81, ZN => n174);
   U194 : NOR2_X1 port map( A1 => n129, A2 => n109, ZN => n81);
   U195 : NAND2_X1 port map( A1 => SH(3), A2 => A(0), ZN => n109);
   U196 : INV_X1 port map( A => n175, ZN => n103);
   U197 : AOI222_X1 port map( A1 => n2, A2 => A(2), B1 => A(1), B2 => n4, C1 =>
                           A(0), C2 => SH(1), ZN => n175);
   U198 : AND2_X1 port map( A1 => SH(3), A2 => n129, ZN => n79);
   U199 : AOI22_X1 port map( A1 => A(9), A2 => n4, B1 => A(10), B2 => n2, ZN =>
                           n176);
   U200 : INV_X1 port map( A => A(7), ZN => n152);
   U201 : INV_X1 port map( A => A(8), ZN => n169);
   U202 : NOR2_X1 port map( A1 => n129, A2 => SH(3), ZN => n74);
   U203 : INV_X1 port map( A => SH(2), ZN => n129);
   U204 : OAI221_X1 port map( B1 => n25, B2 => n171, C1 => n155, C2 => n27, A 
                           => n177, ZN => n104);
   U205 : AOI22_X1 port map( A1 => A(5), A2 => n4, B1 => A(6), B2 => n2, ZN => 
                           n177);
   U206 : NOR2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n31);
   U207 : NOR2_X1 port map( A1 => n178, A2 => SH(1), ZN => n30);
   U208 : INV_X1 port map( A => A(3), ZN => n155);
   U209 : INV_X1 port map( A => A(4), ZN => n171);
   U210 : INV_X1 port map( A => SH(0), ZN => n178);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW01_ash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW01_ash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal SHMAG_3_port, SHMAG_2_port, SHMAG_1_port, SHMAG_0_port, 
      ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, ML_int_1_28_port, 
      ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, ML_int_1_24_port, 
      ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, ML_int_1_20_port, 
      ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, ML_int_1_16_port, 
      ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, ML_int_1_12_port, 
      ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, ML_int_1_8_port, 
      ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, ML_int_1_4_port, 
      ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, ML_int_1_0_port, 
      ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, ML_int_2_28_port, 
      ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, ML_int_2_24_port, 
      ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, ML_int_2_20_port, 
      ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, ML_int_2_16_port, 
      ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, ML_int_2_12_port, 
      ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, ML_int_2_8_port, 
      ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, ML_int_2_4_port, 
      ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, ML_int_2_0_port, 
      ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, ML_int_3_28_port, 
      ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, ML_int_3_24_port, 
      ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, ML_int_3_20_port, 
      ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, ML_int_3_16_port, 
      ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, ML_int_3_12_port, 
      ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, ML_int_3_8_port, 
      ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, ML_int_3_4_port, 
      ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, ML_int_3_0_port, 
      ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, ML_int_4_28_port, 
      ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, ML_int_4_24_port, 
      ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, ML_int_4_20_port, 
      ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, ML_int_4_16_port, 
      ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, ML_int_4_12_port, 
      ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, ML_int_4_8_port, 
      ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, ML_int_4_4_port, 
      ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, ML_int_4_0_port, n1, 
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n1, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n1, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n1, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n1, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n1, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n1, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n1, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n1, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n1, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n1, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n1, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n1, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n2, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n2, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n2, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n2, Z => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => SH(3), Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => SH(3), Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => SH(3), Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => SH(3), Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => SH(3), Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => SH(3), Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => SH(3), Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => SH(3), Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => SH(3), Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => SH(3), Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => SH(3), Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => SH(3), Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => SH(3), Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => SH(3), Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => SH(3), Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => SH(3), Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => SH(3), Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => SH(3), Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => SH(3), Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => SH(3), Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           SH(3), Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           SH(3), Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => SH(2), Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => SH(2), Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => SH(2), Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => SH(2), Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => SH(2), Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => SH(2), Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => SH(2), Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => SH(2), Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => SH(2), Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => SH(2), Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => SH(2), Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => SH(2), Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => SH(2), Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => SH(2), Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => SH(2), Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => SH(2), Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => SH(2), Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => SH(2), Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           SH(2), Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           SH(2), Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           SH(2), Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           SH(2), Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           SH(2), Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           SH(2), Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => SH(1), Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => SH(1), Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => SH(1), Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => SH(1), Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => SH(1), Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => SH(1), Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => SH(1), Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => SH(1), Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => SH(1), Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => SH(1), Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           SH(1), Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           SH(1), Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           SH(1), Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           SH(1), Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           SH(1), Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           SH(1), Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           SH(1), Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           SH(1), Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => SH(0), Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => SH(0), Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => SH(0), Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => SH(0), Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => SH(0), Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => SH(0), Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => SH(0), Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => SH(0), Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => SH(0), Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => SH(0), Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => SH(0), Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => SH(0), Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => SH(0), Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => SH(0), Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => SH(0), Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => SH(0), Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => SH(0), Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => SH(0), Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => SH(0), Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => SH(0), Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => SH(0), Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => SH(0), Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => SH(0), Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => SH(0), Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => SH(0), Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => SH(0), Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => SH(0), Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => SH(0), Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => SH(0), Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => SH(0), Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => SH(0), Z => 
                           ML_int_1_1_port);
   U3 : INV_X1 port map( A => n3, ZN => n1);
   U4 : INV_X1 port map( A => n3, ZN => n2);
   U5 : INV_X1 port map( A => SH(4), ZN => n3);
   U6 : INV_X1 port map( A => SH(4), ZN => n4);
   U7 : INV_X1 port map( A => SH(4), ZN => n5);
   U8 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n5, ZN => B(9));
   U9 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n5, ZN => B(8));
   U10 : NOR2_X1 port map( A1 => n2, A2 => n6, ZN => B(7));
   U11 : NOR2_X1 port map( A1 => n2, A2 => n7, ZN => B(6));
   U12 : NOR2_X1 port map( A1 => n2, A2 => n8, ZN => B(5));
   U13 : NOR2_X1 port map( A1 => n2, A2 => n9, ZN => B(4));
   U14 : NOR2_X1 port map( A1 => n2, A2 => n10, ZN => B(3));
   U15 : NOR2_X1 port map( A1 => n2, A2 => n11, ZN => B(2));
   U16 : NOR2_X1 port map( A1 => n2, A2 => n12, ZN => B(1));
   U17 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n5, ZN => B(15));
   U18 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n4, ZN => B(14));
   U19 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n4, ZN => B(13));
   U20 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n4, ZN => B(12));
   U21 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n4, ZN => B(11));
   U22 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n3, ZN => B(10));
   U23 : NOR2_X1 port map( A1 => n2, A2 => n13, ZN => B(0));
   U24 : INV_X1 port map( A => n6, ZN => ML_int_4_7_port);
   U25 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => SHMAG_3_port, ZN => n6
                           );
   U26 : INV_X1 port map( A => n7, ZN => ML_int_4_6_port);
   U27 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => SHMAG_3_port, ZN => n7
                           );
   U28 : INV_X1 port map( A => n8, ZN => ML_int_4_5_port);
   U29 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => SHMAG_3_port, ZN => n8
                           );
   U30 : INV_X1 port map( A => n9, ZN => ML_int_4_4_port);
   U31 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => SHMAG_3_port, ZN => n9
                           );
   U32 : INV_X1 port map( A => n10, ZN => ML_int_4_3_port);
   U33 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => SHMAG_3_port, ZN => 
                           n10);
   U34 : INV_X1 port map( A => n11, ZN => ML_int_4_2_port);
   U35 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => SHMAG_3_port, ZN => 
                           n11);
   U36 : INV_X1 port map( A => n12, ZN => ML_int_4_1_port);
   U37 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => SHMAG_3_port, ZN => 
                           n12);
   U38 : INV_X1 port map( A => n13, ZN => ML_int_4_0_port);
   U39 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => SHMAG_3_port, ZN => 
                           n13);
   U40 : INV_X1 port map( A => SH(3), ZN => SHMAG_3_port);
   U41 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_3_port);
   U42 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_2_port);
   U43 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_1_port);
   U44 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_0_port);
   U45 : INV_X1 port map( A => SH(2), ZN => SHMAG_2_port);
   U46 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => SHMAG_1_port, ZN => 
                           ML_int_2_1_port);
   U47 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => SHMAG_1_port, ZN => 
                           ML_int_2_0_port);
   U48 : INV_X1 port map( A => SH(1), ZN => SHMAG_1_port);
   U49 : AND2_X1 port map( A1 => A(0), A2 => SHMAG_0_port, ZN => 
                           ML_int_1_0_port);
   U50 : INV_X1 port map( A => SH(0), ZN => SHMAG_0_port);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end DATAPTH_NBIT32_REG_BIT5_DW01_inc_0;

architecture SYN_rpl of DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_7;

architecture SYN_struct of MUX21_GENERIC_NBIT4_7 is

   component MUX21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_28 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_27 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_26 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_25 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_6;

architecture SYN_struct of MUX21_GENERIC_NBIT4_6 is

   component MUX21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_24 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_23 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_22 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_21 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_5;

architecture SYN_struct of MUX21_GENERIC_NBIT4_5 is

   component MUX21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_20 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_19 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_18 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_17 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_4;

architecture SYN_struct of MUX21_GENERIC_NBIT4_4 is

   component MUX21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_16 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_15 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_14 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_13 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_3;

architecture SYN_struct of MUX21_GENERIC_NBIT4_3 is

   component MUX21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_12 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_11 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_10 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_9 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_2;

architecture SYN_struct of MUX21_GENERIC_NBIT4_2 is

   component MUX21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_8 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_7 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_6 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_5 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_1;

architecture SYN_struct of MUX21_GENERIC_NBIT4_1 is

   component MUX21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_4 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_3 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_2 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_1 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_15;

architecture SYN_BEHAVIORAL of RCA_NBIT4_15 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_14;

architecture SYN_BEHAVIORAL of RCA_NBIT4_14 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_13;

architecture SYN_BEHAVIORAL of RCA_NBIT4_13 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_12;

architecture SYN_BEHAVIORAL of RCA_NBIT4_12 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_11;

architecture SYN_BEHAVIORAL of RCA_NBIT4_11 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_10;

architecture SYN_BEHAVIORAL of RCA_NBIT4_10 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_9;

architecture SYN_BEHAVIORAL of RCA_NBIT4_9 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_8;

architecture SYN_BEHAVIORAL of RCA_NBIT4_8 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_7;

architecture SYN_BEHAVIORAL of RCA_NBIT4_7 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_6;

architecture SYN_BEHAVIORAL of RCA_NBIT4_6 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_5;

architecture SYN_BEHAVIORAL of RCA_NBIT4_5 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_4;

architecture SYN_BEHAVIORAL of RCA_NBIT4_4 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_3;

architecture SYN_BEHAVIORAL of RCA_NBIT4_3 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_2;

architecture SYN_BEHAVIORAL of RCA_NBIT4_2 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_1;

architecture SYN_BEHAVIORAL of RCA_NBIT4_1 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_42 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_42;

architecture SYN_behave of P_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_41 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_41;

architecture SYN_behave of P_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_40 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_40;

architecture SYN_behave of P_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_39 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_39;

architecture SYN_behave of P_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_38 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_38;

architecture SYN_behave of P_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_37 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_37;

architecture SYN_behave of P_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_36 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_36;

architecture SYN_behave of P_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_35 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_35;

architecture SYN_behave of P_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_34 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_34;

architecture SYN_behave of P_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_33 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_33;

architecture SYN_behave of P_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_32 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_32;

architecture SYN_behave of P_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_31 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_31;

architecture SYN_behave of P_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_30 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_30;

architecture SYN_behave of P_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_29 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_29;

architecture SYN_behave of P_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_28 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_28;

architecture SYN_behave of P_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_27 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_27;

architecture SYN_behave of P_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_26 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_26;

architecture SYN_behave of P_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_25 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_25;

architecture SYN_behave of P_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_24 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_24;

architecture SYN_behave of P_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_23 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_23;

architecture SYN_behave of P_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_22 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_22;

architecture SYN_behave of P_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_21 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_21;

architecture SYN_behave of P_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_20 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_20;

architecture SYN_behave of P_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_19 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_19;

architecture SYN_behave of P_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_18 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_18;

architecture SYN_behave of P_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_17 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_17;

architecture SYN_behave of P_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_16 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_16;

architecture SYN_behave of P_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_15 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_15;

architecture SYN_behave of P_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_14 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_14;

architecture SYN_behave of P_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_13 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_13;

architecture SYN_behave of P_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_12 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_12;

architecture SYN_behave of P_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_11 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_11;

architecture SYN_behave of P_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_10 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_10;

architecture SYN_behave of P_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_9 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_9;

architecture SYN_behave of P_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_8 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_8;

architecture SYN_behave of P_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_7 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_7;

architecture SYN_behave of P_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_6 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_6;

architecture SYN_behave of P_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_5 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_5;

architecture SYN_behave of P_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_4 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_4;

architecture SYN_behave of P_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_3 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_3;

architecture SYN_behave of P_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_2 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_2;

architecture SYN_behave of P_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_1 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_1;

architecture SYN_behave of P_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_7;

architecture SYN_STRUCTURAL of CSB_NBIT4_7 is

   component MUX21_GENERIC_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1008, n_1009 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1008);
   RCA1 : RCA_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1009);
   MUXCin : MUX21_GENERIC_NBIT4_7 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_6;

architecture SYN_STRUCTURAL of CSB_NBIT4_6 is

   component MUX21_GENERIC_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1010, n_1011 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1010);
   RCA1 : RCA_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1011);
   MUXCin : MUX21_GENERIC_NBIT4_6 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_5;

architecture SYN_STRUCTURAL of CSB_NBIT4_5 is

   component MUX21_GENERIC_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1012, n_1013 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1012);
   RCA1 : RCA_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1013);
   MUXCin : MUX21_GENERIC_NBIT4_5 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_4;

architecture SYN_STRUCTURAL of CSB_NBIT4_4 is

   component MUX21_GENERIC_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1014, n_1015 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1014);
   RCA1 : RCA_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1015);
   MUXCin : MUX21_GENERIC_NBIT4_4 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_3;

architecture SYN_STRUCTURAL of CSB_NBIT4_3 is

   component MUX21_GENERIC_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1016, n_1017 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1016);
   RCA1 : RCA_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1017);
   MUXCin : MUX21_GENERIC_NBIT4_3 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_2;

architecture SYN_STRUCTURAL of CSB_NBIT4_2 is

   component MUX21_GENERIC_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1018, n_1019 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1018);
   RCA1 : RCA_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1019);
   MUXCin : MUX21_GENERIC_NBIT4_2 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_1;

architecture SYN_STRUCTURAL of CSB_NBIT4_1 is

   component MUX21_GENERIC_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1020, n_1021 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1020);
   RCA1 : RCA_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1021);
   MUXCin : MUX21_GENERIC_NBIT4_1 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_42 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_42;

architecture SYN_arch of PG_42 is

   component P_42
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_42
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_42 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_42 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_41 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_41;

architecture SYN_arch of PG_41 is

   component P_41
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_41
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_41 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_41 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_40 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_40;

architecture SYN_arch of PG_40 is

   component P_40
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_40
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_40 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_40 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_39 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_39;

architecture SYN_arch of PG_39 is

   component P_39
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_39
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_39 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_39 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_38 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_38;

architecture SYN_arch of PG_38 is

   component P_38
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_38
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_38 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_38 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_37 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_37;

architecture SYN_arch of PG_37 is

   component P_37
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_37
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_37 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_37 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_36 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_36;

architecture SYN_arch of PG_36 is

   component P_36
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_36
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_36 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_36 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_35 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_35;

architecture SYN_arch of PG_35 is

   component P_35
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_35
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_35 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_35 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_34 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_34;

architecture SYN_arch of PG_34 is

   component P_34
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_34
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_34 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_34 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_33 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_33;

architecture SYN_arch of PG_33 is

   component P_33
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_33
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_33 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_33 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_32 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_32;

architecture SYN_arch of PG_32 is

   component P_32
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_32
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_32 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_32 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_31 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_31;

architecture SYN_arch of PG_31 is

   component P_31
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_31
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_31 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_31 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_30 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_30;

architecture SYN_arch of PG_30 is

   component P_30
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_30
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_30 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_30 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_29 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_29;

architecture SYN_arch of PG_29 is

   component P_29
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_29
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_29 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_29 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_28 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_28;

architecture SYN_arch of PG_28 is

   component P_28
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_28
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_28 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_28 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_27 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_27;

architecture SYN_arch of PG_27 is

   component P_27
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_27
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_27 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_27 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_26 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_26;

architecture SYN_arch of PG_26 is

   component P_26
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_26
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_26 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_26 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_25 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_25;

architecture SYN_arch of PG_25 is

   component P_25
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_25
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_25 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_25 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_24 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_24;

architecture SYN_arch of PG_24 is

   component P_24
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_24
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_24 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_24 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_23 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_23;

architecture SYN_arch of PG_23 is

   component P_23
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_23
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_23 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_23 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_22 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_22;

architecture SYN_arch of PG_22 is

   component P_22
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_22
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_22 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_22 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_21 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_21;

architecture SYN_arch of PG_21 is

   component P_21
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_21
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_21 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_21 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_20 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_20;

architecture SYN_arch of PG_20 is

   component P_20
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_20
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_20 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_20 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_19 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_19;

architecture SYN_arch of PG_19 is

   component P_19
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_19
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_19 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_19 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_18 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_18;

architecture SYN_arch of PG_18 is

   component P_18
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_18
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_18 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_18 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_17 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_17;

architecture SYN_arch of PG_17 is

   component P_17
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_17
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_17 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_17 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_16 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_16;

architecture SYN_arch of PG_16 is

   component P_16
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_16
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_16 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_16 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_15 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_15;

architecture SYN_arch of PG_15 is

   component P_15
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_15
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_15 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_15 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_14 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_14;

architecture SYN_arch of PG_14 is

   component P_14
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_14
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_14 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_14 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_13 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_13;

architecture SYN_arch of PG_13 is

   component P_13
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_13
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_13 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_13 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_12 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_12;

architecture SYN_arch of PG_12 is

   component P_12
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_12
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_12 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_12 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_11 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_11;

architecture SYN_arch of PG_11 is

   component P_11
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_11
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_11 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_11 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_10 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_10;

architecture SYN_arch of PG_10 is

   component P_10
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_10
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_10 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_10 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_9 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_9;

architecture SYN_arch of PG_9 is

   component P_9
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_9
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_9 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_9 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_8 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_8;

architecture SYN_arch of PG_8 is

   component P_8
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_8
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_8 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_8 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_7 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_7;

architecture SYN_arch of PG_7 is

   component P_7
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_7
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_7 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_7 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_6 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_6;

architecture SYN_arch of PG_6 is

   component P_6
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_6
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_6 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_6 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_5 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_5;

architecture SYN_arch of PG_5 is

   component P_5
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_5
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_5 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_5 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_4 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_4;

architecture SYN_arch of PG_4 is

   component P_4
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_4
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_4 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_4 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_3 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_3;

architecture SYN_arch of PG_3 is

   component P_3
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_3
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_3 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_3 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_2 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_2;

architecture SYN_arch of PG_2 is

   component P_2
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_2
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_2 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_2 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_1 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_1;

architecture SYN_arch of PG_1 is

   component P_1
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_1
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_1 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_1 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_52 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_52;

architecture SYN_behave of G_52 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_51 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_51;

architecture SYN_behave of G_51 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_50 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_50;

architecture SYN_behave of G_50 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_49 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_49;

architecture SYN_behave of G_49 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_48 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_48;

architecture SYN_behave of G_48 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_47 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_47;

architecture SYN_behave of G_47 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_46 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_46;

architecture SYN_behave of G_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_45 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_45;

architecture SYN_behave of G_45 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_44 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_44;

architecture SYN_behave of G_44 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_43 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_43;

architecture SYN_behave of G_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_42 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_42;

architecture SYN_behave of G_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_41 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_41;

architecture SYN_behave of G_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_40 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_40;

architecture SYN_behave of G_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_39 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_39;

architecture SYN_behave of G_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_38 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_38;

architecture SYN_behave of G_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_37 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_37;

architecture SYN_behave of G_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_36 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_36;

architecture SYN_behave of G_36 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_35 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_35;

architecture SYN_behave of G_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_34 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_34;

architecture SYN_behave of G_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_33 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_33;

architecture SYN_behave of G_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_32 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_32;

architecture SYN_behave of G_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_31 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_31;

architecture SYN_behave of G_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_30 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_30;

architecture SYN_behave of G_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_29 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_29;

architecture SYN_behave of G_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_28 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_28;

architecture SYN_behave of G_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_27 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_27;

architecture SYN_behave of G_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_26 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_26;

architecture SYN_behave of G_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_25 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_25;

architecture SYN_behave of G_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_24 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_24;

architecture SYN_behave of G_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_23 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_23;

architecture SYN_behave of G_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_22 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_22;

architecture SYN_behave of G_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_21 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_21;

architecture SYN_behave of G_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_20 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_20;

architecture SYN_behave of G_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_19 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_19;

architecture SYN_behave of G_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_18 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_18;

architecture SYN_behave of G_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_17 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_17;

architecture SYN_behave of G_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_16 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_16;

architecture SYN_behave of G_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_15 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_15;

architecture SYN_behave of G_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_14 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_14;

architecture SYN_behave of G_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_13 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_13;

architecture SYN_behave of G_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_12 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_12;

architecture SYN_behave of G_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_11 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_11;

architecture SYN_behave of G_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_10 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_10;

architecture SYN_behave of G_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_9 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_9;

architecture SYN_behave of G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_8 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_8;

architecture SYN_behave of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_7 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_7;

architecture SYN_behave of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_6 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_6;

architecture SYN_behave of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_5 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_5;

architecture SYN_behave of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_4 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_4;

architecture SYN_behave of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_3 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_3;

architecture SYN_behave of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_2 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_2;

architecture SYN_behave of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_1 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_1;

architecture SYN_behave of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_767 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_767;

architecture SYN_ARCH2 of ND2_767 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_766 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_766;

architecture SYN_ARCH2 of ND2_766 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_765 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_765;

architecture SYN_ARCH2 of ND2_765 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_764 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_764;

architecture SYN_ARCH2 of ND2_764 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_763 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_763;

architecture SYN_ARCH2 of ND2_763 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_762 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_762;

architecture SYN_ARCH2 of ND2_762 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_761 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_761;

architecture SYN_ARCH2 of ND2_761 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_760 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_760;

architecture SYN_ARCH2 of ND2_760 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_759 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_759;

architecture SYN_ARCH2 of ND2_759 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_758 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_758;

architecture SYN_ARCH2 of ND2_758 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_757 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_757;

architecture SYN_ARCH2 of ND2_757 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_756 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_756;

architecture SYN_ARCH2 of ND2_756 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_755 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_755;

architecture SYN_ARCH2 of ND2_755 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_754 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_754;

architecture SYN_ARCH2 of ND2_754 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_753 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_753;

architecture SYN_ARCH2 of ND2_753 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_752 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_752;

architecture SYN_ARCH2 of ND2_752 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_751 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_751;

architecture SYN_ARCH2 of ND2_751 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_750 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_750;

architecture SYN_ARCH2 of ND2_750 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_749 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_749;

architecture SYN_ARCH2 of ND2_749 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_748 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_748;

architecture SYN_ARCH2 of ND2_748 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_747 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_747;

architecture SYN_ARCH2 of ND2_747 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_746 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_746;

architecture SYN_ARCH2 of ND2_746 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_745 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_745;

architecture SYN_ARCH2 of ND2_745 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_744 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_744;

architecture SYN_ARCH2 of ND2_744 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_743 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_743;

architecture SYN_ARCH2 of ND2_743 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_742 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_742;

architecture SYN_ARCH2 of ND2_742 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_741 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_741;

architecture SYN_ARCH2 of ND2_741 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_740 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_740;

architecture SYN_ARCH2 of ND2_740 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_739 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_739;

architecture SYN_ARCH2 of ND2_739 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_738 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_738;

architecture SYN_ARCH2 of ND2_738 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_737 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_737;

architecture SYN_ARCH2 of ND2_737 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_736 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_736;

architecture SYN_ARCH2 of ND2_736 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_735 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_735;

architecture SYN_ARCH2 of ND2_735 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_734 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_734;

architecture SYN_ARCH2 of ND2_734 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_733 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_733;

architecture SYN_ARCH2 of ND2_733 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_732 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_732;

architecture SYN_ARCH2 of ND2_732 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_731 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_731;

architecture SYN_ARCH2 of ND2_731 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_730 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_730;

architecture SYN_ARCH2 of ND2_730 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_729 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_729;

architecture SYN_ARCH2 of ND2_729 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_728 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_728;

architecture SYN_ARCH2 of ND2_728 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_727 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_727;

architecture SYN_ARCH2 of ND2_727 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_726 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_726;

architecture SYN_ARCH2 of ND2_726 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_725 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_725;

architecture SYN_ARCH2 of ND2_725 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_724 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_724;

architecture SYN_ARCH2 of ND2_724 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_723 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_723;

architecture SYN_ARCH2 of ND2_723 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_722 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_722;

architecture SYN_ARCH2 of ND2_722 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_721 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_721;

architecture SYN_ARCH2 of ND2_721 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_720 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_720;

architecture SYN_ARCH2 of ND2_720 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_719 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_719;

architecture SYN_ARCH2 of ND2_719 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_718 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_718;

architecture SYN_ARCH2 of ND2_718 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_717 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_717;

architecture SYN_ARCH2 of ND2_717 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_716 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_716;

architecture SYN_ARCH2 of ND2_716 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_715 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_715;

architecture SYN_ARCH2 of ND2_715 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_714 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_714;

architecture SYN_ARCH2 of ND2_714 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_713 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_713;

architecture SYN_ARCH2 of ND2_713 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_712 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_712;

architecture SYN_ARCH2 of ND2_712 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_711 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_711;

architecture SYN_ARCH2 of ND2_711 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_710 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_710;

architecture SYN_ARCH2 of ND2_710 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_709 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_709;

architecture SYN_ARCH2 of ND2_709 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_708 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_708;

architecture SYN_ARCH2 of ND2_708 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_707 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_707;

architecture SYN_ARCH2 of ND2_707 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_706 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_706;

architecture SYN_ARCH2 of ND2_706 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_705 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_705;

architecture SYN_ARCH2 of ND2_705 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_704 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_704;

architecture SYN_ARCH2 of ND2_704 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_703 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_703;

architecture SYN_ARCH2 of ND2_703 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_702 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_702;

architecture SYN_ARCH2 of ND2_702 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_701 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_701;

architecture SYN_ARCH2 of ND2_701 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_700 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_700;

architecture SYN_ARCH2 of ND2_700 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_699 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_699;

architecture SYN_ARCH2 of ND2_699 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_698 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_698;

architecture SYN_ARCH2 of ND2_698 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_697 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_697;

architecture SYN_ARCH2 of ND2_697 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_696 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_696;

architecture SYN_ARCH2 of ND2_696 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_695 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_695;

architecture SYN_ARCH2 of ND2_695 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_694 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_694;

architecture SYN_ARCH2 of ND2_694 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_693 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_693;

architecture SYN_ARCH2 of ND2_693 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_692 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_692;

architecture SYN_ARCH2 of ND2_692 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_691 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_691;

architecture SYN_ARCH2 of ND2_691 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_690 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_690;

architecture SYN_ARCH2 of ND2_690 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_689 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_689;

architecture SYN_ARCH2 of ND2_689 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_688 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_688;

architecture SYN_ARCH2 of ND2_688 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_687 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_687;

architecture SYN_ARCH2 of ND2_687 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_686 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_686;

architecture SYN_ARCH2 of ND2_686 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_685 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_685;

architecture SYN_ARCH2 of ND2_685 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_684 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_684;

architecture SYN_ARCH2 of ND2_684 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_683 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_683;

architecture SYN_ARCH2 of ND2_683 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_682 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_682;

architecture SYN_ARCH2 of ND2_682 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_681 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_681;

architecture SYN_ARCH2 of ND2_681 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_680 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_680;

architecture SYN_ARCH2 of ND2_680 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_679 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_679;

architecture SYN_ARCH2 of ND2_679 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_678 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_678;

architecture SYN_ARCH2 of ND2_678 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_677 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_677;

architecture SYN_ARCH2 of ND2_677 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_676 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_676;

architecture SYN_ARCH2 of ND2_676 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_675 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_675;

architecture SYN_ARCH2 of ND2_675 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_674 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_674;

architecture SYN_ARCH2 of ND2_674 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_673 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_673;

architecture SYN_ARCH2 of ND2_673 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_672 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_672;

architecture SYN_ARCH2 of ND2_672 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_671 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_671;

architecture SYN_ARCH2 of ND2_671 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_670 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_670;

architecture SYN_ARCH2 of ND2_670 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_669 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_669;

architecture SYN_ARCH2 of ND2_669 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_668 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_668;

architecture SYN_ARCH2 of ND2_668 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_667 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_667;

architecture SYN_ARCH2 of ND2_667 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_666 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_666;

architecture SYN_ARCH2 of ND2_666 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_665 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_665;

architecture SYN_ARCH2 of ND2_665 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_664 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_664;

architecture SYN_ARCH2 of ND2_664 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_663 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_663;

architecture SYN_ARCH2 of ND2_663 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_662 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_662;

architecture SYN_ARCH2 of ND2_662 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_661 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_661;

architecture SYN_ARCH2 of ND2_661 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_660 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_660;

architecture SYN_ARCH2 of ND2_660 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_659 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_659;

architecture SYN_ARCH2 of ND2_659 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_658 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_658;

architecture SYN_ARCH2 of ND2_658 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_657 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_657;

architecture SYN_ARCH2 of ND2_657 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_656 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_656;

architecture SYN_ARCH2 of ND2_656 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_655 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_655;

architecture SYN_ARCH2 of ND2_655 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_654 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_654;

architecture SYN_ARCH2 of ND2_654 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_653 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_653;

architecture SYN_ARCH2 of ND2_653 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_652 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_652;

architecture SYN_ARCH2 of ND2_652 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_651 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_651;

architecture SYN_ARCH2 of ND2_651 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_650 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_650;

architecture SYN_ARCH2 of ND2_650 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_649 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_649;

architecture SYN_ARCH2 of ND2_649 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_648 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_648;

architecture SYN_ARCH2 of ND2_648 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_647 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_647;

architecture SYN_ARCH2 of ND2_647 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_646 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_646;

architecture SYN_ARCH2 of ND2_646 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_645 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_645;

architecture SYN_ARCH2 of ND2_645 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_644 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_644;

architecture SYN_ARCH2 of ND2_644 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_643 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_643;

architecture SYN_ARCH2 of ND2_643 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_642 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_642;

architecture SYN_ARCH2 of ND2_642 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_641 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_641;

architecture SYN_ARCH2 of ND2_641 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_640 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_640;

architecture SYN_ARCH2 of ND2_640 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_639 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_639;

architecture SYN_ARCH2 of ND2_639 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_638 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_638;

architecture SYN_ARCH2 of ND2_638 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_637 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_637;

architecture SYN_ARCH2 of ND2_637 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_636 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_636;

architecture SYN_ARCH2 of ND2_636 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_635 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_635;

architecture SYN_ARCH2 of ND2_635 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_634 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_634;

architecture SYN_ARCH2 of ND2_634 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_633 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_633;

architecture SYN_ARCH2 of ND2_633 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_632 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_632;

architecture SYN_ARCH2 of ND2_632 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_631 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_631;

architecture SYN_ARCH2 of ND2_631 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_630 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_630;

architecture SYN_ARCH2 of ND2_630 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_629 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_629;

architecture SYN_ARCH2 of ND2_629 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_628 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_628;

architecture SYN_ARCH2 of ND2_628 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_627 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_627;

architecture SYN_ARCH2 of ND2_627 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_626 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_626;

architecture SYN_ARCH2 of ND2_626 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_625 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_625;

architecture SYN_ARCH2 of ND2_625 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_624 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_624;

architecture SYN_ARCH2 of ND2_624 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_623 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_623;

architecture SYN_ARCH2 of ND2_623 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_622 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_622;

architecture SYN_ARCH2 of ND2_622 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_621 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_621;

architecture SYN_ARCH2 of ND2_621 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_620 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_620;

architecture SYN_ARCH2 of ND2_620 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_619 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_619;

architecture SYN_ARCH2 of ND2_619 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_618 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_618;

architecture SYN_ARCH2 of ND2_618 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_617 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_617;

architecture SYN_ARCH2 of ND2_617 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_616 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_616;

architecture SYN_ARCH2 of ND2_616 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_615 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_615;

architecture SYN_ARCH2 of ND2_615 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_614 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_614;

architecture SYN_ARCH2 of ND2_614 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_613 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_613;

architecture SYN_ARCH2 of ND2_613 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_612 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_612;

architecture SYN_ARCH2 of ND2_612 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_611 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_611;

architecture SYN_ARCH2 of ND2_611 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_610 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_610;

architecture SYN_ARCH2 of ND2_610 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_609 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_609;

architecture SYN_ARCH2 of ND2_609 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_608 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_608;

architecture SYN_ARCH2 of ND2_608 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_607 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_607;

architecture SYN_ARCH2 of ND2_607 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_606 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_606;

architecture SYN_ARCH2 of ND2_606 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_605 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_605;

architecture SYN_ARCH2 of ND2_605 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_604 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_604;

architecture SYN_ARCH2 of ND2_604 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_603 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_603;

architecture SYN_ARCH2 of ND2_603 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_602 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_602;

architecture SYN_ARCH2 of ND2_602 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_601 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_601;

architecture SYN_ARCH2 of ND2_601 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_600 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_600;

architecture SYN_ARCH2 of ND2_600 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_599 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_599;

architecture SYN_ARCH2 of ND2_599 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_598 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_598;

architecture SYN_ARCH2 of ND2_598 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_597 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_597;

architecture SYN_ARCH2 of ND2_597 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_596 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_596;

architecture SYN_ARCH2 of ND2_596 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_595 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_595;

architecture SYN_ARCH2 of ND2_595 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_594 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_594;

architecture SYN_ARCH2 of ND2_594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_593 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_593;

architecture SYN_ARCH2 of ND2_593 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_592 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_592;

architecture SYN_ARCH2 of ND2_592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_591 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_591;

architecture SYN_ARCH2 of ND2_591 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_590 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_590;

architecture SYN_ARCH2 of ND2_590 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_589 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_589;

architecture SYN_ARCH2 of ND2_589 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_588 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_588;

architecture SYN_ARCH2 of ND2_588 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_587 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_587;

architecture SYN_ARCH2 of ND2_587 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_586 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_586;

architecture SYN_ARCH2 of ND2_586 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_585 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_585;

architecture SYN_ARCH2 of ND2_585 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_584 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_584;

architecture SYN_ARCH2 of ND2_584 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_583 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_583;

architecture SYN_ARCH2 of ND2_583 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_582 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_582;

architecture SYN_ARCH2 of ND2_582 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_581 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_581;

architecture SYN_ARCH2 of ND2_581 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_580 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_580;

architecture SYN_ARCH2 of ND2_580 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_579 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_579;

architecture SYN_ARCH2 of ND2_579 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_578 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_578;

architecture SYN_ARCH2 of ND2_578 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_577 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_577;

architecture SYN_ARCH2 of ND2_577 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_576 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_576;

architecture SYN_ARCH2 of ND2_576 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_575 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_575;

architecture SYN_ARCH2 of ND2_575 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_574 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_574;

architecture SYN_ARCH2 of ND2_574 is

   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N1, n1_port : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => N1);
   U2 : INV_X1 port map( A => N1, ZN => n1_port);
   U3 : INV_X8 port map( A => n1_port, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_573 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_573;

architecture SYN_ARCH2 of ND2_573 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_572 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_572;

architecture SYN_ARCH2 of ND2_572 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_571 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_571;

architecture SYN_ARCH2 of ND2_571 is

   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N1, n1_port : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => N1);
   U2 : INV_X1 port map( A => N1, ZN => n1_port);
   U3 : INV_X8 port map( A => n1_port, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_570 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_570;

architecture SYN_ARCH2 of ND2_570 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_569 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_569;

architecture SYN_ARCH2 of ND2_569 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_568 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_568;

architecture SYN_ARCH2 of ND2_568 is

   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N1, n1_port : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => N1);
   U2 : INV_X1 port map( A => N1, ZN => n1_port);
   U3 : INV_X8 port map( A => n1_port, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_567 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_567;

architecture SYN_ARCH2 of ND2_567 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_566 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_566;

architecture SYN_ARCH2 of ND2_566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_565 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_565;

architecture SYN_ARCH2 of ND2_565 is

   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N1, n1_port : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => N1);
   U2 : INV_X1 port map( A => N1, ZN => n1_port);
   U3 : INV_X8 port map( A => n1_port, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_564 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_564;

architecture SYN_ARCH2 of ND2_564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_563 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_563;

architecture SYN_ARCH2 of ND2_563 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_562 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_562;

architecture SYN_ARCH2 of ND2_562 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_561 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_561;

architecture SYN_ARCH2 of ND2_561 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_560 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_560;

architecture SYN_ARCH2 of ND2_560 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_559 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_559;

architecture SYN_ARCH2 of ND2_559 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_558 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_558;

architecture SYN_ARCH2 of ND2_558 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_557 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_557;

architecture SYN_ARCH2 of ND2_557 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_556 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_556;

architecture SYN_ARCH2 of ND2_556 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_555 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_555;

architecture SYN_ARCH2 of ND2_555 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_554 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_554;

architecture SYN_ARCH2 of ND2_554 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_553 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_553;

architecture SYN_ARCH2 of ND2_553 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_552 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_552;

architecture SYN_ARCH2 of ND2_552 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_551 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_551;

architecture SYN_ARCH2 of ND2_551 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_550 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_550;

architecture SYN_ARCH2 of ND2_550 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_549 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_549;

architecture SYN_ARCH2 of ND2_549 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_548 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_548;

architecture SYN_ARCH2 of ND2_548 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_547 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_547;

architecture SYN_ARCH2 of ND2_547 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_546 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_546;

architecture SYN_ARCH2 of ND2_546 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_545 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_545;

architecture SYN_ARCH2 of ND2_545 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_544 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_544;

architecture SYN_ARCH2 of ND2_544 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_543 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_543;

architecture SYN_ARCH2 of ND2_543 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_542 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_542;

architecture SYN_ARCH2 of ND2_542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_541 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_541;

architecture SYN_ARCH2 of ND2_541 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_540 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_540;

architecture SYN_ARCH2 of ND2_540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_539 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_539;

architecture SYN_ARCH2 of ND2_539 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_538 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_538;

architecture SYN_ARCH2 of ND2_538 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_537 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_537;

architecture SYN_ARCH2 of ND2_537 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_536 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_536;

architecture SYN_ARCH2 of ND2_536 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_535 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_535;

architecture SYN_ARCH2 of ND2_535 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_534 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_534;

architecture SYN_ARCH2 of ND2_534 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_533 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_533;

architecture SYN_ARCH2 of ND2_533 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_532 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_532;

architecture SYN_ARCH2 of ND2_532 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_531 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_531;

architecture SYN_ARCH2 of ND2_531 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_530 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_530;

architecture SYN_ARCH2 of ND2_530 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_529 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_529;

architecture SYN_ARCH2 of ND2_529 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_528 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_528;

architecture SYN_ARCH2 of ND2_528 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_527 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_527;

architecture SYN_ARCH2 of ND2_527 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_526 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_526;

architecture SYN_ARCH2 of ND2_526 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_525 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_525;

architecture SYN_ARCH2 of ND2_525 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_524 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_524;

architecture SYN_ARCH2 of ND2_524 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_523 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_523;

architecture SYN_ARCH2 of ND2_523 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_522 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_522;

architecture SYN_ARCH2 of ND2_522 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_521 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_521;

architecture SYN_ARCH2 of ND2_521 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_520 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_520;

architecture SYN_ARCH2 of ND2_520 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_519 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_519;

architecture SYN_ARCH2 of ND2_519 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_518 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_518;

architecture SYN_ARCH2 of ND2_518 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_517 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_517;

architecture SYN_ARCH2 of ND2_517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_516 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_516;

architecture SYN_ARCH2 of ND2_516 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_515 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_515;

architecture SYN_ARCH2 of ND2_515 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_514 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_514;

architecture SYN_ARCH2 of ND2_514 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_513 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_513;

architecture SYN_ARCH2 of ND2_513 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_512 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_512;

architecture SYN_ARCH2 of ND2_512 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_511 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_511;

architecture SYN_ARCH2 of ND2_511 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_510 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_510;

architecture SYN_ARCH2 of ND2_510 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_509 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_509;

architecture SYN_ARCH2 of ND2_509 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_508 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_508;

architecture SYN_ARCH2 of ND2_508 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_507 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_507;

architecture SYN_ARCH2 of ND2_507 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_506 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_506;

architecture SYN_ARCH2 of ND2_506 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_505 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_505;

architecture SYN_ARCH2 of ND2_505 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_504 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_504;

architecture SYN_ARCH2 of ND2_504 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_503 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_503;

architecture SYN_ARCH2 of ND2_503 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_502 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_502;

architecture SYN_ARCH2 of ND2_502 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_501 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_501;

architecture SYN_ARCH2 of ND2_501 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_500 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_500;

architecture SYN_ARCH2 of ND2_500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_499 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_499;

architecture SYN_ARCH2 of ND2_499 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_498 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_498;

architecture SYN_ARCH2 of ND2_498 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_497 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_497;

architecture SYN_ARCH2 of ND2_497 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_496 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_496;

architecture SYN_ARCH2 of ND2_496 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_495 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_495;

architecture SYN_ARCH2 of ND2_495 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_494 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_494;

architecture SYN_ARCH2 of ND2_494 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_493 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_493;

architecture SYN_ARCH2 of ND2_493 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_492 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_492;

architecture SYN_ARCH2 of ND2_492 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_491 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_491;

architecture SYN_ARCH2 of ND2_491 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_490 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_490;

architecture SYN_ARCH2 of ND2_490 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_489 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_489;

architecture SYN_ARCH2 of ND2_489 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_488 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_488;

architecture SYN_ARCH2 of ND2_488 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_487 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_487;

architecture SYN_ARCH2 of ND2_487 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_486 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_486;

architecture SYN_ARCH2 of ND2_486 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_485 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_485;

architecture SYN_ARCH2 of ND2_485 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_484 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_484;

architecture SYN_ARCH2 of ND2_484 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_483 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_483;

architecture SYN_ARCH2 of ND2_483 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_482 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_482;

architecture SYN_ARCH2 of ND2_482 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_481 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_481;

architecture SYN_ARCH2 of ND2_481 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_480 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_480;

architecture SYN_ARCH2 of ND2_480 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_479 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_479;

architecture SYN_ARCH2 of ND2_479 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_478 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_478;

architecture SYN_ARCH2 of ND2_478 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_477 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_477;

architecture SYN_ARCH2 of ND2_477 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_476 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_476;

architecture SYN_ARCH2 of ND2_476 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_475 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_475;

architecture SYN_ARCH2 of ND2_475 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_474 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_474;

architecture SYN_ARCH2 of ND2_474 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_473 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_473;

architecture SYN_ARCH2 of ND2_473 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_472 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_472;

architecture SYN_ARCH2 of ND2_472 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_471 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_471;

architecture SYN_ARCH2 of ND2_471 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_470 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_470;

architecture SYN_ARCH2 of ND2_470 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_469 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_469;

architecture SYN_ARCH2 of ND2_469 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_468 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_468;

architecture SYN_ARCH2 of ND2_468 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_467 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_467;

architecture SYN_ARCH2 of ND2_467 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_466 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_466;

architecture SYN_ARCH2 of ND2_466 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_465 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_465;

architecture SYN_ARCH2 of ND2_465 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_464 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_464;

architecture SYN_ARCH2 of ND2_464 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_463 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_463;

architecture SYN_ARCH2 of ND2_463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_462 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_462;

architecture SYN_ARCH2 of ND2_462 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_461 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_461;

architecture SYN_ARCH2 of ND2_461 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_460 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_460;

architecture SYN_ARCH2 of ND2_460 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_459 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_459;

architecture SYN_ARCH2 of ND2_459 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_458 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_458;

architecture SYN_ARCH2 of ND2_458 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_457 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_457;

architecture SYN_ARCH2 of ND2_457 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_456 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_456;

architecture SYN_ARCH2 of ND2_456 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_455 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_455;

architecture SYN_ARCH2 of ND2_455 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_454 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_454;

architecture SYN_ARCH2 of ND2_454 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_453 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_453;

architecture SYN_ARCH2 of ND2_453 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_452 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_452;

architecture SYN_ARCH2 of ND2_452 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_451 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_451;

architecture SYN_ARCH2 of ND2_451 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_450 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_450;

architecture SYN_ARCH2 of ND2_450 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_449 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_449;

architecture SYN_ARCH2 of ND2_449 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_448 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_448;

architecture SYN_ARCH2 of ND2_448 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_447 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_447;

architecture SYN_ARCH2 of ND2_447 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_446 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_446;

architecture SYN_ARCH2 of ND2_446 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_445 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_445;

architecture SYN_ARCH2 of ND2_445 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_444 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_444;

architecture SYN_ARCH2 of ND2_444 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_443 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_443;

architecture SYN_ARCH2 of ND2_443 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_442 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_442;

architecture SYN_ARCH2 of ND2_442 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_441 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_441;

architecture SYN_ARCH2 of ND2_441 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_440 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_440;

architecture SYN_ARCH2 of ND2_440 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_439 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_439;

architecture SYN_ARCH2 of ND2_439 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_438 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_438;

architecture SYN_ARCH2 of ND2_438 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_437 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_437;

architecture SYN_ARCH2 of ND2_437 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_436 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_436;

architecture SYN_ARCH2 of ND2_436 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_435 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_435;

architecture SYN_ARCH2 of ND2_435 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_434 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_434;

architecture SYN_ARCH2 of ND2_434 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_433 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_433;

architecture SYN_ARCH2 of ND2_433 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_432 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_432;

architecture SYN_ARCH2 of ND2_432 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_431 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_431;

architecture SYN_ARCH2 of ND2_431 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_430 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_430;

architecture SYN_ARCH2 of ND2_430 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_429 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_429;

architecture SYN_ARCH2 of ND2_429 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_428 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_428;

architecture SYN_ARCH2 of ND2_428 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_427 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_427;

architecture SYN_ARCH2 of ND2_427 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_426 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_426;

architecture SYN_ARCH2 of ND2_426 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_425 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_425;

architecture SYN_ARCH2 of ND2_425 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_424 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_424;

architecture SYN_ARCH2 of ND2_424 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_423 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_423;

architecture SYN_ARCH2 of ND2_423 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_422 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_422;

architecture SYN_ARCH2 of ND2_422 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_421 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_421;

architecture SYN_ARCH2 of ND2_421 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_420 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_420;

architecture SYN_ARCH2 of ND2_420 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_419 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_419;

architecture SYN_ARCH2 of ND2_419 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_418 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_418;

architecture SYN_ARCH2 of ND2_418 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_417 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_417;

architecture SYN_ARCH2 of ND2_417 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_416 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_416;

architecture SYN_ARCH2 of ND2_416 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_415 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_415;

architecture SYN_ARCH2 of ND2_415 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_414 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_414;

architecture SYN_ARCH2 of ND2_414 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_413 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_413;

architecture SYN_ARCH2 of ND2_413 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_412 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_412;

architecture SYN_ARCH2 of ND2_412 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_411 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_411;

architecture SYN_ARCH2 of ND2_411 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_410 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_410;

architecture SYN_ARCH2 of ND2_410 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_409 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_409;

architecture SYN_ARCH2 of ND2_409 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_408 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_408;

architecture SYN_ARCH2 of ND2_408 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_407 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_407;

architecture SYN_ARCH2 of ND2_407 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_406 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_406;

architecture SYN_ARCH2 of ND2_406 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_405 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_405;

architecture SYN_ARCH2 of ND2_405 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_404 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_404;

architecture SYN_ARCH2 of ND2_404 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_403 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_403;

architecture SYN_ARCH2 of ND2_403 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_402 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_402;

architecture SYN_ARCH2 of ND2_402 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_401 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_401;

architecture SYN_ARCH2 of ND2_401 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_400 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_400;

architecture SYN_ARCH2 of ND2_400 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_399 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_399;

architecture SYN_ARCH2 of ND2_399 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_398 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_398;

architecture SYN_ARCH2 of ND2_398 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_397 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_397;

architecture SYN_ARCH2 of ND2_397 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_396 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_396;

architecture SYN_ARCH2 of ND2_396 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_395 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_395;

architecture SYN_ARCH2 of ND2_395 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_394 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_394;

architecture SYN_ARCH2 of ND2_394 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_393 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_393;

architecture SYN_ARCH2 of ND2_393 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_392 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_392;

architecture SYN_ARCH2 of ND2_392 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_391 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_391;

architecture SYN_ARCH2 of ND2_391 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_390 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_390;

architecture SYN_ARCH2 of ND2_390 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_389 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_389;

architecture SYN_ARCH2 of ND2_389 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_388 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_388;

architecture SYN_ARCH2 of ND2_388 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_387 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_387;

architecture SYN_ARCH2 of ND2_387 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_386 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_386;

architecture SYN_ARCH2 of ND2_386 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_385 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_385;

architecture SYN_ARCH2 of ND2_385 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_384 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_384;

architecture SYN_ARCH2 of ND2_384 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_383 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_383;

architecture SYN_ARCH2 of ND2_383 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_382 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_382;

architecture SYN_ARCH2 of ND2_382 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_381 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_381;

architecture SYN_ARCH2 of ND2_381 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_380 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_380;

architecture SYN_ARCH2 of ND2_380 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_379 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_379;

architecture SYN_ARCH2 of ND2_379 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_378 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_378;

architecture SYN_ARCH2 of ND2_378 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_377 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_377;

architecture SYN_ARCH2 of ND2_377 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_376 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_376;

architecture SYN_ARCH2 of ND2_376 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_375 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_375;

architecture SYN_ARCH2 of ND2_375 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_374 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_374;

architecture SYN_ARCH2 of ND2_374 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_373 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_373;

architecture SYN_ARCH2 of ND2_373 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_372 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_372;

architecture SYN_ARCH2 of ND2_372 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_371 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_371;

architecture SYN_ARCH2 of ND2_371 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_370 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_370;

architecture SYN_ARCH2 of ND2_370 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_369 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_369;

architecture SYN_ARCH2 of ND2_369 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_368 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_368;

architecture SYN_ARCH2 of ND2_368 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_367 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_367;

architecture SYN_ARCH2 of ND2_367 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_366 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_366;

architecture SYN_ARCH2 of ND2_366 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_365 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_365;

architecture SYN_ARCH2 of ND2_365 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_364 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_364;

architecture SYN_ARCH2 of ND2_364 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_363 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_363;

architecture SYN_ARCH2 of ND2_363 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_362 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_362;

architecture SYN_ARCH2 of ND2_362 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_361 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_361;

architecture SYN_ARCH2 of ND2_361 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_360 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_360;

architecture SYN_ARCH2 of ND2_360 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_359 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_359;

architecture SYN_ARCH2 of ND2_359 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_358 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_358;

architecture SYN_ARCH2 of ND2_358 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_357 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_357;

architecture SYN_ARCH2 of ND2_357 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_356 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_356;

architecture SYN_ARCH2 of ND2_356 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_355 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_355;

architecture SYN_ARCH2 of ND2_355 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_354 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_354;

architecture SYN_ARCH2 of ND2_354 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_353 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_353;

architecture SYN_ARCH2 of ND2_353 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_352 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_352;

architecture SYN_ARCH2 of ND2_352 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_351 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_351;

architecture SYN_ARCH2 of ND2_351 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_350 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_350;

architecture SYN_ARCH2 of ND2_350 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_349 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_349;

architecture SYN_ARCH2 of ND2_349 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_348 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_348;

architecture SYN_ARCH2 of ND2_348 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_347 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_347;

architecture SYN_ARCH2 of ND2_347 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_346 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_346;

architecture SYN_ARCH2 of ND2_346 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_345 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_345;

architecture SYN_ARCH2 of ND2_345 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_344 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_344;

architecture SYN_ARCH2 of ND2_344 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_343 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_343;

architecture SYN_ARCH2 of ND2_343 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_342 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_342;

architecture SYN_ARCH2 of ND2_342 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_341 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_341;

architecture SYN_ARCH2 of ND2_341 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_340 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_340;

architecture SYN_ARCH2 of ND2_340 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_339 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_339;

architecture SYN_ARCH2 of ND2_339 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_338 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_338;

architecture SYN_ARCH2 of ND2_338 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_337 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_337;

architecture SYN_ARCH2 of ND2_337 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_336 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_336;

architecture SYN_ARCH2 of ND2_336 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_335 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_335;

architecture SYN_ARCH2 of ND2_335 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_334 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_334;

architecture SYN_ARCH2 of ND2_334 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_333 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_333;

architecture SYN_ARCH2 of ND2_333 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_332 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_332;

architecture SYN_ARCH2 of ND2_332 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_331 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_331;

architecture SYN_ARCH2 of ND2_331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_330 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_330;

architecture SYN_ARCH2 of ND2_330 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_329 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_329;

architecture SYN_ARCH2 of ND2_329 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_328 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_328;

architecture SYN_ARCH2 of ND2_328 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_327 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_327;

architecture SYN_ARCH2 of ND2_327 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_326 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_326;

architecture SYN_ARCH2 of ND2_326 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_325 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_325;

architecture SYN_ARCH2 of ND2_325 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_324 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_324;

architecture SYN_ARCH2 of ND2_324 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_323 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_323;

architecture SYN_ARCH2 of ND2_323 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_322 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_322;

architecture SYN_ARCH2 of ND2_322 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_321 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_321;

architecture SYN_ARCH2 of ND2_321 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_320 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_320;

architecture SYN_ARCH2 of ND2_320 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_319 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_319;

architecture SYN_ARCH2 of ND2_319 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_318 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_318;

architecture SYN_ARCH2 of ND2_318 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_317 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_317;

architecture SYN_ARCH2 of ND2_317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_316 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_316;

architecture SYN_ARCH2 of ND2_316 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_315 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_315;

architecture SYN_ARCH2 of ND2_315 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_314 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_314;

architecture SYN_ARCH2 of ND2_314 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_313 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_313;

architecture SYN_ARCH2 of ND2_313 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_312 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_312;

architecture SYN_ARCH2 of ND2_312 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_311 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_311;

architecture SYN_ARCH2 of ND2_311 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_310 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_310;

architecture SYN_ARCH2 of ND2_310 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_309 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_309;

architecture SYN_ARCH2 of ND2_309 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_308 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_308;

architecture SYN_ARCH2 of ND2_308 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_307 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_307;

architecture SYN_ARCH2 of ND2_307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_306 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_306;

architecture SYN_ARCH2 of ND2_306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_305 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_305;

architecture SYN_ARCH2 of ND2_305 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_304 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_304;

architecture SYN_ARCH2 of ND2_304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_303 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_303;

architecture SYN_ARCH2 of ND2_303 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_302 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_302;

architecture SYN_ARCH2 of ND2_302 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_301 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_301;

architecture SYN_ARCH2 of ND2_301 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_300 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_300;

architecture SYN_ARCH2 of ND2_300 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_299 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_299;

architecture SYN_ARCH2 of ND2_299 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_298 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_298;

architecture SYN_ARCH2 of ND2_298 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_297 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_297;

architecture SYN_ARCH2 of ND2_297 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_296 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_296;

architecture SYN_ARCH2 of ND2_296 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_295 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_295;

architecture SYN_ARCH2 of ND2_295 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_294 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_294;

architecture SYN_ARCH2 of ND2_294 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_293 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_293;

architecture SYN_ARCH2 of ND2_293 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_292 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_292;

architecture SYN_ARCH2 of ND2_292 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_291 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_291;

architecture SYN_ARCH2 of ND2_291 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_290 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_290;

architecture SYN_ARCH2 of ND2_290 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_289 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_289;

architecture SYN_ARCH2 of ND2_289 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_288 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_288;

architecture SYN_ARCH2 of ND2_288 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_287 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_287;

architecture SYN_ARCH2 of ND2_287 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_286 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_286;

architecture SYN_ARCH2 of ND2_286 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_285 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_285;

architecture SYN_ARCH2 of ND2_285 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_284 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_284;

architecture SYN_ARCH2 of ND2_284 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_283 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_283;

architecture SYN_ARCH2 of ND2_283 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_282 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_282;

architecture SYN_ARCH2 of ND2_282 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_281 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_281;

architecture SYN_ARCH2 of ND2_281 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_280 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_280;

architecture SYN_ARCH2 of ND2_280 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_279 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_279;

architecture SYN_ARCH2 of ND2_279 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_278 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_278;

architecture SYN_ARCH2 of ND2_278 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_277 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_277;

architecture SYN_ARCH2 of ND2_277 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_276 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_276;

architecture SYN_ARCH2 of ND2_276 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_275 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_275;

architecture SYN_ARCH2 of ND2_275 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_274 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_274;

architecture SYN_ARCH2 of ND2_274 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_273 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_273;

architecture SYN_ARCH2 of ND2_273 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_272 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_272;

architecture SYN_ARCH2 of ND2_272 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_271 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_271;

architecture SYN_ARCH2 of ND2_271 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_270 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_270;

architecture SYN_ARCH2 of ND2_270 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_269 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_269;

architecture SYN_ARCH2 of ND2_269 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_268 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_268;

architecture SYN_ARCH2 of ND2_268 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_267 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_267;

architecture SYN_ARCH2 of ND2_267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_266 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_266;

architecture SYN_ARCH2 of ND2_266 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_265 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_265;

architecture SYN_ARCH2 of ND2_265 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_264 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_264;

architecture SYN_ARCH2 of ND2_264 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_263 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_263;

architecture SYN_ARCH2 of ND2_263 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_262 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_262;

architecture SYN_ARCH2 of ND2_262 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_261 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_261;

architecture SYN_ARCH2 of ND2_261 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_260 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_260;

architecture SYN_ARCH2 of ND2_260 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_259 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_259;

architecture SYN_ARCH2 of ND2_259 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_258 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_258;

architecture SYN_ARCH2 of ND2_258 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_257 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_257;

architecture SYN_ARCH2 of ND2_257 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_256 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_256;

architecture SYN_ARCH2 of ND2_256 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_255 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_255;

architecture SYN_ARCH2 of ND2_255 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_254 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_254;

architecture SYN_ARCH2 of ND2_254 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_253 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_253;

architecture SYN_ARCH2 of ND2_253 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_252 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_252;

architecture SYN_ARCH2 of ND2_252 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_251 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_251;

architecture SYN_ARCH2 of ND2_251 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_250 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_250;

architecture SYN_ARCH2 of ND2_250 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_249 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_249;

architecture SYN_ARCH2 of ND2_249 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_248 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_248;

architecture SYN_ARCH2 of ND2_248 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_247 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_247;

architecture SYN_ARCH2 of ND2_247 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_246 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_246;

architecture SYN_ARCH2 of ND2_246 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_245 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_245;

architecture SYN_ARCH2 of ND2_245 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_244 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_244;

architecture SYN_ARCH2 of ND2_244 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_243 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_243;

architecture SYN_ARCH2 of ND2_243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_242 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_242;

architecture SYN_ARCH2 of ND2_242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_241 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_241;

architecture SYN_ARCH2 of ND2_241 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_240 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_240;

architecture SYN_ARCH2 of ND2_240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_239 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_239;

architecture SYN_ARCH2 of ND2_239 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_238 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_238;

architecture SYN_ARCH2 of ND2_238 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_237 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_237;

architecture SYN_ARCH2 of ND2_237 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_236 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_236;

architecture SYN_ARCH2 of ND2_236 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_235 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_235;

architecture SYN_ARCH2 of ND2_235 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_234 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_234;

architecture SYN_ARCH2 of ND2_234 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_233 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_233;

architecture SYN_ARCH2 of ND2_233 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_232 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_232;

architecture SYN_ARCH2 of ND2_232 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_231 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_231;

architecture SYN_ARCH2 of ND2_231 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_230 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_230;

architecture SYN_ARCH2 of ND2_230 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_229 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_229;

architecture SYN_ARCH2 of ND2_229 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_228 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_228;

architecture SYN_ARCH2 of ND2_228 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_227 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_227;

architecture SYN_ARCH2 of ND2_227 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_226 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_226;

architecture SYN_ARCH2 of ND2_226 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_225 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_225;

architecture SYN_ARCH2 of ND2_225 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_224 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_224;

architecture SYN_ARCH2 of ND2_224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_223 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_223;

architecture SYN_ARCH2 of ND2_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_222 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_222;

architecture SYN_ARCH2 of ND2_222 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_221 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_221;

architecture SYN_ARCH2 of ND2_221 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_220 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_220;

architecture SYN_ARCH2 of ND2_220 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_219 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_219;

architecture SYN_ARCH2 of ND2_219 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_218 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_218;

architecture SYN_ARCH2 of ND2_218 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_217 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_217;

architecture SYN_ARCH2 of ND2_217 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_216 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_216;

architecture SYN_ARCH2 of ND2_216 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_215 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_215;

architecture SYN_ARCH2 of ND2_215 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_214 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_214;

architecture SYN_ARCH2 of ND2_214 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_213 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_213;

architecture SYN_ARCH2 of ND2_213 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_212 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_212;

architecture SYN_ARCH2 of ND2_212 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_211 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_211;

architecture SYN_ARCH2 of ND2_211 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_210 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_210;

architecture SYN_ARCH2 of ND2_210 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_209 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_209;

architecture SYN_ARCH2 of ND2_209 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_208 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_208;

architecture SYN_ARCH2 of ND2_208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_207 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_207;

architecture SYN_ARCH2 of ND2_207 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_206 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_206;

architecture SYN_ARCH2 of ND2_206 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_205 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_205;

architecture SYN_ARCH2 of ND2_205 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_204 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_204;

architecture SYN_ARCH2 of ND2_204 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_203 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_203;

architecture SYN_ARCH2 of ND2_203 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_202 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_202;

architecture SYN_ARCH2 of ND2_202 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_201 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_201;

architecture SYN_ARCH2 of ND2_201 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_200 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_200;

architecture SYN_ARCH2 of ND2_200 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_199 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_199;

architecture SYN_ARCH2 of ND2_199 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_198 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_198;

architecture SYN_ARCH2 of ND2_198 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_197 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_197;

architecture SYN_ARCH2 of ND2_197 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_196 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_196;

architecture SYN_ARCH2 of ND2_196 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_195 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_195;

architecture SYN_ARCH2 of ND2_195 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_194 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_194;

architecture SYN_ARCH2 of ND2_194 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_193 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_193;

architecture SYN_ARCH2 of ND2_193 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_192 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_192;

architecture SYN_ARCH2 of ND2_192 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_191;

architecture SYN_ARCH2 of ND2_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_190;

architecture SYN_ARCH2 of ND2_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_189;

architecture SYN_ARCH2 of ND2_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_188;

architecture SYN_ARCH2 of ND2_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_187;

architecture SYN_ARCH2 of ND2_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_186;

architecture SYN_ARCH2 of ND2_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_185;

architecture SYN_ARCH2 of ND2_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_184;

architecture SYN_ARCH2 of ND2_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_183;

architecture SYN_ARCH2 of ND2_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_182;

architecture SYN_ARCH2 of ND2_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_181;

architecture SYN_ARCH2 of ND2_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_180;

architecture SYN_ARCH2 of ND2_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_179;

architecture SYN_ARCH2 of ND2_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_178;

architecture SYN_ARCH2 of ND2_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_177;

architecture SYN_ARCH2 of ND2_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_176;

architecture SYN_ARCH2 of ND2_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_175;

architecture SYN_ARCH2 of ND2_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_174;

architecture SYN_ARCH2 of ND2_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_173;

architecture SYN_ARCH2 of ND2_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_172;

architecture SYN_ARCH2 of ND2_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_171;

architecture SYN_ARCH2 of ND2_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_170;

architecture SYN_ARCH2 of ND2_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_169;

architecture SYN_ARCH2 of ND2_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_168;

architecture SYN_ARCH2 of ND2_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_167;

architecture SYN_ARCH2 of ND2_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_166;

architecture SYN_ARCH2 of ND2_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_165;

architecture SYN_ARCH2 of ND2_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_164;

architecture SYN_ARCH2 of ND2_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_163;

architecture SYN_ARCH2 of ND2_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_162;

architecture SYN_ARCH2 of ND2_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_161;

architecture SYN_ARCH2 of ND2_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_160;

architecture SYN_ARCH2 of ND2_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_159;

architecture SYN_ARCH2 of ND2_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_158;

architecture SYN_ARCH2 of ND2_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_157;

architecture SYN_ARCH2 of ND2_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_156;

architecture SYN_ARCH2 of ND2_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_155;

architecture SYN_ARCH2 of ND2_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_154;

architecture SYN_ARCH2 of ND2_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_153;

architecture SYN_ARCH2 of ND2_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_152;

architecture SYN_ARCH2 of ND2_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_151;

architecture SYN_ARCH2 of ND2_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_150;

architecture SYN_ARCH2 of ND2_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_149;

architecture SYN_ARCH2 of ND2_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_148;

architecture SYN_ARCH2 of ND2_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_147;

architecture SYN_ARCH2 of ND2_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_146;

architecture SYN_ARCH2 of ND2_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_145;

architecture SYN_ARCH2 of ND2_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_144;

architecture SYN_ARCH2 of ND2_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_143;

architecture SYN_ARCH2 of ND2_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_142;

architecture SYN_ARCH2 of ND2_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_141;

architecture SYN_ARCH2 of ND2_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_140;

architecture SYN_ARCH2 of ND2_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_139;

architecture SYN_ARCH2 of ND2_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_138;

architecture SYN_ARCH2 of ND2_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_137;

architecture SYN_ARCH2 of ND2_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_136;

architecture SYN_ARCH2 of ND2_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_135;

architecture SYN_ARCH2 of ND2_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_134;

architecture SYN_ARCH2 of ND2_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_133;

architecture SYN_ARCH2 of ND2_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_132;

architecture SYN_ARCH2 of ND2_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_131;

architecture SYN_ARCH2 of ND2_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_130;

architecture SYN_ARCH2 of ND2_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_129;

architecture SYN_ARCH2 of ND2_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_128;

architecture SYN_ARCH2 of ND2_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_127;

architecture SYN_ARCH2 of ND2_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_126;

architecture SYN_ARCH2 of ND2_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_125;

architecture SYN_ARCH2 of ND2_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_124;

architecture SYN_ARCH2 of ND2_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_123;

architecture SYN_ARCH2 of ND2_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_122;

architecture SYN_ARCH2 of ND2_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_121;

architecture SYN_ARCH2 of ND2_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_120;

architecture SYN_ARCH2 of ND2_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_119;

architecture SYN_ARCH2 of ND2_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_118;

architecture SYN_ARCH2 of ND2_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_117;

architecture SYN_ARCH2 of ND2_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_116;

architecture SYN_ARCH2 of ND2_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_115;

architecture SYN_ARCH2 of ND2_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_114;

architecture SYN_ARCH2 of ND2_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_113;

architecture SYN_ARCH2 of ND2_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_112;

architecture SYN_ARCH2 of ND2_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_111;

architecture SYN_ARCH2 of ND2_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_110;

architecture SYN_ARCH2 of ND2_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_109;

architecture SYN_ARCH2 of ND2_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_108;

architecture SYN_ARCH2 of ND2_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_107;

architecture SYN_ARCH2 of ND2_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_106;

architecture SYN_ARCH2 of ND2_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_105;

architecture SYN_ARCH2 of ND2_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_104;

architecture SYN_ARCH2 of ND2_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_103;

architecture SYN_ARCH2 of ND2_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_102;

architecture SYN_ARCH2 of ND2_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_101;

architecture SYN_ARCH2 of ND2_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_100;

architecture SYN_ARCH2 of ND2_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_99;

architecture SYN_ARCH2 of ND2_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_98;

architecture SYN_ARCH2 of ND2_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_97;

architecture SYN_ARCH2 of ND2_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_96;

architecture SYN_ARCH2 of ND2_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95;

architecture SYN_ARCH2 of ND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94;

architecture SYN_ARCH2 of ND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH2 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH2 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH2 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH2 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH2 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH2 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH2 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH2 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH2 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH2 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH2 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH2 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH2 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH2 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH2 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH2 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH2 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH2 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH2 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH2 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH2 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH2 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH2 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH2 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH2 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH2 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH2 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH2 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH2 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH2 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH2 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH2 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH2 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH2 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH2 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH2 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH2 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH2 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH2 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH2 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH2 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH2 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH2 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH2 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH2 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH2 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH2 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH2 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH2 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH2 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH2 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH2 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH2 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH2 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH2 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH2 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH2 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH2 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH2 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH2 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH2 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH2 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH2 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH2 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH2 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH2 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH2 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH2 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH2 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH2 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH2 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH2 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH2 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH2 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH2 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH2 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH2 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH2 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH2 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH2 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH2 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH2 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH2 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH2 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH2 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH2 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH2 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH2 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH2 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH2 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH2 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH2 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH2 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_255 is

   port( A : in std_logic;  Y : out std_logic);

end IV_255;

architecture SYN_BEHAVIORAL of IV_255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_254 is

   port( A : in std_logic;  Y : out std_logic);

end IV_254;

architecture SYN_BEHAVIORAL of IV_254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_253 is

   port( A : in std_logic;  Y : out std_logic);

end IV_253;

architecture SYN_BEHAVIORAL of IV_253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_252 is

   port( A : in std_logic;  Y : out std_logic);

end IV_252;

architecture SYN_BEHAVIORAL of IV_252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_251 is

   port( A : in std_logic;  Y : out std_logic);

end IV_251;

architecture SYN_BEHAVIORAL of IV_251 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_250 is

   port( A : in std_logic;  Y : out std_logic);

end IV_250;

architecture SYN_BEHAVIORAL of IV_250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_249 is

   port( A : in std_logic;  Y : out std_logic);

end IV_249;

architecture SYN_BEHAVIORAL of IV_249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_248 is

   port( A : in std_logic;  Y : out std_logic);

end IV_248;

architecture SYN_BEHAVIORAL of IV_248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_247 is

   port( A : in std_logic;  Y : out std_logic);

end IV_247;

architecture SYN_BEHAVIORAL of IV_247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_246 is

   port( A : in std_logic;  Y : out std_logic);

end IV_246;

architecture SYN_BEHAVIORAL of IV_246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_245 is

   port( A : in std_logic;  Y : out std_logic);

end IV_245;

architecture SYN_BEHAVIORAL of IV_245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_244 is

   port( A : in std_logic;  Y : out std_logic);

end IV_244;

architecture SYN_BEHAVIORAL of IV_244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_243 is

   port( A : in std_logic;  Y : out std_logic);

end IV_243;

architecture SYN_BEHAVIORAL of IV_243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_242 is

   port( A : in std_logic;  Y : out std_logic);

end IV_242;

architecture SYN_BEHAVIORAL of IV_242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_241 is

   port( A : in std_logic;  Y : out std_logic);

end IV_241;

architecture SYN_BEHAVIORAL of IV_241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_240 is

   port( A : in std_logic;  Y : out std_logic);

end IV_240;

architecture SYN_BEHAVIORAL of IV_240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_239 is

   port( A : in std_logic;  Y : out std_logic);

end IV_239;

architecture SYN_BEHAVIORAL of IV_239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_238 is

   port( A : in std_logic;  Y : out std_logic);

end IV_238;

architecture SYN_BEHAVIORAL of IV_238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_237 is

   port( A : in std_logic;  Y : out std_logic);

end IV_237;

architecture SYN_BEHAVIORAL of IV_237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_236 is

   port( A : in std_logic;  Y : out std_logic);

end IV_236;

architecture SYN_BEHAVIORAL of IV_236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_235 is

   port( A : in std_logic;  Y : out std_logic);

end IV_235;

architecture SYN_BEHAVIORAL of IV_235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_234 is

   port( A : in std_logic;  Y : out std_logic);

end IV_234;

architecture SYN_BEHAVIORAL of IV_234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_233 is

   port( A : in std_logic;  Y : out std_logic);

end IV_233;

architecture SYN_BEHAVIORAL of IV_233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_232 is

   port( A : in std_logic;  Y : out std_logic);

end IV_232;

architecture SYN_BEHAVIORAL of IV_232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_231 is

   port( A : in std_logic;  Y : out std_logic);

end IV_231;

architecture SYN_BEHAVIORAL of IV_231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_230 is

   port( A : in std_logic;  Y : out std_logic);

end IV_230;

architecture SYN_BEHAVIORAL of IV_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_229 is

   port( A : in std_logic;  Y : out std_logic);

end IV_229;

architecture SYN_BEHAVIORAL of IV_229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_228 is

   port( A : in std_logic;  Y : out std_logic);

end IV_228;

architecture SYN_BEHAVIORAL of IV_228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_227 is

   port( A : in std_logic;  Y : out std_logic);

end IV_227;

architecture SYN_BEHAVIORAL of IV_227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_226 is

   port( A : in std_logic;  Y : out std_logic);

end IV_226;

architecture SYN_BEHAVIORAL of IV_226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_225 is

   port( A : in std_logic;  Y : out std_logic);

end IV_225;

architecture SYN_BEHAVIORAL of IV_225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_224 is

   port( A : in std_logic;  Y : out std_logic);

end IV_224;

architecture SYN_BEHAVIORAL of IV_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_223 is

   port( A : in std_logic;  Y : out std_logic);

end IV_223;

architecture SYN_BEHAVIORAL of IV_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_222 is

   port( A : in std_logic;  Y : out std_logic);

end IV_222;

architecture SYN_BEHAVIORAL of IV_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_221 is

   port( A : in std_logic;  Y : out std_logic);

end IV_221;

architecture SYN_BEHAVIORAL of IV_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_220 is

   port( A : in std_logic;  Y : out std_logic);

end IV_220;

architecture SYN_BEHAVIORAL of IV_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_219 is

   port( A : in std_logic;  Y : out std_logic);

end IV_219;

architecture SYN_BEHAVIORAL of IV_219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_218 is

   port( A : in std_logic;  Y : out std_logic);

end IV_218;

architecture SYN_BEHAVIORAL of IV_218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_217 is

   port( A : in std_logic;  Y : out std_logic);

end IV_217;

architecture SYN_BEHAVIORAL of IV_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_216 is

   port( A : in std_logic;  Y : out std_logic);

end IV_216;

architecture SYN_BEHAVIORAL of IV_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_215 is

   port( A : in std_logic;  Y : out std_logic);

end IV_215;

architecture SYN_BEHAVIORAL of IV_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_214 is

   port( A : in std_logic;  Y : out std_logic);

end IV_214;

architecture SYN_BEHAVIORAL of IV_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_213 is

   port( A : in std_logic;  Y : out std_logic);

end IV_213;

architecture SYN_BEHAVIORAL of IV_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_212 is

   port( A : in std_logic;  Y : out std_logic);

end IV_212;

architecture SYN_BEHAVIORAL of IV_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_211 is

   port( A : in std_logic;  Y : out std_logic);

end IV_211;

architecture SYN_BEHAVIORAL of IV_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_210 is

   port( A : in std_logic;  Y : out std_logic);

end IV_210;

architecture SYN_BEHAVIORAL of IV_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_209 is

   port( A : in std_logic;  Y : out std_logic);

end IV_209;

architecture SYN_BEHAVIORAL of IV_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_208 is

   port( A : in std_logic;  Y : out std_logic);

end IV_208;

architecture SYN_BEHAVIORAL of IV_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_207 is

   port( A : in std_logic;  Y : out std_logic);

end IV_207;

architecture SYN_BEHAVIORAL of IV_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_206 is

   port( A : in std_logic;  Y : out std_logic);

end IV_206;

architecture SYN_BEHAVIORAL of IV_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_205 is

   port( A : in std_logic;  Y : out std_logic);

end IV_205;

architecture SYN_BEHAVIORAL of IV_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_204 is

   port( A : in std_logic;  Y : out std_logic);

end IV_204;

architecture SYN_BEHAVIORAL of IV_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_203 is

   port( A : in std_logic;  Y : out std_logic);

end IV_203;

architecture SYN_BEHAVIORAL of IV_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_202 is

   port( A : in std_logic;  Y : out std_logic);

end IV_202;

architecture SYN_BEHAVIORAL of IV_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_201 is

   port( A : in std_logic;  Y : out std_logic);

end IV_201;

architecture SYN_BEHAVIORAL of IV_201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_200 is

   port( A : in std_logic;  Y : out std_logic);

end IV_200;

architecture SYN_BEHAVIORAL of IV_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_199 is

   port( A : in std_logic;  Y : out std_logic);

end IV_199;

architecture SYN_BEHAVIORAL of IV_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_198 is

   port( A : in std_logic;  Y : out std_logic);

end IV_198;

architecture SYN_BEHAVIORAL of IV_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_197 is

   port( A : in std_logic;  Y : out std_logic);

end IV_197;

architecture SYN_BEHAVIORAL of IV_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_196 is

   port( A : in std_logic;  Y : out std_logic);

end IV_196;

architecture SYN_BEHAVIORAL of IV_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_195 is

   port( A : in std_logic;  Y : out std_logic);

end IV_195;

architecture SYN_BEHAVIORAL of IV_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_194 is

   port( A : in std_logic;  Y : out std_logic);

end IV_194;

architecture SYN_BEHAVIORAL of IV_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_193 is

   port( A : in std_logic;  Y : out std_logic);

end IV_193;

architecture SYN_BEHAVIORAL of IV_193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_192 is

   port( A : in std_logic;  Y : out std_logic);

end IV_192;

architecture SYN_BEHAVIORAL of IV_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_191 is

   port( A : in std_logic;  Y : out std_logic);

end IV_191;

architecture SYN_BEHAVIORAL of IV_191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_190 is

   port( A : in std_logic;  Y : out std_logic);

end IV_190;

architecture SYN_BEHAVIORAL of IV_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_189 is

   port( A : in std_logic;  Y : out std_logic);

end IV_189;

architecture SYN_BEHAVIORAL of IV_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_188 is

   port( A : in std_logic;  Y : out std_logic);

end IV_188;

architecture SYN_BEHAVIORAL of IV_188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_187 is

   port( A : in std_logic;  Y : out std_logic);

end IV_187;

architecture SYN_BEHAVIORAL of IV_187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_186 is

   port( A : in std_logic;  Y : out std_logic);

end IV_186;

architecture SYN_BEHAVIORAL of IV_186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_185 is

   port( A : in std_logic;  Y : out std_logic);

end IV_185;

architecture SYN_BEHAVIORAL of IV_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_184 is

   port( A : in std_logic;  Y : out std_logic);

end IV_184;

architecture SYN_BEHAVIORAL of IV_184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_183 is

   port( A : in std_logic;  Y : out std_logic);

end IV_183;

architecture SYN_BEHAVIORAL of IV_183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_182 is

   port( A : in std_logic;  Y : out std_logic);

end IV_182;

architecture SYN_BEHAVIORAL of IV_182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_181 is

   port( A : in std_logic;  Y : out std_logic);

end IV_181;

architecture SYN_BEHAVIORAL of IV_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_180 is

   port( A : in std_logic;  Y : out std_logic);

end IV_180;

architecture SYN_BEHAVIORAL of IV_180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_179 is

   port( A : in std_logic;  Y : out std_logic);

end IV_179;

architecture SYN_BEHAVIORAL of IV_179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_178 is

   port( A : in std_logic;  Y : out std_logic);

end IV_178;

architecture SYN_BEHAVIORAL of IV_178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_177 is

   port( A : in std_logic;  Y : out std_logic);

end IV_177;

architecture SYN_BEHAVIORAL of IV_177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_176 is

   port( A : in std_logic;  Y : out std_logic);

end IV_176;

architecture SYN_BEHAVIORAL of IV_176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_175 is

   port( A : in std_logic;  Y : out std_logic);

end IV_175;

architecture SYN_BEHAVIORAL of IV_175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_174 is

   port( A : in std_logic;  Y : out std_logic);

end IV_174;

architecture SYN_BEHAVIORAL of IV_174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_173 is

   port( A : in std_logic;  Y : out std_logic);

end IV_173;

architecture SYN_BEHAVIORAL of IV_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_172 is

   port( A : in std_logic;  Y : out std_logic);

end IV_172;

architecture SYN_BEHAVIORAL of IV_172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_171 is

   port( A : in std_logic;  Y : out std_logic);

end IV_171;

architecture SYN_BEHAVIORAL of IV_171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_170 is

   port( A : in std_logic;  Y : out std_logic);

end IV_170;

architecture SYN_BEHAVIORAL of IV_170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_169 is

   port( A : in std_logic;  Y : out std_logic);

end IV_169;

architecture SYN_BEHAVIORAL of IV_169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_168 is

   port( A : in std_logic;  Y : out std_logic);

end IV_168;

architecture SYN_BEHAVIORAL of IV_168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_167 is

   port( A : in std_logic;  Y : out std_logic);

end IV_167;

architecture SYN_BEHAVIORAL of IV_167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_166 is

   port( A : in std_logic;  Y : out std_logic);

end IV_166;

architecture SYN_BEHAVIORAL of IV_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_165 is

   port( A : in std_logic;  Y : out std_logic);

end IV_165;

architecture SYN_BEHAVIORAL of IV_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_164 is

   port( A : in std_logic;  Y : out std_logic);

end IV_164;

architecture SYN_BEHAVIORAL of IV_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_163 is

   port( A : in std_logic;  Y : out std_logic);

end IV_163;

architecture SYN_BEHAVIORAL of IV_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_162 is

   port( A : in std_logic;  Y : out std_logic);

end IV_162;

architecture SYN_BEHAVIORAL of IV_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_161 is

   port( A : in std_logic;  Y : out std_logic);

end IV_161;

architecture SYN_BEHAVIORAL of IV_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_160 is

   port( A : in std_logic;  Y : out std_logic);

end IV_160;

architecture SYN_BEHAVIORAL of IV_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_159 is

   port( A : in std_logic;  Y : out std_logic);

end IV_159;

architecture SYN_BEHAVIORAL of IV_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_158 is

   port( A : in std_logic;  Y : out std_logic);

end IV_158;

architecture SYN_BEHAVIORAL of IV_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_157 is

   port( A : in std_logic;  Y : out std_logic);

end IV_157;

architecture SYN_BEHAVIORAL of IV_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_156 is

   port( A : in std_logic;  Y : out std_logic);

end IV_156;

architecture SYN_BEHAVIORAL of IV_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_155 is

   port( A : in std_logic;  Y : out std_logic);

end IV_155;

architecture SYN_BEHAVIORAL of IV_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_154 is

   port( A : in std_logic;  Y : out std_logic);

end IV_154;

architecture SYN_BEHAVIORAL of IV_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_153 is

   port( A : in std_logic;  Y : out std_logic);

end IV_153;

architecture SYN_BEHAVIORAL of IV_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_152 is

   port( A : in std_logic;  Y : out std_logic);

end IV_152;

architecture SYN_BEHAVIORAL of IV_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_151 is

   port( A : in std_logic;  Y : out std_logic);

end IV_151;

architecture SYN_BEHAVIORAL of IV_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_150 is

   port( A : in std_logic;  Y : out std_logic);

end IV_150;

architecture SYN_BEHAVIORAL of IV_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_149 is

   port( A : in std_logic;  Y : out std_logic);

end IV_149;

architecture SYN_BEHAVIORAL of IV_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_148 is

   port( A : in std_logic;  Y : out std_logic);

end IV_148;

architecture SYN_BEHAVIORAL of IV_148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_147 is

   port( A : in std_logic;  Y : out std_logic);

end IV_147;

architecture SYN_BEHAVIORAL of IV_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_146 is

   port( A : in std_logic;  Y : out std_logic);

end IV_146;

architecture SYN_BEHAVIORAL of IV_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_145 is

   port( A : in std_logic;  Y : out std_logic);

end IV_145;

architecture SYN_BEHAVIORAL of IV_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_144 is

   port( A : in std_logic;  Y : out std_logic);

end IV_144;

architecture SYN_BEHAVIORAL of IV_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_143 is

   port( A : in std_logic;  Y : out std_logic);

end IV_143;

architecture SYN_BEHAVIORAL of IV_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_142 is

   port( A : in std_logic;  Y : out std_logic);

end IV_142;

architecture SYN_BEHAVIORAL of IV_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_141 is

   port( A : in std_logic;  Y : out std_logic);

end IV_141;

architecture SYN_BEHAVIORAL of IV_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_140 is

   port( A : in std_logic;  Y : out std_logic);

end IV_140;

architecture SYN_BEHAVIORAL of IV_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_139 is

   port( A : in std_logic;  Y : out std_logic);

end IV_139;

architecture SYN_BEHAVIORAL of IV_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_138 is

   port( A : in std_logic;  Y : out std_logic);

end IV_138;

architecture SYN_BEHAVIORAL of IV_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_137 is

   port( A : in std_logic;  Y : out std_logic);

end IV_137;

architecture SYN_BEHAVIORAL of IV_137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_136 is

   port( A : in std_logic;  Y : out std_logic);

end IV_136;

architecture SYN_BEHAVIORAL of IV_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_135 is

   port( A : in std_logic;  Y : out std_logic);

end IV_135;

architecture SYN_BEHAVIORAL of IV_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_134 is

   port( A : in std_logic;  Y : out std_logic);

end IV_134;

architecture SYN_BEHAVIORAL of IV_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_133 is

   port( A : in std_logic;  Y : out std_logic);

end IV_133;

architecture SYN_BEHAVIORAL of IV_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_132 is

   port( A : in std_logic;  Y : out std_logic);

end IV_132;

architecture SYN_BEHAVIORAL of IV_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_131 is

   port( A : in std_logic;  Y : out std_logic);

end IV_131;

architecture SYN_BEHAVIORAL of IV_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_130 is

   port( A : in std_logic;  Y : out std_logic);

end IV_130;

architecture SYN_BEHAVIORAL of IV_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_129 is

   port( A : in std_logic;  Y : out std_logic);

end IV_129;

architecture SYN_BEHAVIORAL of IV_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_128 is

   port( A : in std_logic;  Y : out std_logic);

end IV_128;

architecture SYN_BEHAVIORAL of IV_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_127 is

   port( A : in std_logic;  Y : out std_logic);

end IV_127;

architecture SYN_BEHAVIORAL of IV_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_126 is

   port( A : in std_logic;  Y : out std_logic);

end IV_126;

architecture SYN_BEHAVIORAL of IV_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_125 is

   port( A : in std_logic;  Y : out std_logic);

end IV_125;

architecture SYN_BEHAVIORAL of IV_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_124 is

   port( A : in std_logic;  Y : out std_logic);

end IV_124;

architecture SYN_BEHAVIORAL of IV_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_123 is

   port( A : in std_logic;  Y : out std_logic);

end IV_123;

architecture SYN_BEHAVIORAL of IV_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_122 is

   port( A : in std_logic;  Y : out std_logic);

end IV_122;

architecture SYN_BEHAVIORAL of IV_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_121 is

   port( A : in std_logic;  Y : out std_logic);

end IV_121;

architecture SYN_BEHAVIORAL of IV_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_120 is

   port( A : in std_logic;  Y : out std_logic);

end IV_120;

architecture SYN_BEHAVIORAL of IV_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_119 is

   port( A : in std_logic;  Y : out std_logic);

end IV_119;

architecture SYN_BEHAVIORAL of IV_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_118 is

   port( A : in std_logic;  Y : out std_logic);

end IV_118;

architecture SYN_BEHAVIORAL of IV_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_117 is

   port( A : in std_logic;  Y : out std_logic);

end IV_117;

architecture SYN_BEHAVIORAL of IV_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_116 is

   port( A : in std_logic;  Y : out std_logic);

end IV_116;

architecture SYN_BEHAVIORAL of IV_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_115 is

   port( A : in std_logic;  Y : out std_logic);

end IV_115;

architecture SYN_BEHAVIORAL of IV_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_114 is

   port( A : in std_logic;  Y : out std_logic);

end IV_114;

architecture SYN_BEHAVIORAL of IV_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_113 is

   port( A : in std_logic;  Y : out std_logic);

end IV_113;

architecture SYN_BEHAVIORAL of IV_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_112 is

   port( A : in std_logic;  Y : out std_logic);

end IV_112;

architecture SYN_BEHAVIORAL of IV_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_111 is

   port( A : in std_logic;  Y : out std_logic);

end IV_111;

architecture SYN_BEHAVIORAL of IV_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_110 is

   port( A : in std_logic;  Y : out std_logic);

end IV_110;

architecture SYN_BEHAVIORAL of IV_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_109 is

   port( A : in std_logic;  Y : out std_logic);

end IV_109;

architecture SYN_BEHAVIORAL of IV_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_108 is

   port( A : in std_logic;  Y : out std_logic);

end IV_108;

architecture SYN_BEHAVIORAL of IV_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_107 is

   port( A : in std_logic;  Y : out std_logic);

end IV_107;

architecture SYN_BEHAVIORAL of IV_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_106 is

   port( A : in std_logic;  Y : out std_logic);

end IV_106;

architecture SYN_BEHAVIORAL of IV_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_105 is

   port( A : in std_logic;  Y : out std_logic);

end IV_105;

architecture SYN_BEHAVIORAL of IV_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_104 is

   port( A : in std_logic;  Y : out std_logic);

end IV_104;

architecture SYN_BEHAVIORAL of IV_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_103 is

   port( A : in std_logic;  Y : out std_logic);

end IV_103;

architecture SYN_BEHAVIORAL of IV_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_102 is

   port( A : in std_logic;  Y : out std_logic);

end IV_102;

architecture SYN_BEHAVIORAL of IV_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_101 is

   port( A : in std_logic;  Y : out std_logic);

end IV_101;

architecture SYN_BEHAVIORAL of IV_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_100 is

   port( A : in std_logic;  Y : out std_logic);

end IV_100;

architecture SYN_BEHAVIORAL of IV_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_99 is

   port( A : in std_logic;  Y : out std_logic);

end IV_99;

architecture SYN_BEHAVIORAL of IV_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_98 is

   port( A : in std_logic;  Y : out std_logic);

end IV_98;

architecture SYN_BEHAVIORAL of IV_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_97 is

   port( A : in std_logic;  Y : out std_logic);

end IV_97;

architecture SYN_BEHAVIORAL of IV_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_96 is

   port( A : in std_logic;  Y : out std_logic);

end IV_96;

architecture SYN_BEHAVIORAL of IV_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_95 is

   port( A : in std_logic;  Y : out std_logic);

end IV_95;

architecture SYN_BEHAVIORAL of IV_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_94 is

   port( A : in std_logic;  Y : out std_logic);

end IV_94;

architecture SYN_BEHAVIORAL of IV_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_93 is

   port( A : in std_logic;  Y : out std_logic);

end IV_93;

architecture SYN_BEHAVIORAL of IV_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_92 is

   port( A : in std_logic;  Y : out std_logic);

end IV_92;

architecture SYN_BEHAVIORAL of IV_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_91 is

   port( A : in std_logic;  Y : out std_logic);

end IV_91;

architecture SYN_BEHAVIORAL of IV_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_90 is

   port( A : in std_logic;  Y : out std_logic);

end IV_90;

architecture SYN_BEHAVIORAL of IV_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_89 is

   port( A : in std_logic;  Y : out std_logic);

end IV_89;

architecture SYN_BEHAVIORAL of IV_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_88 is

   port( A : in std_logic;  Y : out std_logic);

end IV_88;

architecture SYN_BEHAVIORAL of IV_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_87 is

   port( A : in std_logic;  Y : out std_logic);

end IV_87;

architecture SYN_BEHAVIORAL of IV_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_86 is

   port( A : in std_logic;  Y : out std_logic);

end IV_86;

architecture SYN_BEHAVIORAL of IV_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_85 is

   port( A : in std_logic;  Y : out std_logic);

end IV_85;

architecture SYN_BEHAVIORAL of IV_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_84 is

   port( A : in std_logic;  Y : out std_logic);

end IV_84;

architecture SYN_BEHAVIORAL of IV_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_83 is

   port( A : in std_logic;  Y : out std_logic);

end IV_83;

architecture SYN_BEHAVIORAL of IV_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_82 is

   port( A : in std_logic;  Y : out std_logic);

end IV_82;

architecture SYN_BEHAVIORAL of IV_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_81 is

   port( A : in std_logic;  Y : out std_logic);

end IV_81;

architecture SYN_BEHAVIORAL of IV_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_80 is

   port( A : in std_logic;  Y : out std_logic);

end IV_80;

architecture SYN_BEHAVIORAL of IV_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_79 is

   port( A : in std_logic;  Y : out std_logic);

end IV_79;

architecture SYN_BEHAVIORAL of IV_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_78 is

   port( A : in std_logic;  Y : out std_logic);

end IV_78;

architecture SYN_BEHAVIORAL of IV_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_77 is

   port( A : in std_logic;  Y : out std_logic);

end IV_77;

architecture SYN_BEHAVIORAL of IV_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_76 is

   port( A : in std_logic;  Y : out std_logic);

end IV_76;

architecture SYN_BEHAVIORAL of IV_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_75 is

   port( A : in std_logic;  Y : out std_logic);

end IV_75;

architecture SYN_BEHAVIORAL of IV_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_74 is

   port( A : in std_logic;  Y : out std_logic);

end IV_74;

architecture SYN_BEHAVIORAL of IV_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_73 is

   port( A : in std_logic;  Y : out std_logic);

end IV_73;

architecture SYN_BEHAVIORAL of IV_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_72 is

   port( A : in std_logic;  Y : out std_logic);

end IV_72;

architecture SYN_BEHAVIORAL of IV_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_71 is

   port( A : in std_logic;  Y : out std_logic);

end IV_71;

architecture SYN_BEHAVIORAL of IV_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_70 is

   port( A : in std_logic;  Y : out std_logic);

end IV_70;

architecture SYN_BEHAVIORAL of IV_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_69 is

   port( A : in std_logic;  Y : out std_logic);

end IV_69;

architecture SYN_BEHAVIORAL of IV_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_68 is

   port( A : in std_logic;  Y : out std_logic);

end IV_68;

architecture SYN_BEHAVIORAL of IV_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_67 is

   port( A : in std_logic;  Y : out std_logic);

end IV_67;

architecture SYN_BEHAVIORAL of IV_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_66 is

   port( A : in std_logic;  Y : out std_logic);

end IV_66;

architecture SYN_BEHAVIORAL of IV_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_65 is

   port( A : in std_logic;  Y : out std_logic);

end IV_65;

architecture SYN_BEHAVIORAL of IV_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_64 is

   port( A : in std_logic;  Y : out std_logic);

end IV_64;

architecture SYN_BEHAVIORAL of IV_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_255 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_255;

architecture SYN_STRUCTURAL of MUX21_255 is

   component ND2_763
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_764
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_765
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_255
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_255 port map( A => S, Y => SB);
   UND1 : ND2_765 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_764 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_763 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_254 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_254;

architecture SYN_STRUCTURAL of MUX21_254 is

   component ND2_760
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_761
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_762
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_254
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_254 port map( A => S, Y => SB);
   UND1 : ND2_762 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_761 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_760 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_253 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_253;

architecture SYN_STRUCTURAL of MUX21_253 is

   component ND2_757
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_758
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_759
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_253
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_253 port map( A => S, Y => SB);
   UND1 : ND2_759 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_758 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_757 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_252 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_252;

architecture SYN_STRUCTURAL of MUX21_252 is

   component ND2_754
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_755
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_756
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_252
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_252 port map( A => S, Y => SB);
   UND1 : ND2_756 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_755 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_754 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_251 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_251;

architecture SYN_STRUCTURAL of MUX21_251 is

   component ND2_751
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_752
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_753
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_251
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_251 port map( A => S, Y => SB);
   UND1 : ND2_753 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_752 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_751 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_250 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_250;

architecture SYN_STRUCTURAL of MUX21_250 is

   component ND2_748
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_749
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_750
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_250
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_250 port map( A => S, Y => SB);
   UND1 : ND2_750 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_749 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_748 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_249 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_249;

architecture SYN_STRUCTURAL of MUX21_249 is

   component ND2_745
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_746
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_747
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_249
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_249 port map( A => S, Y => SB);
   UND1 : ND2_747 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_746 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_745 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_248 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_248;

architecture SYN_STRUCTURAL of MUX21_248 is

   component ND2_742
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_743
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_744
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_248
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_248 port map( A => S, Y => SB);
   UND1 : ND2_744 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_743 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_742 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_247 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_247;

architecture SYN_STRUCTURAL of MUX21_247 is

   component ND2_739
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_740
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_741
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_247
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_247 port map( A => S, Y => SB);
   UND1 : ND2_741 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_740 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_739 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_246 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_246;

architecture SYN_STRUCTURAL of MUX21_246 is

   component ND2_736
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_737
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_738
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_246
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_246 port map( A => S, Y => SB);
   UND1 : ND2_738 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_737 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_736 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_245 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_245;

architecture SYN_STRUCTURAL of MUX21_245 is

   component ND2_733
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_734
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_735
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_245
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_245 port map( A => S, Y => SB);
   UND1 : ND2_735 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_734 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_733 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_244 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_244;

architecture SYN_STRUCTURAL of MUX21_244 is

   component ND2_730
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_731
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_732
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_244
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_244 port map( A => S, Y => SB);
   UND1 : ND2_732 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_731 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_730 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_243 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_243;

architecture SYN_STRUCTURAL of MUX21_243 is

   component ND2_727
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_728
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_729
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_243
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_243 port map( A => S, Y => SB);
   UND1 : ND2_729 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_728 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_727 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_242 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_242;

architecture SYN_STRUCTURAL of MUX21_242 is

   component ND2_724
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_725
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_726
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_242
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_242 port map( A => S, Y => SB);
   UND1 : ND2_726 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_725 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_724 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_241 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_241;

architecture SYN_STRUCTURAL of MUX21_241 is

   component ND2_721
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_722
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_723
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_241
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_241 port map( A => S, Y => SB);
   UND1 : ND2_723 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_722 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_721 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_240 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_240;

architecture SYN_STRUCTURAL of MUX21_240 is

   component ND2_718
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_719
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_720
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_240
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_240 port map( A => S, Y => SB);
   UND1 : ND2_720 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_719 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_718 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_239 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_239;

architecture SYN_STRUCTURAL of MUX21_239 is

   component ND2_715
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_716
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_717
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_239
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_239 port map( A => S, Y => SB);
   UND1 : ND2_717 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_716 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_715 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_238 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_238;

architecture SYN_STRUCTURAL of MUX21_238 is

   component ND2_712
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_713
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_714
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_238
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_238 port map( A => S, Y => SB);
   UND1 : ND2_714 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_713 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_712 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_237 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_237;

architecture SYN_STRUCTURAL of MUX21_237 is

   component ND2_709
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_710
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_711
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_237
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_237 port map( A => S, Y => SB);
   UND1 : ND2_711 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_710 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_709 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_236 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_236;

architecture SYN_STRUCTURAL of MUX21_236 is

   component ND2_706
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_707
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_708
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_236
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_236 port map( A => S, Y => SB);
   UND1 : ND2_708 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_707 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_706 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_235 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_235;

architecture SYN_STRUCTURAL of MUX21_235 is

   component ND2_703
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_704
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_705
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_235
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_235 port map( A => S, Y => SB);
   UND1 : ND2_705 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_704 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_703 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_234 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_234;

architecture SYN_STRUCTURAL of MUX21_234 is

   component ND2_700
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_701
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_702
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_234
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_234 port map( A => S, Y => SB);
   UND1 : ND2_702 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_701 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_700 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_233 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_233;

architecture SYN_STRUCTURAL of MUX21_233 is

   component ND2_697
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_698
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_699
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_233
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_233 port map( A => S, Y => SB);
   UND1 : ND2_699 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_698 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_697 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_232 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_232;

architecture SYN_STRUCTURAL of MUX21_232 is

   component ND2_694
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_695
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_696
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_232
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_232 port map( A => S, Y => SB);
   UND1 : ND2_696 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_695 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_694 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_231 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_231;

architecture SYN_STRUCTURAL of MUX21_231 is

   component ND2_691
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_692
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_693
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_231
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_231 port map( A => S, Y => SB);
   UND1 : ND2_693 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_692 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_691 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_230 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_230;

architecture SYN_STRUCTURAL of MUX21_230 is

   component ND2_688
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_689
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_690
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_230
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_230 port map( A => S, Y => SB);
   UND1 : ND2_690 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_689 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_688 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_229 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_229;

architecture SYN_STRUCTURAL of MUX21_229 is

   component ND2_685
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_686
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_687
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_229
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_229 port map( A => S, Y => SB);
   UND1 : ND2_687 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_686 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_685 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_228 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_228;

architecture SYN_STRUCTURAL of MUX21_228 is

   component ND2_682
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_683
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_684
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_228
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_228 port map( A => S, Y => SB);
   UND1 : ND2_684 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_683 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_682 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_227 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_227;

architecture SYN_STRUCTURAL of MUX21_227 is

   component ND2_679
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_680
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_681
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_227
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_227 port map( A => S, Y => SB);
   UND1 : ND2_681 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_680 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_679 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_226 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_226;

architecture SYN_STRUCTURAL of MUX21_226 is

   component ND2_676
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_677
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_678
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_226
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_226 port map( A => S, Y => SB);
   UND1 : ND2_678 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_677 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_676 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_225 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_225;

architecture SYN_STRUCTURAL of MUX21_225 is

   component ND2_673
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_674
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_675
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_225
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_225 port map( A => S, Y => SB);
   UND1 : ND2_675 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_674 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_673 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_224 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_224;

architecture SYN_STRUCTURAL of MUX21_224 is

   component ND2_670
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_671
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_672
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_224
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_224 port map( A => S, Y => SB);
   UND1 : ND2_672 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_671 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_670 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_223 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_223;

architecture SYN_STRUCTURAL of MUX21_223 is

   component ND2_667
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_668
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_669
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_223
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_223 port map( A => S, Y => SB);
   UND1 : ND2_669 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_668 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_667 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_222 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_222;

architecture SYN_STRUCTURAL of MUX21_222 is

   component ND2_664
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_665
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_666
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_222
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_222 port map( A => S, Y => SB);
   UND1 : ND2_666 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_665 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_664 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_221 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_221;

architecture SYN_STRUCTURAL of MUX21_221 is

   component ND2_661
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_662
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_663
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_221
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_221 port map( A => S, Y => SB);
   UND1 : ND2_663 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_662 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_661 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_220 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_220;

architecture SYN_STRUCTURAL of MUX21_220 is

   component ND2_658
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_659
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_660
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_220
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_220 port map( A => S, Y => SB);
   UND1 : ND2_660 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_659 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_658 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_219 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_219;

architecture SYN_STRUCTURAL of MUX21_219 is

   component ND2_655
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_656
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_657
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_219
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_219 port map( A => S, Y => SB);
   UND1 : ND2_657 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_656 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_655 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_218 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_218;

architecture SYN_STRUCTURAL of MUX21_218 is

   component ND2_652
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_653
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_654
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_218
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_218 port map( A => S, Y => SB);
   UND1 : ND2_654 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_653 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_652 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_217;

architecture SYN_STRUCTURAL of MUX21_217 is

   component ND2_649
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_650
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_651
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_217
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_217 port map( A => S, Y => SB);
   UND1 : ND2_651 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_650 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_649 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_216;

architecture SYN_STRUCTURAL of MUX21_216 is

   component ND2_646
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_647
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_648
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_216
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_216 port map( A => S, Y => SB);
   UND1 : ND2_648 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_647 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_646 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_215;

architecture SYN_STRUCTURAL of MUX21_215 is

   component ND2_643
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_644
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_645
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_215
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_215 port map( A => S, Y => SB);
   UND1 : ND2_645 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_644 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_643 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_214;

architecture SYN_STRUCTURAL of MUX21_214 is

   component ND2_640
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_641
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_642
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_214
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_214 port map( A => S, Y => SB);
   UND1 : ND2_642 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_641 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_640 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_213;

architecture SYN_STRUCTURAL of MUX21_213 is

   component ND2_637
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_638
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_639
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_213
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_213 port map( A => S, Y => SB);
   UND1 : ND2_639 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_638 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_637 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_212;

architecture SYN_STRUCTURAL of MUX21_212 is

   component ND2_634
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_635
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_636
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_212
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_212 port map( A => S, Y => SB);
   UND1 : ND2_636 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_635 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_634 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_211;

architecture SYN_STRUCTURAL of MUX21_211 is

   component ND2_631
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_632
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_633
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_211
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_211 port map( A => S, Y => SB);
   UND1 : ND2_633 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_632 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_631 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_210;

architecture SYN_STRUCTURAL of MUX21_210 is

   component ND2_628
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_629
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_630
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_210
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_210 port map( A => S, Y => SB);
   UND1 : ND2_630 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_629 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_628 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_209;

architecture SYN_STRUCTURAL of MUX21_209 is

   component ND2_625
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_626
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_627
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_209
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_209 port map( A => S, Y => SB);
   UND1 : ND2_627 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_626 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_625 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_208;

architecture SYN_STRUCTURAL of MUX21_208 is

   component ND2_622
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_623
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_624
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_208
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_208 port map( A => S, Y => SB);
   UND1 : ND2_624 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_623 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_622 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_207;

architecture SYN_STRUCTURAL of MUX21_207 is

   component ND2_619
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_620
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_621
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_207
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_207 port map( A => S, Y => SB);
   UND1 : ND2_621 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_620 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_619 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_206;

architecture SYN_STRUCTURAL of MUX21_206 is

   component ND2_616
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_617
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_618
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_206
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_206 port map( A => S, Y => SB);
   UND1 : ND2_618 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_617 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_616 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_205;

architecture SYN_STRUCTURAL of MUX21_205 is

   component ND2_613
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_614
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_615
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_205
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_205 port map( A => S, Y => SB);
   UND1 : ND2_615 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_614 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_613 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_204;

architecture SYN_STRUCTURAL of MUX21_204 is

   component ND2_610
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_611
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_612
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_204
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_204 port map( A => S, Y => SB);
   UND1 : ND2_612 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_611 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_610 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_203;

architecture SYN_STRUCTURAL of MUX21_203 is

   component ND2_607
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_608
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_609
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_203
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_203 port map( A => S, Y => SB);
   UND1 : ND2_609 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_608 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_607 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_202;

architecture SYN_STRUCTURAL of MUX21_202 is

   component ND2_604
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_605
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_606
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_202
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_202 port map( A => S, Y => SB);
   UND1 : ND2_606 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_605 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_604 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_201;

architecture SYN_STRUCTURAL of MUX21_201 is

   component ND2_601
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_602
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_603
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_201
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_201 port map( A => S, Y => SB);
   UND1 : ND2_603 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_602 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_601 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_200;

architecture SYN_STRUCTURAL of MUX21_200 is

   component ND2_598
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_599
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_600
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_200
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_200 port map( A => S, Y => SB);
   UND1 : ND2_600 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_599 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_598 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_199;

architecture SYN_STRUCTURAL of MUX21_199 is

   component ND2_595
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_596
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_597
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_199
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_199 port map( A => S, Y => SB);
   UND1 : ND2_597 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_596 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_595 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_198;

architecture SYN_STRUCTURAL of MUX21_198 is

   component ND2_592
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_593
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_594
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_198
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_198 port map( A => S, Y => SB);
   UND1 : ND2_594 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_593 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_592 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_197;

architecture SYN_STRUCTURAL of MUX21_197 is

   component ND2_589
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_590
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_591
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_197
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_197 port map( A => S, Y => SB);
   UND1 : ND2_591 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_590 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_589 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_196;

architecture SYN_STRUCTURAL of MUX21_196 is

   component ND2_586
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_587
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_588
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_196
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_196 port map( A => S, Y => SB);
   UND1 : ND2_588 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_587 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_586 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_195;

architecture SYN_STRUCTURAL of MUX21_195 is

   component ND2_583
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_584
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_585
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_195
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_195 port map( A => S, Y => SB);
   UND1 : ND2_585 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_584 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_583 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_194;

architecture SYN_STRUCTURAL of MUX21_194 is

   component ND2_580
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_581
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_582
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_194
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_194 port map( A => S, Y => SB);
   UND1 : ND2_582 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_581 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_580 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_193;

architecture SYN_STRUCTURAL of MUX21_193 is

   component ND2_577
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_578
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_579
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_193
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_193 port map( A => S, Y => SB);
   UND1 : ND2_579 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_578 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_577 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_192;

architecture SYN_STRUCTURAL of MUX21_192 is

   component ND2_574
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_575
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_576
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_192
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_192 port map( A => S, Y => SB);
   UND1 : ND2_576 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_575 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_574 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_191;

architecture SYN_STRUCTURAL of MUX21_191 is

   component ND2_571
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_572
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_573
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_191
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_191 port map( A => S, Y => SB);
   UND1 : ND2_573 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_572 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_571 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_190;

architecture SYN_STRUCTURAL of MUX21_190 is

   component ND2_568
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_569
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_570
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_190
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_190 port map( A => S, Y => SB);
   UND1 : ND2_570 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_569 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_568 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_189;

architecture SYN_STRUCTURAL of MUX21_189 is

   component ND2_565
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_566
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_567
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_189
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_189 port map( A => S, Y => SB);
   UND1 : ND2_567 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_566 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_565 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_188;

architecture SYN_STRUCTURAL of MUX21_188 is

   component ND2_562
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_563
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_564
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_188
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_188 port map( A => S, Y => SB);
   UND1 : ND2_564 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_563 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_562 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_187;

architecture SYN_STRUCTURAL of MUX21_187 is

   component ND2_559
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_560
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_561
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_187
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_187 port map( A => S, Y => SB);
   UND1 : ND2_561 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_560 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_559 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_186;

architecture SYN_STRUCTURAL of MUX21_186 is

   component ND2_556
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_557
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_558
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_186
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_186 port map( A => S, Y => SB);
   UND1 : ND2_558 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_557 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_556 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_185;

architecture SYN_STRUCTURAL of MUX21_185 is

   component ND2_553
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_554
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_555
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_185
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_185 port map( A => S, Y => SB);
   UND1 : ND2_555 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_554 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_553 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_184;

architecture SYN_STRUCTURAL of MUX21_184 is

   component ND2_550
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_551
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_552
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_184
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_184 port map( A => S, Y => SB);
   UND1 : ND2_552 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_551 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_550 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_183;

architecture SYN_STRUCTURAL of MUX21_183 is

   component ND2_547
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_548
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_549
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_183
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_183 port map( A => S, Y => SB);
   UND1 : ND2_549 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_548 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_547 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_182;

architecture SYN_STRUCTURAL of MUX21_182 is

   component ND2_544
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_545
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_546
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_182
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_182 port map( A => S, Y => SB);
   UND1 : ND2_546 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_545 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_544 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_181;

architecture SYN_STRUCTURAL of MUX21_181 is

   component ND2_541
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_542
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_543
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_181
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_181 port map( A => S, Y => SB);
   UND1 : ND2_543 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_542 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_541 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_180;

architecture SYN_STRUCTURAL of MUX21_180 is

   component ND2_538
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_539
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_540
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_180
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_180 port map( A => S, Y => SB);
   UND1 : ND2_540 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_539 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_538 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_179;

architecture SYN_STRUCTURAL of MUX21_179 is

   component ND2_535
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_536
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_537
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_179
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_179 port map( A => S, Y => SB);
   UND1 : ND2_537 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_536 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_535 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_178;

architecture SYN_STRUCTURAL of MUX21_178 is

   component ND2_532
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_533
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_534
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_178
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_178 port map( A => S, Y => SB);
   UND1 : ND2_534 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_533 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_532 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_177;

architecture SYN_STRUCTURAL of MUX21_177 is

   component ND2_529
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_530
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_531
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_177
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_177 port map( A => S, Y => SB);
   UND1 : ND2_531 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_530 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_529 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_176;

architecture SYN_STRUCTURAL of MUX21_176 is

   component ND2_526
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_527
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_528
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_176
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_176 port map( A => S, Y => SB);
   UND1 : ND2_528 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_527 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_526 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_175;

architecture SYN_STRUCTURAL of MUX21_175 is

   component ND2_523
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_524
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_525
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_175
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_175 port map( A => S, Y => SB);
   UND1 : ND2_525 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_524 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_523 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_174;

architecture SYN_STRUCTURAL of MUX21_174 is

   component ND2_520
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_521
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_522
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_174
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_174 port map( A => S, Y => SB);
   UND1 : ND2_522 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_521 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_520 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_173;

architecture SYN_STRUCTURAL of MUX21_173 is

   component ND2_517
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_518
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_519
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_173
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_173 port map( A => S, Y => SB);
   UND1 : ND2_519 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_518 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_517 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_172;

architecture SYN_STRUCTURAL of MUX21_172 is

   component ND2_514
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_515
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_516
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_172
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_172 port map( A => S, Y => SB);
   UND1 : ND2_516 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_515 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_514 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_171;

architecture SYN_STRUCTURAL of MUX21_171 is

   component ND2_511
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_512
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_513
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_171
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_171 port map( A => S, Y => SB);
   UND1 : ND2_513 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_512 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_511 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_170;

architecture SYN_STRUCTURAL of MUX21_170 is

   component ND2_508
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_509
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_510
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_170
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_170 port map( A => S, Y => SB);
   UND1 : ND2_510 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_509 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_508 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_169;

architecture SYN_STRUCTURAL of MUX21_169 is

   component ND2_505
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_506
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_507
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_169
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_169 port map( A => S, Y => SB);
   UND1 : ND2_507 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_506 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_505 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_168;

architecture SYN_STRUCTURAL of MUX21_168 is

   component ND2_502
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_503
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_504
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_168
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_168 port map( A => S, Y => SB);
   UND1 : ND2_504 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_503 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_502 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_167;

architecture SYN_STRUCTURAL of MUX21_167 is

   component ND2_499
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_500
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_501
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_167
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_167 port map( A => S, Y => SB);
   UND1 : ND2_501 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_500 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_499 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_166;

architecture SYN_STRUCTURAL of MUX21_166 is

   component ND2_496
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_497
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_498
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_166
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_166 port map( A => S, Y => SB);
   UND1 : ND2_498 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_497 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_496 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_165;

architecture SYN_STRUCTURAL of MUX21_165 is

   component ND2_493
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_494
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_495
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_165
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_165 port map( A => S, Y => SB);
   UND1 : ND2_495 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_494 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_493 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_164;

architecture SYN_STRUCTURAL of MUX21_164 is

   component ND2_490
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_491
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_492
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_164
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_164 port map( A => S, Y => SB);
   UND1 : ND2_492 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_491 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_490 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_163;

architecture SYN_STRUCTURAL of MUX21_163 is

   component ND2_487
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_488
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_489
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_163
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_163 port map( A => S, Y => SB);
   UND1 : ND2_489 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_488 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_487 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_162;

architecture SYN_STRUCTURAL of MUX21_162 is

   component ND2_484
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_485
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_486
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_162
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_162 port map( A => S, Y => SB);
   UND1 : ND2_486 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_485 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_484 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_161;

architecture SYN_STRUCTURAL of MUX21_161 is

   component ND2_481
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_482
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_483
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_161
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_161 port map( A => S, Y => SB);
   UND1 : ND2_483 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_482 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_481 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_160;

architecture SYN_STRUCTURAL of MUX21_160 is

   component ND2_478
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_479
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_480
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_160
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_160 port map( A => S, Y => SB);
   UND1 : ND2_480 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_479 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_478 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_159;

architecture SYN_STRUCTURAL of MUX21_159 is

   component ND2_475
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_476
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_477
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_159
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_159 port map( A => S, Y => SB);
   UND1 : ND2_477 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_476 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_475 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_158;

architecture SYN_STRUCTURAL of MUX21_158 is

   component ND2_472
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_473
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_474
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_158
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_158 port map( A => S, Y => SB);
   UND1 : ND2_474 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_473 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_472 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_157;

architecture SYN_STRUCTURAL of MUX21_157 is

   component ND2_469
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_470
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_471
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_157
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_157 port map( A => S, Y => SB);
   UND1 : ND2_471 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_470 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_469 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_156;

architecture SYN_STRUCTURAL of MUX21_156 is

   component ND2_466
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_467
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_468
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_156
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_156 port map( A => S, Y => SB);
   UND1 : ND2_468 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_467 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_466 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_155;

architecture SYN_STRUCTURAL of MUX21_155 is

   component ND2_463
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_464
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_465
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_155
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_155 port map( A => S, Y => SB);
   UND1 : ND2_465 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_464 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_463 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_154;

architecture SYN_STRUCTURAL of MUX21_154 is

   component ND2_460
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_461
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_462
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_154
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_154 port map( A => S, Y => SB);
   UND1 : ND2_462 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_461 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_460 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_153;

architecture SYN_STRUCTURAL of MUX21_153 is

   component ND2_457
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_458
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_459
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_153
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_153 port map( A => S, Y => SB);
   UND1 : ND2_459 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_458 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_457 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_152;

architecture SYN_STRUCTURAL of MUX21_152 is

   component ND2_454
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_455
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_456
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_152
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_152 port map( A => S, Y => SB);
   UND1 : ND2_456 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_455 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_454 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_151;

architecture SYN_STRUCTURAL of MUX21_151 is

   component ND2_451
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_452
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_453
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_151
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_151 port map( A => S, Y => SB);
   UND1 : ND2_453 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_452 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_451 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_150;

architecture SYN_STRUCTURAL of MUX21_150 is

   component ND2_448
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_449
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_450
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_150
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_150 port map( A => S, Y => SB);
   UND1 : ND2_450 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_449 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_448 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_149;

architecture SYN_STRUCTURAL of MUX21_149 is

   component ND2_445
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_446
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_447
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_149
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_149 port map( A => S, Y => SB);
   UND1 : ND2_447 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_446 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_445 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_148;

architecture SYN_STRUCTURAL of MUX21_148 is

   component ND2_442
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_443
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_444
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_148
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_148 port map( A => S, Y => SB);
   UND1 : ND2_444 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_443 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_442 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_147;

architecture SYN_STRUCTURAL of MUX21_147 is

   component ND2_439
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_440
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_441
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_147
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_147 port map( A => S, Y => SB);
   UND1 : ND2_441 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_440 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_439 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_146;

architecture SYN_STRUCTURAL of MUX21_146 is

   component ND2_436
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_437
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_438
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_146
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_146 port map( A => S, Y => SB);
   UND1 : ND2_438 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_437 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_436 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_145;

architecture SYN_STRUCTURAL of MUX21_145 is

   component ND2_433
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_434
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_435
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_145
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_145 port map( A => S, Y => SB);
   UND1 : ND2_435 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_434 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_433 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_144;

architecture SYN_STRUCTURAL of MUX21_144 is

   component ND2_430
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_431
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_432
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_144
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_144 port map( A => S, Y => SB);
   UND1 : ND2_432 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_431 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_430 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_143;

architecture SYN_STRUCTURAL of MUX21_143 is

   component ND2_427
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_428
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_429
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_143
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_143 port map( A => S, Y => SB);
   UND1 : ND2_429 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_428 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_427 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_142;

architecture SYN_STRUCTURAL of MUX21_142 is

   component ND2_424
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_425
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_426
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_142
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_142 port map( A => S, Y => SB);
   UND1 : ND2_426 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_425 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_424 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_141;

architecture SYN_STRUCTURAL of MUX21_141 is

   component ND2_421
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_422
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_423
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_141
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_141 port map( A => S, Y => SB);
   UND1 : ND2_423 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_422 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_421 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_140;

architecture SYN_STRUCTURAL of MUX21_140 is

   component ND2_418
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_419
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_420
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_140
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_140 port map( A => S, Y => SB);
   UND1 : ND2_420 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_419 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_418 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_139;

architecture SYN_STRUCTURAL of MUX21_139 is

   component ND2_415
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_416
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_417
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_139
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_139 port map( A => S, Y => SB);
   UND1 : ND2_417 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_416 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_415 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_138;

architecture SYN_STRUCTURAL of MUX21_138 is

   component ND2_412
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_413
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_414
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_138
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_138 port map( A => S, Y => SB);
   UND1 : ND2_414 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_413 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_412 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_137;

architecture SYN_STRUCTURAL of MUX21_137 is

   component ND2_409
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_410
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_411
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_137
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_137 port map( A => S, Y => SB);
   UND1 : ND2_411 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_410 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_409 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_136;

architecture SYN_STRUCTURAL of MUX21_136 is

   component ND2_406
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_407
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_408
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_136
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_136 port map( A => S, Y => SB);
   UND1 : ND2_408 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_407 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_406 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_135;

architecture SYN_STRUCTURAL of MUX21_135 is

   component ND2_403
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_404
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_405
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_135
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_135 port map( A => S, Y => SB);
   UND1 : ND2_405 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_404 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_403 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_134;

architecture SYN_STRUCTURAL of MUX21_134 is

   component ND2_400
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_401
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_402
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_134
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_134 port map( A => S, Y => SB);
   UND1 : ND2_402 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_401 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_400 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_133;

architecture SYN_STRUCTURAL of MUX21_133 is

   component ND2_397
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_398
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_399
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_133
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_133 port map( A => S, Y => SB);
   UND1 : ND2_399 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_398 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_397 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_132;

architecture SYN_STRUCTURAL of MUX21_132 is

   component ND2_394
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_395
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_396
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_132
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_132 port map( A => S, Y => SB);
   UND1 : ND2_396 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_395 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_394 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_131;

architecture SYN_STRUCTURAL of MUX21_131 is

   component ND2_391
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_392
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_393
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_131
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_131 port map( A => S, Y => SB);
   UND1 : ND2_393 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_392 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_391 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_130;

architecture SYN_STRUCTURAL of MUX21_130 is

   component ND2_388
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_389
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_390
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_130
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_130 port map( A => S, Y => SB);
   UND1 : ND2_390 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_389 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_388 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_129;

architecture SYN_STRUCTURAL of MUX21_129 is

   component ND2_385
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_386
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_387
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_129
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_129 port map( A => S, Y => SB);
   UND1 : ND2_387 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_386 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_385 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_128;

architecture SYN_STRUCTURAL of MUX21_128 is

   component ND2_382
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_383
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_384
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_128
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_128 port map( A => S, Y => SB);
   UND1 : ND2_384 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_383 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_382 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_127 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_127;

architecture SYN_STRUCTURAL of MUX21_127 is

   component ND2_379
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_380
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_381
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_127
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_127 port map( A => S, Y => SB);
   UND1 : ND2_381 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_380 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_379 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_126 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_126;

architecture SYN_STRUCTURAL of MUX21_126 is

   component ND2_376
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_377
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_378
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_126
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_126 port map( A => S, Y => SB);
   UND1 : ND2_378 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_377 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_376 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_125 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_125;

architecture SYN_STRUCTURAL of MUX21_125 is

   component ND2_373
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_374
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_375
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_125
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_125 port map( A => S, Y => SB);
   UND1 : ND2_375 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_374 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_373 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_124 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_124;

architecture SYN_STRUCTURAL of MUX21_124 is

   component ND2_370
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_371
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_372
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_124
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_124 port map( A => S, Y => SB);
   UND1 : ND2_372 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_371 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_370 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_123 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_123;

architecture SYN_STRUCTURAL of MUX21_123 is

   component ND2_367
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_368
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_369
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_123
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_123 port map( A => S, Y => SB);
   UND1 : ND2_369 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_368 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_367 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_122 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_122;

architecture SYN_STRUCTURAL of MUX21_122 is

   component ND2_364
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_365
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_366
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_122
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_122 port map( A => S, Y => SB);
   UND1 : ND2_366 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_365 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_364 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_121 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_121;

architecture SYN_STRUCTURAL of MUX21_121 is

   component ND2_361
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_362
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_363
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_121
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_121 port map( A => S, Y => SB);
   UND1 : ND2_363 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_362 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_361 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_120 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_120;

architecture SYN_STRUCTURAL of MUX21_120 is

   component ND2_358
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_359
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_360
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_120
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_120 port map( A => S, Y => SB);
   UND1 : ND2_360 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_359 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_358 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_119 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_119;

architecture SYN_STRUCTURAL of MUX21_119 is

   component ND2_355
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_356
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_357
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_119
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_119 port map( A => S, Y => SB);
   UND1 : ND2_357 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_356 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_355 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_118 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_118;

architecture SYN_STRUCTURAL of MUX21_118 is

   component ND2_352
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_353
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_354
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_118
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_118 port map( A => S, Y => SB);
   UND1 : ND2_354 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_353 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_352 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_117 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_117;

architecture SYN_STRUCTURAL of MUX21_117 is

   component ND2_349
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_350
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_351
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_117
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_117 port map( A => S, Y => SB);
   UND1 : ND2_351 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_350 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_349 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_116 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_116;

architecture SYN_STRUCTURAL of MUX21_116 is

   component ND2_346
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_347
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_348
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_116
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_116 port map( A => S, Y => SB);
   UND1 : ND2_348 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_347 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_346 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_115 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_115;

architecture SYN_STRUCTURAL of MUX21_115 is

   component ND2_343
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_344
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_345
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_115
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_115 port map( A => S, Y => SB);
   UND1 : ND2_345 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_344 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_343 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_114 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_114;

architecture SYN_STRUCTURAL of MUX21_114 is

   component ND2_340
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_341
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_342
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_114
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_114 port map( A => S, Y => SB);
   UND1 : ND2_342 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_341 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_340 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_113 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_113;

architecture SYN_STRUCTURAL of MUX21_113 is

   component ND2_337
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_338
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_339
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_113
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_113 port map( A => S, Y => SB);
   UND1 : ND2_339 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_338 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_337 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_112 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_112;

architecture SYN_STRUCTURAL of MUX21_112 is

   component ND2_334
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_335
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_336
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_112
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_112 port map( A => S, Y => SB);
   UND1 : ND2_336 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_335 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_334 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_111 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_111;

architecture SYN_STRUCTURAL of MUX21_111 is

   component ND2_331
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_332
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_333
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_111
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_111 port map( A => S, Y => SB);
   UND1 : ND2_333 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_332 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_331 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_110 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_110;

architecture SYN_STRUCTURAL of MUX21_110 is

   component ND2_328
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_329
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_330
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_110
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_110 port map( A => S, Y => SB);
   UND1 : ND2_330 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_329 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_328 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_109 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_109;

architecture SYN_STRUCTURAL of MUX21_109 is

   component ND2_325
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_326
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_327
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_109
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_109 port map( A => S, Y => SB);
   UND1 : ND2_327 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_326 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_325 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_108 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_108;

architecture SYN_STRUCTURAL of MUX21_108 is

   component ND2_322
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_323
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_324
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_108
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_108 port map( A => S, Y => SB);
   UND1 : ND2_324 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_323 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_322 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_107 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_107;

architecture SYN_STRUCTURAL of MUX21_107 is

   component ND2_319
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_320
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_321
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_107
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_107 port map( A => S, Y => SB);
   UND1 : ND2_321 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_320 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_319 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_106 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_106;

architecture SYN_STRUCTURAL of MUX21_106 is

   component ND2_316
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_317
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_318
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_106
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_106 port map( A => S, Y => SB);
   UND1 : ND2_318 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_317 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_316 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_105 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_105;

architecture SYN_STRUCTURAL of MUX21_105 is

   component ND2_313
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_314
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_315
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_105
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_105 port map( A => S, Y => SB);
   UND1 : ND2_315 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_314 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_313 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_104 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_104;

architecture SYN_STRUCTURAL of MUX21_104 is

   component ND2_310
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_311
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_312
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_104
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_104 port map( A => S, Y => SB);
   UND1 : ND2_312 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_311 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_310 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_103 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_103;

architecture SYN_STRUCTURAL of MUX21_103 is

   component ND2_307
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_308
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_309
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_103
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_103 port map( A => S, Y => SB);
   UND1 : ND2_309 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_308 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_307 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_102 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_102;

architecture SYN_STRUCTURAL of MUX21_102 is

   component ND2_304
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_305
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_306
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_102
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_102 port map( A => S, Y => SB);
   UND1 : ND2_306 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_305 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_304 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_101 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_101;

architecture SYN_STRUCTURAL of MUX21_101 is

   component ND2_301
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_302
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_303
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_101
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_101 port map( A => S, Y => SB);
   UND1 : ND2_303 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_302 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_301 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_100 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_100;

architecture SYN_STRUCTURAL of MUX21_100 is

   component ND2_298
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_299
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_300
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_100
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_100 port map( A => S, Y => SB);
   UND1 : ND2_300 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_299 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_298 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_99 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_99;

architecture SYN_STRUCTURAL of MUX21_99 is

   component ND2_295
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_296
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_297
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_99
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_99 port map( A => S, Y => SB);
   UND1 : ND2_297 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_296 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_295 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_98 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_98;

architecture SYN_STRUCTURAL of MUX21_98 is

   component ND2_292
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_293
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_294
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_98
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_98 port map( A => S, Y => SB);
   UND1 : ND2_294 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_293 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_292 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_97 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_97;

architecture SYN_STRUCTURAL of MUX21_97 is

   component ND2_289
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_290
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_291
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_97
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_97 port map( A => S, Y => SB);
   UND1 : ND2_291 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_290 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_289 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_96 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_96;

architecture SYN_STRUCTURAL of MUX21_96 is

   component ND2_286
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_287
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_288
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_96
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_96 port map( A => S, Y => SB);
   UND1 : ND2_288 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_287 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_286 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_95 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_95;

architecture SYN_STRUCTURAL of MUX21_95 is

   component ND2_283
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_284
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_285
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_95
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_95 port map( A => S, Y => SB);
   UND1 : ND2_285 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_284 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_283 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_94 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_94;

architecture SYN_STRUCTURAL of MUX21_94 is

   component ND2_280
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_281
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_282
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_94
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_94 port map( A => S, Y => SB);
   UND1 : ND2_282 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_281 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_280 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_93 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_93;

architecture SYN_STRUCTURAL of MUX21_93 is

   component ND2_277
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_278
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_279
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_93
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_93 port map( A => S, Y => SB);
   UND1 : ND2_279 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_278 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_277 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_92 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_92;

architecture SYN_STRUCTURAL of MUX21_92 is

   component ND2_274
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_275
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_276
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_92
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_92 port map( A => S, Y => SB);
   UND1 : ND2_276 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_275 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_274 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_91 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_91;

architecture SYN_STRUCTURAL of MUX21_91 is

   component ND2_271
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_272
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_273
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_91
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_91 port map( A => S, Y => SB);
   UND1 : ND2_273 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_272 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_271 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_90 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_90;

architecture SYN_STRUCTURAL of MUX21_90 is

   component ND2_268
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_269
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_270
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_90
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_90 port map( A => S, Y => SB);
   UND1 : ND2_270 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_269 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_268 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_89 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_89;

architecture SYN_STRUCTURAL of MUX21_89 is

   component ND2_265
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_266
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_267
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_89
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_89 port map( A => S, Y => SB);
   UND1 : ND2_267 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_266 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_265 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_88 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_88;

architecture SYN_STRUCTURAL of MUX21_88 is

   component ND2_262
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_263
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_264
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_88
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_88 port map( A => S, Y => SB);
   UND1 : ND2_264 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_263 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_262 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_87 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_87;

architecture SYN_STRUCTURAL of MUX21_87 is

   component ND2_259
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_260
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_261
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_87
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_87 port map( A => S, Y => SB);
   UND1 : ND2_261 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_260 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_259 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_86 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_86;

architecture SYN_STRUCTURAL of MUX21_86 is

   component ND2_256
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_257
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_258
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_86
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_86 port map( A => S, Y => SB);
   UND1 : ND2_258 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_257 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_256 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_85 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_85;

architecture SYN_STRUCTURAL of MUX21_85 is

   component ND2_253
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_254
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_255
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_85
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_85 port map( A => S, Y => SB);
   UND1 : ND2_255 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_254 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_253 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_84 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_84;

architecture SYN_STRUCTURAL of MUX21_84 is

   component ND2_250
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_251
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_252
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_84
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_84 port map( A => S, Y => SB);
   UND1 : ND2_252 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_251 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_250 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_83 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_83;

architecture SYN_STRUCTURAL of MUX21_83 is

   component ND2_247
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_248
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_249
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_83
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_83 port map( A => S, Y => SB);
   UND1 : ND2_249 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_248 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_247 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_82 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_82;

architecture SYN_STRUCTURAL of MUX21_82 is

   component ND2_244
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_245
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_246
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_82
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_82 port map( A => S, Y => SB);
   UND1 : ND2_246 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_245 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_244 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_81 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_81;

architecture SYN_STRUCTURAL of MUX21_81 is

   component ND2_241
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_242
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_243
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_81
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_81 port map( A => S, Y => SB);
   UND1 : ND2_243 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_242 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_241 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_80 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_80;

architecture SYN_STRUCTURAL of MUX21_80 is

   component ND2_238
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_239
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_240
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_80
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_80 port map( A => S, Y => SB);
   UND1 : ND2_240 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_239 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_238 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_79 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_79;

architecture SYN_STRUCTURAL of MUX21_79 is

   component ND2_235
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_236
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_237
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_79
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_79 port map( A => S, Y => SB);
   UND1 : ND2_237 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_236 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_235 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_78 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_78;

architecture SYN_STRUCTURAL of MUX21_78 is

   component ND2_232
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_233
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_234
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_78
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_78 port map( A => S, Y => SB);
   UND1 : ND2_234 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_233 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_232 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_77 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_77;

architecture SYN_STRUCTURAL of MUX21_77 is

   component ND2_229
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_230
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_231
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_77
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_77 port map( A => S, Y => SB);
   UND1 : ND2_231 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_230 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_229 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_76 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_76;

architecture SYN_STRUCTURAL of MUX21_76 is

   component ND2_226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_76
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_76 port map( A => S, Y => SB);
   UND1 : ND2_228 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_227 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_226 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_75 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_75;

architecture SYN_STRUCTURAL of MUX21_75 is

   component ND2_223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_75
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_75 port map( A => S, Y => SB);
   UND1 : ND2_225 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_224 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_223 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_74 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_74;

architecture SYN_STRUCTURAL of MUX21_74 is

   component ND2_220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_74
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_74 port map( A => S, Y => SB);
   UND1 : ND2_222 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_221 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_220 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_73 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_73;

architecture SYN_STRUCTURAL of MUX21_73 is

   component ND2_217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_73
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_73 port map( A => S, Y => SB);
   UND1 : ND2_219 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_218 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_217 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_72 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_72;

architecture SYN_STRUCTURAL of MUX21_72 is

   component ND2_214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_72
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_72 port map( A => S, Y => SB);
   UND1 : ND2_216 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_215 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_214 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_71 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_71;

architecture SYN_STRUCTURAL of MUX21_71 is

   component ND2_211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_71
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_71 port map( A => S, Y => SB);
   UND1 : ND2_213 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_212 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_211 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_70 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_70;

architecture SYN_STRUCTURAL of MUX21_70 is

   component ND2_208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_70
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_70 port map( A => S, Y => SB);
   UND1 : ND2_210 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_209 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_208 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_69 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_69;

architecture SYN_STRUCTURAL of MUX21_69 is

   component ND2_205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_69
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_69 port map( A => S, Y => SB);
   UND1 : ND2_207 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_206 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_205 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_68 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_68;

architecture SYN_STRUCTURAL of MUX21_68 is

   component ND2_202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_68
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_68 port map( A => S, Y => SB);
   UND1 : ND2_204 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_203 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_202 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_67 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_67;

architecture SYN_STRUCTURAL of MUX21_67 is

   component ND2_199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_67
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_67 port map( A => S, Y => SB);
   UND1 : ND2_201 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_200 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_199 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_66 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_66;

architecture SYN_STRUCTURAL of MUX21_66 is

   component ND2_196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_66
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_66 port map( A => S, Y => SB);
   UND1 : ND2_198 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_197 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_196 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_65 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_65;

architecture SYN_STRUCTURAL of MUX21_65 is

   component ND2_193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_65
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_65 port map( A => S, Y => SB);
   UND1 : ND2_195 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_194 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_193 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_64 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_64;

architecture SYN_STRUCTURAL of MUX21_64 is

   component ND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_64
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_64 port map( A => S, Y => SB);
   UND1 : ND2_192 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_191 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_190 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_63 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_63;

architecture SYN_STRUCTURAL of MUX21_63 is

   component ND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_63 port map( A => S, Y => SB);
   UND1 : ND2_189 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_188 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_187 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_62 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_62;

architecture SYN_STRUCTURAL of MUX21_62 is

   component ND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_62 port map( A => S, Y => SB);
   UND1 : ND2_186 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_185 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_184 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_61 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_61;

architecture SYN_STRUCTURAL of MUX21_61 is

   component ND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_61 port map( A => S, Y => SB);
   UND1 : ND2_183 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_182 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_181 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_60;

architecture SYN_STRUCTURAL of MUX21_60 is

   component ND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_60 port map( A => S, Y => SB);
   UND1 : ND2_180 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_179 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_178 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_59;

architecture SYN_STRUCTURAL of MUX21_59 is

   component ND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_59 port map( A => S, Y => SB);
   UND1 : ND2_177 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_176 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_175 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_58;

architecture SYN_STRUCTURAL of MUX21_58 is

   component ND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_58 port map( A => S, Y => SB);
   UND1 : ND2_174 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_173 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_172 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_57;

architecture SYN_STRUCTURAL of MUX21_57 is

   component ND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_57 port map( A => S, Y => SB);
   UND1 : ND2_171 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_170 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_169 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_56;

architecture SYN_STRUCTURAL of MUX21_56 is

   component ND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_56 port map( A => S, Y => SB);
   UND1 : ND2_168 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_167 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_166 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_55;

architecture SYN_STRUCTURAL of MUX21_55 is

   component ND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_55 port map( A => S, Y => SB);
   UND1 : ND2_165 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_164 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_163 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_54;

architecture SYN_STRUCTURAL of MUX21_54 is

   component ND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_54 port map( A => S, Y => SB);
   UND1 : ND2_162 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_161 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_160 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_53;

architecture SYN_STRUCTURAL of MUX21_53 is

   component ND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_53 port map( A => S, Y => SB);
   UND1 : ND2_159 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_158 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_157 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_52;

architecture SYN_STRUCTURAL of MUX21_52 is

   component ND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_52 port map( A => S, Y => SB);
   UND1 : ND2_156 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_155 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_154 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_51;

architecture SYN_STRUCTURAL of MUX21_51 is

   component ND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_51 port map( A => S, Y => SB);
   UND1 : ND2_153 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_152 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_151 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_50;

architecture SYN_STRUCTURAL of MUX21_50 is

   component ND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_50 port map( A => S, Y => SB);
   UND1 : ND2_150 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_149 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_148 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_49;

architecture SYN_STRUCTURAL of MUX21_49 is

   component ND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_49 port map( A => S, Y => SB);
   UND1 : ND2_147 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_146 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_145 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_48;

architecture SYN_STRUCTURAL of MUX21_48 is

   component ND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_48 port map( A => S, Y => SB);
   UND1 : ND2_144 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_143 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_142 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_47;

architecture SYN_STRUCTURAL of MUX21_47 is

   component ND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_47 port map( A => S, Y => SB);
   UND1 : ND2_141 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_140 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_139 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_46;

architecture SYN_STRUCTURAL of MUX21_46 is

   component ND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_46 port map( A => S, Y => SB);
   UND1 : ND2_138 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_137 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_136 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_45;

architecture SYN_STRUCTURAL of MUX21_45 is

   component ND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_45 port map( A => S, Y => SB);
   UND1 : ND2_135 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_134 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_133 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_44;

architecture SYN_STRUCTURAL of MUX21_44 is

   component ND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_44 port map( A => S, Y => SB);
   UND1 : ND2_132 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_131 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_130 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_43;

architecture SYN_STRUCTURAL of MUX21_43 is

   component ND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_43 port map( A => S, Y => SB);
   UND1 : ND2_129 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_128 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_127 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_42;

architecture SYN_STRUCTURAL of MUX21_42 is

   component ND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_42 port map( A => S, Y => SB);
   UND1 : ND2_126 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_125 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_124 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_41;

architecture SYN_STRUCTURAL of MUX21_41 is

   component ND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_41 port map( A => S, Y => SB);
   UND1 : ND2_123 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_122 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_121 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_40;

architecture SYN_STRUCTURAL of MUX21_40 is

   component ND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_40 port map( A => S, Y => SB);
   UND1 : ND2_120 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_119 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_118 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_39;

architecture SYN_STRUCTURAL of MUX21_39 is

   component ND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_39 port map( A => S, Y => SB);
   UND1 : ND2_117 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_116 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_115 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_38;

architecture SYN_STRUCTURAL of MUX21_38 is

   component ND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_38 port map( A => S, Y => SB);
   UND1 : ND2_114 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_113 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_112 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_37;

architecture SYN_STRUCTURAL of MUX21_37 is

   component ND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_37 port map( A => S, Y => SB);
   UND1 : ND2_111 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_110 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_109 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_36;

architecture SYN_STRUCTURAL of MUX21_36 is

   component ND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_36 port map( A => S, Y => SB);
   UND1 : ND2_108 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_107 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_106 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_35;

architecture SYN_STRUCTURAL of MUX21_35 is

   component ND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_35 port map( A => S, Y => SB);
   UND1 : ND2_105 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_104 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_103 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_34;

architecture SYN_STRUCTURAL of MUX21_34 is

   component ND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_34 port map( A => S, Y => SB);
   UND1 : ND2_102 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_101 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_100 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_33;

architecture SYN_STRUCTURAL of MUX21_33 is

   component ND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_33 port map( A => S, Y => SB);
   UND1 : ND2_99 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_98 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_97 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_32;

architecture SYN_STRUCTURAL of MUX21_32 is

   component ND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_32 port map( A => S, Y => SB);
   UND1 : ND2_96 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31;

architecture SYN_STRUCTURAL of MUX21_31 is

   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31 port map( A => S, Y => SB);
   UND1 : ND2_93 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_92 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_91 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30;

architecture SYN_STRUCTURAL of MUX21_30 is

   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30 port map( A => S, Y => SB);
   UND1 : ND2_90 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_89 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_88 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_29;

architecture SYN_STRUCTURAL of MUX21_29 is

   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_29 port map( A => S, Y => SB);
   UND1 : ND2_87 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_86 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_85 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_28;

architecture SYN_STRUCTURAL of MUX21_28 is

   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_28 port map( A => S, Y => SB);
   UND1 : ND2_84 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_83 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_82 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_27;

architecture SYN_STRUCTURAL_architecture of MUX21_27 is

   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_27 port map( A => S, Y => SB);
   UND1 : ND2_81 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_80 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_79 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_26;

architecture SYN_STRUCTURAL_architecture2 of MUX21_26 is

   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_26 port map( A => S, Y => SB);
   UND1 : ND2_78 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_77 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_76 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_25;

architecture SYN_STRUCTURAL_architecture3 of MUX21_25 is

   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_25 port map( A => S, Y => SB);
   UND1 : ND2_75 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_74 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_73 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_24;

architecture SYN_STRUCTURAL of MUX21_24 is

   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_24 port map( A => S, Y => SB);
   UND1 : ND2_72 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_71 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_70 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_23;

architecture SYN_STRUCTURAL_architecture of MUX21_23 is

   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_23 port map( A => S, Y => SB);
   UND1 : ND2_69 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_68 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_67 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_22;

architecture SYN_STRUCTURAL_architecture2 of MUX21_22 is

   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_22 port map( A => S, Y => SB);
   UND1 : ND2_66 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_65 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_64 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_21;

architecture SYN_STRUCTURAL_architecture3 of MUX21_21 is

   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_21 port map( A => S, Y => SB);
   UND1 : ND2_63 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_62 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_61 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_20;

architecture SYN_STRUCTURAL of MUX21_20 is

   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_20 port map( A => S, Y => SB);
   UND1 : ND2_60 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_59 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_58 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_19;

architecture SYN_STRUCTURAL_architecture of MUX21_19 is

   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_19 port map( A => S, Y => SB);
   UND1 : ND2_57 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_56 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_55 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_18;

architecture SYN_STRUCTURAL_architecture2 of MUX21_18 is

   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_18 port map( A => S, Y => SB);
   UND1 : ND2_54 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_53 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_52 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_17;

architecture SYN_STRUCTURAL_architecture3 of MUX21_17 is

   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_17 port map( A => S, Y => SB);
   UND1 : ND2_51 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_50 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_49 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_16;

architecture SYN_STRUCTURAL of MUX21_16 is

   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_16 port map( A => S, Y => SB);
   UND1 : ND2_48 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_47 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_46 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_15;

architecture SYN_STRUCTURAL_architecture of MUX21_15 is

   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_15 port map( A => S, Y => SB);
   UND1 : ND2_45 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_44 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_43 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_14;

architecture SYN_STRUCTURAL_architecture2 of MUX21_14 is

   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_14 port map( A => S, Y => SB);
   UND1 : ND2_42 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_41 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_40 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_13;

architecture SYN_STRUCTURAL_architecture3 of MUX21_13 is

   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_13 port map( A => S, Y => SB);
   UND1 : ND2_39 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_38 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_37 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_12;

architecture SYN_STRUCTURAL of MUX21_12 is

   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_12 port map( A => S, Y => SB);
   UND1 : ND2_36 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_35 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_34 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_11;

architecture SYN_STRUCTURAL_architecture of MUX21_11 is

   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_11 port map( A => S, Y => SB);
   UND1 : ND2_33 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_32 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_31 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_10;

architecture SYN_STRUCTURAL_architecture2 of MUX21_10 is

   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_10 port map( A => S, Y => SB);
   UND1 : ND2_30 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_29 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_28 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_9;

architecture SYN_STRUCTURAL_architecture3 of MUX21_9 is

   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_9 port map( A => S, Y => SB);
   UND1 : ND2_27 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_26 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_25 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_8;

architecture SYN_STRUCTURAL of MUX21_8 is

   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_8 port map( A => S, Y => SB);
   UND1 : ND2_24 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_23 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_22 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_7;

architecture SYN_STRUCTURAL_architecture of MUX21_7 is

   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_7 port map( A => S, Y => SB);
   UND1 : ND2_21 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_20 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_19 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_6;

architecture SYN_STRUCTURAL_architecture2 of MUX21_6 is

   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_6 port map( A => S, Y => SB);
   UND1 : ND2_18 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_17 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_16 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_5;

architecture SYN_STRUCTURAL_architecture3 of MUX21_5 is

   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_5 port map( A => S, Y => SB);
   UND1 : ND2_15 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_14 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_13 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_4;

architecture SYN_STRUCTURAL of MUX21_4 is

   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_4 port map( A => S, Y => SB);
   UND1 : ND2_12 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_11 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_10 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_3;

architecture SYN_STRUCTURAL_architecture of MUX21_3 is

   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_3 port map( A => S, Y => SB);
   UND1 : ND2_9 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_8 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_7 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_2;

architecture SYN_STRUCTURAL_architecture2 of MUX21_2 is

   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_2 port map( A => S, Y => SB);
   UND1 : ND2_6 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_5 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_4 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_1;

architecture SYN_STRUCTURAL_architecture3 of MUX21_1 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_1 port map( A => S, Y => SB);
   UND1 : ND2_3 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_2 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT6_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 downto 
         0);  Q : out std_logic_vector (5 downto 0));

end regFFD_NBIT6_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT6_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
      n33, n34, n35, n36 : std_logic;

begin
   
   Q_reg_5_inst : DFFR_X1 port map( D => n19, CK => CK, RN => RESET, Q => Q(5),
                           QN => n25);
   Q_reg_4_inst : DFFR_X1 port map( D => n20, CK => CK, RN => RESET, Q => Q(4),
                           QN => n26);
   Q_reg_3_inst : DFFR_X1 port map( D => n21, CK => CK, RN => RESET, Q => Q(3),
                           QN => n27);
   Q_reg_2_inst : DFFR_X1 port map( D => n22, CK => CK, RN => RESET, Q => Q(2),
                           QN => n28);
   Q_reg_1_inst : DFFR_X1 port map( D => n23, CK => CK, RN => RESET, Q => Q(1),
                           QN => n29);
   Q_reg_0_inst : DFFR_X1 port map( D => n24, CK => CK, RN => RESET, Q => Q(0),
                           QN => n30);
   U2 : OAI21_X1 port map( B1 => n30, B2 => ENABLE, A => n36, ZN => n24);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n36);
   U4 : OAI21_X1 port map( B1 => n29, B2 => ENABLE, A => n35, ZN => n23);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n35);
   U6 : OAI21_X1 port map( B1 => n28, B2 => ENABLE, A => n34, ZN => n22);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n34);
   U8 : OAI21_X1 port map( B1 => n27, B2 => ENABLE, A => n33, ZN => n21);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n33);
   U10 : OAI21_X1 port map( B1 => n26, B2 => ENABLE, A => n32, ZN => n20);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n32);
   U12 : OAI21_X1 port map( B1 => n25, B2 => ENABLE, A => n31, ZN => n19);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n31);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_2 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_2;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n16, CK => CK, RN => RESET, Q => Q(4),
                           QN => n21);
   Q_reg_3_inst : DFFR_X1 port map( D => n17, CK => CK, RN => RESET, Q => Q(3),
                           QN => n22);
   Q_reg_2_inst : DFFR_X1 port map( D => n18, CK => CK, RN => RESET, Q => Q(2),
                           QN => n23);
   Q_reg_1_inst : DFFR_X1 port map( D => n19, CK => CK, RN => RESET, Q => Q(1),
                           QN => n24);
   Q_reg_0_inst : DFFR_X1 port map( D => n20, CK => CK, RN => RESET, Q => Q(0),
                           QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => ENABLE, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => ENABLE, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => ENABLE, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => ENABLE, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => ENABLE, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n26);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n16, CK => CK, RN => RESET, Q => Q(4),
                           QN => n21);
   Q_reg_3_inst : DFFR_X1 port map( D => n17, CK => CK, RN => RESET, Q => Q(3),
                           QN => n22);
   Q_reg_2_inst : DFFR_X1 port map( D => n18, CK => CK, RN => RESET, Q => Q(2),
                           QN => n23);
   Q_reg_1_inst : DFFR_X1 port map( D => n19, CK => CK, RN => RESET, Q => Q(1),
                           QN => n24);
   Q_reg_0_inst : DFFR_X1 port map( D => n20, CK => CK, RN => RESET, Q => Q(0),
                           QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => ENABLE, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => ENABLE, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => ENABLE, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => ENABLE, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => ENABLE, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n26);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_7 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_7;

architecture SYN_SYNC_BHV of FF_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n5, n6, n7, n8, n_1022 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1022);
   U3 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => n5);
   U4 : INV_X1 port map( A => RESET, ZN => n7);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n6, ZN => n8)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n6);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_6 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_6;

architecture SYN_SYNC_BHV of FF_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n5, n6, n7, n8, n_1023 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1023);
   U3 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => n5);
   U4 : INV_X1 port map( A => RESET, ZN => n7);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n6, ZN => n8)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n6);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_5 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_5;

architecture SYN_SYNC_BHV of FF_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n5, n6, n7, n8, n_1024 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1024);
   U3 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => n5);
   U4 : INV_X1 port map( A => RESET, ZN => n7);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n6, ZN => n8)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n6);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_4 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_4;

architecture SYN_SYNC_BHV of FF_4 is

   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal Q_port, n2, n4, n5, n_1025 : std_logic;

begin
   Q <= Q_port;
   
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n4, ZN => n5)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n4);
   Q_reg : SDFF_X1 port map( D => RESET, SI => n2, SE => n5, CK => CLK, Q => 
                           Q_port, QN => n_1025);
   n2 <= '0';

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_3 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_3;

architecture SYN_SYNC_BHV of FF_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n5, n6, n7, n8, n_1026 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1026);
   U3 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => n5);
   U4 : INV_X1 port map( A => RESET, ZN => n7);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n6, ZN => n8)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n6);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_2 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_2;

architecture SYN_SYNC_BHV of FF_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n5, n6, n7, n8, n_1027 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1027);
   U3 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => n5);
   U4 : INV_X1 port map( A => RESET, ZN => n7);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n6, ZN => n8)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n6);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_1 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_1;

architecture SYN_SYNC_BHV of FF_1 is

   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n11, n5, Q_port, n7, n8, n9, n10, n_1028 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n7, CK => CLK, Q => n11, QN => n_1028);
   U3 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n7);
   U4 : INV_X1 port map( A => RESET, ZN => n9);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n8, ZN => n10
                           );
   U6 : INV_X1 port map( A => EN, ZN => n8);
   U7 : INV_X1 port map( A => n11, ZN => n5);
   U8 : INV_X4 port map( A => n5, ZN => Q_port);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_6;

architecture SYN_struct of MUX21_GENERIC_NBIT32_6 is

   component MUX21_193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_218
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_219
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_220
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_221
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_222
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_223
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_224
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_224 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_223 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_222 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_221 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_220 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_219 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_218 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_217 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_216 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_215 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_214 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_213 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_212 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_211 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_210 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_209 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_208 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_207 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_206 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_205 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_204 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_203 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_202 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_201 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_200 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_199 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_198 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_197 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_196 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_195 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_194 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_193 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_5;

architecture SYN_struct of MUX21_GENERIC_NBIT32_5 is

   component MUX21_161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_192 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_191 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_190 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_189 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_188 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_187 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_186 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_185 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_184 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_183 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_182 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_181 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_180 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_179 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_178 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_177 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_176 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_175 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_174 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_173 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_172 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_171 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_170 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_169 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_168 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_167 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_166 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_165 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_164 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_163 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_162 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_161 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_4;

architecture SYN_struct of MUX21_GENERIC_NBIT32_4 is

   component MUX21_129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_160 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_159 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_158 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_157 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_156 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_155 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_154 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_153 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_152 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_151 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_150 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_149 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_148 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_147 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_146 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_145 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_144 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_143 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_142 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_141 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_140 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_139 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_138 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_137 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_136 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_135 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_134 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_133 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_132 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_131 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_130 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_129 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_3;

architecture SYN_struct of MUX21_GENERIC_NBIT32_3 is

   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_97
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_98
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_99
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_100
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_101
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_102
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_103
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_104
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_105
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_106
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_107
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_108
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_109
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_110
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_111
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_112
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_113
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_114
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_115
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_116
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_117
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_118
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_119
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_120
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_121
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_122
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_123
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_124
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_125
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_126
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_127
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   gen1_0 : MUX21_128 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   gen1_1 : MUX21_127 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   gen1_2 : MUX21_126 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   gen1_3 : MUX21_125 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   gen1_4 : MUX21_124 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   gen1_5 : MUX21_123 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   gen1_6 : MUX21_122 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   gen1_7 : MUX21_121 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   gen1_8 : MUX21_120 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   gen1_9 : MUX21_119 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   gen1_10 : MUX21_118 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   gen1_11 : MUX21_117 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   gen1_12 : MUX21_116 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   gen1_13 : MUX21_115 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   gen1_14 : MUX21_114 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   gen1_15 : MUX21_113 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   gen1_16 : MUX21_112 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   gen1_17 : MUX21_111 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   gen1_18 : MUX21_110 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   gen1_19 : MUX21_109 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   gen1_20 : MUX21_108 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   gen1_21 : MUX21_107 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   gen1_22 : MUX21_106 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   gen1_23 : MUX21_105 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   gen1_24 : MUX21_104 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   gen1_25 : MUX21_103 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   gen1_26 : MUX21_102 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   gen1_27 : MUX21_101 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   gen1_28 : MUX21_100 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   gen1_29 : MUX21_99 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   gen1_30 : MUX21_98 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   gen1_31 : MUX21_97 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : CLKBUF_X3 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X3 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X3 port map( A => SEL, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_2;

architecture SYN_struct of MUX21_GENERIC_NBIT32_2 is

   component MUX21_65
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_66
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_67
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_68
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_69
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_70
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_71
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_72
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_73
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_74
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_75
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_76
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_77
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_78
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_79
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_80
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_81
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_82
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_83
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_84
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_85
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_86
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_87
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_88
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_89
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_90
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_91
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_92
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_93
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_94
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_95
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_96
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_96 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_95 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_94 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_93 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_92 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_91 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_90 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_89 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_88 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_87 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_86 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_85 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_84 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_83 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_82 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_81 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_80 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_79 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_78 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_77 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_76 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_75 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_74 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_73 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_72 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_71 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_70 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_69 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_68 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_67 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_66 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_65 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_1;

architecture SYN_struct of MUX21_GENERIC_NBIT32_1 is

   component MUX21_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_61
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_62
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_63
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_64
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_64 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_63 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_62 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_61 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_60 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_59 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_58 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_57 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_56 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_55 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_54 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_53 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_52 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_51 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_50 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_49 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_48 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_47 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_46 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_45 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_44 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_43 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_42 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_41 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_40 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_39 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_38 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_37 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_36 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_35 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_34 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_33 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_18 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_18;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_17 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_17;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_16 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_16;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_15 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_15;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_14 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_14;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_13 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_13;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_12 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_12;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_11 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_11;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n163);
   U2 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U4 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U6 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U8 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U10 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U12 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U14 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U16 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U18 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U20 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U22 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U24 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U26 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U28 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U30 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U32 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U34 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U36 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U38 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U40 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U42 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U44 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U46 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U48 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U50 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U52 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U54 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U56 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U58 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U60 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U62 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U64 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);
   Q_reg_31_inst : SDFFR_X1 port map( D => n98, SI => n99, SE => n97, CK => CK,
                           RN => RESET, Q => Q(31), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n137);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n135);
   U66 : INV_X1 port map( A => n100, ZN => n97);
   n98 <= '1';
   n99 <= '0';

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_10 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_10;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_9 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_9;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_8 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_8;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_7 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_7;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_6 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_6;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_5 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_5;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_4 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_4;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_3 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_3;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_2 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_2;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192 : 
      std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n97, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n129);
   Q_reg_30_inst : DFFR_X1 port map( D => n98, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n99, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n131);
   Q_reg_28_inst : DFFR_X1 port map( D => n100, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n132);
   Q_reg_27_inst : DFFR_X1 port map( D => n101, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n133);
   Q_reg_26_inst : DFFR_X1 port map( D => n102, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n134);
   Q_reg_25_inst : DFFR_X1 port map( D => n103, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n135);
   Q_reg_24_inst : DFFR_X1 port map( D => n104, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n136);
   Q_reg_23_inst : DFFR_X1 port map( D => n105, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n137);
   Q_reg_22_inst : DFFR_X1 port map( D => n106, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n138);
   Q_reg_21_inst : DFFR_X1 port map( D => n107, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n139);
   Q_reg_20_inst : DFFR_X1 port map( D => n108, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n140);
   Q_reg_19_inst : DFFR_X1 port map( D => n109, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n141);
   Q_reg_18_inst : DFFR_X1 port map( D => n110, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n142);
   Q_reg_17_inst : DFFR_X1 port map( D => n111, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n143);
   Q_reg_16_inst : DFFR_X1 port map( D => n112, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n144);
   Q_reg_15_inst : DFFR_X1 port map( D => n113, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n145);
   Q_reg_14_inst : DFFR_X1 port map( D => n114, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n146);
   Q_reg_13_inst : DFFR_X1 port map( D => n115, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n147);
   Q_reg_12_inst : DFFR_X1 port map( D => n116, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n148);
   Q_reg_11_inst : DFFR_X1 port map( D => n117, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n149);
   Q_reg_10_inst : DFFR_X1 port map( D => n118, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n150);
   Q_reg_9_inst : DFFR_X1 port map( D => n119, CK => CK, RN => RESET, Q => Q(9)
                           , QN => n151);
   Q_reg_8_inst : DFFR_X1 port map( D => n120, CK => CK, RN => RESET, Q => Q(8)
                           , QN => n152);
   Q_reg_7_inst : DFFR_X1 port map( D => n121, CK => CK, RN => RESET, Q => Q(7)
                           , QN => n153);
   Q_reg_6_inst : DFFR_X1 port map( D => n122, CK => CK, RN => RESET, Q => Q(6)
                           , QN => n154);
   Q_reg_5_inst : DFFR_X1 port map( D => n123, CK => CK, RN => RESET, Q => Q(5)
                           , QN => n155);
   Q_reg_4_inst : DFFR_X1 port map( D => n124, CK => CK, RN => RESET, Q => Q(4)
                           , QN => n156);
   Q_reg_3_inst : DFFR_X1 port map( D => n125, CK => CK, RN => RESET, Q => Q(3)
                           , QN => n157);
   Q_reg_2_inst : DFFR_X1 port map( D => n126, CK => CK, RN => RESET, Q => Q(2)
                           , QN => n158);
   Q_reg_1_inst : DFFR_X1 port map( D => n127, CK => CK, RN => RESET, Q => Q(1)
                           , QN => n159);
   Q_reg_0_inst : DFFR_X1 port map( D => n128, CK => CK, RN => RESET, Q => Q(0)
                           , QN => n160);
   U2 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n192);
   U4 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n191);
   U6 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n190);
   U8 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n189);
   U10 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n188);
   U12 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n187);
   U14 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n186);
   U16 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n185);
   U18 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n184);
   U20 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n183);
   U22 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n182);
   U24 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n181);
   U26 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n180);
   U28 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n179);
   U30 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n178);
   U32 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n177);
   U34 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n176);
   U36 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n175);
   U38 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n174);
   U40 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n173);
   U42 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n172);
   U44 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n171);
   U46 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n170);
   U48 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n169);
   U50 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n168);
   U52 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n167);
   U54 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n166);
   U56 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n165);
   U58 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n164);
   U60 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n163, ZN => n99);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n163);
   U62 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n162, ZN => n98);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n162);
   U64 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n161, ZN => n97);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n161);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_0;

architecture SYN_struct of MUX21_GENERIC_NBIT4_0 is

   component MUX21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_32 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_31 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_30 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_29 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_0;

architecture SYN_BEHAVIORAL of RCA_NBIT4_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_0 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_0;

architecture SYN_behave of P_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_0;

architecture SYN_STRUCTURAL of CSB_NBIT4_0 is

   component MUX21_GENERIC_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1029, n_1030 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1029);
   RCA1 : RCA_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1030);
   MUXCin : MUX21_GENERIC_NBIT4_0 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_0 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_0;

architecture SYN_arch of PG_0 is

   component P_0
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_43
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_43 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_0 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_0 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_0;

architecture SYN_behave of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n1);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_STRUCTURAL of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component CSB_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_0 : CSB_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), S(2) 
                           => S(2), S(1) => S(1), S(0) => S(0));
   CSBI_1 : CSB_NBIT4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5), 
                           A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1) => 
                           B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), S(2) 
                           => S(6), S(1) => S(5), S(0) => S(4));
   CSBI_2 : CSB_NBIT4_6 port map( A(3) => A(11), A(2) => A(10), A(1) => A(9), 
                           A(0) => A(8), B(3) => B(11), B(2) => B(10), B(1) => 
                           B(9), B(0) => B(8), Ci => Ci(2), S(3) => S(11), S(2)
                           => S(10), S(1) => S(9), S(0) => S(8));
   CSBI_3 : CSB_NBIT4_5 port map( A(3) => A(15), A(2) => A(14), A(1) => A(13), 
                           A(0) => A(12), B(3) => B(15), B(2) => B(14), B(1) =>
                           B(13), B(0) => B(12), Ci => Ci(3), S(3) => S(15), 
                           S(2) => S(14), S(1) => S(13), S(0) => S(12));
   CSBI_4 : CSB_NBIT4_4 port map( A(3) => A(19), A(2) => A(18), A(1) => A(17), 
                           A(0) => A(16), B(3) => B(19), B(2) => B(18), B(1) =>
                           B(17), B(0) => B(16), Ci => Ci(4), S(3) => S(19), 
                           S(2) => S(18), S(1) => S(17), S(0) => S(16));
   CSBI_5 : CSB_NBIT4_3 port map( A(3) => A(23), A(2) => A(22), A(1) => A(21), 
                           A(0) => A(20), B(3) => B(23), B(2) => B(22), B(1) =>
                           B(21), B(0) => B(20), Ci => Ci(5), S(3) => S(23), 
                           S(2) => S(22), S(1) => S(21), S(0) => S(20));
   CSBI_6 : CSB_NBIT4_2 port map( A(3) => A(27), A(2) => A(26), A(1) => A(25), 
                           A(0) => A(24), B(3) => B(27), B(2) => B(26), B(1) =>
                           B(25), B(0) => B(24), Ci => Ci(6), S(3) => S(27), 
                           S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CSBI_7 : CSB_NBIT4_1 port map( A(3) => A(31), A(2) => A(30), A(1) => A(29), 
                           A(0) => A(28), B(3) => B(31), B(2) => B(30), B(1) =>
                           B(29), B(0) => B(28), Ci => Ci(7), S(3) => S(31), 
                           S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_arch of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 is

   component G_44
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_45
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_46
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_47
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_1
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_2
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_48
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_49
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_3
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_4
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_5
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_50
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_6
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_7
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_8
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_9
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_10
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_11
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_12
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_51
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_13
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_14
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_15
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_16
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_17
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_18
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_19
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_20
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_21
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_22
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_23
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_24
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_25
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_26
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_27
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_28
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_29
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_30
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_31
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_32
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_33
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_34
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_35
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_36
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_37
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_38
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_39
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_40
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_41
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_42
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_52
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_0
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_0
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port,
      Co_2_port, Co_1_port, Co_0_port, gi_32_4_port, gi_32_3_port, gi_32_2_port
      , gi_32_1_port, gi_32_0_port, gi_31_0_port, gi_30_0_port, gi_29_0_port, 
      gi_28_4_port, gi_28_2_port, gi_28_1_port, gi_28_0_port, gi_27_0_port, 
      gi_26_0_port, gi_25_0_port, gi_24_3_port, gi_24_2_port, gi_24_1_port, 
      gi_24_0_port, gi_23_0_port, gi_22_0_port, gi_21_0_port, gi_20_2_port, 
      gi_20_1_port, gi_20_0_port, gi_19_0_port, gi_18_0_port, gi_17_0_port, 
      gi_16_3_port, gi_16_2_port, gi_16_1_port, gi_16_0_port, gi_15_0_port, 
      gi_14_0_port, gi_13_0_port, gi_12_2_port, gi_12_1_port, gi_12_0_port, 
      gi_11_0_port, gi_10_0_port, gi_9_0_port, gi_8_2_port, gi_8_1_port, 
      gi_8_0_port, gi_7_0_port, gi_6_0_port, gi_5_0_port, gi_4_1_port, 
      gi_4_0_port, gi_3_0_port, gi_2_1_port, gi_2_0_port, gi_1_0_port, 
      gi_0_0_port, pi_32_4_port, pi_32_3_port, pi_32_2_port, pi_32_1_port, 
      pi_32_0_port, pi_31_0_port, pi_30_0_port, pi_29_0_port, pi_28_4_port, 
      pi_28_2_port, pi_28_1_port, pi_28_0_port, pi_27_0_port, pi_26_0_port, 
      pi_25_0_port, pi_24_3_port, pi_24_2_port, pi_24_1_port, pi_24_0_port, 
      pi_23_0_port, pi_22_0_port, pi_21_0_port, pi_20_2_port, pi_20_1_port, 
      pi_20_0_port, pi_19_0_port, pi_18_0_port, pi_17_0_port, pi_16_3_port, 
      pi_16_2_port, pi_16_1_port, pi_16_0_port, pi_15_0_port, pi_14_0_port, 
      pi_13_0_port, pi_12_2_port, pi_12_1_port, pi_12_0_port, pi_11_0_port, 
      pi_10_0_port, pi_9_0_port, pi_8_2_port, pi_8_1_port, pi_8_0_port, 
      pi_7_0_port, pi_6_0_port, pi_5_0_port, pi_4_1_port, pi_4_0_port, 
      pi_3_0_port, pi_2_0_port, pi_0_0_port, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   X_Logic0_port <= '0';
   U2 : XOR2_X1 port map( A => B(8), B => A(8), Z => pi_9_0_port);
   U3 : XOR2_X1 port map( A => B(7), B => A(7), Z => pi_8_0_port);
   U4 : XOR2_X1 port map( A => B(6), B => A(6), Z => pi_7_0_port);
   U5 : XOR2_X1 port map( A => B(5), B => A(5), Z => pi_6_0_port);
   U6 : XOR2_X1 port map( A => B(4), B => A(4), Z => pi_5_0_port);
   U7 : XOR2_X1 port map( A => B(3), B => A(3), Z => pi_4_0_port);
   U8 : XOR2_X1 port map( A => B(2), B => A(2), Z => pi_3_0_port);
   U9 : XOR2_X1 port map( A => B(31), B => A(31), Z => pi_32_0_port);
   U10 : XOR2_X1 port map( A => B(30), B => A(30), Z => pi_31_0_port);
   U11 : XOR2_X1 port map( A => B(29), B => A(29), Z => pi_30_0_port);
   U12 : XOR2_X1 port map( A => B(1), B => A(1), Z => pi_2_0_port);
   U13 : XOR2_X1 port map( A => B(28), B => A(28), Z => pi_29_0_port);
   U14 : XOR2_X1 port map( A => B(27), B => A(27), Z => pi_28_0_port);
   U15 : XOR2_X1 port map( A => B(26), B => A(26), Z => pi_27_0_port);
   U16 : XOR2_X1 port map( A => B(25), B => A(25), Z => pi_26_0_port);
   U17 : XOR2_X1 port map( A => B(24), B => A(24), Z => pi_25_0_port);
   U18 : XOR2_X1 port map( A => B(23), B => A(23), Z => pi_24_0_port);
   U19 : XOR2_X1 port map( A => B(22), B => A(22), Z => pi_23_0_port);
   U20 : XOR2_X1 port map( A => B(21), B => A(21), Z => pi_22_0_port);
   U21 : XOR2_X1 port map( A => B(20), B => A(20), Z => pi_21_0_port);
   U22 : XOR2_X1 port map( A => B(19), B => A(19), Z => pi_20_0_port);
   U23 : XOR2_X1 port map( A => B(18), B => A(18), Z => pi_19_0_port);
   U24 : XOR2_X1 port map( A => B(17), B => A(17), Z => pi_18_0_port);
   U25 : XOR2_X1 port map( A => B(16), B => A(16), Z => pi_17_0_port);
   U26 : XOR2_X1 port map( A => B(15), B => A(15), Z => pi_16_0_port);
   U27 : XOR2_X1 port map( A => B(14), B => A(14), Z => pi_15_0_port);
   U28 : XOR2_X1 port map( A => B(13), B => A(13), Z => pi_14_0_port);
   U29 : XOR2_X1 port map( A => B(12), B => A(12), Z => pi_13_0_port);
   U30 : XOR2_X1 port map( A => B(11), B => A(11), Z => pi_12_0_port);
   U31 : XOR2_X1 port map( A => B(10), B => A(10), Z => pi_11_0_port);
   U32 : XOR2_X1 port map( A => B(9), B => A(9), Z => pi_10_0_port);
   U33 : XOR2_X1 port map( A => B(0), B => A(0), Z => pi_0_0_port);
   U34 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => gi_9_0_port);
   U35 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => gi_8_0_port);
   U36 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => gi_7_0_port);
   U37 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => gi_6_0_port);
   U38 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => gi_5_0_port);
   U39 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => gi_4_0_port);
   U40 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => gi_3_0_port);
   U41 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => gi_32_0_port);
   U42 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => gi_31_0_port);
   U43 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => gi_30_0_port);
   U44 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => gi_2_0_port);
   U45 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => gi_29_0_port);
   U46 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => gi_28_0_port);
   U47 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => gi_27_0_port);
   U48 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => gi_26_0_port);
   U49 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => gi_25_0_port);
   U50 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => gi_24_0_port);
   U51 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => gi_23_0_port);
   U52 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => gi_22_0_port);
   U53 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => gi_21_0_port);
   U54 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => gi_20_0_port);
   U55 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => gi_19_0_port);
   U56 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => gi_18_0_port);
   U57 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => gi_17_0_port);
   U58 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => gi_16_0_port);
   U59 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => gi_15_0_port);
   U60 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => gi_14_0_port);
   U61 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => gi_13_0_port);
   U62 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => gi_12_0_port);
   U63 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => gi_11_0_port);
   U64 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => gi_10_0_port);
   U65 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => gi_0_0_port);
   g_port0_0_1 : G_0 port map( G1 => gi_0_0_port, P => pi_0_0_port, G2 => Cin, 
                           Co => gi_1_0_port);
   pg_port2_1_1 : PG_0 port map( G1 => gi_1_0_port, P1 => X_Logic0_port, G2 => 
                           gi_0_0_port, P2 => pi_0_0_port, gout => n_1031, pout
                           => n_1032);
   g_port1_1_2 : G_52 port map( G1 => gi_2_0_port, P => pi_2_0_port, G2 => 
                           gi_1_0_port, Co => gi_2_1_port);
   pg_port2_1_3 : PG_42 port map( G1 => gi_3_0_port, P1 => pi_3_0_port, G2 => 
                           gi_2_0_port, P2 => pi_2_0_port, gout => n_1033, pout
                           => n_1034);
   pg_port2_1_4 : PG_41 port map( G1 => gi_4_0_port, P1 => pi_4_0_port, G2 => 
                           gi_3_0_port, P2 => pi_3_0_port, gout => gi_4_1_port,
                           pout => pi_4_1_port);
   pg_port2_1_5 : PG_40 port map( G1 => gi_5_0_port, P1 => pi_5_0_port, G2 => 
                           gi_4_0_port, P2 => pi_4_0_port, gout => n_1035, pout
                           => n_1036);
   pg_port2_1_6 : PG_39 port map( G1 => gi_6_0_port, P1 => pi_6_0_port, G2 => 
                           gi_5_0_port, P2 => pi_5_0_port, gout => n_1037, pout
                           => n_1038);
   pg_port2_1_7 : PG_38 port map( G1 => gi_7_0_port, P1 => pi_7_0_port, G2 => 
                           gi_6_0_port, P2 => pi_6_0_port, gout => n_1039, pout
                           => n_1040);
   pg_port2_1_8 : PG_37 port map( G1 => gi_8_0_port, P1 => pi_8_0_port, G2 => 
                           gi_7_0_port, P2 => pi_7_0_port, gout => gi_8_1_port,
                           pout => pi_8_1_port);
   pg_port2_1_9 : PG_36 port map( G1 => gi_9_0_port, P1 => pi_9_0_port, G2 => 
                           gi_8_0_port, P2 => pi_8_0_port, gout => n_1041, pout
                           => n_1042);
   pg_port2_1_10 : PG_35 port map( G1 => gi_10_0_port, P1 => pi_10_0_port, G2 
                           => gi_9_0_port, P2 => pi_9_0_port, gout => n_1043, 
                           pout => n_1044);
   pg_port2_1_11 : PG_34 port map( G1 => gi_11_0_port, P1 => pi_11_0_port, G2 
                           => gi_10_0_port, P2 => pi_10_0_port, gout => n_1045,
                           pout => n_1046);
   pg_port2_1_12 : PG_33 port map( G1 => gi_12_0_port, P1 => pi_12_0_port, G2 
                           => gi_11_0_port, P2 => pi_11_0_port, gout => 
                           gi_12_1_port, pout => pi_12_1_port);
   pg_port2_1_13 : PG_32 port map( G1 => gi_13_0_port, P1 => pi_13_0_port, G2 
                           => gi_12_0_port, P2 => pi_12_0_port, gout => n_1047,
                           pout => n_1048);
   pg_port2_1_14 : PG_31 port map( G1 => gi_14_0_port, P1 => pi_14_0_port, G2 
                           => gi_13_0_port, P2 => pi_13_0_port, gout => n_1049,
                           pout => n_1050);
   pg_port2_1_15 : PG_30 port map( G1 => gi_15_0_port, P1 => pi_15_0_port, G2 
                           => gi_14_0_port, P2 => pi_14_0_port, gout => n_1051,
                           pout => n_1052);
   pg_port2_1_16 : PG_29 port map( G1 => gi_16_0_port, P1 => pi_16_0_port, G2 
                           => gi_15_0_port, P2 => pi_15_0_port, gout => 
                           gi_16_1_port, pout => pi_16_1_port);
   pg_port2_1_17 : PG_28 port map( G1 => gi_17_0_port, P1 => pi_17_0_port, G2 
                           => gi_16_0_port, P2 => pi_16_0_port, gout => n_1053,
                           pout => n_1054);
   pg_port2_1_18 : PG_27 port map( G1 => gi_18_0_port, P1 => pi_18_0_port, G2 
                           => gi_17_0_port, P2 => pi_17_0_port, gout => n_1055,
                           pout => n_1056);
   pg_port2_1_19 : PG_26 port map( G1 => gi_19_0_port, P1 => pi_19_0_port, G2 
                           => gi_18_0_port, P2 => pi_18_0_port, gout => n_1057,
                           pout => n_1058);
   pg_port2_1_20 : PG_25 port map( G1 => gi_20_0_port, P1 => pi_20_0_port, G2 
                           => gi_19_0_port, P2 => pi_19_0_port, gout => 
                           gi_20_1_port, pout => pi_20_1_port);
   pg_port2_1_21 : PG_24 port map( G1 => gi_21_0_port, P1 => pi_21_0_port, G2 
                           => gi_20_0_port, P2 => pi_20_0_port, gout => n_1059,
                           pout => n_1060);
   pg_port2_1_22 : PG_23 port map( G1 => gi_22_0_port, P1 => pi_22_0_port, G2 
                           => gi_21_0_port, P2 => pi_21_0_port, gout => n_1061,
                           pout => n_1062);
   pg_port2_1_23 : PG_22 port map( G1 => gi_23_0_port, P1 => pi_23_0_port, G2 
                           => gi_22_0_port, P2 => pi_22_0_port, gout => n_1063,
                           pout => n_1064);
   pg_port2_1_24 : PG_21 port map( G1 => gi_24_0_port, P1 => pi_24_0_port, G2 
                           => gi_23_0_port, P2 => pi_23_0_port, gout => 
                           gi_24_1_port, pout => pi_24_1_port);
   pg_port2_1_25 : PG_20 port map( G1 => gi_25_0_port, P1 => pi_25_0_port, G2 
                           => gi_24_0_port, P2 => pi_24_0_port, gout => n_1065,
                           pout => n_1066);
   pg_port2_1_26 : PG_19 port map( G1 => gi_26_0_port, P1 => pi_26_0_port, G2 
                           => gi_25_0_port, P2 => pi_25_0_port, gout => n_1067,
                           pout => n_1068);
   pg_port2_1_27 : PG_18 port map( G1 => gi_27_0_port, P1 => pi_27_0_port, G2 
                           => gi_26_0_port, P2 => pi_26_0_port, gout => n_1069,
                           pout => n_1070);
   pg_port2_1_28 : PG_17 port map( G1 => gi_28_0_port, P1 => pi_28_0_port, G2 
                           => gi_27_0_port, P2 => pi_27_0_port, gout => 
                           gi_28_1_port, pout => pi_28_1_port);
   pg_port2_1_29 : PG_16 port map( G1 => gi_29_0_port, P1 => pi_29_0_port, G2 
                           => gi_28_0_port, P2 => pi_28_0_port, gout => n_1071,
                           pout => n_1072);
   pg_port2_1_30 : PG_15 port map( G1 => gi_30_0_port, P1 => pi_30_0_port, G2 
                           => gi_29_0_port, P2 => pi_29_0_port, gout => n_1073,
                           pout => n_1074);
   pg_port2_1_31 : PG_14 port map( G1 => gi_31_0_port, P1 => pi_31_0_port, G2 
                           => gi_30_0_port, P2 => pi_30_0_port, gout => n_1075,
                           pout => n_1076);
   pg_port2_1_32 : PG_13 port map( G1 => gi_32_0_port, P1 => pi_32_0_port, G2 
                           => gi_31_0_port, P2 => pi_31_0_port, gout => 
                           gi_32_1_port, pout => pi_32_1_port);
   g_port_0 : G_51 port map( G1 => gi_4_1_port, P => pi_4_1_port, G2 => 
                           gi_2_1_port, Co => Co_0_port);
   pg_port2_0_1_2 : PG_12 port map( G1 => gi_8_1_port, P1 => pi_8_1_port, G2 =>
                           gi_4_1_port, P2 => pi_4_1_port, gout => gi_8_2_port,
                           pout => pi_8_2_port);
   pg_port2_0_2_3 : PG_11 port map( G1 => gi_12_1_port, P1 => pi_12_1_port, G2 
                           => gi_8_1_port, P2 => pi_8_1_port, gout => 
                           gi_12_2_port, pout => pi_12_2_port);
   pg_port2_0_3_4 : PG_10 port map( G1 => gi_16_1_port, P1 => pi_16_1_port, G2 
                           => gi_12_1_port, P2 => pi_12_1_port, gout => 
                           gi_16_2_port, pout => pi_16_2_port);
   pg_port2_0_4_5 : PG_9 port map( G1 => gi_20_1_port, P1 => pi_20_1_port, G2 
                           => gi_16_1_port, P2 => pi_16_1_port, gout => 
                           gi_20_2_port, pout => pi_20_2_port);
   pg_port2_0_5_6 : PG_8 port map( G1 => gi_24_1_port, P1 => pi_24_1_port, G2 
                           => gi_20_1_port, P2 => pi_20_1_port, gout => 
                           gi_24_2_port, pout => pi_24_2_port);
   pg_port2_0_6_7 : PG_7 port map( G1 => gi_28_1_port, P1 => pi_28_1_port, G2 
                           => gi_24_1_port, P2 => pi_24_1_port, gout => 
                           gi_28_2_port, pout => pi_28_2_port);
   pg_port2_0_7_8 : PG_6 port map( G1 => gi_32_1_port, P1 => pi_32_1_port, G2 
                           => gi_28_1_port, P2 => pi_28_1_port, gout => 
                           gi_32_2_port, pout => pi_32_2_port);
   g_port_1_2 : G_50 port map( G1 => gi_8_2_port, P => pi_8_2_port, G2 => 
                           Co_0_port, Co => Co_1_port);
   pg_port2_1_1_4 : PG_5 port map( G1 => gi_16_2_port, P1 => pi_16_2_port, G2 
                           => gi_12_2_port, P2 => pi_12_2_port, gout => 
                           gi_16_3_port, pout => pi_16_3_port);
   pg_port2_1_2_6 : PG_4 port map( G1 => gi_24_2_port, P1 => pi_24_2_port, G2 
                           => gi_20_2_port, P2 => pi_20_2_port, gout => 
                           gi_24_3_port, pout => pi_24_3_port);
   pg_port2_1_3_8 : PG_3 port map( G1 => gi_32_2_port, P1 => pi_32_2_port, G2 
                           => gi_28_2_port, P2 => pi_28_2_port, gout => 
                           gi_32_3_port, pout => pi_32_3_port);
   g_port_2_3 : G_49 port map( G1 => gi_12_2_port, P => pi_12_2_port, G2 => 
                           Co_1_port, Co => Co_2_port);
   g_port_2_4 : G_48 port map( G1 => gi_16_3_port, P => pi_16_3_port, G2 => 
                           Co_1_port, Co => Co_3_port);
   pg_port2_2_1_7 : PG_2 port map( G1 => gi_28_2_port, P1 => pi_28_2_port, G2 
                           => gi_24_3_port, P2 => pi_24_3_port, gout => 
                           gi_28_4_port, pout => pi_28_4_port);
   pg_port2_2_1_8 : PG_1 port map( G1 => gi_32_3_port, P1 => pi_32_3_port, G2 
                           => gi_24_3_port, P2 => pi_24_3_port, gout => 
                           gi_32_4_port, pout => pi_32_4_port);
   g_port_3_5 : G_47 port map( G1 => gi_20_2_port, P => pi_20_2_port, G2 => 
                           Co_3_port, Co => Co_4_port);
   g_port_3_6 : G_46 port map( G1 => gi_24_3_port, P => pi_24_3_port, G2 => 
                           Co_3_port, Co => Co_5_port);
   g_port_3_7 : G_45 port map( G1 => gi_28_4_port, P => pi_28_4_port, G2 => 
                           Co_3_port, Co => Co_6_port);
   g_port_3_8 : G_44 port map( G1 => gi_32_4_port, P => pi_32_4_port, G2 => 
                           Co_3_port, Co => Co_7_port);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0;

architecture SYN_ARCH2 of ND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P4_ADDER_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4_ADDER_NBIT32;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32 is

   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal Cout_gen_6_port, Cout_gen_5_port, Cout_gen_4_port, Cout_gen_3_port, 
      Cout_gen_2_port, Cout_gen_1_port, Cout_gen_0_port : std_logic;

begin
   
   carry_logic : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 port map( A(31) => 
                           A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           Cin => Cin, Co(7) => Cout, Co(6) => Cout_gen_6_port,
                           Co(5) => Cout_gen_5_port, Co(4) => Cout_gen_4_port, 
                           Co(3) => Cout_gen_3_port, Co(2) => Cout_gen_2_port, 
                           Co(1) => Cout_gen_1_port, Co(0) => Cout_gen_0_port);
   sum_logic : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31),
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           Cout_gen_6_port, Ci(6) => Cout_gen_5_port, Ci(5) => 
                           Cout_gen_4_port, Ci(4) => Cout_gen_3_port, Ci(3) => 
                           Cout_gen_2_port, Ci(2) => Cout_gen_1_port, Ci(1) => 
                           Cout_gen_0_port, Ci(0) => Cin, S(31) => S(31), S(30)
                           => S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
         downto 0);  LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE : in std_logic;  
         OUTPUT : out std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32;

architecture SYN_BEHAVIORAL of SHIFTER_GENERIC_N32 is

   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_lbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sla_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, 
      N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35
      , N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, 
      N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64
      , N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109, N110, N111,
      N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, 
      N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, 
      N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, 
      N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N202, N203, N204, 
      N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, 
      N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, 
      N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, 
      N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, 
      N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, 
      N265, n13_port, n14_port, n15_port, n16_port, n17_port, n18_port, 
      n19_port, n20_port, n21_port, n22_port, n23_port, n24_port, n25_port, 
      n26_port, n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, 
      n33_port, n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, 
      n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, 
      n47_port, n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, 
      n54_port, n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, 
      n61_port, n62_port, n63_port, n64_port, n65_port, n66_port, n67_port, 
      n68_port, n69_port, n70_port, n71, n72, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n1 : 
      std_logic;

begin
   
   n13_port <= '0';
   n14_port <= '0';
   n15_port <= '0';
   n16_port <= '0';
   n17_port <= '0';
   n18_port <= '0';
   U13 : NAND2_X1 port map( A1 => n19_port, A2 => n20_port, ZN => OUTPUT(9));
   U14 : AOI222_X1 port map( A1 => N211, A2 => n21_port, B1 => N114, B2 => 
                           n22_port, C1 => N146, C2 => n23_port, ZN => n20_port
                           );
   U15 : AOI222_X1 port map( A1 => N48, A2 => n24_port, B1 => N243, B2 => 
                           n25_port, C1 => N16, C2 => n26_port, ZN => n19_port)
                           ;
   U16 : NAND2_X1 port map( A1 => n27_port, A2 => n28_port, ZN => OUTPUT(8));
   U17 : AOI222_X1 port map( A1 => N210, A2 => n21_port, B1 => N113, B2 => 
                           n22_port, C1 => N145, C2 => n23_port, ZN => n28_port
                           );
   U18 : AOI222_X1 port map( A1 => N47, A2 => n24_port, B1 => N242, B2 => 
                           n25_port, C1 => N15, C2 => n26_port, ZN => n27_port)
                           ;
   U19 : NAND2_X1 port map( A1 => n29_port, A2 => n30_port, ZN => OUTPUT(7));
   U20 : AOI222_X1 port map( A1 => N209, A2 => n21_port, B1 => N112, B2 => 
                           n22_port, C1 => N144, C2 => n23_port, ZN => n30_port
                           );
   U21 : AOI222_X1 port map( A1 => N46, A2 => n24_port, B1 => N241, B2 => 
                           n25_port, C1 => N14, C2 => n26_port, ZN => n29_port)
                           ;
   U22 : NAND2_X1 port map( A1 => n31_port, A2 => n32_port, ZN => OUTPUT(6));
   U23 : AOI222_X1 port map( A1 => N208, A2 => n21_port, B1 => N111, B2 => 
                           n22_port, C1 => N143, C2 => n23_port, ZN => n32_port
                           );
   U24 : AOI222_X1 port map( A1 => N45, A2 => n24_port, B1 => N240, B2 => 
                           n25_port, C1 => N13, C2 => n26_port, ZN => n31_port)
                           ;
   U25 : NAND2_X1 port map( A1 => n33_port, A2 => n34_port, ZN => OUTPUT(5));
   U26 : AOI222_X1 port map( A1 => N207, A2 => n21_port, B1 => N110, B2 => 
                           n22_port, C1 => N142, C2 => n23_port, ZN => n34_port
                           );
   U27 : AOI222_X1 port map( A1 => N44, A2 => n24_port, B1 => N239, B2 => 
                           n25_port, C1 => N12, C2 => n26_port, ZN => n33_port)
                           ;
   U28 : NAND2_X1 port map( A1 => n35_port, A2 => n36_port, ZN => OUTPUT(4));
   U29 : AOI222_X1 port map( A1 => N206, A2 => n21_port, B1 => N109, B2 => 
                           n22_port, C1 => N141, C2 => n23_port, ZN => n36_port
                           );
   U30 : AOI222_X1 port map( A1 => N43, A2 => n24_port, B1 => N238, B2 => 
                           n25_port, C1 => N11, C2 => n26_port, ZN => n35_port)
                           ;
   U31 : NAND2_X1 port map( A1 => n37_port, A2 => n38_port, ZN => OUTPUT(3));
   U32 : AOI222_X1 port map( A1 => N205, A2 => n21_port, B1 => N108, B2 => 
                           n22_port, C1 => N140, C2 => n23_port, ZN => n38_port
                           );
   U33 : AOI222_X1 port map( A1 => N42, A2 => n24_port, B1 => N237, B2 => 
                           n25_port, C1 => N10, C2 => n26_port, ZN => n37_port)
                           ;
   U34 : NAND2_X1 port map( A1 => n39_port, A2 => n40_port, ZN => OUTPUT(31));
   U35 : AOI222_X1 port map( A1 => N233, A2 => n21_port, B1 => N136, B2 => 
                           n22_port, C1 => N168, C2 => n23_port, ZN => n40_port
                           );
   U36 : AOI222_X1 port map( A1 => N70, A2 => n24_port, B1 => N265, B2 => 
                           n25_port, C1 => N38, C2 => n26_port, ZN => n39_port)
                           ;
   U37 : NAND2_X1 port map( A1 => n41_port, A2 => n42_port, ZN => OUTPUT(30));
   U38 : AOI222_X1 port map( A1 => N232, A2 => n21_port, B1 => N135, B2 => 
                           n22_port, C1 => N167, C2 => n23_port, ZN => n42_port
                           );
   U39 : AOI222_X1 port map( A1 => N69, A2 => n24_port, B1 => N264, B2 => 
                           n25_port, C1 => N37, C2 => n26_port, ZN => n41_port)
                           ;
   U40 : NAND2_X1 port map( A1 => n43_port, A2 => n44_port, ZN => OUTPUT(2));
   U41 : AOI222_X1 port map( A1 => N204, A2 => n21_port, B1 => N107, B2 => 
                           n22_port, C1 => N139, C2 => n23_port, ZN => n44_port
                           );
   U42 : AOI222_X1 port map( A1 => N41, A2 => n24_port, B1 => N236, B2 => 
                           n25_port, C1 => N9, C2 => n26_port, ZN => n43_port);
   U43 : NAND2_X1 port map( A1 => n45_port, A2 => n46_port, ZN => OUTPUT(29));
   U44 : AOI222_X1 port map( A1 => N231, A2 => n21_port, B1 => N134, B2 => 
                           n22_port, C1 => N166, C2 => n23_port, ZN => n46_port
                           );
   U45 : AOI222_X1 port map( A1 => N68, A2 => n24_port, B1 => N263, B2 => 
                           n25_port, C1 => N36, C2 => n26_port, ZN => n45_port)
                           ;
   U46 : NAND2_X1 port map( A1 => n47_port, A2 => n48_port, ZN => OUTPUT(28));
   U47 : AOI222_X1 port map( A1 => N230, A2 => n21_port, B1 => N133, B2 => 
                           n22_port, C1 => N165, C2 => n23_port, ZN => n48_port
                           );
   U48 : AOI222_X1 port map( A1 => N67, A2 => n24_port, B1 => N262, B2 => 
                           n25_port, C1 => N35, C2 => n26_port, ZN => n47_port)
                           ;
   U49 : NAND2_X1 port map( A1 => n49_port, A2 => n50_port, ZN => OUTPUT(27));
   U50 : AOI222_X1 port map( A1 => N229, A2 => n21_port, B1 => N132, B2 => 
                           n22_port, C1 => N164, C2 => n23_port, ZN => n50_port
                           );
   U51 : AOI222_X1 port map( A1 => N66, A2 => n24_port, B1 => N261, B2 => 
                           n25_port, C1 => N34, C2 => n26_port, ZN => n49_port)
                           ;
   U52 : NAND2_X1 port map( A1 => n51_port, A2 => n52_port, ZN => OUTPUT(26));
   U53 : AOI222_X1 port map( A1 => N228, A2 => n21_port, B1 => N131, B2 => 
                           n22_port, C1 => N163, C2 => n23_port, ZN => n52_port
                           );
   U54 : AOI222_X1 port map( A1 => N65, A2 => n24_port, B1 => N260, B2 => 
                           n25_port, C1 => N33, C2 => n26_port, ZN => n51_port)
                           ;
   U55 : NAND2_X1 port map( A1 => n53_port, A2 => n54_port, ZN => OUTPUT(25));
   U56 : AOI222_X1 port map( A1 => N227, A2 => n21_port, B1 => N130, B2 => 
                           n22_port, C1 => N162, C2 => n23_port, ZN => n54_port
                           );
   U57 : AOI222_X1 port map( A1 => N64, A2 => n24_port, B1 => N259, B2 => 
                           n25_port, C1 => N32, C2 => n26_port, ZN => n53_port)
                           ;
   U58 : NAND2_X1 port map( A1 => n55_port, A2 => n56_port, ZN => OUTPUT(24));
   U59 : AOI222_X1 port map( A1 => N226, A2 => n21_port, B1 => N129, B2 => 
                           n22_port, C1 => N161, C2 => n23_port, ZN => n56_port
                           );
   U60 : AOI222_X1 port map( A1 => N63, A2 => n24_port, B1 => N258, B2 => 
                           n25_port, C1 => N31, C2 => n26_port, ZN => n55_port)
                           ;
   U61 : NAND2_X1 port map( A1 => n57_port, A2 => n58_port, ZN => OUTPUT(23));
   U62 : AOI222_X1 port map( A1 => N225, A2 => n21_port, B1 => N128, B2 => 
                           n22_port, C1 => N160, C2 => n23_port, ZN => n58_port
                           );
   U63 : AOI222_X1 port map( A1 => N62, A2 => n24_port, B1 => N257, B2 => 
                           n25_port, C1 => N30, C2 => n26_port, ZN => n57_port)
                           ;
   U64 : NAND2_X1 port map( A1 => n59_port, A2 => n60_port, ZN => OUTPUT(22));
   U65 : AOI222_X1 port map( A1 => N224, A2 => n21_port, B1 => N127, B2 => 
                           n22_port, C1 => N159, C2 => n23_port, ZN => n60_port
                           );
   U66 : AOI222_X1 port map( A1 => N61, A2 => n24_port, B1 => N256, B2 => 
                           n25_port, C1 => N29, C2 => n26_port, ZN => n59_port)
                           ;
   U67 : NAND2_X1 port map( A1 => n61_port, A2 => n62_port, ZN => OUTPUT(21));
   U68 : AOI222_X1 port map( A1 => N223, A2 => n21_port, B1 => N126, B2 => 
                           n22_port, C1 => N158, C2 => n23_port, ZN => n62_port
                           );
   U69 : AOI222_X1 port map( A1 => N60, A2 => n24_port, B1 => N255, B2 => 
                           n25_port, C1 => N28, C2 => n26_port, ZN => n61_port)
                           ;
   U70 : NAND2_X1 port map( A1 => n63_port, A2 => n64_port, ZN => OUTPUT(20));
   U71 : AOI222_X1 port map( A1 => N222, A2 => n21_port, B1 => N125, B2 => 
                           n22_port, C1 => N157, C2 => n23_port, ZN => n64_port
                           );
   U72 : AOI222_X1 port map( A1 => N59, A2 => n24_port, B1 => N254, B2 => 
                           n25_port, C1 => N27, C2 => n26_port, ZN => n63_port)
                           ;
   U73 : NAND2_X1 port map( A1 => n65_port, A2 => n66_port, ZN => OUTPUT(1));
   U74 : AOI222_X1 port map( A1 => N203, A2 => n21_port, B1 => N106, B2 => 
                           n22_port, C1 => N138, C2 => n23_port, ZN => n66_port
                           );
   U75 : AOI222_X1 port map( A1 => N40, A2 => n24_port, B1 => N235, B2 => 
                           n25_port, C1 => N8, C2 => n26_port, ZN => n65_port);
   U76 : NAND2_X1 port map( A1 => n67_port, A2 => n68_port, ZN => OUTPUT(19));
   U77 : AOI222_X1 port map( A1 => N221, A2 => n21_port, B1 => N124, B2 => 
                           n22_port, C1 => N156, C2 => n23_port, ZN => n68_port
                           );
   U78 : AOI222_X1 port map( A1 => N58, A2 => n24_port, B1 => N253, B2 => 
                           n25_port, C1 => N26, C2 => n26_port, ZN => n67_port)
                           ;
   U79 : NAND2_X1 port map( A1 => n69_port, A2 => n70_port, ZN => OUTPUT(18));
   U80 : AOI222_X1 port map( A1 => N220, A2 => n21_port, B1 => N123, B2 => 
                           n22_port, C1 => N155, C2 => n23_port, ZN => n70_port
                           );
   U81 : AOI222_X1 port map( A1 => N57, A2 => n24_port, B1 => N252, B2 => 
                           n25_port, C1 => N25, C2 => n26_port, ZN => n69_port)
                           ;
   U82 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => OUTPUT(17));
   U83 : AOI222_X1 port map( A1 => N219, A2 => n21_port, B1 => N122, B2 => 
                           n22_port, C1 => N154, C2 => n23_port, ZN => n72);
   U84 : AOI222_X1 port map( A1 => N56, A2 => n24_port, B1 => N251, B2 => 
                           n25_port, C1 => N24, C2 => n26_port, ZN => n71);
   U85 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => OUTPUT(16));
   U86 : AOI222_X1 port map( A1 => N218, A2 => n21_port, B1 => N121, B2 => 
                           n22_port, C1 => N153, C2 => n23_port, ZN => n74);
   U87 : AOI222_X1 port map( A1 => N55, A2 => n24_port, B1 => N250, B2 => 
                           n25_port, C1 => N23, C2 => n26_port, ZN => n73);
   U88 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => OUTPUT(15));
   U89 : AOI222_X1 port map( A1 => N217, A2 => n21_port, B1 => N120, B2 => 
                           n22_port, C1 => N152, C2 => n23_port, ZN => n76);
   U90 : AOI222_X1 port map( A1 => N54, A2 => n24_port, B1 => N249, B2 => 
                           n25_port, C1 => N22, C2 => n26_port, ZN => n75);
   U91 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => OUTPUT(14));
   U92 : AOI222_X1 port map( A1 => N216, A2 => n21_port, B1 => N119, B2 => 
                           n22_port, C1 => N151, C2 => n23_port, ZN => n78);
   U93 : AOI222_X1 port map( A1 => N53, A2 => n24_port, B1 => N248, B2 => 
                           n25_port, C1 => N21, C2 => n26_port, ZN => n77);
   U94 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => OUTPUT(13));
   U95 : AOI222_X1 port map( A1 => N215, A2 => n21_port, B1 => N118, B2 => 
                           n22_port, C1 => N150, C2 => n23_port, ZN => n80);
   U96 : AOI222_X1 port map( A1 => N52, A2 => n24_port, B1 => N247, B2 => 
                           n25_port, C1 => N20, C2 => n26_port, ZN => n79);
   U97 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => OUTPUT(12));
   U98 : AOI222_X1 port map( A1 => N214, A2 => n21_port, B1 => N117, B2 => 
                           n22_port, C1 => N149, C2 => n23_port, ZN => n82);
   U99 : AOI222_X1 port map( A1 => N51, A2 => n24_port, B1 => N246, B2 => 
                           n25_port, C1 => N19, C2 => n26_port, ZN => n81);
   U100 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => OUTPUT(11));
   U101 : AOI222_X1 port map( A1 => N213, A2 => n21_port, B1 => N116, B2 => 
                           n22_port, C1 => N148, C2 => n23_port, ZN => n84);
   U102 : AOI222_X1 port map( A1 => N50, A2 => n24_port, B1 => N245, B2 => 
                           n25_port, C1 => N18, C2 => n26_port, ZN => n83);
   U103 : NAND2_X1 port map( A1 => n85, A2 => n86, ZN => OUTPUT(10));
   U104 : AOI222_X1 port map( A1 => N212, A2 => n21_port, B1 => N115, B2 => 
                           n22_port, C1 => N147, C2 => n23_port, ZN => n86);
   U105 : AOI222_X1 port map( A1 => N49, A2 => n24_port, B1 => N244, B2 => 
                           n25_port, C1 => N17, C2 => n26_port, ZN => n85);
   U106 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => OUTPUT(0));
   U107 : AOI222_X1 port map( A1 => N202, A2 => n21_port, B1 => N105, B2 => 
                           n22_port, C1 => N137, C2 => n23_port, ZN => n88);
   U111 : NOR2_X1 port map( A1 => n92, A2 => LOGIC_ARITH, ZN => n91);
   U112 : INV_X1 port map( A => SHIFT_ROTATE, ZN => n92);
   U113 : AOI222_X1 port map( A1 => N39, A2 => n24_port, B1 => N234, B2 => 
                           n25_port, C1 => N7, C2 => n26_port, ZN => n87);
   U116 : AND2_X1 port map( A1 => LOGIC_ARITH, A2 => SHIFT_ROTATE, ZN => n89);
   U118 : INV_X1 port map( A => LEFT_RIGHT, ZN => n90);
   sll_49 : SHIFTER_GENERIC_N32_DW01_ash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n13_port, SH(4) =>
                           n1, SH(3) => B(3), SH(2) => B(2), SH(1) => B(1), 
                           SH(0) => B(0), SH_TC => n13_port, B(31) => N265, 
                           B(30) => N264, B(29) => N263, B(28) => N262, B(27) 
                           => N261, B(26) => N260, B(25) => N259, B(24) => N258
                           , B(23) => N257, B(22) => N256, B(21) => N255, B(20)
                           => N254, B(19) => N253, B(18) => N252, B(17) => N251
                           , B(16) => N250, B(15) => N249, B(14) => N248, B(13)
                           => N247, B(12) => N246, B(11) => N245, B(10) => N244
                           , B(9) => N243, B(8) => N242, B(7) => N241, B(6) => 
                           N240, B(5) => N239, B(4) => N238, B(3) => N237, B(2)
                           => N236, B(1) => N235, B(0) => N234);
   sla_47 : SHIFTER_GENERIC_N32_DW_sla_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n1, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n14_port, B(31) => N233, B(30) => N232, B(29) => 
                           N231, B(28) => N230, B(27) => N229, B(26) => N228, 
                           B(25) => N227, B(24) => N226, B(23) => N225, B(22) 
                           => N224, B(21) => N223, B(20) => N222, B(19) => N221
                           , B(18) => N220, B(17) => N219, B(16) => N218, B(15)
                           => N217, B(14) => N216, B(13) => N215, B(12) => N214
                           , B(11) => N213, B(10) => N212, B(9) => N211, B(8) 
                           => N210, B(7) => N209, B(6) => N208, B(5) => N207, 
                           B(4) => N206, B(3) => N205, B(2) => N204, B(1) => 
                           N203, B(0) => N202);
   srl_42 : SHIFTER_GENERIC_N32_DW_rash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n15_port, SH(4) =>
                           n1, SH(3) => B(3), SH(2) => B(2), SH(1) => B(1), 
                           SH(0) => B(0), SH_TC => n15_port, B(31) => N168, 
                           B(30) => N167, B(29) => N166, B(28) => N165, B(27) 
                           => N164, B(26) => N163, B(25) => N162, B(24) => N161
                           , B(23) => N160, B(22) => N159, B(21) => N158, B(20)
                           => N157, B(19) => N156, B(18) => N155, B(17) => N154
                           , B(16) => N153, B(15) => N152, B(14) => N151, B(13)
                           => N150, B(12) => N149, B(11) => N148, B(10) => N147
                           , B(9) => N146, B(8) => N145, B(7) => N144, B(6) => 
                           N143, B(5) => N142, B(4) => N141, B(3) => N140, B(2)
                           => N139, B(1) => N138, B(0) => N137);
   sra_40 : SHIFTER_GENERIC_N32_DW_sra_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n1, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n16_port, B(31) => N136, B(30) => N135, B(29) => 
                           N134, B(28) => N133, B(27) => N132, B(26) => N131, 
                           B(25) => N130, B(24) => N129, B(23) => N128, B(22) 
                           => N127, B(21) => N126, B(20) => N125, B(19) => N124
                           , B(18) => N123, B(17) => N122, B(16) => N121, B(15)
                           => N120, B(14) => N119, B(13) => N118, B(12) => N117
                           , B(11) => N116, B(10) => N115, B(9) => N114, B(8) 
                           => N113, B(7) => N112, B(6) => N111, B(5) => N110, 
                           B(4) => N109, B(3) => N108, B(2) => N107, B(1) => 
                           N106, B(0) => N105);
   rol_33 : SHIFTER_GENERIC_N32_DW_lbsh_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n1, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n17_port, B(31) => N70, B(30) => N69, B(29) => 
                           N68, B(28) => N67, B(27) => N66, B(26) => N65, B(25)
                           => N64, B(24) => N63, B(23) => N62, B(22) => N61, 
                           B(21) => N60, B(20) => N59, B(19) => N58, B(18) => 
                           N57, B(17) => N56, B(16) => N55, B(15) => N54, B(14)
                           => N53, B(13) => N52, B(12) => N51, B(11) => N50, 
                           B(10) => N49, B(9) => N48, B(8) => N47, B(7) => N46,
                           B(6) => N45, B(5) => N44, B(4) => N43, B(3) => N42, 
                           B(2) => N41, B(1) => N40, B(0) => N39);
   ror_31 : SHIFTER_GENERIC_N32_DW_rbsh_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n1, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n18_port, B(31) => N38, B(30) => N37, B(29) => 
                           N36, B(28) => N35, B(27) => N34, B(26) => N33, B(25)
                           => N32, B(24) => N31, B(23) => N30, B(22) => N29, 
                           B(21) => N28, B(20) => N27, B(19) => N26, B(18) => 
                           N25, B(17) => N24, B(16) => N23, B(15) => N22, B(14)
                           => N21, B(13) => N20, B(12) => N19, B(11) => N18, 
                           B(10) => N17, B(9) => N16, B(8) => N15, B(7) => N14,
                           B(6) => N13, B(5) => N12, B(4) => N11, B(3) => N10, 
                           B(2) => N9, B(1) => N8, B(0) => N7);
   U5 : AND2_X2 port map( A1 => n89, A2 => n90, ZN => n23_port);
   U6 : AND2_X2 port map( A1 => n91, A2 => n90, ZN => n22_port);
   U7 : AND2_X2 port map( A1 => LEFT_RIGHT, A2 => n89, ZN => n25_port);
   U8 : AND2_X2 port map( A1 => LEFT_RIGHT, A2 => n91, ZN => n21_port);
   U9 : NOR2_X4 port map( A1 => n90, A2 => SHIFT_ROTATE, ZN => n24_port);
   U10 : NOR2_X4 port map( A1 => LEFT_RIGHT, A2 => SHIFT_ROTATE, ZN => n26_port
                           );
   U108 : BUF_X4 port map( A => B(4), Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity comparator is

   port( DATA1 : in std_logic_vector (31 downto 0);  DATA2i : in std_logic;  
         tipo : in std_logic_vector (0 to 5);  OUTALU : out std_logic_vector 
         (31 downto 0));

end comparator;

architecture SYN_Architectural of comparator is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N57, N58, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49 : std_logic;

begin
   
   OUTALU_reg_0_inst : DLH_X1 port map( G => N57, D => N58, Q => OUTALU(0));
   OUTALU(1) <= '0';
   OUTALU(2) <= '0';
   OUTALU(3) <= '0';
   OUTALU(4) <= '0';
   OUTALU(5) <= '0';
   OUTALU(6) <= '0';
   OUTALU(7) <= '0';
   OUTALU(8) <= '0';
   OUTALU(9) <= '0';
   OUTALU(10) <= '0';
   OUTALU(11) <= '0';
   OUTALU(12) <= '0';
   OUTALU(13) <= '0';
   OUTALU(14) <= '0';
   OUTALU(15) <= '0';
   OUTALU(16) <= '0';
   OUTALU(17) <= '0';
   OUTALU(18) <= '0';
   OUTALU(19) <= '0';
   OUTALU(20) <= '0';
   OUTALU(21) <= '0';
   OUTALU(22) <= '0';
   OUTALU(23) <= '0';
   OUTALU(24) <= '0';
   OUTALU(25) <= '0';
   OUTALU(26) <= '0';
   OUTALU(27) <= '0';
   OUTALU(28) <= '0';
   OUTALU(29) <= '0';
   OUTALU(30) <= '0';
   OUTALU(31) <= '0';
   U33 : OAI211_X1 port map( C1 => n1, C2 => n2, A => n3, B => n4, ZN => N58);
   U34 : AOI22_X1 port map( A1 => n5, A2 => n2, B1 => n6, B2 => n7, ZN => n4);
   U35 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n10, ZN => n3);
   U36 : INV_X1 port map( A => DATA2i, ZN => n2);
   U37 : AOI21_X1 port map( B1 => n11, B2 => n7, A => n12, ZN => n1);
   U38 : INV_X1 port map( A => n10, ZN => n7);
   U39 : NOR2_X1 port map( A1 => n13, A2 => n14, ZN => n10);
   U40 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n14);
   U41 : NOR4_X1 port map( A1 => DATA1(23), A2 => DATA1(22), A3 => DATA1(21), 
                           A4 => DATA1(20), ZN => n18);
   U42 : NOR4_X1 port map( A1 => DATA1(1), A2 => DATA1(19), A3 => DATA1(18), A4
                           => DATA1(17), ZN => n17);
   U43 : NOR4_X1 port map( A1 => DATA1(16), A2 => DATA1(15), A3 => DATA1(14), 
                           A4 => DATA1(13), ZN => n16);
   U44 : NOR4_X1 port map( A1 => DATA1(12), A2 => DATA1(11), A3 => DATA1(10), 
                           A4 => DATA1(0), ZN => n15);
   U45 : NAND4_X1 port map( A1 => n19, A2 => n20, A3 => n21, A4 => n22, ZN => 
                           n13);
   U46 : NOR4_X1 port map( A1 => DATA1(9), A2 => DATA1(8), A3 => DATA1(7), A4 
                           => DATA1(6), ZN => n22);
   U47 : NOR4_X1 port map( A1 => DATA1(5), A2 => DATA1(4), A3 => DATA1(3), A4 
                           => DATA1(31), ZN => n21);
   U48 : NOR4_X1 port map( A1 => DATA1(30), A2 => DATA1(2), A3 => DATA1(29), A4
                           => DATA1(28), ZN => n20);
   U49 : NOR4_X1 port map( A1 => DATA1(27), A2 => DATA1(26), A3 => DATA1(25), 
                           A4 => DATA1(24), ZN => n19);
   U50 : OR4_X1 port map( A1 => n6, A2 => n5, A3 => n23, A4 => n11, ZN => N57);
   U51 : OAI21_X1 port map( B1 => n24, B2 => n25, A => n26, ZN => n11);
   U52 : INV_X1 port map( A => n27, ZN => n26);
   U53 : AOI21_X1 port map( B1 => n28, B2 => n29, A => n30, ZN => n27);
   U54 : OR2_X1 port map( A1 => n8, A2 => n12, ZN => n23);
   U55 : OAI221_X1 port map( B1 => n31, B2 => n28, C1 => n25, C2 => n32, A => 
                           n33, ZN => n12);
   U56 : INV_X1 port map( A => n34, ZN => n33);
   U57 : AOI211_X1 port map( C1 => n29, C2 => n35, A => n36, B => n37, ZN => 
                           n34);
   U58 : NAND4_X1 port map( A1 => tipo(0), A2 => tipo(1), A3 => n38, A4 => n39,
                           ZN => n28);
   U59 : INV_X1 port map( A => tipo(3), ZN => n38);
   U60 : OAI21_X1 port map( B1 => n40, B2 => n30, A => n41, ZN => n8);
   U61 : NAND4_X1 port map( A1 => tipo(1), A2 => tipo(3), A3 => n42, A4 => n43,
                           ZN => n41);
   U62 : INV_X1 port map( A => n25, ZN => n43);
   U63 : NOR2_X1 port map( A1 => tipo(0), A2 => n39, ZN => n42);
   U64 : OAI221_X1 port map( B1 => n44, B2 => n45, C1 => n24, C2 => n31, A => 
                           n46, ZN => n5);
   U65 : INV_X1 port map( A => n9, ZN => n46);
   U66 : OAI22_X1 port map( A1 => n31, A2 => n32, B1 => n25, B2 => n35, ZN => 
                           n9);
   U67 : NAND2_X1 port map( A1 => tipo(4), A2 => n37, ZN => n25);
   U68 : AND2_X1 port map( A1 => n40, A2 => n29, ZN => n24);
   U69 : NAND3_X1 port map( A1 => n47, A2 => n39, A3 => tipo(0), ZN => n29);
   U70 : NAND3_X1 port map( A1 => tipo(2), A2 => n47, A3 => tipo(0), ZN => n40)
                           ;
   U71 : NAND2_X1 port map( A1 => tipo(5), A2 => tipo(3), ZN => n45);
   U72 : NAND3_X1 port map( A1 => tipo(2), A2 => n48, A3 => tipo(4), ZN => n44)
                           ;
   U73 : XNOR2_X1 port map( A => n49, B => tipo(1), ZN => n48);
   U74 : OAI22_X1 port map( A1 => n35, A2 => n31, B1 => n32, B2 => n30, ZN => 
                           n6);
   U75 : NAND2_X1 port map( A1 => n37, A2 => n36, ZN => n30);
   U76 : INV_X1 port map( A => tipo(5), ZN => n37);
   U77 : NAND4_X1 port map( A1 => tipo(1), A2 => tipo(3), A3 => n39, A4 => n49,
                           ZN => n32);
   U78 : INV_X1 port map( A => tipo(2), ZN => n39);
   U79 : NAND2_X1 port map( A1 => tipo(5), A2 => n36, ZN => n31);
   U80 : INV_X1 port map( A => tipo(4), ZN => n36);
   U81 : NAND3_X1 port map( A1 => n47, A2 => n49, A3 => tipo(2), ZN => n35);
   U82 : INV_X1 port map( A => tipo(0), ZN => n49);
   U83 : NOR2_X1 port map( A1 => tipo(1), A2 => tipo(3), ZN => n47);

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity logic_N32 is

   port( FUNC : in std_logic_vector (0 to 5);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUT_ALU : out std_logic_vector (31 
         downto 0));

end logic_N32;

architecture SYN_Architectural of logic_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n25, n141, n142, n143, n144 : std_logic;

begin
   
   U2 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           OUT_ALU(9));
   U3 : AOI21_X1 port map( B1 => n5, B2 => n2, A => n143, ZN => n3);
   U4 : INV_X1 port map( A => DATA2(9), ZN => n2);
   U5 : AOI221_X1 port map( B1 => n5, B2 => n4, C1 => n141, C2 => DATA1(9), A 
                           => n143, ZN => n1);
   U6 : INV_X1 port map( A => DATA1(9), ZN => n4);
   U7 : OAI22_X1 port map( A1 => n8, A2 => n9, B1 => n10, B2 => n11, ZN => 
                           OUT_ALU(8));
   U8 : AOI21_X1 port map( B1 => n5, B2 => n9, A => n143, ZN => n10);
   U9 : INV_X1 port map( A => DATA2(8), ZN => n9);
   U10 : AOI221_X1 port map( B1 => n5, B2 => n11, C1 => DATA1(8), C2 => n141, A
                           => n143, ZN => n8);
   U11 : INV_X1 port map( A => DATA1(8), ZN => n11);
   U12 : OAI22_X1 port map( A1 => n12, A2 => n13, B1 => n14, B2 => n15, ZN => 
                           OUT_ALU(7));
   U13 : AOI21_X1 port map( B1 => n5, B2 => n13, A => n143, ZN => n14);
   U14 : INV_X1 port map( A => DATA2(7), ZN => n13);
   U15 : AOI221_X1 port map( B1 => n5, B2 => n15, C1 => DATA1(7), C2 => n141, A
                           => n143, ZN => n12);
   U16 : INV_X1 port map( A => DATA1(7), ZN => n15);
   U17 : OAI22_X1 port map( A1 => n16, A2 => n17, B1 => n18, B2 => n19, ZN => 
                           OUT_ALU(6));
   U18 : AOI21_X1 port map( B1 => n5, B2 => n17, A => n143, ZN => n18);
   U19 : INV_X1 port map( A => DATA2(6), ZN => n17);
   U20 : AOI221_X1 port map( B1 => n5, B2 => n19, C1 => DATA1(6), C2 => n141, A
                           => n143, ZN => n16);
   U21 : INV_X1 port map( A => DATA1(6), ZN => n19);
   U22 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => n22, B2 => n23, ZN => 
                           OUT_ALU(5));
   U23 : AOI21_X1 port map( B1 => n5, B2 => n21, A => n143, ZN => n22);
   U24 : INV_X1 port map( A => DATA2(5), ZN => n21);
   U25 : AOI221_X1 port map( B1 => n5, B2 => n23, C1 => DATA1(5), C2 => n141, A
                           => n143, ZN => n20);
   U26 : INV_X1 port map( A => DATA1(5), ZN => n23);
   U27 : OAI22_X1 port map( A1 => n24, A2 => n144, B1 => n26, B2 => n27, ZN => 
                           OUT_ALU(4));
   U28 : AOI21_X1 port map( B1 => n5, B2 => n144, A => n143, ZN => n26);
   U30 : AOI221_X1 port map( B1 => n5, B2 => n27, C1 => DATA1(4), C2 => n141, A
                           => n143, ZN => n24);
   U31 : INV_X1 port map( A => DATA1(4), ZN => n27);
   U32 : OAI22_X1 port map( A1 => n28, A2 => n29, B1 => n30, B2 => n31, ZN => 
                           OUT_ALU(3));
   U33 : AOI21_X1 port map( B1 => n5, B2 => n29, A => n143, ZN => n30);
   U34 : INV_X1 port map( A => DATA2(3), ZN => n29);
   U35 : AOI221_X1 port map( B1 => n5, B2 => n31, C1 => DATA1(3), C2 => n141, A
                           => n143, ZN => n28);
   U36 : INV_X1 port map( A => DATA1(3), ZN => n31);
   U37 : OAI22_X1 port map( A1 => n32, A2 => n33, B1 => n34, B2 => n35, ZN => 
                           OUT_ALU(31));
   U38 : AOI21_X1 port map( B1 => n5, B2 => n33, A => n143, ZN => n34);
   U39 : INV_X1 port map( A => DATA2(31), ZN => n33);
   U40 : AOI221_X1 port map( B1 => n5, B2 => n35, C1 => DATA1(31), C2 => n141, 
                           A => n143, ZN => n32);
   U41 : INV_X1 port map( A => DATA1(31), ZN => n35);
   U42 : OAI22_X1 port map( A1 => n36, A2 => n37, B1 => n38, B2 => n39, ZN => 
                           OUT_ALU(30));
   U43 : AOI21_X1 port map( B1 => n5, B2 => n37, A => n143, ZN => n38);
   U44 : INV_X1 port map( A => DATA2(30), ZN => n37);
   U45 : AOI221_X1 port map( B1 => n5, B2 => n39, C1 => DATA1(30), C2 => n141, 
                           A => n143, ZN => n36);
   U46 : INV_X1 port map( A => DATA1(30), ZN => n39);
   U47 : OAI22_X1 port map( A1 => n40, A2 => n41, B1 => n42, B2 => n43, ZN => 
                           OUT_ALU(2));
   U48 : AOI21_X1 port map( B1 => n5, B2 => n41, A => n143, ZN => n42);
   U49 : INV_X1 port map( A => DATA2(2), ZN => n41);
   U50 : AOI221_X1 port map( B1 => n5, B2 => n43, C1 => DATA1(2), C2 => n141, A
                           => n143, ZN => n40);
   U51 : INV_X1 port map( A => DATA1(2), ZN => n43);
   U52 : OAI22_X1 port map( A1 => n44, A2 => n45, B1 => n46, B2 => n47, ZN => 
                           OUT_ALU(29));
   U53 : AOI21_X1 port map( B1 => n5, B2 => n45, A => n143, ZN => n46);
   U54 : INV_X1 port map( A => DATA2(29), ZN => n45);
   U55 : AOI221_X1 port map( B1 => n5, B2 => n47, C1 => DATA1(29), C2 => n141, 
                           A => n143, ZN => n44);
   U56 : INV_X1 port map( A => DATA1(29), ZN => n47);
   U57 : OAI22_X1 port map( A1 => n48, A2 => n49, B1 => n50, B2 => n51, ZN => 
                           OUT_ALU(28));
   U58 : AOI21_X1 port map( B1 => n5, B2 => n49, A => n143, ZN => n50);
   U59 : INV_X1 port map( A => DATA2(28), ZN => n49);
   U60 : AOI221_X1 port map( B1 => n5, B2 => n51, C1 => DATA1(28), C2 => n141, 
                           A => n143, ZN => n48);
   U61 : INV_X1 port map( A => DATA1(28), ZN => n51);
   U62 : OAI22_X1 port map( A1 => n52, A2 => n53, B1 => n54, B2 => n55, ZN => 
                           OUT_ALU(27));
   U63 : AOI21_X1 port map( B1 => n5, B2 => n53, A => n143, ZN => n54);
   U64 : INV_X1 port map( A => DATA2(27), ZN => n53);
   U65 : AOI221_X1 port map( B1 => n5, B2 => n55, C1 => DATA1(27), C2 => n141, 
                           A => n143, ZN => n52);
   U66 : INV_X1 port map( A => DATA1(27), ZN => n55);
   U67 : OAI22_X1 port map( A1 => n56, A2 => n57, B1 => n58, B2 => n59, ZN => 
                           OUT_ALU(26));
   U68 : AOI21_X1 port map( B1 => n5, B2 => n57, A => n143, ZN => n58);
   U69 : INV_X1 port map( A => DATA2(26), ZN => n57);
   U70 : AOI221_X1 port map( B1 => n5, B2 => n59, C1 => DATA1(26), C2 => n141, 
                           A => n143, ZN => n56);
   U71 : INV_X1 port map( A => DATA1(26), ZN => n59);
   U72 : OAI22_X1 port map( A1 => n60, A2 => n61, B1 => n62, B2 => n63, ZN => 
                           OUT_ALU(25));
   U73 : AOI21_X1 port map( B1 => n5, B2 => n61, A => n143, ZN => n62);
   U74 : INV_X1 port map( A => DATA2(25), ZN => n61);
   U75 : AOI221_X1 port map( B1 => n5, B2 => n63, C1 => DATA1(25), C2 => n141, 
                           A => n143, ZN => n60);
   U76 : INV_X1 port map( A => DATA1(25), ZN => n63);
   U77 : OAI22_X1 port map( A1 => n64, A2 => n65, B1 => n66, B2 => n67, ZN => 
                           OUT_ALU(24));
   U78 : AOI21_X1 port map( B1 => n5, B2 => n65, A => n143, ZN => n66);
   U79 : INV_X1 port map( A => DATA2(24), ZN => n65);
   U80 : AOI221_X1 port map( B1 => n5, B2 => n67, C1 => DATA1(24), C2 => n141, 
                           A => n143, ZN => n64);
   U81 : INV_X1 port map( A => DATA1(24), ZN => n67);
   U82 : OAI22_X1 port map( A1 => n68, A2 => n69, B1 => n70, B2 => n71, ZN => 
                           OUT_ALU(23));
   U83 : AOI21_X1 port map( B1 => n5, B2 => n69, A => n143, ZN => n70);
   U84 : INV_X1 port map( A => DATA2(23), ZN => n69);
   U85 : AOI221_X1 port map( B1 => n5, B2 => n71, C1 => DATA1(23), C2 => n141, 
                           A => n143, ZN => n68);
   U86 : INV_X1 port map( A => DATA1(23), ZN => n71);
   U87 : OAI22_X1 port map( A1 => n72, A2 => n73, B1 => n74, B2 => n75, ZN => 
                           OUT_ALU(22));
   U88 : AOI21_X1 port map( B1 => n5, B2 => n73, A => n143, ZN => n74);
   U89 : INV_X1 port map( A => DATA2(22), ZN => n73);
   U90 : AOI221_X1 port map( B1 => n5, B2 => n75, C1 => DATA1(22), C2 => n141, 
                           A => n143, ZN => n72);
   U91 : INV_X1 port map( A => DATA1(22), ZN => n75);
   U92 : OAI22_X1 port map( A1 => n76, A2 => n77, B1 => n78, B2 => n79, ZN => 
                           OUT_ALU(21));
   U93 : AOI21_X1 port map( B1 => n5, B2 => n77, A => n143, ZN => n78);
   U94 : INV_X1 port map( A => DATA2(21), ZN => n77);
   U95 : AOI221_X1 port map( B1 => n5, B2 => n79, C1 => DATA1(21), C2 => n141, 
                           A => n143, ZN => n76);
   U96 : INV_X1 port map( A => DATA1(21), ZN => n79);
   U97 : OAI22_X1 port map( A1 => n80, A2 => n81, B1 => n82, B2 => n83, ZN => 
                           OUT_ALU(20));
   U98 : AOI21_X1 port map( B1 => n5, B2 => n81, A => n143, ZN => n82);
   U99 : INV_X1 port map( A => DATA2(20), ZN => n81);
   U100 : AOI221_X1 port map( B1 => n5, B2 => n83, C1 => DATA1(20), C2 => n141,
                           A => n143, ZN => n80);
   U101 : INV_X1 port map( A => DATA1(20), ZN => n83);
   U102 : OAI22_X1 port map( A1 => n84, A2 => n85, B1 => n86, B2 => n87, ZN => 
                           OUT_ALU(1));
   U103 : AOI21_X1 port map( B1 => n5, B2 => n85, A => n143, ZN => n86);
   U104 : INV_X1 port map( A => DATA2(1), ZN => n85);
   U105 : AOI221_X1 port map( B1 => n5, B2 => n87, C1 => DATA1(1), C2 => n141, 
                           A => n143, ZN => n84);
   U106 : INV_X1 port map( A => DATA1(1), ZN => n87);
   U107 : OAI22_X1 port map( A1 => n88, A2 => n89, B1 => n90, B2 => n91, ZN => 
                           OUT_ALU(19));
   U108 : AOI21_X1 port map( B1 => n5, B2 => n89, A => n143, ZN => n90);
   U109 : INV_X1 port map( A => DATA2(19), ZN => n89);
   U110 : AOI221_X1 port map( B1 => n5, B2 => n91, C1 => DATA1(19), C2 => n141,
                           A => n143, ZN => n88);
   U111 : INV_X1 port map( A => DATA1(19), ZN => n91);
   U112 : OAI22_X1 port map( A1 => n92, A2 => n93, B1 => n94, B2 => n95, ZN => 
                           OUT_ALU(18));
   U113 : AOI21_X1 port map( B1 => n5, B2 => n93, A => n143, ZN => n94);
   U114 : INV_X1 port map( A => DATA2(18), ZN => n93);
   U115 : AOI221_X1 port map( B1 => n5, B2 => n95, C1 => DATA1(18), C2 => n141,
                           A => n143, ZN => n92);
   U116 : INV_X1 port map( A => DATA1(18), ZN => n95);
   U117 : OAI22_X1 port map( A1 => n96, A2 => n97, B1 => n98, B2 => n99, ZN => 
                           OUT_ALU(17));
   U118 : AOI21_X1 port map( B1 => n5, B2 => n97, A => n143, ZN => n98);
   U119 : INV_X1 port map( A => DATA2(17), ZN => n97);
   U120 : AOI221_X1 port map( B1 => n5, B2 => n99, C1 => DATA1(17), C2 => n141,
                           A => n143, ZN => n96);
   U121 : INV_X1 port map( A => DATA1(17), ZN => n99);
   U122 : OAI22_X1 port map( A1 => n100, A2 => n101, B1 => n102, B2 => n103, ZN
                           => OUT_ALU(16));
   U123 : AOI21_X1 port map( B1 => n5, B2 => n101, A => n143, ZN => n102);
   U124 : INV_X1 port map( A => DATA2(16), ZN => n101);
   U125 : AOI221_X1 port map( B1 => n5, B2 => n103, C1 => DATA1(16), C2 => n141
                           , A => n143, ZN => n100);
   U126 : INV_X1 port map( A => DATA1(16), ZN => n103);
   U127 : OAI22_X1 port map( A1 => n104, A2 => n105, B1 => n106, B2 => n107, ZN
                           => OUT_ALU(15));
   U128 : AOI21_X1 port map( B1 => n5, B2 => n105, A => n143, ZN => n106);
   U129 : INV_X1 port map( A => DATA2(15), ZN => n105);
   U130 : AOI221_X1 port map( B1 => n5, B2 => n107, C1 => DATA1(15), C2 => n141
                           , A => n143, ZN => n104);
   U131 : INV_X1 port map( A => DATA1(15), ZN => n107);
   U132 : OAI22_X1 port map( A1 => n108, A2 => n109, B1 => n110, B2 => n111, ZN
                           => OUT_ALU(14));
   U133 : AOI21_X1 port map( B1 => n5, B2 => n109, A => n143, ZN => n110);
   U134 : INV_X1 port map( A => DATA2(14), ZN => n109);
   U135 : AOI221_X1 port map( B1 => n5, B2 => n111, C1 => DATA1(14), C2 => n141
                           , A => n143, ZN => n108);
   U136 : INV_X1 port map( A => DATA1(14), ZN => n111);
   U137 : OAI22_X1 port map( A1 => n112, A2 => n113, B1 => n114, B2 => n115, ZN
                           => OUT_ALU(13));
   U138 : AOI21_X1 port map( B1 => n5, B2 => n113, A => n143, ZN => n114);
   U139 : INV_X1 port map( A => DATA2(13), ZN => n113);
   U140 : AOI221_X1 port map( B1 => n5, B2 => n115, C1 => DATA1(13), C2 => n141
                           , A => n143, ZN => n112);
   U141 : INV_X1 port map( A => DATA1(13), ZN => n115);
   U142 : OAI22_X1 port map( A1 => n116, A2 => n117, B1 => n118, B2 => n119, ZN
                           => OUT_ALU(12));
   U143 : AOI21_X1 port map( B1 => n5, B2 => n117, A => n143, ZN => n118);
   U144 : INV_X1 port map( A => DATA2(12), ZN => n117);
   U145 : AOI221_X1 port map( B1 => n5, B2 => n119, C1 => DATA1(12), C2 => n141
                           , A => n143, ZN => n116);
   U146 : INV_X1 port map( A => DATA1(12), ZN => n119);
   U147 : OAI22_X1 port map( A1 => n120, A2 => n121, B1 => n122, B2 => n123, ZN
                           => OUT_ALU(11));
   U148 : AOI21_X1 port map( B1 => n5, B2 => n121, A => n143, ZN => n122);
   U149 : INV_X1 port map( A => DATA2(11), ZN => n121);
   U150 : AOI221_X1 port map( B1 => n5, B2 => n123, C1 => DATA1(11), C2 => n141
                           , A => n143, ZN => n120);
   U151 : INV_X1 port map( A => DATA1(11), ZN => n123);
   U152 : OAI22_X1 port map( A1 => n124, A2 => n125, B1 => n126, B2 => n127, ZN
                           => OUT_ALU(10));
   U153 : AOI21_X1 port map( B1 => n5, B2 => n125, A => n143, ZN => n126);
   U154 : INV_X1 port map( A => DATA2(10), ZN => n125);
   U155 : AOI221_X1 port map( B1 => n5, B2 => n127, C1 => DATA1(10), C2 => n141
                           , A => n143, ZN => n124);
   U156 : INV_X1 port map( A => DATA1(10), ZN => n127);
   U157 : OAI22_X1 port map( A1 => n128, A2 => n129, B1 => n130, B2 => n131, ZN
                           => OUT_ALU(0));
   U158 : AOI21_X1 port map( B1 => n5, B2 => n129, A => n143, ZN => n130);
   U159 : INV_X1 port map( A => DATA2(0), ZN => n129);
   U160 : AOI221_X1 port map( B1 => n5, B2 => n131, C1 => DATA1(0), C2 => n141,
                           A => n143, ZN => n128);
   U161 : OAI21_X1 port map( B1 => FUNC(5), B2 => n132, A => n133, ZN => n6);
   U162 : OR3_X1 port map( A1 => n134, A2 => FUNC(2), A3 => n135, ZN => n133);
   U163 : AOI21_X1 port map( B1 => n135, B2 => FUNC(2), A => n134, ZN => n7);
   U164 : NAND4_X1 port map( A1 => FUNC(3), A2 => FUNC(4), A3 => n136, A4 => 
                           n137, ZN => n134);
   U165 : INV_X1 port map( A => FUNC(0), ZN => n137);
   U166 : INV_X1 port map( A => DATA1(0), ZN => n131);
   U168 : NAND4_X1 port map( A1 => FUNC(2), A2 => n139, A3 => n135, A4 => n136,
                           ZN => n138);
   U169 : INV_X1 port map( A => FUNC(1), ZN => n136);
   U170 : INV_X1 port map( A => FUNC(5), ZN => n135);
   U171 : NAND3_X1 port map( A1 => n139, A2 => n140, A3 => FUNC(1), ZN => n132)
                           ;
   U172 : INV_X1 port map( A => FUNC(2), ZN => n140);
   U173 : NOR3_X1 port map( A1 => FUNC(3), A2 => FUNC(0), A3 => FUNC(4), ZN => 
                           n139);
   U29 : INV_X1 port map( A => n7, ZN => n25);
   U167 : INV_X2 port map( A => n25, ZN => n141);
   U174 : NAND2_X4 port map( A1 => n132, A2 => n138, ZN => n5);
   U175 : INV_X1 port map( A => n6, ZN => n142);
   U176 : INV_X4 port map( A => n142, ZN => n143);
   U177 : INV_X1 port map( A => DATA2(4), ZN => n144);

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in26_N_out32 is

   port( IR_out : in std_logic_vector (25 downto 0);  signed_val : in std_logic
         ;  Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in26_N_out32;

architecture SYN_BHV of sign_eval_N_in26_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal Immediate_31, n1 : std_logic;

begin
   Immediate <= ( Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, IR_out(25), IR_out(24), IR_out(23), 
      IR_out(22), IR_out(21), IR_out(20), IR_out(19), IR_out(18), IR_out(17), 
      IR_out(16), IR_out(15), IR_out(14), IR_out(13), IR_out(12), IR_out(11), 
      IR_out(10), IR_out(9), IR_out(8), IR_out(7), IR_out(6), IR_out(5), 
      IR_out(4), IR_out(3), IR_out(2), IR_out(1), IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n1, ZN => Immediate_31);
   U2 : INV_X1 port map( A => IR_out(25), ZN => n1);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in16_N_out32 is

   port( IR_out : in std_logic_vector (15 downto 0);  signed_val : in std_logic
         ;  Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in16_N_out32;

architecture SYN_BHV of sign_eval_N_in16_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal Immediate_31, n1 : std_logic;

begin
   Immediate <= ( Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, IR_out(15), IR_out(14), IR_out(13), 
      IR_out(12), IR_out(11), IR_out(10), IR_out(9), IR_out(8), IR_out(7), 
      IR_out(6), IR_out(5), IR_out(4), IR_out(3), IR_out(2), IR_out(1), 
      IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n1, ZN => Immediate_31);
   U2 : INV_X1 port map( A => IR_out(15), ZN => n1);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in5_N_out32 is

   port( IR_out : in std_logic_vector (4 downto 0);  signed_val : in std_logic;
         Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in5_N_out32;

architecture SYN_BHV of sign_eval_N_in5_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal Immediate_31, n1 : std_logic;

begin
   Immediate <= ( Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, Immediate_31, Immediate_31, Immediate_31, 
      Immediate_31, Immediate_31, Immediate_31, IR_out(4), IR_out(3), IR_out(2)
      , IR_out(1), IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n1, ZN => Immediate_31);
   U2 : INV_X1 port map( A => IR_out(4), ZN => n1);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0;

architecture SYN_STRUCTURAL of MUX21_0 is

   component ND2_766
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_767
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0 port map( A => S, Y => SB);
   UND1 : ND2_0 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_767 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_766 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity load_data is

   port( data_in : in std_logic_vector (31 downto 0);  signed_val, load_op : in
         std_logic;  load_type : in std_logic_vector (1 downto 0);  data_out : 
         out std_logic_vector (31 downto 0));

end load_data;

architecture SYN_bhv_load of load_data is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
      N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64
      , N65, N66, N67, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30 : std_logic;

begin
   
   data_out_reg_31_inst : DLH_X1 port map( G => load_op, D => N67, Q => 
                           data_out(31));
   data_out_reg_30_inst : DLH_X1 port map( G => load_op, D => N66, Q => 
                           data_out(30));
   data_out_reg_29_inst : DLH_X1 port map( G => load_op, D => N65, Q => 
                           data_out(29));
   data_out_reg_28_inst : DLH_X1 port map( G => load_op, D => N64, Q => 
                           data_out(28));
   data_out_reg_27_inst : DLH_X1 port map( G => load_op, D => N63, Q => 
                           data_out(27));
   data_out_reg_26_inst : DLH_X1 port map( G => load_op, D => N62, Q => 
                           data_out(26));
   data_out_reg_25_inst : DLH_X1 port map( G => load_op, D => N61, Q => 
                           data_out(25));
   data_out_reg_24_inst : DLH_X1 port map( G => load_op, D => N60, Q => 
                           data_out(24));
   data_out_reg_23_inst : DLH_X1 port map( G => load_op, D => N59, Q => 
                           data_out(23));
   data_out_reg_22_inst : DLH_X1 port map( G => load_op, D => N58, Q => 
                           data_out(22));
   data_out_reg_21_inst : DLH_X1 port map( G => load_op, D => N57, Q => 
                           data_out(21));
   data_out_reg_20_inst : DLH_X1 port map( G => load_op, D => N56, Q => 
                           data_out(20));
   data_out_reg_19_inst : DLH_X1 port map( G => load_op, D => N55, Q => 
                           data_out(19));
   data_out_reg_18_inst : DLH_X1 port map( G => load_op, D => N54, Q => 
                           data_out(18));
   data_out_reg_17_inst : DLH_X1 port map( G => load_op, D => N53, Q => 
                           data_out(17));
   data_out_reg_16_inst : DLH_X1 port map( G => load_op, D => N52, Q => 
                           data_out(16));
   data_out_reg_15_inst : DLH_X1 port map( G => load_op, D => N51, Q => 
                           data_out(15));
   data_out_reg_14_inst : DLH_X1 port map( G => load_op, D => N50, Q => 
                           data_out(14));
   data_out_reg_13_inst : DLH_X1 port map( G => load_op, D => N49, Q => 
                           data_out(13));
   data_out_reg_12_inst : DLH_X1 port map( G => load_op, D => N48, Q => 
                           data_out(12));
   data_out_reg_11_inst : DLH_X1 port map( G => load_op, D => N47, Q => 
                           data_out(11));
   data_out_reg_10_inst : DLH_X1 port map( G => load_op, D => N46, Q => 
                           data_out(10));
   data_out_reg_9_inst : DLH_X1 port map( G => load_op, D => N45, Q => 
                           data_out(9));
   data_out_reg_8_inst : DLH_X1 port map( G => load_op, D => N44, Q => 
                           data_out(8));
   data_out_reg_7_inst : DLH_X1 port map( G => load_op, D => N43, Q => 
                           data_out(7));
   data_out_reg_6_inst : DLH_X1 port map( G => load_op, D => N42, Q => 
                           data_out(6));
   data_out_reg_5_inst : DLH_X1 port map( G => load_op, D => N41, Q => 
                           data_out(5));
   data_out_reg_4_inst : DLH_X1 port map( G => load_op, D => N40, Q => 
                           data_out(4));
   data_out_reg_3_inst : DLH_X1 port map( G => load_op, D => N39, Q => 
                           data_out(3));
   data_out_reg_2_inst : DLH_X1 port map( G => load_op, D => N38, Q => 
                           data_out(2));
   data_out_reg_1_inst : DLH_X1 port map( G => load_op, D => N37, Q => 
                           data_out(1));
   data_out_reg_0_inst : DLH_X1 port map( G => load_op, D => N36, Q => 
                           data_out(0));
   U2 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => N67);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N66);
   U4 : NAND2_X1 port map( A1 => data_in(30), A2 => n5, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n3, A2 => n6, ZN => N65);
   U6 : NAND2_X1 port map( A1 => data_in(29), A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n3, A2 => n7, ZN => N64);
   U8 : NAND2_X1 port map( A1 => data_in(28), A2 => n5, ZN => n7);
   U9 : NAND2_X1 port map( A1 => n3, A2 => n8, ZN => N63);
   U10 : NAND2_X1 port map( A1 => data_in(27), A2 => n5, ZN => n8);
   U11 : NAND2_X1 port map( A1 => n3, A2 => n9, ZN => N62);
   U12 : NAND2_X1 port map( A1 => data_in(26), A2 => n5, ZN => n9);
   U13 : NAND2_X1 port map( A1 => n3, A2 => n10, ZN => N61);
   U14 : NAND2_X1 port map( A1 => data_in(25), A2 => n5, ZN => n10);
   U15 : NAND2_X1 port map( A1 => n3, A2 => n11, ZN => N60);
   U16 : NAND2_X1 port map( A1 => data_in(24), A2 => n5, ZN => n11);
   U17 : NAND2_X1 port map( A1 => n3, A2 => n12, ZN => N59);
   U18 : NAND2_X1 port map( A1 => data_in(23), A2 => n5, ZN => n12);
   U19 : NAND2_X1 port map( A1 => n3, A2 => n13, ZN => N58);
   U20 : NAND2_X1 port map( A1 => data_in(22), A2 => n5, ZN => n13);
   U21 : NAND2_X1 port map( A1 => n3, A2 => n14, ZN => N57);
   U22 : NAND2_X1 port map( A1 => data_in(21), A2 => n5, ZN => n14);
   U23 : NAND2_X1 port map( A1 => n3, A2 => n15, ZN => N56);
   U24 : NAND2_X1 port map( A1 => data_in(20), A2 => n5, ZN => n15);
   U25 : NAND2_X1 port map( A1 => n3, A2 => n16, ZN => N55);
   U26 : NAND2_X1 port map( A1 => data_in(19), A2 => n5, ZN => n16);
   U27 : NAND2_X1 port map( A1 => n3, A2 => n17, ZN => N54);
   U28 : NAND2_X1 port map( A1 => data_in(18), A2 => n5, ZN => n17);
   U29 : NAND2_X1 port map( A1 => n3, A2 => n18, ZN => N53);
   U30 : NAND2_X1 port map( A1 => data_in(17), A2 => n5, ZN => n18);
   U31 : NAND2_X1 port map( A1 => n3, A2 => n19, ZN => N52);
   U32 : NAND2_X1 port map( A1 => data_in(16), A2 => n5, ZN => n19);
   U33 : INV_X1 port map( A => n1, ZN => n5);
   U34 : NAND2_X1 port map( A1 => load_type(1), A2 => load_type(0), ZN => n1);
   U35 : NAND2_X1 port map( A1 => n3, A2 => n20, ZN => N51);
   U36 : NAND2_X1 port map( A1 => data_in(15), A2 => load_type(0), ZN => n20);
   U37 : NAND2_X1 port map( A1 => n3, A2 => n21, ZN => N50);
   U38 : NAND2_X1 port map( A1 => data_in(14), A2 => load_type(0), ZN => n21);
   U39 : NAND2_X1 port map( A1 => n3, A2 => n22, ZN => N49);
   U40 : NAND2_X1 port map( A1 => data_in(13), A2 => load_type(0), ZN => n22);
   U41 : NAND2_X1 port map( A1 => n3, A2 => n23, ZN => N48);
   U42 : NAND2_X1 port map( A1 => data_in(12), A2 => load_type(0), ZN => n23);
   U43 : NAND2_X1 port map( A1 => n3, A2 => n24, ZN => N47);
   U44 : NAND2_X1 port map( A1 => data_in(11), A2 => load_type(0), ZN => n24);
   U45 : NAND2_X1 port map( A1 => n3, A2 => n25, ZN => N46);
   U46 : NAND2_X1 port map( A1 => data_in(10), A2 => load_type(0), ZN => n25);
   U47 : NAND2_X1 port map( A1 => n3, A2 => n26, ZN => N45);
   U48 : NAND2_X1 port map( A1 => data_in(9), A2 => load_type(0), ZN => n26);
   U49 : NAND2_X1 port map( A1 => n3, A2 => n27, ZN => N44);
   U50 : NAND2_X1 port map( A1 => data_in(8), A2 => load_type(0), ZN => n27);
   U51 : OR3_X1 port map( A1 => signed_val, A2 => n2, A3 => n28, ZN => n3);
   U52 : INV_X1 port map( A => data_in(31), ZN => n2);
   U53 : AND2_X1 port map( A1 => data_in(7), A2 => n29, ZN => N43);
   U54 : AND2_X1 port map( A1 => data_in(6), A2 => n29, ZN => N42);
   U55 : AND2_X1 port map( A1 => data_in(5), A2 => n29, ZN => N41);
   U56 : AND2_X1 port map( A1 => data_in(4), A2 => n29, ZN => N40);
   U57 : AND2_X1 port map( A1 => data_in(3), A2 => n29, ZN => N39);
   U58 : AND2_X1 port map( A1 => data_in(2), A2 => n29, ZN => N38);
   U59 : AND2_X1 port map( A1 => data_in(1), A2 => n29, ZN => N37);
   U60 : AND2_X1 port map( A1 => data_in(0), A2 => n29, ZN => N36);
   U61 : NAND2_X1 port map( A1 => n30, A2 => n28, ZN => n29);
   U62 : OR2_X1 port map( A1 => load_type(1), A2 => load_type(0), ZN => n28);
   U63 : INV_X1 port map( A => load_type(0), ZN => n30);

end SYN_bhv_load;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity COND_BT_NBIT32 is

   port( ZERO_BIT, OPCODE_0, branch_op : in std_logic;  con_sign : out 
         std_logic);

end COND_BT_NBIT32;

architecture SYN_BHV of COND_BT_NBIT32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => branch_op, A2 => n1, ZN => con_sign);
   U3 : XOR2_X1 port map( A => ZERO_BIT, B => OPCODE_0, Z => n1);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity zero_eval_NBIT32 is

   port( input : in std_logic_vector (31 downto 0);  res : out std_logic);

end zero_eval_NBIT32;

architecture SYN_bhv of zero_eval_NBIT32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => res);
   U2 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => n2);
   U3 : NOR4_X1 port map( A1 => input(23), A2 => input(22), A3 => input(21), A4
                           => input(20), ZN => n6);
   U4 : NOR4_X1 port map( A1 => input(1), A2 => input(19), A3 => input(18), A4 
                           => input(17), ZN => n5);
   U5 : NOR4_X1 port map( A1 => input(16), A2 => input(15), A3 => input(14), A4
                           => input(13), ZN => n4);
   U6 : NOR4_X1 port map( A1 => input(12), A2 => input(11), A3 => input(10), A4
                           => input(0), ZN => n3);
   U7 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => n9, A4 => n10, ZN => n1);
   U8 : NOR4_X1 port map( A1 => input(9), A2 => input(8), A3 => input(7), A4 =>
                           input(6), ZN => n10);
   U9 : NOR4_X1 port map( A1 => input(5), A2 => input(4), A3 => input(3), A4 =>
                           input(31), ZN => n9);
   U10 : NOR4_X1 port map( A1 => input(30), A2 => input(2), A3 => input(29), A4
                           => input(28), ZN => n8);
   U11 : NOR4_X1 port map( A1 => input(27), A2 => input(26), A3 => input(25), 
                           A4 => input(24), ZN => n7);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ALU_N32 is

   port( CLK : in std_logic;  FUNC : in std_logic_vector (0 to 5);  DATA1, 
         DATA2 : in std_logic_vector (31 downto 0);  OUT_ALU : out 
         std_logic_vector (31 downto 0));

end ALU_N32;

architecture SYN_Architectural of ALU_N32 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component P4_ADDER_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component SHIFTER_GENERIC_N32
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
            downto 0);  LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE : in std_logic;  
            OUTPUT : out std_logic_vector (31 downto 0));
   end component;
   
   component comparator
      port( DATA1 : in std_logic_vector (31 downto 0);  DATA2i : in std_logic; 
            tipo : in std_logic_vector (0 to 5);  OUTALU : out std_logic_vector
            (31 downto 0));
   end component;
   
   component logic_N32
      port( FUNC : in std_logic_vector (0 to 5);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUT_ALU : out std_logic_vector (31
            downto 0));
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal OUTPUT_alu_i_31_port, OUTPUT_alu_i_30_port, OUTPUT_alu_i_29_port, 
      OUTPUT_alu_i_28_port, OUTPUT_alu_i_27_port, OUTPUT_alu_i_26_port, 
      OUTPUT_alu_i_25_port, OUTPUT_alu_i_24_port, OUTPUT_alu_i_23_port, 
      OUTPUT_alu_i_22_port, OUTPUT_alu_i_21_port, OUTPUT_alu_i_20_port, 
      OUTPUT_alu_i_19_port, OUTPUT_alu_i_18_port, OUTPUT_alu_i_17_port, 
      OUTPUT_alu_i_16_port, OUTPUT_alu_i_15_port, OUTPUT_alu_i_14_port, 
      OUTPUT_alu_i_13_port, OUTPUT_alu_i_12_port, OUTPUT_alu_i_11_port, 
      OUTPUT_alu_i_10_port, OUTPUT_alu_i_9_port, OUTPUT_alu_i_8_port, 
      OUTPUT_alu_i_7_port, OUTPUT_alu_i_6_port, OUTPUT_alu_i_5_port, 
      OUTPUT_alu_i_4_port, OUTPUT_alu_i_3_port, OUTPUT_alu_i_2_port, 
      OUTPUT_alu_i_1_port, OUTPUT_alu_i_0_port, OUTPUT4_31_port, 
      OUTPUT4_30_port, OUTPUT4_29_port, OUTPUT4_28_port, OUTPUT4_27_port, 
      OUTPUT4_26_port, OUTPUT4_25_port, OUTPUT4_24_port, OUTPUT4_23_port, 
      OUTPUT4_22_port, OUTPUT4_21_port, OUTPUT4_20_port, OUTPUT4_19_port, 
      OUTPUT4_18_port, OUTPUT4_17_port, OUTPUT4_16_port, OUTPUT4_15_port, 
      OUTPUT4_14_port, OUTPUT4_13_port, OUTPUT4_12_port, OUTPUT4_11_port, 
      OUTPUT4_10_port, OUTPUT4_9_port, OUTPUT4_8_port, OUTPUT4_7_port, 
      OUTPUT4_6_port, OUTPUT4_5_port, OUTPUT4_4_port, OUTPUT4_3_port, 
      OUTPUT4_2_port, OUTPUT4_1_port, OUTPUT4_0_port, OUTPUT2_31_port, 
      OUTPUT2_30_port, OUTPUT2_29_port, OUTPUT2_28_port, OUTPUT2_27_port, 
      OUTPUT2_26_port, OUTPUT2_25_port, OUTPUT2_24_port, OUTPUT2_23_port, 
      OUTPUT2_22_port, OUTPUT2_21_port, OUTPUT2_20_port, OUTPUT2_19_port, 
      OUTPUT2_18_port, OUTPUT2_17_port, OUTPUT2_16_port, OUTPUT2_15_port, 
      OUTPUT2_14_port, OUTPUT2_13_port, OUTPUT2_12_port, OUTPUT2_11_port, 
      OUTPUT2_10_port, OUTPUT2_9_port, OUTPUT2_8_port, OUTPUT2_7_port, 
      OUTPUT2_6_port, OUTPUT2_5_port, OUTPUT2_4_port, OUTPUT2_3_port, 
      OUTPUT2_2_port, OUTPUT2_1_port, OUTPUT2_0_port, Cout_i, OUTPUT3_0_port, 
      LOGIC_ARITH_i, LEFT_RIGHT_i, SHIFT_ROTATE_i, OUTPUT1_31_port, 
      OUTPUT1_30_port, OUTPUT1_29_port, OUTPUT1_28_port, OUTPUT1_27_port, 
      OUTPUT1_26_port, OUTPUT1_25_port, OUTPUT1_24_port, OUTPUT1_23_port, 
      OUTPUT1_22_port, OUTPUT1_21_port, OUTPUT1_20_port, OUTPUT1_19_port, 
      OUTPUT1_18_port, OUTPUT1_17_port, OUTPUT1_16_port, OUTPUT1_15_port, 
      OUTPUT1_14_port, OUTPUT1_13_port, OUTPUT1_12_port, OUTPUT1_11_port, 
      OUTPUT1_10_port, OUTPUT1_9_port, OUTPUT1_8_port, OUTPUT1_7_port, 
      OUTPUT1_6_port, OUTPUT1_5_port, OUTPUT1_4_port, OUTPUT1_3_port, 
      OUTPUT1_2_port, OUTPUT1_1_port, OUTPUT1_0_port, data1i_31_port, 
      data1i_30_port, data1i_29_port, data1i_28_port, data1i_27_port, 
      data1i_26_port, data1i_25_port, data1i_24_port, data1i_23_port, 
      data1i_22_port, data1i_21_port, data1i_20_port, data1i_19_port, 
      data1i_18_port, data1i_17_port, data1i_16_port, data1i_15_port, 
      data1i_14_port, data1i_13_port, data1i_12_port, data1i_11_port, 
      data1i_10_port, data1i_9_port, data1i_8_port, data1i_7_port, 
      data1i_6_port, data1i_5_port, data1i_4_port, data1i_3_port, data1i_2_port
      , data1i_1_port, data1i_0_port, data2i_31_port, data2i_30_port, 
      data2i_29_port, data2i_28_port, data2i_27_port, data2i_26_port, 
      data2i_25_port, data2i_24_port, data2i_23_port, data2i_22_port, 
      data2i_21_port, data2i_20_port, data2i_19_port, data2i_18_port, 
      data2i_17_port, data2i_16_port, data2i_15_port, data2i_14_port, 
      data2i_13_port, data2i_12_port, data2i_11_port, data2i_10_port, 
      data2i_9_port, data2i_8_port, data2i_7_port, data2i_6_port, data2i_5_port
      , data2i_4_port, data2i_3_port, data2i_2_port, data2i_1_port, 
      data2i_0_port, Cin_i, N139, N140, N141, N142, N143, N144, N145, N146, 
      N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, 
      N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, 
      N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, 
      N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, 
      N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, 
      N207, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
      n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102
      , n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139_port, n140_port, n141_port, n142_port, n143_port, n144_port, 
      n145_port, n146_port, n147_port, n148_port, n149_port, n150_port, 
      n151_port, n152_port, n153_port, n154_port, n155_port, n156_port, 
      n157_port, n158_port, n159_port, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139 : std_logic;

begin
   
   Cin_i_reg : DLH_X1 port map( G => n155_port, D => N140, Q => Cin_i);
   data2i_reg_31_inst : DLH_X1 port map( G => n155_port, D => N205, Q => 
                           data2i_31_port);
   data2i_reg_30_inst : DLH_X1 port map( G => n155_port, D => N204, Q => 
                           data2i_30_port);
   data2i_reg_29_inst : DLH_X1 port map( G => n155_port, D => N203, Q => 
                           data2i_29_port);
   data2i_reg_28_inst : DLH_X1 port map( G => n155_port, D => N202, Q => 
                           data2i_28_port);
   data2i_reg_27_inst : DLH_X1 port map( G => n155_port, D => N201, Q => 
                           data2i_27_port);
   data2i_reg_26_inst : DLH_X1 port map( G => n155_port, D => N200, Q => 
                           data2i_26_port);
   data2i_reg_25_inst : DLH_X1 port map( G => n155_port, D => N199, Q => 
                           data2i_25_port);
   data2i_reg_24_inst : DLH_X1 port map( G => n155_port, D => N198, Q => 
                           data2i_24_port);
   data2i_reg_23_inst : DLH_X1 port map( G => n155_port, D => N197, Q => 
                           data2i_23_port);
   data2i_reg_22_inst : DLH_X1 port map( G => n155_port, D => N196, Q => 
                           data2i_22_port);
   data2i_reg_21_inst : DLH_X1 port map( G => n155_port, D => N195, Q => 
                           data2i_21_port);
   data2i_reg_20_inst : DLH_X1 port map( G => n155_port, D => N194, Q => 
                           data2i_20_port);
   data2i_reg_19_inst : DLH_X1 port map( G => n155_port, D => N193, Q => 
                           data2i_19_port);
   data2i_reg_18_inst : DLH_X1 port map( G => n155_port, D => N192, Q => 
                           data2i_18_port);
   data2i_reg_17_inst : DLH_X1 port map( G => n155_port, D => N191, Q => 
                           data2i_17_port);
   data2i_reg_16_inst : DLH_X1 port map( G => n155_port, D => N190, Q => 
                           data2i_16_port);
   data2i_reg_15_inst : DLH_X1 port map( G => n155_port, D => N189, Q => 
                           data2i_15_port);
   data2i_reg_14_inst : DLH_X1 port map( G => n155_port, D => N188, Q => 
                           data2i_14_port);
   data2i_reg_13_inst : DLH_X1 port map( G => n155_port, D => N187, Q => 
                           data2i_13_port);
   data2i_reg_12_inst : DLH_X1 port map( G => n155_port, D => N186, Q => 
                           data2i_12_port);
   data2i_reg_11_inst : DLH_X1 port map( G => n155_port, D => N185, Q => 
                           data2i_11_port);
   data2i_reg_10_inst : DLH_X1 port map( G => n155_port, D => N184, Q => 
                           data2i_10_port);
   data2i_reg_9_inst : DLH_X1 port map( G => n155_port, D => N183, Q => 
                           data2i_9_port);
   data2i_reg_8_inst : DLH_X1 port map( G => n155_port, D => N182, Q => 
                           data2i_8_port);
   data2i_reg_7_inst : DLH_X1 port map( G => n155_port, D => N181, Q => 
                           data2i_7_port);
   data2i_reg_6_inst : DLH_X1 port map( G => n155_port, D => N180, Q => 
                           data2i_6_port);
   data2i_reg_5_inst : DLH_X1 port map( G => n155_port, D => N179, Q => 
                           data2i_5_port);
   data2i_reg_4_inst : DLH_X1 port map( G => n155_port, D => N178, Q => 
                           data2i_4_port);
   data2i_reg_3_inst : DLH_X1 port map( G => n155_port, D => N177, Q => 
                           data2i_3_port);
   data2i_reg_2_inst : DLH_X1 port map( G => n155_port, D => N176, Q => 
                           data2i_2_port);
   data2i_reg_1_inst : DLH_X1 port map( G => n155_port, D => N175, Q => 
                           data2i_1_port);
   data2i_reg_0_inst : DLH_X1 port map( G => n155_port, D => N174, Q => 
                           data2i_0_port);
   data1i_reg_31_inst : DLH_X1 port map( G => n155_port, D => DATA1(31), Q => 
                           data1i_31_port);
   data1i_reg_30_inst : DLH_X1 port map( G => n155_port, D => DATA1(30), Q => 
                           data1i_30_port);
   data1i_reg_29_inst : DLH_X1 port map( G => n155_port, D => DATA1(29), Q => 
                           data1i_29_port);
   data1i_reg_28_inst : DLH_X1 port map( G => n155_port, D => DATA1(28), Q => 
                           data1i_28_port);
   data1i_reg_27_inst : DLH_X1 port map( G => n155_port, D => DATA1(27), Q => 
                           data1i_27_port);
   data1i_reg_26_inst : DLH_X1 port map( G => n155_port, D => DATA1(26), Q => 
                           data1i_26_port);
   data1i_reg_25_inst : DLH_X1 port map( G => n155_port, D => DATA1(25), Q => 
                           data1i_25_port);
   data1i_reg_24_inst : DLH_X1 port map( G => n155_port, D => DATA1(24), Q => 
                           data1i_24_port);
   data1i_reg_23_inst : DLH_X1 port map( G => n155_port, D => DATA1(23), Q => 
                           data1i_23_port);
   data1i_reg_22_inst : DLH_X1 port map( G => n155_port, D => DATA1(22), Q => 
                           data1i_22_port);
   data1i_reg_21_inst : DLH_X1 port map( G => n155_port, D => DATA1(21), Q => 
                           data1i_21_port);
   data1i_reg_20_inst : DLH_X1 port map( G => n155_port, D => DATA1(20), Q => 
                           data1i_20_port);
   data1i_reg_19_inst : DLH_X1 port map( G => n155_port, D => DATA1(19), Q => 
                           data1i_19_port);
   data1i_reg_18_inst : DLH_X1 port map( G => n155_port, D => DATA1(18), Q => 
                           data1i_18_port);
   data1i_reg_17_inst : DLH_X1 port map( G => n155_port, D => DATA1(17), Q => 
                           data1i_17_port);
   data1i_reg_16_inst : DLH_X1 port map( G => n155_port, D => DATA1(16), Q => 
                           data1i_16_port);
   data1i_reg_15_inst : DLH_X1 port map( G => n155_port, D => DATA1(15), Q => 
                           data1i_15_port);
   data1i_reg_14_inst : DLH_X1 port map( G => n155_port, D => DATA1(14), Q => 
                           data1i_14_port);
   data1i_reg_13_inst : DLH_X1 port map( G => n155_port, D => DATA1(13), Q => 
                           data1i_13_port);
   data1i_reg_12_inst : DLH_X1 port map( G => n155_port, D => DATA1(12), Q => 
                           data1i_12_port);
   data1i_reg_11_inst : DLH_X1 port map( G => n155_port, D => DATA1(11), Q => 
                           data1i_11_port);
   data1i_reg_10_inst : DLH_X1 port map( G => n155_port, D => DATA1(10), Q => 
                           data1i_10_port);
   data1i_reg_9_inst : DLH_X1 port map( G => n155_port, D => DATA1(9), Q => 
                           data1i_9_port);
   data1i_reg_8_inst : DLH_X1 port map( G => n155_port, D => DATA1(8), Q => 
                           data1i_8_port);
   data1i_reg_7_inst : DLH_X1 port map( G => n155_port, D => DATA1(7), Q => 
                           data1i_7_port);
   data1i_reg_6_inst : DLH_X1 port map( G => n155_port, D => DATA1(6), Q => 
                           data1i_6_port);
   data1i_reg_5_inst : DLH_X1 port map( G => n155_port, D => DATA1(5), Q => 
                           data1i_5_port);
   data1i_reg_4_inst : DLH_X1 port map( G => n155_port, D => DATA1(4), Q => 
                           data1i_4_port);
   data1i_reg_3_inst : DLH_X1 port map( G => n155_port, D => DATA1(3), Q => 
                           data1i_3_port);
   data1i_reg_2_inst : DLH_X1 port map( G => n155_port, D => DATA1(2), Q => 
                           data1i_2_port);
   data1i_reg_1_inst : DLH_X1 port map( G => n155_port, D => DATA1(1), Q => 
                           data1i_1_port);
   data1i_reg_0_inst : DLH_X1 port map( G => n155_port, D => DATA1(0), Q => 
                           data1i_0_port);
   LOGIC_ARITH_i_reg : DLH_X1 port map( G => n159_port, D => N207, Q => 
                           LOGIC_ARITH_i);
   LEFT_RIGHT_i_reg : DLH_X1 port map( G => n159_port, D => N207, Q => 
                           LEFT_RIGHT_i);
   OUTPUT_alu_i_reg_0_inst : DLH_X1 port map( G => N141, D => N142, Q => 
                           OUTPUT_alu_i_0_port);
   OUT_ALU_reg_0_inst : DFF_X1 port map( D => OUTPUT_alu_i_0_port, CK => CLK, Q
                           => OUT_ALU(0), QN => n_1077);
   OUTPUT_alu_i_reg_1_inst : DLH_X1 port map( G => N141, D => N143, Q => 
                           OUTPUT_alu_i_1_port);
   OUT_ALU_reg_1_inst : DFF_X1 port map( D => OUTPUT_alu_i_1_port, CK => CLK, Q
                           => OUT_ALU(1), QN => n_1078);
   OUTPUT_alu_i_reg_2_inst : DLH_X1 port map( G => N141, D => N144, Q => 
                           OUTPUT_alu_i_2_port);
   OUT_ALU_reg_2_inst : DFF_X1 port map( D => OUTPUT_alu_i_2_port, CK => CLK, Q
                           => OUT_ALU(2), QN => n_1079);
   OUTPUT_alu_i_reg_3_inst : DLH_X1 port map( G => N141, D => N145, Q => 
                           OUTPUT_alu_i_3_port);
   OUT_ALU_reg_3_inst : DFF_X1 port map( D => OUTPUT_alu_i_3_port, CK => CLK, Q
                           => OUT_ALU(3), QN => n_1080);
   OUTPUT_alu_i_reg_4_inst : DLH_X1 port map( G => N141, D => N146, Q => 
                           OUTPUT_alu_i_4_port);
   OUT_ALU_reg_4_inst : DFF_X1 port map( D => OUTPUT_alu_i_4_port, CK => CLK, Q
                           => OUT_ALU(4), QN => n_1081);
   OUTPUT_alu_i_reg_5_inst : DLH_X1 port map( G => N141, D => N147, Q => 
                           OUTPUT_alu_i_5_port);
   OUT_ALU_reg_5_inst : DFF_X1 port map( D => OUTPUT_alu_i_5_port, CK => CLK, Q
                           => OUT_ALU(5), QN => n_1082);
   OUTPUT_alu_i_reg_6_inst : DLH_X1 port map( G => N141, D => N148, Q => 
                           OUTPUT_alu_i_6_port);
   OUT_ALU_reg_6_inst : DFF_X1 port map( D => OUTPUT_alu_i_6_port, CK => CLK, Q
                           => OUT_ALU(6), QN => n_1083);
   OUTPUT_alu_i_reg_7_inst : DLH_X1 port map( G => N141, D => N149, Q => 
                           OUTPUT_alu_i_7_port);
   OUT_ALU_reg_7_inst : DFF_X1 port map( D => OUTPUT_alu_i_7_port, CK => CLK, Q
                           => OUT_ALU(7), QN => n_1084);
   OUTPUT_alu_i_reg_8_inst : DLH_X1 port map( G => N141, D => N150, Q => 
                           OUTPUT_alu_i_8_port);
   OUT_ALU_reg_8_inst : DFF_X1 port map( D => OUTPUT_alu_i_8_port, CK => CLK, Q
                           => OUT_ALU(8), QN => n_1085);
   OUTPUT_alu_i_reg_9_inst : DLH_X1 port map( G => N141, D => N151, Q => 
                           OUTPUT_alu_i_9_port);
   OUT_ALU_reg_9_inst : DFF_X1 port map( D => OUTPUT_alu_i_9_port, CK => CLK, Q
                           => OUT_ALU(9), QN => n_1086);
   OUTPUT_alu_i_reg_10_inst : DLH_X1 port map( G => N141, D => N152, Q => 
                           OUTPUT_alu_i_10_port);
   OUT_ALU_reg_10_inst : DFF_X1 port map( D => OUTPUT_alu_i_10_port, CK => CLK,
                           Q => OUT_ALU(10), QN => n_1087);
   OUTPUT_alu_i_reg_11_inst : DLH_X1 port map( G => N141, D => N153, Q => 
                           OUTPUT_alu_i_11_port);
   OUT_ALU_reg_11_inst : DFF_X1 port map( D => OUTPUT_alu_i_11_port, CK => CLK,
                           Q => OUT_ALU(11), QN => n_1088);
   OUTPUT_alu_i_reg_12_inst : DLH_X1 port map( G => N141, D => N154, Q => 
                           OUTPUT_alu_i_12_port);
   OUT_ALU_reg_12_inst : DFF_X1 port map( D => OUTPUT_alu_i_12_port, CK => CLK,
                           Q => OUT_ALU(12), QN => n_1089);
   OUTPUT_alu_i_reg_13_inst : DLH_X1 port map( G => N141, D => N155, Q => 
                           OUTPUT_alu_i_13_port);
   OUT_ALU_reg_13_inst : DFF_X1 port map( D => OUTPUT_alu_i_13_port, CK => CLK,
                           Q => OUT_ALU(13), QN => n_1090);
   OUTPUT_alu_i_reg_14_inst : DLH_X1 port map( G => N141, D => N156, Q => 
                           OUTPUT_alu_i_14_port);
   OUT_ALU_reg_14_inst : DFF_X1 port map( D => OUTPUT_alu_i_14_port, CK => CLK,
                           Q => OUT_ALU(14), QN => n_1091);
   OUTPUT_alu_i_reg_15_inst : DLH_X1 port map( G => N141, D => N157, Q => 
                           OUTPUT_alu_i_15_port);
   OUT_ALU_reg_15_inst : DFF_X1 port map( D => OUTPUT_alu_i_15_port, CK => CLK,
                           Q => OUT_ALU(15), QN => n_1092);
   OUTPUT_alu_i_reg_16_inst : DLH_X1 port map( G => N141, D => N158, Q => 
                           OUTPUT_alu_i_16_port);
   OUT_ALU_reg_16_inst : DFF_X1 port map( D => OUTPUT_alu_i_16_port, CK => CLK,
                           Q => OUT_ALU(16), QN => n_1093);
   OUTPUT_alu_i_reg_17_inst : DLH_X1 port map( G => N141, D => N159, Q => 
                           OUTPUT_alu_i_17_port);
   OUT_ALU_reg_17_inst : DFF_X1 port map( D => OUTPUT_alu_i_17_port, CK => CLK,
                           Q => OUT_ALU(17), QN => n_1094);
   OUTPUT_alu_i_reg_18_inst : DLH_X1 port map( G => N141, D => N160, Q => 
                           OUTPUT_alu_i_18_port);
   OUT_ALU_reg_18_inst : DFF_X1 port map( D => OUTPUT_alu_i_18_port, CK => CLK,
                           Q => OUT_ALU(18), QN => n_1095);
   OUTPUT_alu_i_reg_19_inst : DLH_X1 port map( G => N141, D => N161, Q => 
                           OUTPUT_alu_i_19_port);
   OUT_ALU_reg_19_inst : DFF_X1 port map( D => OUTPUT_alu_i_19_port, CK => CLK,
                           Q => OUT_ALU(19), QN => n_1096);
   OUTPUT_alu_i_reg_20_inst : DLH_X1 port map( G => N141, D => N162, Q => 
                           OUTPUT_alu_i_20_port);
   OUT_ALU_reg_20_inst : DFF_X1 port map( D => OUTPUT_alu_i_20_port, CK => CLK,
                           Q => OUT_ALU(20), QN => n_1097);
   OUTPUT_alu_i_reg_21_inst : DLH_X1 port map( G => N141, D => N163, Q => 
                           OUTPUT_alu_i_21_port);
   OUT_ALU_reg_21_inst : DFF_X1 port map( D => OUTPUT_alu_i_21_port, CK => CLK,
                           Q => OUT_ALU(21), QN => n_1098);
   OUTPUT_alu_i_reg_22_inst : DLH_X1 port map( G => N141, D => N164, Q => 
                           OUTPUT_alu_i_22_port);
   OUT_ALU_reg_22_inst : DFF_X1 port map( D => OUTPUT_alu_i_22_port, CK => CLK,
                           Q => OUT_ALU(22), QN => n_1099);
   OUTPUT_alu_i_reg_23_inst : DLH_X1 port map( G => N141, D => N165, Q => 
                           OUTPUT_alu_i_23_port);
   OUT_ALU_reg_23_inst : DFF_X1 port map( D => OUTPUT_alu_i_23_port, CK => CLK,
                           Q => OUT_ALU(23), QN => n_1100);
   OUTPUT_alu_i_reg_24_inst : DLH_X1 port map( G => N141, D => N166, Q => 
                           OUTPUT_alu_i_24_port);
   OUT_ALU_reg_24_inst : DFF_X1 port map( D => OUTPUT_alu_i_24_port, CK => CLK,
                           Q => OUT_ALU(24), QN => n_1101);
   OUTPUT_alu_i_reg_25_inst : DLH_X1 port map( G => N141, D => N167, Q => 
                           OUTPUT_alu_i_25_port);
   OUT_ALU_reg_25_inst : DFF_X1 port map( D => OUTPUT_alu_i_25_port, CK => CLK,
                           Q => OUT_ALU(25), QN => n_1102);
   OUTPUT_alu_i_reg_26_inst : DLH_X1 port map( G => N141, D => N168, Q => 
                           OUTPUT_alu_i_26_port);
   OUT_ALU_reg_26_inst : DFF_X1 port map( D => OUTPUT_alu_i_26_port, CK => CLK,
                           Q => OUT_ALU(26), QN => n_1103);
   OUTPUT_alu_i_reg_27_inst : DLH_X1 port map( G => N141, D => N169, Q => 
                           OUTPUT_alu_i_27_port);
   OUT_ALU_reg_27_inst : DFF_X1 port map( D => OUTPUT_alu_i_27_port, CK => CLK,
                           Q => OUT_ALU(27), QN => n_1104);
   OUTPUT_alu_i_reg_28_inst : DLH_X1 port map( G => N141, D => N170, Q => 
                           OUTPUT_alu_i_28_port);
   OUT_ALU_reg_28_inst : DFF_X1 port map( D => OUTPUT_alu_i_28_port, CK => CLK,
                           Q => OUT_ALU(28), QN => n_1105);
   OUTPUT_alu_i_reg_29_inst : DLH_X1 port map( G => N141, D => N171, Q => 
                           OUTPUT_alu_i_29_port);
   OUT_ALU_reg_29_inst : DFF_X1 port map( D => OUTPUT_alu_i_29_port, CK => CLK,
                           Q => OUT_ALU(29), QN => n_1106);
   OUTPUT_alu_i_reg_30_inst : DLH_X1 port map( G => N141, D => N172, Q => 
                           OUTPUT_alu_i_30_port);
   OUT_ALU_reg_30_inst : DFF_X1 port map( D => OUTPUT_alu_i_30_port, CK => CLK,
                           Q => OUT_ALU(30), QN => n_1107);
   OUTPUT_alu_i_reg_31_inst : DLH_X1 port map( G => N141, D => N173, Q => 
                           OUTPUT_alu_i_31_port);
   OUT_ALU_reg_31_inst : DFF_X1 port map( D => OUTPUT_alu_i_31_port, CK => CLK,
                           Q => OUT_ALU(31), QN => n_1108);
   SHIFT_ROTATE_i <= '1';
   U4 : INV_X1 port map( A => n1, ZN => N207);
   U5 : OAI22_X1 port map( A1 => DATA2(31), A2 => n157_port, B1 => n3, B2 => n4
                           , ZN => N205);
   U6 : INV_X1 port map( A => DATA2(31), ZN => n4);
   U7 : OAI22_X1 port map( A1 => DATA2(30), A2 => n157_port, B1 => n3, B2 => n5
                           , ZN => N204);
   U8 : INV_X1 port map( A => DATA2(30), ZN => n5);
   U9 : OAI22_X1 port map( A1 => DATA2(29), A2 => n157_port, B1 => n3, B2 => n6
                           , ZN => N203);
   U10 : INV_X1 port map( A => DATA2(29), ZN => n6);
   U11 : OAI22_X1 port map( A1 => DATA2(28), A2 => n157_port, B1 => n3, B2 => 
                           n7, ZN => N202);
   U12 : INV_X1 port map( A => DATA2(28), ZN => n7);
   U13 : OAI22_X1 port map( A1 => DATA2(27), A2 => n157_port, B1 => n3, B2 => 
                           n8, ZN => N201);
   U14 : INV_X1 port map( A => DATA2(27), ZN => n8);
   U15 : OAI22_X1 port map( A1 => DATA2(26), A2 => n157_port, B1 => n3, B2 => 
                           n9, ZN => N200);
   U16 : INV_X1 port map( A => DATA2(26), ZN => n9);
   U17 : OAI22_X1 port map( A1 => DATA2(25), A2 => n157_port, B1 => n3, B2 => 
                           n10, ZN => N199);
   U18 : INV_X1 port map( A => DATA2(25), ZN => n10);
   U19 : OAI22_X1 port map( A1 => DATA2(24), A2 => n157_port, B1 => n3, B2 => 
                           n11, ZN => N198);
   U20 : INV_X1 port map( A => DATA2(24), ZN => n11);
   U21 : OAI22_X1 port map( A1 => DATA2(23), A2 => n157_port, B1 => n3, B2 => 
                           n12, ZN => N197);
   U22 : INV_X1 port map( A => DATA2(23), ZN => n12);
   U23 : OAI22_X1 port map( A1 => DATA2(22), A2 => n157_port, B1 => n3, B2 => 
                           n13, ZN => N196);
   U24 : INV_X1 port map( A => DATA2(22), ZN => n13);
   U25 : OAI22_X1 port map( A1 => DATA2(21), A2 => n157_port, B1 => n3, B2 => 
                           n14, ZN => N195);
   U26 : INV_X1 port map( A => DATA2(21), ZN => n14);
   U27 : OAI22_X1 port map( A1 => DATA2(20), A2 => n157_port, B1 => n3, B2 => 
                           n15, ZN => N194);
   U28 : INV_X1 port map( A => DATA2(20), ZN => n15);
   U29 : OAI22_X1 port map( A1 => DATA2(19), A2 => n157_port, B1 => n3, B2 => 
                           n16, ZN => N193);
   U30 : INV_X1 port map( A => DATA2(19), ZN => n16);
   U31 : OAI22_X1 port map( A1 => DATA2(18), A2 => n157_port, B1 => n3, B2 => 
                           n17, ZN => N192);
   U32 : INV_X1 port map( A => DATA2(18), ZN => n17);
   U33 : OAI22_X1 port map( A1 => DATA2(17), A2 => n157_port, B1 => n3, B2 => 
                           n18, ZN => N191);
   U34 : INV_X1 port map( A => DATA2(17), ZN => n18);
   U35 : OAI22_X1 port map( A1 => DATA2(16), A2 => n157_port, B1 => n3, B2 => 
                           n19, ZN => N190);
   U36 : INV_X1 port map( A => DATA2(16), ZN => n19);
   U37 : OAI22_X1 port map( A1 => DATA2(15), A2 => n157_port, B1 => n3, B2 => 
                           n20, ZN => N189);
   U38 : INV_X1 port map( A => DATA2(15), ZN => n20);
   U39 : OAI22_X1 port map( A1 => DATA2(14), A2 => n157_port, B1 => n3, B2 => 
                           n21, ZN => N188);
   U40 : INV_X1 port map( A => DATA2(14), ZN => n21);
   U41 : OAI22_X1 port map( A1 => DATA2(13), A2 => n157_port, B1 => n3, B2 => 
                           n22, ZN => N187);
   U42 : INV_X1 port map( A => DATA2(13), ZN => n22);
   U43 : OAI22_X1 port map( A1 => DATA2(12), A2 => n157_port, B1 => n3, B2 => 
                           n23, ZN => N186);
   U44 : INV_X1 port map( A => DATA2(12), ZN => n23);
   U45 : OAI22_X1 port map( A1 => DATA2(11), A2 => n157_port, B1 => n3, B2 => 
                           n24, ZN => N185);
   U46 : INV_X1 port map( A => DATA2(11), ZN => n24);
   U47 : OAI22_X1 port map( A1 => DATA2(10), A2 => n157_port, B1 => n3, B2 => 
                           n25, ZN => N184);
   U48 : INV_X1 port map( A => DATA2(10), ZN => n25);
   U49 : OAI22_X1 port map( A1 => DATA2(9), A2 => n157_port, B1 => n3, B2 => 
                           n26, ZN => N183);
   U50 : INV_X1 port map( A => DATA2(9), ZN => n26);
   U51 : OAI22_X1 port map( A1 => DATA2(8), A2 => n157_port, B1 => n3, B2 => 
                           n27, ZN => N182);
   U52 : INV_X1 port map( A => DATA2(8), ZN => n27);
   U53 : OAI22_X1 port map( A1 => DATA2(7), A2 => n157_port, B1 => n3, B2 => 
                           n28, ZN => N181);
   U54 : INV_X1 port map( A => DATA2(7), ZN => n28);
   U55 : OAI22_X1 port map( A1 => DATA2(6), A2 => n157_port, B1 => n3, B2 => 
                           n29, ZN => N180);
   U56 : INV_X1 port map( A => DATA2(6), ZN => n29);
   U57 : OAI22_X1 port map( A1 => DATA2(5), A2 => n157_port, B1 => n3, B2 => 
                           n30, ZN => N179);
   U58 : INV_X1 port map( A => DATA2(5), ZN => n30);
   U59 : OAI22_X1 port map( A1 => DATA2(4), A2 => n157_port, B1 => n3, B2 => 
                           n31, ZN => N178);
   U60 : INV_X1 port map( A => DATA2(4), ZN => n31);
   U61 : OAI22_X1 port map( A1 => DATA2(3), A2 => n157_port, B1 => n3, B2 => 
                           n32, ZN => N177);
   U62 : INV_X1 port map( A => DATA2(3), ZN => n32);
   U63 : OAI22_X1 port map( A1 => DATA2(2), A2 => n157_port, B1 => n3, B2 => 
                           n33, ZN => N176);
   U64 : INV_X1 port map( A => DATA2(2), ZN => n33);
   U65 : OAI22_X1 port map( A1 => DATA2(1), A2 => n157_port, B1 => n3, B2 => 
                           n34, ZN => N175);
   U66 : INV_X1 port map( A => DATA2(1), ZN => n34);
   U67 : OAI22_X1 port map( A1 => DATA2(0), A2 => n157_port, B1 => n3, B2 => 
                           n35, ZN => N174);
   U68 : INV_X1 port map( A => DATA2(0), ZN => n35);
   U70 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => N173);
   U71 : AOI22_X1 port map( A1 => OUTPUT2_31_port, A2 => n39, B1 => 
                           OUTPUT4_31_port, B2 => n153_port, ZN => n38);
   U73 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => N172);
   U74 : AOI22_X1 port map( A1 => OUTPUT2_30_port, A2 => n39, B1 => 
                           OUTPUT4_30_port, B2 => n153_port, ZN => n43);
   U76 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => N171);
   U77 : AOI22_X1 port map( A1 => OUTPUT2_29_port, A2 => n39, B1 => 
                           OUTPUT4_29_port, B2 => n153_port, ZN => n45);
   U79 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => N170);
   U80 : AOI22_X1 port map( A1 => OUTPUT2_28_port, A2 => n39, B1 => 
                           OUTPUT4_28_port, B2 => n153_port, ZN => n47);
   U82 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => N169);
   U83 : AOI22_X1 port map( A1 => OUTPUT2_27_port, A2 => n39, B1 => 
                           OUTPUT4_27_port, B2 => n153_port, ZN => n49);
   U85 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => N168);
   U86 : AOI22_X1 port map( A1 => OUTPUT2_26_port, A2 => n39, B1 => 
                           OUTPUT4_26_port, B2 => n153_port, ZN => n51);
   U88 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => N167);
   U89 : AOI22_X1 port map( A1 => OUTPUT2_25_port, A2 => n39, B1 => 
                           OUTPUT4_25_port, B2 => n153_port, ZN => n53);
   U91 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => N166);
   U92 : AOI22_X1 port map( A1 => OUTPUT2_24_port, A2 => n39, B1 => 
                           OUTPUT4_24_port, B2 => n153_port, ZN => n55);
   U94 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => N165);
   U95 : AOI22_X1 port map( A1 => OUTPUT2_23_port, A2 => n39, B1 => 
                           OUTPUT4_23_port, B2 => n153_port, ZN => n57);
   U97 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N164);
   U98 : AOI22_X1 port map( A1 => OUTPUT2_22_port, A2 => n39, B1 => 
                           OUTPUT4_22_port, B2 => n153_port, ZN => n59);
   U100 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N163);
   U101 : AOI22_X1 port map( A1 => OUTPUT2_21_port, A2 => n39, B1 => 
                           OUTPUT4_21_port, B2 => n153_port, ZN => n61);
   U103 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N162);
   U104 : AOI22_X1 port map( A1 => OUTPUT2_20_port, A2 => n39, B1 => 
                           OUTPUT4_20_port, B2 => n153_port, ZN => n63);
   U106 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N161);
   U107 : AOI22_X1 port map( A1 => OUTPUT2_19_port, A2 => n39, B1 => 
                           OUTPUT4_19_port, B2 => n153_port, ZN => n65);
   U109 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N160);
   U110 : AOI22_X1 port map( A1 => OUTPUT2_18_port, A2 => n39, B1 => 
                           OUTPUT4_18_port, B2 => n153_port, ZN => n67);
   U112 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N159);
   U113 : AOI22_X1 port map( A1 => OUTPUT2_17_port, A2 => n39, B1 => 
                           OUTPUT4_17_port, B2 => n153_port, ZN => n69);
   U115 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N158);
   U116 : AOI22_X1 port map( A1 => OUTPUT2_16_port, A2 => n39, B1 => 
                           OUTPUT4_16_port, B2 => n153_port, ZN => n71);
   U118 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => N157);
   U119 : AOI22_X1 port map( A1 => OUTPUT2_15_port, A2 => n39, B1 => 
                           OUTPUT4_15_port, B2 => n153_port, ZN => n73);
   U121 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => N156);
   U122 : AOI22_X1 port map( A1 => OUTPUT2_14_port, A2 => n39, B1 => 
                           OUTPUT4_14_port, B2 => n153_port, ZN => n75);
   U124 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => N155);
   U125 : AOI22_X1 port map( A1 => OUTPUT2_13_port, A2 => n39, B1 => 
                           OUTPUT4_13_port, B2 => n153_port, ZN => n77);
   U127 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => N154);
   U128 : AOI22_X1 port map( A1 => OUTPUT2_12_port, A2 => n39, B1 => 
                           OUTPUT4_12_port, B2 => n153_port, ZN => n79);
   U130 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => N153);
   U131 : AOI22_X1 port map( A1 => OUTPUT2_11_port, A2 => n39, B1 => 
                           OUTPUT4_11_port, B2 => n153_port, ZN => n81);
   U133 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => N152);
   U134 : AOI22_X1 port map( A1 => OUTPUT2_10_port, A2 => n39, B1 => 
                           OUTPUT4_10_port, B2 => n153_port, ZN => n83);
   U136 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => N151);
   U137 : AOI22_X1 port map( A1 => OUTPUT2_9_port, A2 => n39, B1 => 
                           OUTPUT4_9_port, B2 => n153_port, ZN => n85);
   U139 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => N150);
   U140 : AOI22_X1 port map( A1 => OUTPUT2_8_port, A2 => n39, B1 => 
                           OUTPUT4_8_port, B2 => n153_port, ZN => n87);
   U142 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => N149);
   U143 : AOI22_X1 port map( A1 => OUTPUT2_7_port, A2 => n39, B1 => 
                           OUTPUT4_7_port, B2 => n153_port, ZN => n89);
   U145 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => N148);
   U146 : AOI22_X1 port map( A1 => OUTPUT2_6_port, A2 => n39, B1 => 
                           OUTPUT4_6_port, B2 => n153_port, ZN => n91);
   U148 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => N147);
   U149 : AOI22_X1 port map( A1 => OUTPUT2_5_port, A2 => n39, B1 => 
                           OUTPUT4_5_port, B2 => n153_port, ZN => n93);
   U151 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => N146);
   U152 : AOI22_X1 port map( A1 => OUTPUT2_4_port, A2 => n39, B1 => 
                           OUTPUT4_4_port, B2 => n153_port, ZN => n95);
   U154 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => N145);
   U155 : AOI22_X1 port map( A1 => OUTPUT2_3_port, A2 => n39, B1 => 
                           OUTPUT4_3_port, B2 => n153_port, ZN => n97);
   U157 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => N144);
   U158 : AOI22_X1 port map( A1 => OUTPUT2_2_port, A2 => n39, B1 => 
                           OUTPUT4_2_port, B2 => n153_port, ZN => n99);
   U160 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => N143);
   U161 : AOI22_X1 port map( A1 => OUTPUT2_1_port, A2 => n39, B1 => 
                           OUTPUT4_1_port, B2 => n153_port, ZN => n101);
   U163 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => N142);
   U164 : AOI22_X1 port map( A1 => OUTPUT2_0_port, A2 => n39, B1 => 
                           OUTPUT4_0_port, B2 => n153_port, ZN => n103);
   U165 : AOI22_X1 port map( A1 => OUTPUT3_0_port, A2 => n41, B1 => 
                           OUTPUT1_0_port, B2 => n159_port, ZN => n102);
   U166 : OR3_X1 port map( A1 => n155_port, A2 => n159_port, A3 => n153_port, 
                           ZN => N141);
   U167 : OAI221_X1 port map( B1 => n104, B2 => n105, C1 => n106, C2 => n107, A
                           => n108, ZN => n40);
   U168 : INV_X1 port map( A => n109, ZN => n108);
   U169 : OAI22_X1 port map( A1 => n110, A2 => n111, B1 => n112, B2 => n113, ZN
                           => n109);
   U170 : INV_X1 port map( A => n114, ZN => n111);
   U171 : OAI211_X1 port map( C1 => n115, C2 => n116, A => n117, B => n1, ZN =>
                           N206);
   U172 : NAND2_X1 port map( A1 => n118, A2 => n119, ZN => n1);
   U173 : OAI21_X1 port map( B1 => n120, B2 => n119, A => n121, ZN => n117);
   U174 : NAND2_X1 port map( A1 => n122, A2 => n112, ZN => n119);
   U175 : NAND2_X1 port map( A1 => n123, A2 => n124, ZN => n112);
   U176 : NOR3_X1 port map( A1 => n125, A2 => FUNC(2), A3 => n126, ZN => n120);
   U177 : INV_X1 port map( A => n157_port, ZN => N140);
   U178 : NOR3_X1 port map( A1 => n127, A2 => n128, A3 => n41, ZN => n2);
   U179 : OR2_X1 port map( A1 => n39, A2 => n41, ZN => N139);
   U180 : OAI221_X1 port map( B1 => n116, B2 => n105, C1 => n106, C2 => n129, A
                           => n130, ZN => n41);
   U181 : AOI221_X1 port map( B1 => n131, B2 => n114, C1 => n132, C2 => n133, A
                           => n134, ZN => n130);
   U182 : NOR3_X1 port map( A1 => n135, A2 => n113, A3 => n136, ZN => n134);
   U183 : NAND2_X1 port map( A1 => n137, A2 => n138, ZN => n132);
   U184 : NAND2_X1 port map( A1 => n106, A2 => n139_port, ZN => n114);
   U185 : OAI211_X1 port map( C1 => n136, C2 => n126, A => n105, B => n115, ZN 
                           => n131);
   U186 : INV_X1 port map( A => n140_port, ZN => n126);
   U187 : NAND2_X1 port map( A1 => n141_port, A2 => n142_port, ZN => n105);
   U189 : OAI221_X1 port map( B1 => n113, B2 => n107, C1 => n116, C2 => n122, A
                           => n143_port, ZN => n36);
   U190 : AOI222_X1 port map( A1 => n144_port, A2 => n133, B1 => n121, B2 => 
                           n145_port, C1 => n146_port, C2 => n147_port, ZN => 
                           n143_port);
   U191 : NAND4_X1 port map( A1 => n110, A2 => n148_port, A3 => n115, A4 => 
                           n122, ZN => n147_port);
   U192 : NAND2_X1 port map( A1 => n149_port, A2 => n124, ZN => n115);
   U193 : NAND3_X1 port map( A1 => n138, A2 => n137, A3 => n148_port, ZN => 
                           n145_port);
   U194 : NAND3_X1 port map( A1 => n124, A2 => n150_port, A3 => FUNC(3), ZN => 
                           n137);
   U195 : NAND2_X1 port map( A1 => n141_port, A2 => n140_port, ZN => n138);
   U196 : INV_X1 port map( A => n106, ZN => n121);
   U197 : NAND2_X1 port map( A1 => FUNC(5), A2 => FUNC(4), ZN => n106);
   U198 : NAND2_X1 port map( A1 => n113, A2 => n139_port, ZN => n133);
   U199 : INV_X1 port map( A => n129, ZN => n144_port);
   U200 : NAND2_X1 port map( A1 => n149_port, A2 => n140_port, ZN => n129);
   U201 : NOR2_X1 port map( A1 => n135, A2 => FUNC(1), ZN => n140_port);
   U202 : NAND2_X1 port map( A1 => n142_port, A2 => n123, ZN => n122);
   U203 : INV_X1 port map( A => n136, ZN => n123);
   U204 : NAND2_X1 port map( A1 => n150_port, A2 => n125, ZN => n136);
   U205 : AND2_X1 port map( A1 => n116, A2 => n104, ZN => n113);
   U206 : INV_X1 port map( A => n146_port, ZN => n104);
   U207 : NOR2_X1 port map( A1 => FUNC(4), A2 => FUNC(5), ZN => n146_port);
   U208 : AOI21_X1 port map( B1 => n110, B2 => n148_port, A => n116, ZN => n128
                           );
   U209 : NAND2_X1 port map( A1 => FUNC(5), A2 => n151_port, ZN => n116);
   U210 : NAND3_X1 port map( A1 => n142_port, A2 => n150_port, A3 => FUNC(3), 
                           ZN => n110);
   U211 : AOI21_X1 port map( B1 => n148_port, B2 => n107, A => n139_port, ZN =>
                           n127);
   U212 : INV_X1 port map( A => n118, ZN => n139_port);
   U213 : NOR2_X1 port map( A1 => n151_port, A2 => FUNC(5), ZN => n118);
   U214 : INV_X1 port map( A => FUNC(4), ZN => n151_port);
   U215 : NAND2_X1 port map( A1 => n149_port, A2 => n142_port, ZN => n107);
   U216 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n142_port);
   U217 : NOR2_X1 port map( A1 => n150_port, A2 => n125, ZN => n149_port);
   U218 : INV_X1 port map( A => FUNC(3), ZN => n125);
   U219 : NAND2_X1 port map( A1 => n141_port, A2 => n124, ZN => n148_port);
   U220 : AND2_X1 port map( A1 => FUNC(1), A2 => n135, ZN => n124);
   U221 : INV_X1 port map( A => FUNC(0), ZN => n135);
   U222 : NOR2_X1 port map( A1 => n150_port, A2 => FUNC(3), ZN => n141_port);
   U223 : INV_X1 port map( A => FUNC(2), ZN => n150_port);
   log : logic_N32 port map( FUNC(0) => FUNC(0), FUNC(1) => FUNC(1), FUNC(2) =>
                           FUNC(2), FUNC(3) => FUNC(3), FUNC(4) => FUNC(4), 
                           FUNC(5) => FUNC(5), DATA1(31) => DATA1(31), 
                           DATA1(30) => DATA1(30), DATA1(29) => DATA1(29), 
                           DATA1(28) => DATA1(28), DATA1(27) => DATA1(27), 
                           DATA1(26) => DATA1(26), DATA1(25) => DATA1(25), 
                           DATA1(24) => DATA1(24), DATA1(23) => DATA1(23), 
                           DATA1(22) => DATA1(22), DATA1(21) => DATA1(21), 
                           DATA1(20) => DATA1(20), DATA1(19) => DATA1(19), 
                           DATA1(18) => DATA1(18), DATA1(17) => DATA1(17), 
                           DATA1(16) => DATA1(16), DATA1(15) => DATA1(15), 
                           DATA1(14) => DATA1(14), DATA1(13) => DATA1(13), 
                           DATA1(12) => DATA1(12), DATA1(11) => DATA1(11), 
                           DATA1(10) => DATA1(10), DATA1(9) => DATA1(9), 
                           DATA1(8) => DATA1(8), DATA1(7) => DATA1(7), DATA1(6)
                           => DATA1(6), DATA1(5) => DATA1(5), DATA1(4) => 
                           DATA1(4), DATA1(3) => DATA1(3), DATA1(2) => DATA1(2)
                           , DATA1(1) => DATA1(1), DATA1(0) => DATA1(0), 
                           DATA2(31) => DATA2(31), DATA2(30) => DATA2(30), 
                           DATA2(29) => DATA2(29), DATA2(28) => DATA2(28), 
                           DATA2(27) => DATA2(27), DATA2(26) => DATA2(26), 
                           DATA2(25) => DATA2(25), DATA2(24) => DATA2(24), 
                           DATA2(23) => DATA2(23), DATA2(22) => DATA2(22), 
                           DATA2(21) => DATA2(21), DATA2(20) => DATA2(20), 
                           DATA2(19) => DATA2(19), DATA2(18) => DATA2(18), 
                           DATA2(17) => DATA2(17), DATA2(16) => DATA2(16), 
                           DATA2(15) => DATA2(15), DATA2(14) => DATA2(14), 
                           DATA2(13) => DATA2(13), DATA2(12) => DATA2(12), 
                           DATA2(11) => DATA2(11), DATA2(10) => DATA2(10), 
                           DATA2(9) => DATA2(9), DATA2(8) => DATA2(8), DATA2(7)
                           => DATA2(7), DATA2(6) => DATA2(6), DATA2(5) => 
                           DATA2(5), DATA2(4) => DATA2(4), DATA2(3) => DATA2(3)
                           , DATA2(2) => DATA2(2), DATA2(1) => DATA2(1), 
                           DATA2(0) => DATA2(0), OUT_ALU(31) => OUTPUT4_31_port
                           , OUT_ALU(30) => OUTPUT4_30_port, OUT_ALU(29) => 
                           OUTPUT4_29_port, OUT_ALU(28) => OUTPUT4_28_port, 
                           OUT_ALU(27) => OUTPUT4_27_port, OUT_ALU(26) => 
                           OUTPUT4_26_port, OUT_ALU(25) => OUTPUT4_25_port, 
                           OUT_ALU(24) => OUTPUT4_24_port, OUT_ALU(23) => 
                           OUTPUT4_23_port, OUT_ALU(22) => OUTPUT4_22_port, 
                           OUT_ALU(21) => OUTPUT4_21_port, OUT_ALU(20) => 
                           OUTPUT4_20_port, OUT_ALU(19) => OUTPUT4_19_port, 
                           OUT_ALU(18) => OUTPUT4_18_port, OUT_ALU(17) => 
                           OUTPUT4_17_port, OUT_ALU(16) => OUTPUT4_16_port, 
                           OUT_ALU(15) => OUTPUT4_15_port, OUT_ALU(14) => 
                           OUTPUT4_14_port, OUT_ALU(13) => OUTPUT4_13_port, 
                           OUT_ALU(12) => OUTPUT4_12_port, OUT_ALU(11) => 
                           OUTPUT4_11_port, OUT_ALU(10) => OUTPUT4_10_port, 
                           OUT_ALU(9) => OUTPUT4_9_port, OUT_ALU(8) => 
                           OUTPUT4_8_port, OUT_ALU(7) => OUTPUT4_7_port, 
                           OUT_ALU(6) => OUTPUT4_6_port, OUT_ALU(5) => 
                           OUTPUT4_5_port, OUT_ALU(4) => OUTPUT4_4_port, 
                           OUT_ALU(3) => OUTPUT4_3_port, OUT_ALU(2) => 
                           OUTPUT4_2_port, OUT_ALU(1) => OUTPUT4_1_port, 
                           OUT_ALU(0) => OUTPUT4_0_port);
   comp : comparator port map( DATA1(31) => OUTPUT2_31_port, DATA1(30) => 
                           OUTPUT2_30_port, DATA1(29) => OUTPUT2_29_port, 
                           DATA1(28) => OUTPUT2_28_port, DATA1(27) => 
                           OUTPUT2_27_port, DATA1(26) => OUTPUT2_26_port, 
                           DATA1(25) => OUTPUT2_25_port, DATA1(24) => 
                           OUTPUT2_24_port, DATA1(23) => OUTPUT2_23_port, 
                           DATA1(22) => OUTPUT2_22_port, DATA1(21) => 
                           OUTPUT2_21_port, DATA1(20) => OUTPUT2_20_port, 
                           DATA1(19) => OUTPUT2_19_port, DATA1(18) => 
                           OUTPUT2_18_port, DATA1(17) => OUTPUT2_17_port, 
                           DATA1(16) => OUTPUT2_16_port, DATA1(15) => 
                           OUTPUT2_15_port, DATA1(14) => OUTPUT2_14_port, 
                           DATA1(13) => OUTPUT2_13_port, DATA1(12) => 
                           OUTPUT2_12_port, DATA1(11) => OUTPUT2_11_port, 
                           DATA1(10) => OUTPUT2_10_port, DATA1(9) => 
                           OUTPUT2_9_port, DATA1(8) => OUTPUT2_8_port, DATA1(7)
                           => OUTPUT2_7_port, DATA1(6) => OUTPUT2_6_port, 
                           DATA1(5) => OUTPUT2_5_port, DATA1(4) => 
                           OUTPUT2_4_port, DATA1(3) => OUTPUT2_3_port, DATA1(2)
                           => OUTPUT2_2_port, DATA1(1) => OUTPUT2_1_port, 
                           DATA1(0) => OUTPUT2_0_port, DATA2i => Cout_i, 
                           tipo(0) => FUNC(0), tipo(1) => FUNC(1), tipo(2) => 
                           FUNC(2), tipo(3) => FUNC(3), tipo(4) => FUNC(4), 
                           tipo(5) => FUNC(5), OUTALU(31) => n_1109, OUTALU(30)
                           => n_1110, OUTALU(29) => n_1111, OUTALU(28) => 
                           n_1112, OUTALU(27) => n_1113, OUTALU(26) => n_1114, 
                           OUTALU(25) => n_1115, OUTALU(24) => n_1116, 
                           OUTALU(23) => n_1117, OUTALU(22) => n_1118, 
                           OUTALU(21) => n_1119, OUTALU(20) => n_1120, 
                           OUTALU(19) => n_1121, OUTALU(18) => n_1122, 
                           OUTALU(17) => n_1123, OUTALU(16) => n_1124, 
                           OUTALU(15) => n_1125, OUTALU(14) => n_1126, 
                           OUTALU(13) => n_1127, OUTALU(12) => n_1128, 
                           OUTALU(11) => n_1129, OUTALU(10) => n_1130, 
                           OUTALU(9) => n_1131, OUTALU(8) => n_1132, OUTALU(7) 
                           => n_1133, OUTALU(6) => n_1134, OUTALU(5) => n_1135,
                           OUTALU(4) => n_1136, OUTALU(3) => n_1137, OUTALU(2) 
                           => n_1138, OUTALU(1) => n_1139, OUTALU(0) => 
                           OUTPUT3_0_port);
   shifter : SHIFTER_GENERIC_N32 port map( A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28), 
                           A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), B(4) => 
                           DATA2(4), B(3) => DATA2(3), B(2) => DATA2(2), B(1) 
                           => DATA2(1), B(0) => DATA2(0), LOGIC_ARITH => 
                           LOGIC_ARITH_i, LEFT_RIGHT => LEFT_RIGHT_i, 
                           SHIFT_ROTATE => SHIFT_ROTATE_i, OUTPUT(31) => 
                           OUTPUT1_31_port, OUTPUT(30) => OUTPUT1_30_port, 
                           OUTPUT(29) => OUTPUT1_29_port, OUTPUT(28) => 
                           OUTPUT1_28_port, OUTPUT(27) => OUTPUT1_27_port, 
                           OUTPUT(26) => OUTPUT1_26_port, OUTPUT(25) => 
                           OUTPUT1_25_port, OUTPUT(24) => OUTPUT1_24_port, 
                           OUTPUT(23) => OUTPUT1_23_port, OUTPUT(22) => 
                           OUTPUT1_22_port, OUTPUT(21) => OUTPUT1_21_port, 
                           OUTPUT(20) => OUTPUT1_20_port, OUTPUT(19) => 
                           OUTPUT1_19_port, OUTPUT(18) => OUTPUT1_18_port, 
                           OUTPUT(17) => OUTPUT1_17_port, OUTPUT(16) => 
                           OUTPUT1_16_port, OUTPUT(15) => OUTPUT1_15_port, 
                           OUTPUT(14) => OUTPUT1_14_port, OUTPUT(13) => 
                           OUTPUT1_13_port, OUTPUT(12) => OUTPUT1_12_port, 
                           OUTPUT(11) => OUTPUT1_11_port, OUTPUT(10) => 
                           OUTPUT1_10_port, OUTPUT(9) => OUTPUT1_9_port, 
                           OUTPUT(8) => OUTPUT1_8_port, OUTPUT(7) => 
                           OUTPUT1_7_port, OUTPUT(6) => OUTPUT1_6_port, 
                           OUTPUT(5) => OUTPUT1_5_port, OUTPUT(4) => 
                           OUTPUT1_4_port, OUTPUT(3) => OUTPUT1_3_port, 
                           OUTPUT(2) => OUTPUT1_2_port, OUTPUT(1) => 
                           OUTPUT1_1_port, OUTPUT(0) => OUTPUT1_0_port);
   adder : P4_ADDER_NBIT32 port map( A(31) => data1i_31_port, A(30) => 
                           data1i_30_port, A(29) => data1i_29_port, A(28) => 
                           data1i_28_port, A(27) => data1i_27_port, A(26) => 
                           data1i_26_port, A(25) => data1i_25_port, A(24) => 
                           data1i_24_port, A(23) => data1i_23_port, A(22) => 
                           data1i_22_port, A(21) => data1i_21_port, A(20) => 
                           data1i_20_port, A(19) => data1i_19_port, A(18) => 
                           data1i_18_port, A(17) => data1i_17_port, A(16) => 
                           data1i_16_port, A(15) => data1i_15_port, A(14) => 
                           data1i_14_port, A(13) => data1i_13_port, A(12) => 
                           data1i_12_port, A(11) => data1i_11_port, A(10) => 
                           data1i_10_port, A(9) => data1i_9_port, A(8) => 
                           data1i_8_port, A(7) => data1i_7_port, A(6) => 
                           data1i_6_port, A(5) => data1i_5_port, A(4) => 
                           data1i_4_port, A(3) => data1i_3_port, A(2) => 
                           data1i_2_port, A(1) => data1i_1_port, A(0) => 
                           data1i_0_port, B(31) => data2i_31_port, B(30) => 
                           data2i_30_port, B(29) => data2i_29_port, B(28) => 
                           data2i_28_port, B(27) => data2i_27_port, B(26) => 
                           data2i_26_port, B(25) => data2i_25_port, B(24) => 
                           data2i_24_port, B(23) => data2i_23_port, B(22) => 
                           data2i_22_port, B(21) => data2i_21_port, B(20) => 
                           data2i_20_port, B(19) => data2i_19_port, B(18) => 
                           data2i_18_port, B(17) => data2i_17_port, B(16) => 
                           data2i_16_port, B(15) => data2i_15_port, B(14) => 
                           data2i_14_port, B(13) => data2i_13_port, B(12) => 
                           data2i_12_port, B(11) => data2i_11_port, B(10) => 
                           data2i_10_port, B(9) => data2i_9_port, B(8) => 
                           data2i_8_port, B(7) => data2i_7_port, B(6) => 
                           data2i_6_port, B(5) => data2i_5_port, B(4) => 
                           data2i_4_port, B(3) => data2i_3_port, B(2) => 
                           data2i_2_port, B(1) => data2i_1_port, B(0) => 
                           data2i_0_port, Cin => Cin_i, S(31) => 
                           OUTPUT2_31_port, S(30) => OUTPUT2_30_port, S(29) => 
                           OUTPUT2_29_port, S(28) => OUTPUT2_28_port, S(27) => 
                           OUTPUT2_27_port, S(26) => OUTPUT2_26_port, S(25) => 
                           OUTPUT2_25_port, S(24) => OUTPUT2_24_port, S(23) => 
                           OUTPUT2_23_port, S(22) => OUTPUT2_22_port, S(21) => 
                           OUTPUT2_21_port, S(20) => OUTPUT2_20_port, S(19) => 
                           OUTPUT2_19_port, S(18) => OUTPUT2_18_port, S(17) => 
                           OUTPUT2_17_port, S(16) => OUTPUT2_16_port, S(15) => 
                           OUTPUT2_15_port, S(14) => OUTPUT2_14_port, S(13) => 
                           OUTPUT2_13_port, S(12) => OUTPUT2_12_port, S(11) => 
                           OUTPUT2_11_port, S(10) => OUTPUT2_10_port, S(9) => 
                           OUTPUT2_9_port, S(8) => OUTPUT2_8_port, S(7) => 
                           OUTPUT2_7_port, S(6) => OUTPUT2_6_port, S(5) => 
                           OUTPUT2_5_port, S(4) => OUTPUT2_4_port, S(3) => 
                           OUTPUT2_3_port, S(2) => OUTPUT2_2_port, S(1) => 
                           OUTPUT2_1_port, S(0) => OUTPUT2_0_port, Cout => 
                           Cout_i);
   U69 : INV_X2 port map( A => n36, ZN => n3);
   U72 : OR3_X2 port map( A1 => n127, A2 => n128, A3 => n36, ZN => n39);
   U75 : INV_X1 port map( A => n40, ZN => n152_port);
   U78 : INV_X2 port map( A => n152_port, ZN => n153_port);
   U81 : INV_X1 port map( A => N139, ZN => n154_port);
   U84 : INV_X2 port map( A => n154_port, ZN => n155_port);
   U87 : INV_X1 port map( A => n2, ZN => n156_port);
   U90 : INV_X2 port map( A => n156_port, ZN => n157_port);
   U93 : INV_X1 port map( A => N206, ZN => n158_port);
   U96 : INV_X4 port map( A => n158_port, ZN => n159_port);
   U99 : NAND2_X2 port map( A1 => OUTPUT1_31_port, A2 => n159_port, ZN => n37);
   U102 : NAND2_X2 port map( A1 => OUTPUT1_30_port, A2 => n159_port, ZN => n42)
                           ;
   U105 : NAND2_X2 port map( A1 => OUTPUT1_29_port, A2 => n159_port, ZN => n44)
                           ;
   U108 : NAND2_X2 port map( A1 => OUTPUT1_28_port, A2 => n159_port, ZN => n46)
                           ;
   U111 : NAND2_X2 port map( A1 => OUTPUT1_27_port, A2 => n159_port, ZN => n48)
                           ;
   U114 : NAND2_X2 port map( A1 => OUTPUT1_26_port, A2 => n159_port, ZN => n50)
                           ;
   U117 : NAND2_X2 port map( A1 => OUTPUT1_25_port, A2 => n159_port, ZN => n52)
                           ;
   U120 : NAND2_X2 port map( A1 => OUTPUT1_24_port, A2 => n159_port, ZN => n54)
                           ;
   U123 : NAND2_X2 port map( A1 => OUTPUT1_23_port, A2 => n159_port, ZN => n56)
                           ;
   U126 : NAND2_X2 port map( A1 => OUTPUT1_22_port, A2 => n159_port, ZN => n58)
                           ;
   U129 : NAND2_X2 port map( A1 => OUTPUT1_21_port, A2 => n159_port, ZN => n60)
                           ;
   U132 : NAND2_X2 port map( A1 => OUTPUT1_20_port, A2 => n159_port, ZN => n62)
                           ;
   U135 : NAND2_X2 port map( A1 => OUTPUT1_19_port, A2 => n159_port, ZN => n64)
                           ;
   U138 : NAND2_X2 port map( A1 => OUTPUT1_18_port, A2 => n159_port, ZN => n66)
                           ;
   U141 : NAND2_X2 port map( A1 => OUTPUT1_17_port, A2 => n159_port, ZN => n68)
                           ;
   U144 : NAND2_X2 port map( A1 => OUTPUT1_16_port, A2 => n159_port, ZN => n70)
                           ;
   U147 : NAND2_X2 port map( A1 => OUTPUT1_15_port, A2 => n159_port, ZN => n72)
                           ;
   U150 : NAND2_X2 port map( A1 => OUTPUT1_14_port, A2 => n159_port, ZN => n74)
                           ;
   U153 : NAND2_X2 port map( A1 => OUTPUT1_13_port, A2 => n159_port, ZN => n76)
                           ;
   U156 : NAND2_X2 port map( A1 => OUTPUT1_12_port, A2 => n159_port, ZN => n78)
                           ;
   U159 : NAND2_X2 port map( A1 => OUTPUT1_11_port, A2 => n159_port, ZN => n80)
                           ;
   U162 : NAND2_X2 port map( A1 => OUTPUT1_10_port, A2 => n159_port, ZN => n82)
                           ;
   U188 : NAND2_X2 port map( A1 => OUTPUT1_9_port, A2 => n159_port, ZN => n84);
   U224 : NAND2_X2 port map( A1 => OUTPUT1_8_port, A2 => n159_port, ZN => n86);
   U225 : NAND2_X2 port map( A1 => OUTPUT1_7_port, A2 => n159_port, ZN => n88);
   U226 : NAND2_X2 port map( A1 => OUTPUT1_6_port, A2 => n159_port, ZN => n90);
   U227 : NAND2_X2 port map( A1 => OUTPUT1_5_port, A2 => n159_port, ZN => n92);
   U228 : NAND2_X2 port map( A1 => OUTPUT1_4_port, A2 => n159_port, ZN => n94);
   U229 : NAND2_X2 port map( A1 => OUTPUT1_3_port, A2 => n159_port, ZN => n96);
   U230 : NAND2_X2 port map( A1 => OUTPUT1_2_port, A2 => n159_port, ZN => n98);
   U231 : NAND2_X2 port map( A1 => OUTPUT1_1_port, A2 => n159_port, ZN => n100)
                           ;

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT6_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 downto 
         0);  Q : out std_logic_vector (5 downto 0));

end regFFD_NBIT6_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT6_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   Q_reg_5_inst : DFFR_X1 port map( D => n18, CK => CK, RN => RESET, Q => Q(5),
                           QN => n12);
   Q_reg_4_inst : DFFR_X1 port map( D => n17, CK => CK, RN => RESET, Q => Q(4),
                           QN => n11);
   Q_reg_3_inst : DFFR_X1 port map( D => n16, CK => CK, RN => RESET, Q => Q(3),
                           QN => n10);
   Q_reg_2_inst : DFFR_X1 port map( D => n15, CK => CK, RN => RESET, Q => Q(2),
                           QN => n9);
   Q_reg_1_inst : DFFR_X1 port map( D => n14, CK => CK, RN => RESET, Q => Q(1),
                           QN => n8);
   Q_reg_0_inst : DFFR_X1 port map( D => n13, CK => CK, RN => RESET, Q => Q(0),
                           QN => n7);
   U2 : OAI21_X1 port map( B1 => n7, B2 => ENABLE, A => n1, ZN => n13);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n8, B2 => ENABLE, A => n2, ZN => n14);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n9, B2 => ENABLE, A => n3, ZN => n15);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n10, B2 => ENABLE, A => n4, ZN => n16);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n4);
   U10 : OAI21_X1 port map( B1 => n11, B2 => ENABLE, A => n5, ZN => n17);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n5);
   U12 : OAI21_X1 port map( B1 => n12, B2 => ENABLE, A => n6, ZN => n18);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n6);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15 : 
      std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n15, CK => CK, RN => RESET, Q => Q(4),
                           QN => n10);
   Q_reg_3_inst : DFFR_X1 port map( D => n14, CK => CK, RN => RESET, Q => Q(3),
                           QN => n9);
   Q_reg_2_inst : DFFR_X1 port map( D => n13, CK => CK, RN => RESET, Q => Q(2),
                           QN => n8);
   Q_reg_1_inst : DFFR_X1 port map( D => n12, CK => CK, RN => RESET, Q => Q(1),
                           QN => n7);
   Q_reg_0_inst : DFFR_X1 port map( D => n11, CK => CK, RN => RESET, Q => Q(0),
                           QN => n6);
   U2 : OAI21_X1 port map( B1 => n6, B2 => ENABLE, A => n1, ZN => n11);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n7, B2 => ENABLE, A => n2, ZN => n12);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n8, B2 => ENABLE, A => n3, ZN => n13);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n9, B2 => ENABLE, A => n4, ZN => n14);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n4);
   U10 : OAI21_X1 port map( B1 => n10, B2 => ENABLE, A => n5, ZN => n15);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n5);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_0 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_0;

architecture SYN_SYNC_BHV of FF_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n3, n4, n_1140 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n4, CK => CLK, Q => Q_port, QN => n_1140);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => n4);
   U4 : INV_X1 port map( A => RESET, ZN => n2);
   U5 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n3, ZN => n1)
                           ;
   U6 : INV_X1 port map( A => EN, ZN => n3);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0);  wr_signal : in std_logic);

end register_file;

architecture SYN_A of register_file is

   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal REGISTERS_2_31_port, REGISTERS_2_30_port, REGISTERS_2_29_port, 
      REGISTERS_2_28_port, REGISTERS_2_27_port, REGISTERS_2_26_port, 
      REGISTERS_2_25_port, REGISTERS_2_24_port, REGISTERS_2_23_port, 
      REGISTERS_2_22_port, REGISTERS_2_21_port, REGISTERS_2_20_port, 
      REGISTERS_2_19_port, REGISTERS_2_18_port, REGISTERS_2_17_port, 
      REGISTERS_2_16_port, REGISTERS_2_15_port, REGISTERS_2_14_port, 
      REGISTERS_2_13_port, REGISTERS_2_12_port, REGISTERS_2_11_port, 
      REGISTERS_2_10_port, REGISTERS_2_9_port, REGISTERS_2_8_port, 
      REGISTERS_2_7_port, REGISTERS_2_6_port, REGISTERS_2_5_port, 
      REGISTERS_2_4_port, REGISTERS_2_3_port, REGISTERS_2_2_port, 
      REGISTERS_2_1_port, REGISTERS_2_0_port, REGISTERS_3_31_port, 
      REGISTERS_3_30_port, REGISTERS_3_29_port, REGISTERS_3_28_port, 
      REGISTERS_3_27_port, REGISTERS_3_26_port, REGISTERS_3_25_port, 
      REGISTERS_3_24_port, REGISTERS_3_23_port, REGISTERS_3_22_port, 
      REGISTERS_3_21_port, REGISTERS_3_20_port, REGISTERS_3_19_port, 
      REGISTERS_3_18_port, REGISTERS_3_17_port, REGISTERS_3_16_port, 
      REGISTERS_3_15_port, REGISTERS_3_14_port, REGISTERS_3_13_port, 
      REGISTERS_3_12_port, REGISTERS_3_11_port, REGISTERS_3_10_port, 
      REGISTERS_3_9_port, REGISTERS_3_8_port, REGISTERS_3_7_port, 
      REGISTERS_3_6_port, REGISTERS_3_5_port, REGISTERS_3_4_port, 
      REGISTERS_3_3_port, REGISTERS_3_2_port, REGISTERS_3_1_port, 
      REGISTERS_3_0_port, REGISTERS_6_31_port, REGISTERS_6_30_port, 
      REGISTERS_6_29_port, REGISTERS_6_28_port, REGISTERS_6_27_port, 
      REGISTERS_6_26_port, REGISTERS_6_25_port, REGISTERS_6_24_port, 
      REGISTERS_6_23_port, REGISTERS_6_22_port, REGISTERS_6_21_port, 
      REGISTERS_6_20_port, REGISTERS_6_19_port, REGISTERS_6_18_port, 
      REGISTERS_6_17_port, REGISTERS_6_16_port, REGISTERS_6_15_port, 
      REGISTERS_6_14_port, REGISTERS_6_13_port, REGISTERS_6_12_port, 
      REGISTERS_6_11_port, REGISTERS_6_10_port, REGISTERS_6_9_port, 
      REGISTERS_6_8_port, REGISTERS_6_7_port, REGISTERS_6_6_port, 
      REGISTERS_6_5_port, REGISTERS_6_4_port, REGISTERS_6_3_port, 
      REGISTERS_6_2_port, REGISTERS_6_1_port, REGISTERS_6_0_port, 
      REGISTERS_7_31_port, REGISTERS_7_30_port, REGISTERS_7_29_port, 
      REGISTERS_7_28_port, REGISTERS_7_27_port, REGISTERS_7_26_port, 
      REGISTERS_7_25_port, REGISTERS_7_24_port, REGISTERS_7_23_port, 
      REGISTERS_7_22_port, REGISTERS_7_21_port, REGISTERS_7_20_port, 
      REGISTERS_7_19_port, REGISTERS_7_18_port, REGISTERS_7_17_port, 
      REGISTERS_7_16_port, REGISTERS_7_15_port, REGISTERS_7_14_port, 
      REGISTERS_7_13_port, REGISTERS_7_12_port, REGISTERS_7_11_port, 
      REGISTERS_7_10_port, REGISTERS_7_9_port, REGISTERS_7_8_port, 
      REGISTERS_7_7_port, REGISTERS_7_6_port, REGISTERS_7_5_port, 
      REGISTERS_7_4_port, REGISTERS_7_3_port, REGISTERS_7_2_port, 
      REGISTERS_7_1_port, REGISTERS_7_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_14_31_port, REGISTERS_14_30_port, REGISTERS_14_29_port, 
      REGISTERS_14_28_port, REGISTERS_14_27_port, REGISTERS_14_26_port, 
      REGISTERS_14_25_port, REGISTERS_14_24_port, REGISTERS_14_23_port, 
      REGISTERS_14_22_port, REGISTERS_14_21_port, REGISTERS_14_20_port, 
      REGISTERS_14_19_port, REGISTERS_14_18_port, REGISTERS_14_17_port, 
      REGISTERS_14_16_port, REGISTERS_14_15_port, REGISTERS_14_14_port, 
      REGISTERS_14_13_port, REGISTERS_14_12_port, REGISTERS_14_11_port, 
      REGISTERS_14_10_port, REGISTERS_14_9_port, REGISTERS_14_8_port, 
      REGISTERS_14_7_port, REGISTERS_14_6_port, REGISTERS_14_5_port, 
      REGISTERS_14_4_port, REGISTERS_14_3_port, REGISTERS_14_2_port, 
      REGISTERS_14_1_port, REGISTERS_14_0_port, REGISTERS_15_31_port, 
      REGISTERS_15_30_port, REGISTERS_15_29_port, REGISTERS_15_28_port, 
      REGISTERS_15_27_port, REGISTERS_15_26_port, REGISTERS_15_25_port, 
      REGISTERS_15_24_port, REGISTERS_15_23_port, REGISTERS_15_22_port, 
      REGISTERS_15_21_port, REGISTERS_15_20_port, REGISTERS_15_19_port, 
      REGISTERS_15_18_port, REGISTERS_15_17_port, REGISTERS_15_16_port, 
      REGISTERS_15_15_port, REGISTERS_15_14_port, REGISTERS_15_13_port, 
      REGISTERS_15_12_port, REGISTERS_15_11_port, REGISTERS_15_10_port, 
      REGISTERS_15_9_port, REGISTERS_15_8_port, REGISTERS_15_7_port, 
      REGISTERS_15_6_port, REGISTERS_15_5_port, REGISTERS_15_4_port, 
      REGISTERS_15_3_port, REGISTERS_15_2_port, REGISTERS_15_1_port, 
      REGISTERS_15_0_port, REGISTERS_18_31_port, REGISTERS_18_30_port, 
      REGISTERS_18_29_port, REGISTERS_18_28_port, REGISTERS_18_27_port, 
      REGISTERS_18_26_port, REGISTERS_18_25_port, REGISTERS_18_24_port, 
      REGISTERS_18_23_port, REGISTERS_18_22_port, REGISTERS_18_21_port, 
      REGISTERS_18_20_port, REGISTERS_18_19_port, REGISTERS_18_18_port, 
      REGISTERS_18_17_port, REGISTERS_18_16_port, REGISTERS_18_15_port, 
      REGISTERS_18_14_port, REGISTERS_18_13_port, REGISTERS_18_12_port, 
      REGISTERS_18_11_port, REGISTERS_18_10_port, REGISTERS_18_9_port, 
      REGISTERS_18_8_port, REGISTERS_18_7_port, REGISTERS_18_6_port, 
      REGISTERS_18_5_port, REGISTERS_18_4_port, REGISTERS_18_3_port, 
      REGISTERS_18_2_port, REGISTERS_18_1_port, REGISTERS_18_0_port, 
      REGISTERS_19_31_port, REGISTERS_19_30_port, REGISTERS_19_29_port, 
      REGISTERS_19_28_port, REGISTERS_19_27_port, REGISTERS_19_26_port, 
      REGISTERS_19_25_port, REGISTERS_19_24_port, REGISTERS_19_23_port, 
      REGISTERS_19_22_port, REGISTERS_19_21_port, REGISTERS_19_20_port, 
      REGISTERS_19_19_port, REGISTERS_19_18_port, REGISTERS_19_17_port, 
      REGISTERS_19_16_port, REGISTERS_19_15_port, REGISTERS_19_14_port, 
      REGISTERS_19_13_port, REGISTERS_19_12_port, REGISTERS_19_11_port, 
      REGISTERS_19_10_port, REGISTERS_19_9_port, REGISTERS_19_8_port, 
      REGISTERS_19_7_port, REGISTERS_19_6_port, REGISTERS_19_5_port, 
      REGISTERS_19_4_port, REGISTERS_19_3_port, REGISTERS_19_2_port, 
      REGISTERS_19_1_port, REGISTERS_19_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_26_31_port, REGISTERS_26_30_port, REGISTERS_26_29_port, 
      REGISTERS_26_28_port, REGISTERS_26_27_port, REGISTERS_26_26_port, 
      REGISTERS_26_25_port, REGISTERS_26_24_port, REGISTERS_26_23_port, 
      REGISTERS_26_22_port, REGISTERS_26_21_port, REGISTERS_26_20_port, 
      REGISTERS_26_19_port, REGISTERS_26_18_port, REGISTERS_26_17_port, 
      REGISTERS_26_16_port, REGISTERS_26_15_port, REGISTERS_26_14_port, 
      REGISTERS_26_13_port, REGISTERS_26_12_port, REGISTERS_26_11_port, 
      REGISTERS_26_10_port, REGISTERS_26_9_port, REGISTERS_26_8_port, 
      REGISTERS_26_7_port, REGISTERS_26_6_port, REGISTERS_26_5_port, 
      REGISTERS_26_4_port, REGISTERS_26_3_port, REGISTERS_26_2_port, 
      REGISTERS_26_1_port, REGISTERS_26_0_port, REGISTERS_27_31_port, 
      REGISTERS_27_30_port, REGISTERS_27_29_port, REGISTERS_27_28_port, 
      REGISTERS_27_27_port, REGISTERS_27_26_port, REGISTERS_27_25_port, 
      REGISTERS_27_24_port, REGISTERS_27_23_port, REGISTERS_27_22_port, 
      REGISTERS_27_21_port, REGISTERS_27_20_port, REGISTERS_27_19_port, 
      REGISTERS_27_18_port, REGISTERS_27_17_port, REGISTERS_27_16_port, 
      REGISTERS_27_15_port, REGISTERS_27_14_port, REGISTERS_27_13_port, 
      REGISTERS_27_12_port, REGISTERS_27_11_port, REGISTERS_27_10_port, 
      REGISTERS_27_9_port, REGISTERS_27_8_port, REGISTERS_27_7_port, 
      REGISTERS_27_6_port, REGISTERS_27_5_port, REGISTERS_27_4_port, 
      REGISTERS_27_3_port, REGISTERS_27_2_port, REGISTERS_27_1_port, 
      REGISTERS_27_0_port, REGISTERS_28_31_port, REGISTERS_28_30_port, 
      REGISTERS_28_29_port, REGISTERS_28_28_port, REGISTERS_28_27_port, 
      REGISTERS_28_26_port, REGISTERS_28_25_port, REGISTERS_28_24_port, 
      REGISTERS_28_23_port, REGISTERS_28_22_port, REGISTERS_28_21_port, 
      REGISTERS_28_20_port, REGISTERS_28_19_port, REGISTERS_28_18_port, 
      REGISTERS_28_17_port, REGISTERS_28_16_port, REGISTERS_28_15_port, 
      REGISTERS_28_14_port, REGISTERS_28_13_port, REGISTERS_28_12_port, 
      REGISTERS_28_11_port, REGISTERS_28_10_port, REGISTERS_28_9_port, 
      REGISTERS_28_8_port, REGISTERS_28_7_port, REGISTERS_28_6_port, 
      REGISTERS_28_5_port, REGISTERS_28_4_port, REGISTERS_28_3_port, 
      REGISTERS_28_2_port, REGISTERS_28_1_port, REGISTERS_28_0_port, 
      REGISTERS_29_31_port, REGISTERS_29_30_port, REGISTERS_29_29_port, 
      REGISTERS_29_28_port, REGISTERS_29_27_port, REGISTERS_29_26_port, 
      REGISTERS_29_25_port, REGISTERS_29_24_port, REGISTERS_29_23_port, 
      REGISTERS_29_22_port, REGISTERS_29_21_port, REGISTERS_29_20_port, 
      REGISTERS_29_19_port, REGISTERS_29_18_port, REGISTERS_29_17_port, 
      REGISTERS_29_16_port, REGISTERS_29_15_port, REGISTERS_29_14_port, 
      REGISTERS_29_13_port, REGISTERS_29_12_port, REGISTERS_29_11_port, 
      REGISTERS_29_10_port, REGISTERS_29_9_port, REGISTERS_29_8_port, 
      REGISTERS_29_7_port, REGISTERS_29_6_port, REGISTERS_29_5_port, 
      REGISTERS_29_4_port, REGISTERS_29_3_port, REGISTERS_29_2_port, 
      REGISTERS_29_1_port, REGISTERS_29_0_port, N286, N287, N288, N289, N290, 
      N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, 
      N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, 
      N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, 
      N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, 
      N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, 
      N351, N352, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286_port, n287_port, n288_port, n289_port, 
      n290_port, n291_port, n292_port, n293_port, n294_port, n295_port, 
      n296_port, n297_port, n298_port, n299_port, n300_port, n301_port, 
      n302_port, n303_port, n304_port, n305_port, n306_port, n307_port, 
      n308_port, n309_port, n310_port, n311_port, n312_port, n313_port, 
      n314_port, n315_port, n316_port, n317_port, n318_port, n319_port, 
      n320_port, n321_port, n322_port, n323_port, n324_port, n325_port, 
      n326_port, n327_port, n328_port, n329_port, n330_port, n331_port, 
      n332_port, n333_port, n334_port, n335_port, n336_port, n337_port, 
      n338_port, n339_port, n340_port, n341_port, n342_port, n343_port, 
      n344_port, n345_port, n346_port, n347_port, n348_port, n349_port, 
      n350_port, n351_port, n352_port, n353, n354, n355, n356, n357, n358, n359
      , n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, 
      n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
      n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, 
      n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, 
      n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, 
      n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, 
      n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
      n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, 
      n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, 
      n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, 
      n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, 
      n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
      n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
      n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, 
      n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, 
      n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, 
      n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
      n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, 
      n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, 
      n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
      n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
      n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
      n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
      n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, 
      n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, 
      n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, 
      n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
      n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, 
      n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
      n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, 
      n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
      n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
      n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, 
      n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, 
      n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, 
      n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, 
      n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
      n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, 
      n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
      n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, 
      n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
      n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
      n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, 
      n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
      n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, 
      n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, 
      n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
      n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, 
      n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, 
      n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
      n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
      n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
      n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
      n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
      n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
      n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
      n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, 
      n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, 
      n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
      n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
      n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, 
      n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
      n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
      n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, 
      n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
      n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
      n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
      n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, 
      n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, 
      n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
      n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
      n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, 
      n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, 
      n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
      n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
      n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, 
      n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, 
      n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
      n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
      n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, 
      n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
      n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
      n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
      n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, 
      n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
      n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
      n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
      n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, 
      n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, 
      n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
      n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
      n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, 
      n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, 
      n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
      n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
      n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, 
      n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, 
      n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, 
      n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
      n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, 
      n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, 
      n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
      n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
      n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
      n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, 
      n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, 
      n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, 
      n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, 
      n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, 
      n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
      n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
      n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
      n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, 
      n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
      n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, 
      n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
      n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, 
      n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, 
      n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, 
      n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
      n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, 
      n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, 
      n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
      n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
      n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, 
      n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, 
      n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, 
      n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
      n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, 
      n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, 
      n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, 
      n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
      n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
      n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, 
      n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
      n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
      n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
      n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, 
      n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
      n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, 
      n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, 
      n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, 
      n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
      n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, 
      n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, 
      n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, 
      n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
      n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, 
      n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, 
      n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, 
      n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, 
      n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
      n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, 
      n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, 
      n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, 
      n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, 
      n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, 
      n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, 
      n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
      n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
      n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, 
      n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, 
      n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, 
      n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, 
      n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, 
      n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
      n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, 
      n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, 
      n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, 
      n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, 
      n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
      n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
      n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
      n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
      n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
      n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, 
      n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
      n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
      n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
      n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
      n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
      n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
      n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
      n3417, n3418, n3419, n3420, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, 
      n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, 
      n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, 
      n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, 
      n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, 
      n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, 
      n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, 
      n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, 
      n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, 
      n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, 
      n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, 
      n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, 
      n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, 
      n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, 
      n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, 
      n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, 
      n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, 
      n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, 
      n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, 
      n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, 
      n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, 
      n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, 
      n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, 
      n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, 
      n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, 
      n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, 
      n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, 
      n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, 
      n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, 
      n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, 
      n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, 
      n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, 
      n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, 
      n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, 
      n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, 
      n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, 
      n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, 
      n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, 
      n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, 
      n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, 
      n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, 
      n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, 
      n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, 
      n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, 
      n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, 
      n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, 
      n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, 
      n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, 
      n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, 
      n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, 
      n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, 
      n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, 
      n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, 
      n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, 
      n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, 
      n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, 
      n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, 
      n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, 
      n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, 
      n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, 
      n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, 
      n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, 
      n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, 
      n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, 
      n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, 
      n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, 
      n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, 
      n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, 
      n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, 
      n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, 
      n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, 
      n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, 
      n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, 
      n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, 
      n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, 
      n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, 
      n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, 
      n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, 
      n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, 
      n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, 
      n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, 
      n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, 
      n_2163, n_2164 : std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFFR_X1 port map( D => n3420, CK => CLK, RN => 
                           RESET, Q => n_1141, QN => n1138);
   REGISTERS_reg_0_30_inst : DFFR_X1 port map( D => n3419, CK => CLK, RN => 
                           RESET, Q => n_1142, QN => n1137);
   REGISTERS_reg_0_29_inst : DFFR_X1 port map( D => n3418, CK => CLK, RN => 
                           RESET, Q => n_1143, QN => n1136);
   REGISTERS_reg_0_28_inst : DFFR_X1 port map( D => n3417, CK => CLK, RN => 
                           RESET, Q => n_1144, QN => n1135);
   REGISTERS_reg_0_27_inst : DFFR_X1 port map( D => n3416, CK => CLK, RN => 
                           RESET, Q => n_1145, QN => n1134);
   REGISTERS_reg_0_26_inst : DFFR_X1 port map( D => n3415, CK => CLK, RN => 
                           RESET, Q => n_1146, QN => n1133);
   REGISTERS_reg_0_25_inst : DFFR_X1 port map( D => n3414, CK => CLK, RN => 
                           RESET, Q => n_1147, QN => n1132);
   REGISTERS_reg_0_24_inst : DFFR_X1 port map( D => n3413, CK => CLK, RN => 
                           RESET, Q => n_1148, QN => n1131);
   REGISTERS_reg_0_23_inst : DFFR_X1 port map( D => n3412, CK => CLK, RN => 
                           RESET, Q => n_1149, QN => n1130);
   REGISTERS_reg_0_22_inst : DFFR_X1 port map( D => n3411, CK => CLK, RN => 
                           RESET, Q => n_1150, QN => n1129);
   REGISTERS_reg_0_21_inst : DFFR_X1 port map( D => n3410, CK => CLK, RN => 
                           RESET, Q => n_1151, QN => n1128);
   REGISTERS_reg_0_20_inst : DFFR_X1 port map( D => n3409, CK => CLK, RN => 
                           RESET, Q => n_1152, QN => n1127);
   REGISTERS_reg_0_19_inst : DFFR_X1 port map( D => n3408, CK => CLK, RN => 
                           RESET, Q => n_1153, QN => n1126);
   REGISTERS_reg_0_18_inst : DFFR_X1 port map( D => n3407, CK => CLK, RN => 
                           RESET, Q => n_1154, QN => n1125);
   REGISTERS_reg_0_17_inst : DFFR_X1 port map( D => n3406, CK => CLK, RN => 
                           RESET, Q => n_1155, QN => n1124);
   REGISTERS_reg_0_16_inst : DFFR_X1 port map( D => n3405, CK => CLK, RN => 
                           RESET, Q => n_1156, QN => n1123);
   REGISTERS_reg_0_15_inst : DFFR_X1 port map( D => n3404, CK => CLK, RN => 
                           RESET, Q => n_1157, QN => n1122);
   REGISTERS_reg_0_14_inst : DFFR_X1 port map( D => n3403, CK => CLK, RN => 
                           RESET, Q => n_1158, QN => n1121);
   REGISTERS_reg_0_13_inst : DFFR_X1 port map( D => n3402, CK => CLK, RN => 
                           RESET, Q => n_1159, QN => n1120);
   REGISTERS_reg_0_12_inst : DFFR_X1 port map( D => n3401, CK => CLK, RN => 
                           RESET, Q => n_1160, QN => n1119);
   REGISTERS_reg_0_11_inst : DFFR_X1 port map( D => n3400, CK => CLK, RN => 
                           RESET, Q => n_1161, QN => n1118);
   REGISTERS_reg_0_10_inst : DFFR_X1 port map( D => n3399, CK => CLK, RN => 
                           RESET, Q => n_1162, QN => n1117);
   REGISTERS_reg_0_9_inst : DFFR_X1 port map( D => n3398, CK => CLK, RN => 
                           RESET, Q => n_1163, QN => n1116);
   REGISTERS_reg_0_8_inst : DFFR_X1 port map( D => n3397, CK => CLK, RN => 
                           RESET, Q => n_1164, QN => n1115);
   REGISTERS_reg_0_7_inst : DFFR_X1 port map( D => n3396, CK => CLK, RN => 
                           RESET, Q => n_1165, QN => n1114);
   REGISTERS_reg_0_6_inst : DFFR_X1 port map( D => n3395, CK => CLK, RN => 
                           RESET, Q => n_1166, QN => n1113);
   REGISTERS_reg_0_5_inst : DFFR_X1 port map( D => n3394, CK => CLK, RN => 
                           RESET, Q => n_1167, QN => n1112);
   REGISTERS_reg_0_4_inst : DFFR_X1 port map( D => n3393, CK => CLK, RN => 
                           RESET, Q => n_1168, QN => n1111);
   REGISTERS_reg_0_3_inst : DFFR_X1 port map( D => n3392, CK => CLK, RN => 
                           RESET, Q => n_1169, QN => n1110);
   REGISTERS_reg_0_2_inst : DFFR_X1 port map( D => n3391, CK => CLK, RN => 
                           RESET, Q => n_1170, QN => n1109);
   REGISTERS_reg_0_1_inst : DFFR_X1 port map( D => n3390, CK => CLK, RN => 
                           RESET, Q => n_1171, QN => n1108);
   REGISTERS_reg_0_0_inst : DFFR_X1 port map( D => n3389, CK => CLK, RN => 
                           RESET, Q => n_1172, QN => n1107);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n3388, CK => CLK, RN => 
                           RESET, Q => n_1173, QN => n1104);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n3387, CK => CLK, RN => 
                           RESET, Q => n_1174, QN => n1103);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n3386, CK => CLK, RN => 
                           RESET, Q => n_1175, QN => n1102);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n3385, CK => CLK, RN => 
                           RESET, Q => n_1176, QN => n1101);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n3384, CK => CLK, RN => 
                           RESET, Q => n_1177, QN => n1100);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n3383, CK => CLK, RN => 
                           RESET, Q => n_1178, QN => n1099);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n3382, CK => CLK, RN => 
                           RESET, Q => n_1179, QN => n1098);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n3381, CK => CLK, RN => 
                           RESET, Q => n_1180, QN => n1097);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n3380, CK => CLK, RN => 
                           RESET, Q => n_1181, QN => n1096);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n3379, CK => CLK, RN => 
                           RESET, Q => n_1182, QN => n1095);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n3378, CK => CLK, RN => 
                           RESET, Q => n_1183, QN => n1094);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n3377, CK => CLK, RN => 
                           RESET, Q => n_1184, QN => n1093);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n3376, CK => CLK, RN => 
                           RESET, Q => n_1185, QN => n1092);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n3375, CK => CLK, RN => 
                           RESET, Q => n_1186, QN => n1091);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n3374, CK => CLK, RN => 
                           RESET, Q => n_1187, QN => n1090);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n3373, CK => CLK, RN => 
                           RESET, Q => n_1188, QN => n1089);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n3372, CK => CLK, RN => 
                           RESET, Q => n_1189, QN => n1088);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n3371, CK => CLK, RN => 
                           RESET, Q => n_1190, QN => n1087);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n3370, CK => CLK, RN => 
                           RESET, Q => n_1191, QN => n1086);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n3369, CK => CLK, RN => 
                           RESET, Q => n_1192, QN => n1085);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n3368, CK => CLK, RN => 
                           RESET, Q => n_1193, QN => n1084);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n3367, CK => CLK, RN => 
                           RESET, Q => n_1194, QN => n1083);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n3366, CK => CLK, RN => 
                           RESET, Q => n_1195, QN => n1082);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n3365, CK => CLK, RN => 
                           RESET, Q => n_1196, QN => n1081);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n3364, CK => CLK, RN => 
                           RESET, Q => n_1197, QN => n1080);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n3363, CK => CLK, RN => 
                           RESET, Q => n_1198, QN => n1079);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n3362, CK => CLK, RN => 
                           RESET, Q => n_1199, QN => n1078);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n3361, CK => CLK, RN => 
                           RESET, Q => n_1200, QN => n1077);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n3360, CK => CLK, RN => 
                           RESET, Q => n_1201, QN => n1076);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n3359, CK => CLK, RN => 
                           RESET, Q => n_1202, QN => n1075);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n3358, CK => CLK, RN => 
                           RESET, Q => n_1203, QN => n1074);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n3357, CK => CLK, RN => 
                           RESET, Q => n_1204, QN => n1073);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n3356, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_31_port, QN => n_1205);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n3355, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_30_port, QN => n_1206);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n3354, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_29_port, QN => n_1207);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n3353, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_28_port, QN => n_1208);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n3352, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_27_port, QN => n_1209);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n3351, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_26_port, QN => n_1210);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n3350, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_25_port, QN => n_1211);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n3349, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_24_port, QN => n_1212);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n3348, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_23_port, QN => n_1213);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n3347, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_22_port, QN => n_1214);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n3346, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_21_port, QN => n_1215);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n3345, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_20_port, QN => n_1216);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n3344, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_19_port, QN => n_1217);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n3343, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_18_port, QN => n_1218);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n3342, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_17_port, QN => n_1219);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n3341, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_16_port, QN => n_1220);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n3340, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_15_port, QN => n_1221);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n3339, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_14_port, QN => n_1222);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n3338, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_13_port, QN => n_1223);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n3337, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_12_port, QN => n_1224);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n3336, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_11_port, QN => n_1225);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n3335, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_10_port, QN => n_1226);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n3334, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_9_port, QN => n_1227);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n3333, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_8_port, QN => n_1228);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n3332, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_7_port, QN => n_1229);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n3331, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_6_port, QN => n_1230);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n3330, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_5_port, QN => n_1231);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n3329, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_4_port, QN => n_1232);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n3328, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_3_port, QN => n_1233);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n3327, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_2_port, QN => n_1234);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n3326, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_1_port, QN => n_1235);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n3325, CK => CLK, RN => 
                           RESET, Q => REGISTERS_2_0_port, QN => n_1236);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n3324, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_31_port, QN => n_1237);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n3323, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_30_port, QN => n_1238);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n3322, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_29_port, QN => n_1239);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n3321, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_28_port, QN => n_1240);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n3320, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_27_port, QN => n_1241);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n3319, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_26_port, QN => n_1242);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n3318, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_25_port, QN => n_1243);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n3317, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_24_port, QN => n_1244);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n3316, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_23_port, QN => n_1245);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n3315, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_22_port, QN => n_1246);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n3314, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_21_port, QN => n_1247);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n3313, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_20_port, QN => n_1248);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n3312, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_19_port, QN => n_1249);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n3311, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_18_port, QN => n_1250);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n3310, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_17_port, QN => n_1251);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n3309, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_16_port, QN => n_1252);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n3308, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_15_port, QN => n_1253);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n3307, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_14_port, QN => n_1254);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n3306, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_13_port, QN => n_1255);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n3305, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_12_port, QN => n_1256);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n3304, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_11_port, QN => n_1257);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n3303, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_10_port, QN => n_1258);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n3302, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_9_port, QN => n_1259);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n3301, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_8_port, QN => n_1260);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n3300, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_7_port, QN => n_1261);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n3299, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_6_port, QN => n_1262);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n3298, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_5_port, QN => n_1263);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n3297, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_4_port, QN => n_1264);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n3296, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_3_port, QN => n_1265);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n3295, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_2_port, QN => n_1266);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n3294, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_1_port, QN => n_1267);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n3293, CK => CLK, RN => 
                           RESET, Q => REGISTERS_3_0_port, QN => n_1268);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n3292, CK => CLK, RN => 
                           RESET, Q => n_1269, QN => n1002);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n3291, CK => CLK, RN => 
                           RESET, Q => n_1270, QN => n1001);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n3290, CK => CLK, RN => 
                           RESET, Q => n_1271, QN => n1000);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n3289, CK => CLK, RN => 
                           RESET, Q => n_1272, QN => n999);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n3288, CK => CLK, RN => 
                           RESET, Q => n_1273, QN => n998);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n3287, CK => CLK, RN => 
                           RESET, Q => n_1274, QN => n997);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n3286, CK => CLK, RN => 
                           RESET, Q => n_1275, QN => n996);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n3285, CK => CLK, RN => 
                           RESET, Q => n_1276, QN => n995);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n3284, CK => CLK, RN => 
                           RESET, Q => n_1277, QN => n994);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n3283, CK => CLK, RN => 
                           RESET, Q => n_1278, QN => n993);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n3282, CK => CLK, RN => 
                           RESET, Q => n_1279, QN => n992);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n3281, CK => CLK, RN => 
                           RESET, Q => n_1280, QN => n991);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n3280, CK => CLK, RN => 
                           RESET, Q => n_1281, QN => n990);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n3279, CK => CLK, RN => 
                           RESET, Q => n_1282, QN => n989);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n3278, CK => CLK, RN => 
                           RESET, Q => n_1283, QN => n988);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n3277, CK => CLK, RN => 
                           RESET, Q => n_1284, QN => n987);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n3276, CK => CLK, RN => 
                           RESET, Q => n_1285, QN => n986);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n3275, CK => CLK, RN => 
                           RESET, Q => n_1286, QN => n985);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n3274, CK => CLK, RN => 
                           RESET, Q => n_1287, QN => n984);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n3273, CK => CLK, RN => 
                           RESET, Q => n_1288, QN => n983);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n3272, CK => CLK, RN => 
                           RESET, Q => n_1289, QN => n982);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n3271, CK => CLK, RN => 
                           RESET, Q => n_1290, QN => n981);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n3270, CK => CLK, RN => 
                           RESET, Q => n_1291, QN => n980);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n3269, CK => CLK, RN => 
                           RESET, Q => n_1292, QN => n979);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n3268, CK => CLK, RN => 
                           RESET, Q => n_1293, QN => n978);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n3267, CK => CLK, RN => 
                           RESET, Q => n_1294, QN => n977);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n3266, CK => CLK, RN => 
                           RESET, Q => n_1295, QN => n976);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n3265, CK => CLK, RN => 
                           RESET, Q => n_1296, QN => n975);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n3264, CK => CLK, RN => 
                           RESET, Q => n_1297, QN => n974);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n3263, CK => CLK, RN => 
                           RESET, Q => n_1298, QN => n973);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n3262, CK => CLK, RN => 
                           RESET, Q => n_1299, QN => n972);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n3261, CK => CLK, RN => 
                           RESET, Q => n_1300, QN => n971);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n3260, CK => CLK, RN => 
                           RESET, Q => n_1301, QN => n968);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n3259, CK => CLK, RN => 
                           RESET, Q => n_1302, QN => n967);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n3258, CK => CLK, RN => 
                           RESET, Q => n_1303, QN => n966);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n3257, CK => CLK, RN => 
                           RESET, Q => n_1304, QN => n965);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n3256, CK => CLK, RN => 
                           RESET, Q => n_1305, QN => n964);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n3255, CK => CLK, RN => 
                           RESET, Q => n_1306, QN => n963);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n3254, CK => CLK, RN => 
                           RESET, Q => n_1307, QN => n962);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n3253, CK => CLK, RN => 
                           RESET, Q => n_1308, QN => n961);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n3252, CK => CLK, RN => 
                           RESET, Q => n_1309, QN => n960);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n3251, CK => CLK, RN => 
                           RESET, Q => n_1310, QN => n959);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n3250, CK => CLK, RN => 
                           RESET, Q => n_1311, QN => n958);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n3249, CK => CLK, RN => 
                           RESET, Q => n_1312, QN => n957);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n3248, CK => CLK, RN => 
                           RESET, Q => n_1313, QN => n956);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n3247, CK => CLK, RN => 
                           RESET, Q => n_1314, QN => n955);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n3246, CK => CLK, RN => 
                           RESET, Q => n_1315, QN => n954);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n3245, CK => CLK, RN => 
                           RESET, Q => n_1316, QN => n953);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n3244, CK => CLK, RN => 
                           RESET, Q => n_1317, QN => n952);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n3243, CK => CLK, RN => 
                           RESET, Q => n_1318, QN => n951);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n3242, CK => CLK, RN => 
                           RESET, Q => n_1319, QN => n950);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n3241, CK => CLK, RN => 
                           RESET, Q => n_1320, QN => n949);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n3240, CK => CLK, RN => 
                           RESET, Q => n_1321, QN => n948);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n3239, CK => CLK, RN => 
                           RESET, Q => n_1322, QN => n947);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n3238, CK => CLK, RN => 
                           RESET, Q => n_1323, QN => n946);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n3237, CK => CLK, RN => 
                           RESET, Q => n_1324, QN => n945);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n3236, CK => CLK, RN => 
                           RESET, Q => n_1325, QN => n944);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n3235, CK => CLK, RN => 
                           RESET, Q => n_1326, QN => n943);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n3234, CK => CLK, RN => 
                           RESET, Q => n_1327, QN => n942);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n3233, CK => CLK, RN => 
                           RESET, Q => n_1328, QN => n941);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n3232, CK => CLK, RN => 
                           RESET, Q => n_1329, QN => n940);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n3231, CK => CLK, RN => 
                           RESET, Q => n_1330, QN => n939);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n3230, CK => CLK, RN => 
                           RESET, Q => n_1331, QN => n938);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n3229, CK => CLK, RN => 
                           RESET, Q => n_1332, QN => n937);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n3228, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_31_port, QN => n_1333);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n3227, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_30_port, QN => n_1334);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n3226, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_29_port, QN => n_1335);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n3225, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_28_port, QN => n_1336);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n3224, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_27_port, QN => n_1337);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n3223, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_26_port, QN => n_1338);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n3222, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_25_port, QN => n_1339);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n3221, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_24_port, QN => n_1340);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n3220, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_23_port, QN => n_1341);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n3219, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_22_port, QN => n_1342);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n3218, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_21_port, QN => n_1343);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n3217, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_20_port, QN => n_1344);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n3216, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_19_port, QN => n_1345);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n3215, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_18_port, QN => n_1346);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n3214, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_17_port, QN => n_1347);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n3213, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_16_port, QN => n_1348);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n3212, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_15_port, QN => n_1349);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n3211, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_14_port, QN => n_1350);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n3210, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_13_port, QN => n_1351);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n3209, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_12_port, QN => n_1352);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n3208, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_11_port, QN => n_1353);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n3207, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_10_port, QN => n_1354);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n3206, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_9_port, QN => n_1355);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n3205, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_8_port, QN => n_1356);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n3204, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_7_port, QN => n_1357);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n3203, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_6_port, QN => n_1358);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n3202, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_5_port, QN => n_1359);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n3201, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_4_port, QN => n_1360);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n3200, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_3_port, QN => n_1361);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n3199, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_2_port, QN => n_1362);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n3198, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_1_port, QN => n_1363);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n3197, CK => CLK, RN => 
                           RESET, Q => REGISTERS_6_0_port, QN => n_1364);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n3196, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_31_port, QN => n_1365);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n3195, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_30_port, QN => n_1366);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n3194, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_29_port, QN => n_1367);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n3193, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_28_port, QN => n_1368);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n3192, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_27_port, QN => n_1369);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n3191, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_26_port, QN => n_1370);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n3190, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_25_port, QN => n_1371);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n3189, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_24_port, QN => n_1372);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n3188, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_23_port, QN => n_1373);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n3187, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_22_port, QN => n_1374);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n3186, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_21_port, QN => n_1375);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n3185, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_20_port, QN => n_1376);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n3184, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_19_port, QN => n_1377);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n3183, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_18_port, QN => n_1378);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n3182, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_17_port, QN => n_1379);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n3181, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_16_port, QN => n_1380);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n3180, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_15_port, QN => n_1381);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n3179, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_14_port, QN => n_1382);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n3178, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_13_port, QN => n_1383);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n3177, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_12_port, QN => n_1384);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n3176, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_11_port, QN => n_1385);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n3175, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_10_port, QN => n_1386);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n3174, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_9_port, QN => n_1387);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n3173, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_8_port, QN => n_1388);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n3172, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_7_port, QN => n_1389);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n3171, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_6_port, QN => n_1390);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n3170, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_5_port, QN => n_1391);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n3169, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_4_port, QN => n_1392);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n3168, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_3_port, QN => n_1393);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n3167, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_2_port, QN => n_1394);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n3166, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_1_port, QN => n_1395);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n3165, CK => CLK, RN => 
                           RESET, Q => REGISTERS_7_0_port, QN => n_1396);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n3164, CK => CLK, RN => 
                           RESET, Q => n_1397, QN => n861);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n3163, CK => CLK, RN => 
                           RESET, Q => n_1398, QN => n860);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n3162, CK => CLK, RN => 
                           RESET, Q => n_1399, QN => n859);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n3161, CK => CLK, RN => 
                           RESET, Q => n_1400, QN => n858);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n3160, CK => CLK, RN => 
                           RESET, Q => n_1401, QN => n857);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n3159, CK => CLK, RN => 
                           RESET, Q => n_1402, QN => n856);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n3158, CK => CLK, RN => 
                           RESET, Q => n_1403, QN => n855);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n3157, CK => CLK, RN => 
                           RESET, Q => n_1404, QN => n854);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n3156, CK => CLK, RN => 
                           RESET, Q => n_1405, QN => n853);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n3155, CK => CLK, RN => 
                           RESET, Q => n_1406, QN => n852);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n3154, CK => CLK, RN => 
                           RESET, Q => n_1407, QN => n851);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n3153, CK => CLK, RN => 
                           RESET, Q => n_1408, QN => n850);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n3152, CK => CLK, RN => 
                           RESET, Q => n_1409, QN => n849);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n3151, CK => CLK, RN => 
                           RESET, Q => n_1410, QN => n848);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n3150, CK => CLK, RN => 
                           RESET, Q => n_1411, QN => n847);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n3149, CK => CLK, RN => 
                           RESET, Q => n_1412, QN => n846);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n3148, CK => CLK, RN => 
                           RESET, Q => n_1413, QN => n845);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n3147, CK => CLK, RN => 
                           RESET, Q => n_1414, QN => n844);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n3146, CK => CLK, RN => 
                           RESET, Q => n_1415, QN => n843);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n3145, CK => CLK, RN => 
                           RESET, Q => n_1416, QN => n842);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n3144, CK => CLK, RN => 
                           RESET, Q => n_1417, QN => n841);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n3143, CK => CLK, RN => 
                           RESET, Q => n_1418, QN => n840);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n3142, CK => CLK, RN => 
                           RESET, Q => n_1419, QN => n839);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n3141, CK => CLK, RN => 
                           RESET, Q => n_1420, QN => n838);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n3140, CK => CLK, RN => 
                           RESET, Q => n_1421, QN => n837);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n3139, CK => CLK, RN => 
                           RESET, Q => n_1422, QN => n836);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n3138, CK => CLK, RN => 
                           RESET, Q => n_1423, QN => n835);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n3137, CK => CLK, RN => 
                           RESET, Q => n_1424, QN => n834);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n3136, CK => CLK, RN => 
                           RESET, Q => n_1425, QN => n833);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n3135, CK => CLK, RN => 
                           RESET, Q => n_1426, QN => n832);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n3134, CK => CLK, RN => 
                           RESET, Q => n_1427, QN => n831);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n3133, CK => CLK, RN => 
                           RESET, Q => n_1428, QN => n830);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n3132, CK => CLK, RN => 
                           RESET, Q => n_1429, QN => n827);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n3131, CK => CLK, RN => 
                           RESET, Q => n_1430, QN => n826);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n3130, CK => CLK, RN => 
                           RESET, Q => n_1431, QN => n825);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n3129, CK => CLK, RN => 
                           RESET, Q => n_1432, QN => n824);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n3128, CK => CLK, RN => 
                           RESET, Q => n_1433, QN => n823);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n3127, CK => CLK, RN => 
                           RESET, Q => n_1434, QN => n822);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n3126, CK => CLK, RN => 
                           RESET, Q => n_1435, QN => n821);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n3125, CK => CLK, RN => 
                           RESET, Q => n_1436, QN => n820);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n3124, CK => CLK, RN => 
                           RESET, Q => n_1437, QN => n819);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n3123, CK => CLK, RN => 
                           RESET, Q => n_1438, QN => n818);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n3122, CK => CLK, RN => 
                           RESET, Q => n_1439, QN => n817);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n3121, CK => CLK, RN => 
                           RESET, Q => n_1440, QN => n816);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n3120, CK => CLK, RN => 
                           RESET, Q => n_1441, QN => n815);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n3119, CK => CLK, RN => 
                           RESET, Q => n_1442, QN => n814);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n3118, CK => CLK, RN => 
                           RESET, Q => n_1443, QN => n813);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n3117, CK => CLK, RN => 
                           RESET, Q => n_1444, QN => n812);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n3116, CK => CLK, RN => 
                           RESET, Q => n_1445, QN => n811);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n3115, CK => CLK, RN => 
                           RESET, Q => n_1446, QN => n810);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n3114, CK => CLK, RN => 
                           RESET, Q => n_1447, QN => n809);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n3113, CK => CLK, RN => 
                           RESET, Q => n_1448, QN => n808);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n3112, CK => CLK, RN => 
                           RESET, Q => n_1449, QN => n807);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n3111, CK => CLK, RN => 
                           RESET, Q => n_1450, QN => n806);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n3110, CK => CLK, RN => 
                           RESET, Q => n_1451, QN => n805);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n3109, CK => CLK, RN => 
                           RESET, Q => n_1452, QN => n804);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n3108, CK => CLK, RN => 
                           RESET, Q => n_1453, QN => n803);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n3107, CK => CLK, RN => 
                           RESET, Q => n_1454, QN => n802);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n3106, CK => CLK, RN => 
                           RESET, Q => n_1455, QN => n801);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n3105, CK => CLK, RN => 
                           RESET, Q => n_1456, QN => n800);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n3104, CK => CLK, RN => 
                           RESET, Q => n_1457, QN => n799);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n3103, CK => CLK, RN => 
                           RESET, Q => n_1458, QN => n798);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n3102, CK => CLK, RN => 
                           RESET, Q => n_1459, QN => n797);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n3101, CK => CLK, RN => 
                           RESET, Q => n_1460, QN => n796);
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n3100, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_31_port, QN => n_1461);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n3099, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_30_port, QN => n_1462);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n3098, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_29_port, QN => n_1463);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n3097, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_28_port, QN => n_1464);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n3096, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_27_port, QN => n_1465);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n3095, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_26_port, QN => n_1466);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n3094, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_25_port, QN => n_1467);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n3093, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_24_port, QN => n_1468);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n3092, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_23_port, QN => n_1469);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n3091, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_22_port, QN => n_1470);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n3090, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_21_port, QN => n_1471);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n3089, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_20_port, QN => n_1472);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n3088, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_19_port, QN => n_1473);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n3087, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_18_port, QN => n_1474);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n3086, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_17_port, QN => n_1475);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n3085, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_16_port, QN => n_1476);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n3084, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_15_port, QN => n_1477);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n3083, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_14_port, QN => n_1478);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n3082, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_13_port, QN => n_1479);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n3081, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_12_port, QN => n_1480);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n3080, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_11_port, QN => n_1481);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n3079, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_10_port, QN => n_1482);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n3078, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_9_port, QN => n_1483);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n3077, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_8_port, QN => n_1484);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n3076, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_7_port, QN => n_1485);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n3075, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_6_port, QN => n_1486);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n3074, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_5_port, QN => n_1487);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n3073, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_4_port, QN => n_1488);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n3072, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_3_port, QN => n_1489);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n3071, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_2_port, QN => n_1490);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n3070, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_1_port, QN => n_1491);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n3069, CK => CLK, RN => 
                           RESET, Q => REGISTERS_10_0_port, QN => n_1492);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n3068, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_31_port, QN => n_1493);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n3067, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_30_port, QN => n_1494);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n3066, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_29_port, QN => n_1495);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n3065, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_28_port, QN => n_1496);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n3064, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_27_port, QN => n_1497);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n3063, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_26_port, QN => n_1498);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n3062, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_25_port, QN => n_1499);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n3061, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_24_port, QN => n_1500);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n3060, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_23_port, QN => n_1501);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n3059, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_22_port, QN => n_1502);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n3058, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_21_port, QN => n_1503);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n3057, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_20_port, QN => n_1504);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n3056, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_19_port, QN => n_1505);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n3055, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_18_port, QN => n_1506);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n3054, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_17_port, QN => n_1507);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n3053, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_16_port, QN => n_1508);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n3052, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_15_port, QN => n_1509);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n3051, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_14_port, QN => n_1510);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n3050, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_13_port, QN => n_1511);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n3049, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_12_port, QN => n_1512);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n3048, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_11_port, QN => n_1513);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n3047, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_10_port, QN => n_1514);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n3046, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_9_port, QN => n_1515);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n3045, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_8_port, QN => n_1516);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n3044, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_7_port, QN => n_1517);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n3043, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_6_port, QN => n_1518);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n3042, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_5_port, QN => n_1519);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n3041, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_4_port, QN => n_1520);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n3040, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_3_port, QN => n_1521);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n3039, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_2_port, QN => n_1522);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n3038, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_1_port, QN => n_1523);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n3037, CK => CLK, RN => 
                           RESET, Q => REGISTERS_11_0_port, QN => n_1524);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n3036, CK => CLK, RN => 
                           RESET, Q => n_1525, QN => n725);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n3035, CK => CLK, RN => 
                           RESET, Q => n_1526, QN => n724);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n3034, CK => CLK, RN => 
                           RESET, Q => n_1527, QN => n723);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n3033, CK => CLK, RN => 
                           RESET, Q => n_1528, QN => n722);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n3032, CK => CLK, RN => 
                           RESET, Q => n_1529, QN => n721);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n3031, CK => CLK, RN => 
                           RESET, Q => n_1530, QN => n720);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n3030, CK => CLK, RN => 
                           RESET, Q => n_1531, QN => n719);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n3029, CK => CLK, RN => 
                           RESET, Q => n_1532, QN => n718);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n3028, CK => CLK, RN => 
                           RESET, Q => n_1533, QN => n717);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n3027, CK => CLK, RN => 
                           RESET, Q => n_1534, QN => n716);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n3026, CK => CLK, RN => 
                           RESET, Q => n_1535, QN => n715);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n3025, CK => CLK, RN => 
                           RESET, Q => n_1536, QN => n714);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n3024, CK => CLK, RN => 
                           RESET, Q => n_1537, QN => n713);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n3023, CK => CLK, RN => 
                           RESET, Q => n_1538, QN => n712);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n3022, CK => CLK, RN => 
                           RESET, Q => n_1539, QN => n711);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n3021, CK => CLK, RN => 
                           RESET, Q => n_1540, QN => n710);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n3020, CK => CLK, RN => 
                           RESET, Q => n_1541, QN => n709);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n3019, CK => CLK, RN => 
                           RESET, Q => n_1542, QN => n708);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n3018, CK => CLK, RN => 
                           RESET, Q => n_1543, QN => n707);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n3017, CK => CLK, RN => 
                           RESET, Q => n_1544, QN => n706);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n3016, CK => CLK, RN => 
                           RESET, Q => n_1545, QN => n705);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n3015, CK => CLK, RN => 
                           RESET, Q => n_1546, QN => n704);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n3014, CK => CLK, RN => 
                           RESET, Q => n_1547, QN => n703);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n3013, CK => CLK, RN => 
                           RESET, Q => n_1548, QN => n702);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n3012, CK => CLK, RN => 
                           RESET, Q => n_1549, QN => n701);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n3011, CK => CLK, RN => 
                           RESET, Q => n_1550, QN => n700);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n3010, CK => CLK, RN => 
                           RESET, Q => n_1551, QN => n699);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n3009, CK => CLK, RN => 
                           RESET, Q => n_1552, QN => n698);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n3008, CK => CLK, RN => 
                           RESET, Q => n_1553, QN => n697);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n3007, CK => CLK, RN => 
                           RESET, Q => n_1554, QN => n696);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n3006, CK => CLK, RN => 
                           RESET, Q => n_1555, QN => n695);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n3005, CK => CLK, RN => 
                           RESET, Q => n_1556, QN => n694);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n3004, CK => CLK, RN => 
                           RESET, Q => n_1557, QN => n691);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n3003, CK => CLK, RN => 
                           RESET, Q => n_1558, QN => n690);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n3002, CK => CLK, RN => 
                           RESET, Q => n_1559, QN => n689);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n3001, CK => CLK, RN => 
                           RESET, Q => n_1560, QN => n688);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n3000, CK => CLK, RN => 
                           RESET, Q => n_1561, QN => n687);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n2999, CK => CLK, RN => 
                           RESET, Q => n_1562, QN => n686);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n2998, CK => CLK, RN => 
                           RESET, Q => n_1563, QN => n685);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n2997, CK => CLK, RN => 
                           RESET, Q => n_1564, QN => n684);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n2996, CK => CLK, RN => 
                           RESET, Q => n_1565, QN => n683);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n2995, CK => CLK, RN => 
                           RESET, Q => n_1566, QN => n682);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n2994, CK => CLK, RN => 
                           RESET, Q => n_1567, QN => n681);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n2993, CK => CLK, RN => 
                           RESET, Q => n_1568, QN => n680);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n2992, CK => CLK, RN => 
                           RESET, Q => n_1569, QN => n679);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n2991, CK => CLK, RN => 
                           RESET, Q => n_1570, QN => n678);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n2990, CK => CLK, RN => 
                           RESET, Q => n_1571, QN => n677);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n2989, CK => CLK, RN => 
                           RESET, Q => n_1572, QN => n676);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n2988, CK => CLK, RN => 
                           RESET, Q => n_1573, QN => n675);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n2987, CK => CLK, RN => 
                           RESET, Q => n_1574, QN => n674);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n2986, CK => CLK, RN => 
                           RESET, Q => n_1575, QN => n673);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n2985, CK => CLK, RN => 
                           RESET, Q => n_1576, QN => n672);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n2984, CK => CLK, RN => 
                           RESET, Q => n_1577, QN => n671);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n2983, CK => CLK, RN => 
                           RESET, Q => n_1578, QN => n670);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n2982, CK => CLK, RN => 
                           RESET, Q => n_1579, QN => n669);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n2981, CK => CLK, RN => 
                           RESET, Q => n_1580, QN => n668);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n2980, CK => CLK, RN => 
                           RESET, Q => n_1581, QN => n667);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n2979, CK => CLK, RN => 
                           RESET, Q => n_1582, QN => n666);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n2978, CK => CLK, RN => 
                           RESET, Q => n_1583, QN => n665);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n2977, CK => CLK, RN => 
                           RESET, Q => n_1584, QN => n664);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n2976, CK => CLK, RN => 
                           RESET, Q => n_1585, QN => n663);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n2975, CK => CLK, RN => 
                           RESET, Q => n_1586, QN => n662);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n2974, CK => CLK, RN => 
                           RESET, Q => n_1587, QN => n661);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n2973, CK => CLK, RN => 
                           RESET, Q => n_1588, QN => n660);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n2972, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_31_port, QN => n_1589);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n2971, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_30_port, QN => n_1590);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n2970, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_29_port, QN => n_1591);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n2969, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_28_port, QN => n_1592);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n2968, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_27_port, QN => n_1593);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n2967, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_26_port, QN => n_1594);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n2966, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_25_port, QN => n_1595);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n2965, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_24_port, QN => n_1596);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n2964, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_23_port, QN => n_1597);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n2963, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_22_port, QN => n_1598);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n2962, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_21_port, QN => n_1599);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n2961, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_20_port, QN => n_1600);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n2960, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_19_port, QN => n_1601);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n2959, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_18_port, QN => n_1602);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n2958, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_17_port, QN => n_1603);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n2957, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_16_port, QN => n_1604);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n2956, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_15_port, QN => n_1605);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n2955, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_14_port, QN => n_1606);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n2954, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_13_port, QN => n_1607);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n2953, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_12_port, QN => n_1608);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n2952, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_11_port, QN => n_1609);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n2951, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_10_port, QN => n_1610);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n2950, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_9_port, QN => n_1611);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n2949, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_8_port, QN => n_1612);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n2948, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_7_port, QN => n_1613);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n2947, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_6_port, QN => n_1614);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n2946, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_5_port, QN => n_1615);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n2945, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_4_port, QN => n_1616);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n2944, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_3_port, QN => n_1617);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n2943, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_2_port, QN => n_1618);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n2942, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_1_port, QN => n_1619);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n2941, CK => CLK, RN => 
                           RESET, Q => REGISTERS_14_0_port, QN => n_1620);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n2940, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_31_port, QN => n_1621);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n2939, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_30_port, QN => n_1622);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n2938, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_29_port, QN => n_1623);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n2937, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_28_port, QN => n_1624);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n2936, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_27_port, QN => n_1625);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n2935, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_26_port, QN => n_1626);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n2934, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_25_port, QN => n_1627);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n2933, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_24_port, QN => n_1628);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n2932, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_23_port, QN => n_1629);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n2931, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_22_port, QN => n_1630);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n2930, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_21_port, QN => n_1631);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n2929, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_20_port, QN => n_1632);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n2928, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_19_port, QN => n_1633);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n2927, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_18_port, QN => n_1634);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n2926, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_17_port, QN => n_1635);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n2925, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_16_port, QN => n_1636);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n2924, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_15_port, QN => n_1637);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n2923, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_14_port, QN => n_1638);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n2922, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_13_port, QN => n_1639);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n2921, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_12_port, QN => n_1640);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n2920, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_11_port, QN => n_1641);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n2919, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_10_port, QN => n_1642);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n2918, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_9_port, QN => n_1643);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n2917, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_8_port, QN => n_1644);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n2916, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_7_port, QN => n_1645);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n2915, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_6_port, QN => n_1646);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n2914, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_5_port, QN => n_1647);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n2913, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_4_port, QN => n_1648);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n2912, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_3_port, QN => n_1649);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n2911, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_2_port, QN => n_1650);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n2910, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_1_port, QN => n_1651);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n2909, CK => CLK, RN => 
                           RESET, Q => REGISTERS_15_0_port, QN => n_1652);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n2908, CK => CLK, RN => 
                           RESET, Q => n_1653, QN => n587);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n2907, CK => CLK, RN => 
                           RESET, Q => n_1654, QN => n586);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n2906, CK => CLK, RN => 
                           RESET, Q => n_1655, QN => n585);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n2905, CK => CLK, RN => 
                           RESET, Q => n_1656, QN => n584);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n2904, CK => CLK, RN => 
                           RESET, Q => n_1657, QN => n583);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n2903, CK => CLK, RN => 
                           RESET, Q => n_1658, QN => n582);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n2902, CK => CLK, RN => 
                           RESET, Q => n_1659, QN => n581);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n2901, CK => CLK, RN => 
                           RESET, Q => n_1660, QN => n580);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n2900, CK => CLK, RN => 
                           RESET, Q => n_1661, QN => n579);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n2899, CK => CLK, RN => 
                           RESET, Q => n_1662, QN => n578);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n2898, CK => CLK, RN => 
                           RESET, Q => n_1663, QN => n577);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n2897, CK => CLK, RN => 
                           RESET, Q => n_1664, QN => n576);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n2896, CK => CLK, RN => 
                           RESET, Q => n_1665, QN => n575);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n2895, CK => CLK, RN => 
                           RESET, Q => n_1666, QN => n574);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n2894, CK => CLK, RN => 
                           RESET, Q => n_1667, QN => n573);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n2893, CK => CLK, RN => 
                           RESET, Q => n_1668, QN => n572);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n2892, CK => CLK, RN => 
                           RESET, Q => n_1669, QN => n571);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n2891, CK => CLK, RN => 
                           RESET, Q => n_1670, QN => n570);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n2890, CK => CLK, RN => 
                           RESET, Q => n_1671, QN => n569);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n2889, CK => CLK, RN => 
                           RESET, Q => n_1672, QN => n568);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n2888, CK => CLK, RN => 
                           RESET, Q => n_1673, QN => n567);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n2887, CK => CLK, RN => 
                           RESET, Q => n_1674, QN => n566);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n2886, CK => CLK, RN => 
                           RESET, Q => n_1675, QN => n565);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n2885, CK => CLK, RN => 
                           RESET, Q => n_1676, QN => n564);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n2884, CK => CLK, RN => 
                           RESET, Q => n_1677, QN => n563);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n2883, CK => CLK, RN => 
                           RESET, Q => n_1678, QN => n562);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n2882, CK => CLK, RN => 
                           RESET, Q => n_1679, QN => n561);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n2881, CK => CLK, RN => 
                           RESET, Q => n_1680, QN => n560);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n2880, CK => CLK, RN => 
                           RESET, Q => n_1681, QN => n559);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n2879, CK => CLK, RN => 
                           RESET, Q => n_1682, QN => n558);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n2878, CK => CLK, RN => 
                           RESET, Q => n_1683, QN => n557);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n2877, CK => CLK, RN => 
                           RESET, Q => n_1684, QN => n556);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n2876, CK => CLK, RN => 
                           RESET, Q => n_1685, QN => n553);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n2875, CK => CLK, RN => 
                           RESET, Q => n_1686, QN => n552);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n2874, CK => CLK, RN => 
                           RESET, Q => n_1687, QN => n551);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n2873, CK => CLK, RN => 
                           RESET, Q => n_1688, QN => n550);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n2872, CK => CLK, RN => 
                           RESET, Q => n_1689, QN => n549);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n2871, CK => CLK, RN => 
                           RESET, Q => n_1690, QN => n548);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n2870, CK => CLK, RN => 
                           RESET, Q => n_1691, QN => n547);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n2869, CK => CLK, RN => 
                           RESET, Q => n_1692, QN => n546);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n2868, CK => CLK, RN => 
                           RESET, Q => n_1693, QN => n545);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n2867, CK => CLK, RN => 
                           RESET, Q => n_1694, QN => n544);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n2866, CK => CLK, RN => 
                           RESET, Q => n_1695, QN => n543);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n2865, CK => CLK, RN => 
                           RESET, Q => n_1696, QN => n542);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n2864, CK => CLK, RN => 
                           RESET, Q => n_1697, QN => n541);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n2863, CK => CLK, RN => 
                           RESET, Q => n_1698, QN => n540);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n2862, CK => CLK, RN => 
                           RESET, Q => n_1699, QN => n539);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n2861, CK => CLK, RN => 
                           RESET, Q => n_1700, QN => n538);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n2860, CK => CLK, RN => 
                           RESET, Q => n_1701, QN => n537);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n2859, CK => CLK, RN => 
                           RESET, Q => n_1702, QN => n536);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n2858, CK => CLK, RN => 
                           RESET, Q => n_1703, QN => n535);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n2857, CK => CLK, RN => 
                           RESET, Q => n_1704, QN => n534);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n2856, CK => CLK, RN => 
                           RESET, Q => n_1705, QN => n533);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n2855, CK => CLK, RN => 
                           RESET, Q => n_1706, QN => n532);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n2854, CK => CLK, RN => 
                           RESET, Q => n_1707, QN => n531);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n2853, CK => CLK, RN => 
                           RESET, Q => n_1708, QN => n530);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n2852, CK => CLK, RN => 
                           RESET, Q => n_1709, QN => n529);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n2851, CK => CLK, RN => 
                           RESET, Q => n_1710, QN => n528);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n2850, CK => CLK, RN => 
                           RESET, Q => n_1711, QN => n527);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n2849, CK => CLK, RN => 
                           RESET, Q => n_1712, QN => n526);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n2848, CK => CLK, RN => 
                           RESET, Q => n_1713, QN => n525);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n2847, CK => CLK, RN => 
                           RESET, Q => n_1714, QN => n524);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n2846, CK => CLK, RN => 
                           RESET, Q => n_1715, QN => n523);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n2845, CK => CLK, RN => 
                           RESET, Q => n_1716, QN => n522);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n2844, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_31_port, QN => n_1717);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n2843, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_30_port, QN => n_1718);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n2842, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_29_port, QN => n_1719);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n2841, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_28_port, QN => n_1720);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n2840, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_27_port, QN => n_1721);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n2839, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_26_port, QN => n_1722);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n2838, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_25_port, QN => n_1723);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n2837, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_24_port, QN => n_1724);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n2836, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_23_port, QN => n_1725);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n2835, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_22_port, QN => n_1726);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n2834, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_21_port, QN => n_1727);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n2833, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_20_port, QN => n_1728);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n2832, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_19_port, QN => n_1729);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n2831, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_18_port, QN => n_1730);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n2830, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_17_port, QN => n_1731);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n2829, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_16_port, QN => n_1732);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n2828, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_15_port, QN => n_1733);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n2827, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_14_port, QN => n_1734);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n2826, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_13_port, QN => n_1735);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n2825, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_12_port, QN => n_1736);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n2824, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_11_port, QN => n_1737);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n2823, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_10_port, QN => n_1738);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n2822, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_9_port, QN => n_1739);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n2821, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_8_port, QN => n_1740);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n2820, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_7_port, QN => n_1741);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n2819, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_6_port, QN => n_1742);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n2818, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_5_port, QN => n_1743);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n2817, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_4_port, QN => n_1744);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n2816, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_3_port, QN => n_1745);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n2815, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_2_port, QN => n_1746);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n2814, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_1_port, QN => n_1747);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n2813, CK => CLK, RN => 
                           RESET, Q => REGISTERS_18_0_port, QN => n_1748);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n2812, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_31_port, QN => n_1749);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n2811, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_30_port, QN => n_1750);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n2810, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_29_port, QN => n_1751);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n2809, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_28_port, QN => n_1752);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n2808, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_27_port, QN => n_1753);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n2807, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_26_port, QN => n_1754);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n2806, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_25_port, QN => n_1755);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n2805, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_24_port, QN => n_1756);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n2804, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_23_port, QN => n_1757);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n2803, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_22_port, QN => n_1758);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n2802, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_21_port, QN => n_1759);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n2801, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_20_port, QN => n_1760);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n2800, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_19_port, QN => n_1761);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n2799, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_18_port, QN => n_1762);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n2798, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_17_port, QN => n_1763);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n2797, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_16_port, QN => n_1764);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n2796, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_15_port, QN => n_1765);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n2795, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_14_port, QN => n_1766);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n2794, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_13_port, QN => n_1767);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n2793, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_12_port, QN => n_1768);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n2792, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_11_port, QN => n_1769);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n2791, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_10_port, QN => n_1770);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n2790, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_9_port, QN => n_1771);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n2789, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_8_port, QN => n_1772);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n2788, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_7_port, QN => n_1773);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n2787, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_6_port, QN => n_1774);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n2786, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_5_port, QN => n_1775);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n2785, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_4_port, QN => n_1776);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n2784, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_3_port, QN => n_1777);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n2783, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_2_port, QN => n_1778);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n2782, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_1_port, QN => n_1779);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n2781, CK => CLK, RN => 
                           RESET, Q => REGISTERS_19_0_port, QN => n_1780);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n2780, CK => CLK, RN => 
                           RESET, Q => n_1781, QN => n451);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n2779, CK => CLK, RN => 
                           RESET, Q => n_1782, QN => n450);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n2778, CK => CLK, RN => 
                           RESET, Q => n_1783, QN => n449);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n2777, CK => CLK, RN => 
                           RESET, Q => n_1784, QN => n448);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n2776, CK => CLK, RN => 
                           RESET, Q => n_1785, QN => n447);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n2775, CK => CLK, RN => 
                           RESET, Q => n_1786, QN => n446);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n2774, CK => CLK, RN => 
                           RESET, Q => n_1787, QN => n445);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n2773, CK => CLK, RN => 
                           RESET, Q => n_1788, QN => n444);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n2772, CK => CLK, RN => 
                           RESET, Q => n_1789, QN => n443);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n2771, CK => CLK, RN => 
                           RESET, Q => n_1790, QN => n442);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n2770, CK => CLK, RN => 
                           RESET, Q => n_1791, QN => n441);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n2769, CK => CLK, RN => 
                           RESET, Q => n_1792, QN => n440);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n2768, CK => CLK, RN => 
                           RESET, Q => n_1793, QN => n439);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n2767, CK => CLK, RN => 
                           RESET, Q => n_1794, QN => n438);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n2766, CK => CLK, RN => 
                           RESET, Q => n_1795, QN => n437);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n2765, CK => CLK, RN => 
                           RESET, Q => n_1796, QN => n436);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n2764, CK => CLK, RN => 
                           RESET, Q => n_1797, QN => n435);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n2763, CK => CLK, RN => 
                           RESET, Q => n_1798, QN => n434);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n2762, CK => CLK, RN => 
                           RESET, Q => n_1799, QN => n433);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n2761, CK => CLK, RN => 
                           RESET, Q => n_1800, QN => n432);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n2760, CK => CLK, RN => 
                           RESET, Q => n_1801, QN => n431);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n2759, CK => CLK, RN => 
                           RESET, Q => n_1802, QN => n430);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n2758, CK => CLK, RN => 
                           RESET, Q => n_1803, QN => n429);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n2757, CK => CLK, RN => 
                           RESET, Q => n_1804, QN => n428);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n2756, CK => CLK, RN => 
                           RESET, Q => n_1805, QN => n427);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n2755, CK => CLK, RN => 
                           RESET, Q => n_1806, QN => n426);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n2754, CK => CLK, RN => 
                           RESET, Q => n_1807, QN => n425);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n2753, CK => CLK, RN => 
                           RESET, Q => n_1808, QN => n424);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n2752, CK => CLK, RN => 
                           RESET, Q => n_1809, QN => n423);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n2751, CK => CLK, RN => 
                           RESET, Q => n_1810, QN => n422);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n2750, CK => CLK, RN => 
                           RESET, Q => n_1811, QN => n421);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n2749, CK => CLK, RN => 
                           RESET, Q => n_1812, QN => n420);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n2748, CK => CLK, RN => 
                           RESET, Q => n_1813, QN => n417);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n2747, CK => CLK, RN => 
                           RESET, Q => n_1814, QN => n416);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n2746, CK => CLK, RN => 
                           RESET, Q => n_1815, QN => n415);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n2745, CK => CLK, RN => 
                           RESET, Q => n_1816, QN => n414);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n2744, CK => CLK, RN => 
                           RESET, Q => n_1817, QN => n413);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n2743, CK => CLK, RN => 
                           RESET, Q => n_1818, QN => n412);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n2742, CK => CLK, RN => 
                           RESET, Q => n_1819, QN => n411);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n2741, CK => CLK, RN => 
                           RESET, Q => n_1820, QN => n410);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n2740, CK => CLK, RN => 
                           RESET, Q => n_1821, QN => n409);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n2739, CK => CLK, RN => 
                           RESET, Q => n_1822, QN => n408);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n2738, CK => CLK, RN => 
                           RESET, Q => n_1823, QN => n407);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n2737, CK => CLK, RN => 
                           RESET, Q => n_1824, QN => n406);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n2736, CK => CLK, RN => 
                           RESET, Q => n_1825, QN => n405);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n2735, CK => CLK, RN => 
                           RESET, Q => n_1826, QN => n404);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n2734, CK => CLK, RN => 
                           RESET, Q => n_1827, QN => n403);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n2733, CK => CLK, RN => 
                           RESET, Q => n_1828, QN => n402);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n2732, CK => CLK, RN => 
                           RESET, Q => n_1829, QN => n401);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n2731, CK => CLK, RN => 
                           RESET, Q => n_1830, QN => n400);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n2730, CK => CLK, RN => 
                           RESET, Q => n_1831, QN => n399);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n2729, CK => CLK, RN => 
                           RESET, Q => n_1832, QN => n398);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n2728, CK => CLK, RN => 
                           RESET, Q => n_1833, QN => n397);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n2727, CK => CLK, RN => 
                           RESET, Q => n_1834, QN => n396);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n2726, CK => CLK, RN => 
                           RESET, Q => n_1835, QN => n395);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n2725, CK => CLK, RN => 
                           RESET, Q => n_1836, QN => n394);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n2724, CK => CLK, RN => 
                           RESET, Q => n_1837, QN => n393);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n2723, CK => CLK, RN => 
                           RESET, Q => n_1838, QN => n392);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n2722, CK => CLK, RN => 
                           RESET, Q => n_1839, QN => n391);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n2721, CK => CLK, RN => 
                           RESET, Q => n_1840, QN => n390);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n2720, CK => CLK, RN => 
                           RESET, Q => n_1841, QN => n389);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n2719, CK => CLK, RN => 
                           RESET, Q => n_1842, QN => n388);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n2718, CK => CLK, RN => 
                           RESET, Q => n_1843, QN => n387);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n2717, CK => CLK, RN => 
                           RESET, Q => n_1844, QN => n386);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n2716, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_31_port, QN => n_1845);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n2715, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_30_port, QN => n_1846);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n2714, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_29_port, QN => n_1847);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n2713, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_28_port, QN => n_1848);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n2712, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_27_port, QN => n_1849);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n2711, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_26_port, QN => n_1850);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n2710, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_25_port, QN => n_1851);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n2709, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_24_port, QN => n_1852);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n2708, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_23_port, QN => n_1853);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n2707, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_22_port, QN => n_1854);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n2706, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_21_port, QN => n_1855);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n2705, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_20_port, QN => n_1856);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n2704, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_19_port, QN => n_1857);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n2703, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_18_port, QN => n_1858);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n2702, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_17_port, QN => n_1859);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n2701, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_16_port, QN => n_1860);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n2700, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_15_port, QN => n_1861);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n2699, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_14_port, QN => n_1862);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n2698, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_13_port, QN => n_1863);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n2697, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_12_port, QN => n_1864);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n2696, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_11_port, QN => n_1865);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n2695, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_10_port, QN => n_1866);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n2694, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_9_port, QN => n_1867);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n2693, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_8_port, QN => n_1868);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n2692, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_7_port, QN => n_1869);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n2691, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_6_port, QN => n_1870);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n2690, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_5_port, QN => n_1871);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n2689, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_4_port, QN => n_1872);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n2688, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_3_port, QN => n_1873);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n2687, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_2_port, QN => n_1874);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n2686, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_1_port, QN => n_1875);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n2685, CK => CLK, RN => 
                           RESET, Q => REGISTERS_22_0_port, QN => n_1876);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n2684, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_31_port, QN => n_1877);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n2683, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_30_port, QN => n_1878);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n2682, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_29_port, QN => n_1879);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n2681, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_28_port, QN => n_1880);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n2680, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_27_port, QN => n_1881);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n2679, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_26_port, QN => n_1882);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n2678, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_25_port, QN => n_1883);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n2677, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_24_port, QN => n_1884);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n2676, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_23_port, QN => n_1885);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n2675, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_22_port, QN => n_1886);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n2674, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_21_port, QN => n_1887);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n2673, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_20_port, QN => n_1888);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n2672, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_19_port, QN => n_1889);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n2671, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_18_port, QN => n_1890);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n2670, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_17_port, QN => n_1891);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n2669, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_16_port, QN => n_1892);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n2668, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_15_port, QN => n_1893);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n2667, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_14_port, QN => n_1894);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n2666, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_13_port, QN => n_1895);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n2665, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_12_port, QN => n_1896);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n2664, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_11_port, QN => n_1897);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n2663, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_10_port, QN => n_1898);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n2662, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_9_port, QN => n_1899);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n2661, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_8_port, QN => n_1900);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n2660, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_7_port, QN => n_1901);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n2659, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_6_port, QN => n_1902);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n2658, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_5_port, QN => n_1903);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n2657, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_4_port, QN => n_1904);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n2656, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_3_port, QN => n_1905);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n2655, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_2_port, QN => n_1906);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n2654, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_1_port, QN => n_1907);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n2653, CK => CLK, RN => 
                           RESET, Q => REGISTERS_23_0_port, QN => n_1908);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n2652, CK => CLK, RN => 
                           RESET, Q => n_1909, QN => n312_port);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n2651, CK => CLK, RN => 
                           RESET, Q => n_1910, QN => n311_port);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n2650, CK => CLK, RN => 
                           RESET, Q => n_1911, QN => n310_port);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n2649, CK => CLK, RN => 
                           RESET, Q => n_1912, QN => n309_port);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n2648, CK => CLK, RN => 
                           RESET, Q => n_1913, QN => n308_port);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n2647, CK => CLK, RN => 
                           RESET, Q => n_1914, QN => n307_port);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n2646, CK => CLK, RN => 
                           RESET, Q => n_1915, QN => n306_port);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n2645, CK => CLK, RN => 
                           RESET, Q => n_1916, QN => n305_port);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n2644, CK => CLK, RN => 
                           RESET, Q => n_1917, QN => n304_port);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n2643, CK => CLK, RN => 
                           RESET, Q => n_1918, QN => n303_port);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n2642, CK => CLK, RN => 
                           RESET, Q => n_1919, QN => n302_port);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n2641, CK => CLK, RN => 
                           RESET, Q => n_1920, QN => n301_port);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n2640, CK => CLK, RN => 
                           RESET, Q => n_1921, QN => n300_port);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n2639, CK => CLK, RN => 
                           RESET, Q => n_1922, QN => n299_port);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n2638, CK => CLK, RN => 
                           RESET, Q => n_1923, QN => n298_port);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n2637, CK => CLK, RN => 
                           RESET, Q => n_1924, QN => n297_port);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n2636, CK => CLK, RN => 
                           RESET, Q => n_1925, QN => n296_port);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n2635, CK => CLK, RN => 
                           RESET, Q => n_1926, QN => n295_port);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n2634, CK => CLK, RN => 
                           RESET, Q => n_1927, QN => n294_port);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n2633, CK => CLK, RN => 
                           RESET, Q => n_1928, QN => n293_port);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n2632, CK => CLK, RN => 
                           RESET, Q => n_1929, QN => n292_port);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n2631, CK => CLK, RN => 
                           RESET, Q => n_1930, QN => n291_port);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n2630, CK => CLK, RN => 
                           RESET, Q => n_1931, QN => n290_port);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n2629, CK => CLK, RN => 
                           RESET, Q => n_1932, QN => n289_port);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n2628, CK => CLK, RN => 
                           RESET, Q => n_1933, QN => n288_port);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n2627, CK => CLK, RN => 
                           RESET, Q => n_1934, QN => n287_port);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n2626, CK => CLK, RN => 
                           RESET, Q => n_1935, QN => n286_port);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n2625, CK => CLK, RN => 
                           RESET, Q => n_1936, QN => n285);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n2624, CK => CLK, RN => 
                           RESET, Q => n_1937, QN => n284);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n2623, CK => CLK, RN => 
                           RESET, Q => n_1938, QN => n283);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n2622, CK => CLK, RN => 
                           RESET, Q => n_1939, QN => n282);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n2621, CK => CLK, RN => 
                           RESET, Q => n_1940, QN => n281);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n2620, CK => CLK, RN => 
                           RESET, Q => n_1941, QN => n277);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n2619, CK => CLK, RN => 
                           RESET, Q => n_1942, QN => n276);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n2618, CK => CLK, RN => 
                           RESET, Q => n_1943, QN => n275);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n2617, CK => CLK, RN => 
                           RESET, Q => n_1944, QN => n274);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n2616, CK => CLK, RN => 
                           RESET, Q => n_1945, QN => n273);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n2615, CK => CLK, RN => 
                           RESET, Q => n_1946, QN => n272);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n2614, CK => CLK, RN => 
                           RESET, Q => n_1947, QN => n271);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n2613, CK => CLK, RN => 
                           RESET, Q => n_1948, QN => n270);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n2612, CK => CLK, RN => 
                           RESET, Q => n_1949, QN => n269);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n2611, CK => CLK, RN => 
                           RESET, Q => n_1950, QN => n268);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n2610, CK => CLK, RN => 
                           RESET, Q => n_1951, QN => n267);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n2609, CK => CLK, RN => 
                           RESET, Q => n_1952, QN => n266);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n2608, CK => CLK, RN => 
                           RESET, Q => n_1953, QN => n265);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n2607, CK => CLK, RN => 
                           RESET, Q => n_1954, QN => n264);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n2606, CK => CLK, RN => 
                           RESET, Q => n_1955, QN => n263);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n2605, CK => CLK, RN => 
                           RESET, Q => n_1956, QN => n262);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n2604, CK => CLK, RN => 
                           RESET, Q => n_1957, QN => n261);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n2603, CK => CLK, RN => 
                           RESET, Q => n_1958, QN => n260);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n2602, CK => CLK, RN => 
                           RESET, Q => n_1959, QN => n259);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n2601, CK => CLK, RN => 
                           RESET, Q => n_1960, QN => n258);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n2600, CK => CLK, RN => 
                           RESET, Q => n_1961, QN => n257);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n2599, CK => CLK, RN => 
                           RESET, Q => n_1962, QN => n256);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n2598, CK => CLK, RN => 
                           RESET, Q => n_1963, QN => n255);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n2597, CK => CLK, RN => 
                           RESET, Q => n_1964, QN => n254);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n2596, CK => CLK, RN => 
                           RESET, Q => n_1965, QN => n253);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n2595, CK => CLK, RN => 
                           RESET, Q => n_1966, QN => n252);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n2594, CK => CLK, RN => 
                           RESET, Q => n_1967, QN => n251);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n2593, CK => CLK, RN => 
                           RESET, Q => n_1968, QN => n250);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n2592, CK => CLK, RN => 
                           RESET, Q => n_1969, QN => n249);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n2591, CK => CLK, RN => 
                           RESET, Q => n_1970, QN => n248);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n2590, CK => CLK, RN => 
                           RESET, Q => n_1971, QN => n247);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n2589, CK => CLK, RN => 
                           RESET, Q => n_1972, QN => n246);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n2588, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_31_port, QN => n_1973);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n2587, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_30_port, QN => n_1974);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n2586, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_29_port, QN => n_1975);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n2585, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_28_port, QN => n_1976);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n2584, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_27_port, QN => n_1977);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n2583, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_26_port, QN => n_1978);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n2582, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_25_port, QN => n_1979);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n2581, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_24_port, QN => n_1980);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n2580, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_23_port, QN => n_1981);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n2579, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_22_port, QN => n_1982);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n2578, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_21_port, QN => n_1983);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n2577, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_20_port, QN => n_1984);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n2576, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_19_port, QN => n_1985);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n2575, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_18_port, QN => n_1986);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n2574, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_17_port, QN => n_1987);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n2573, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_16_port, QN => n_1988);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n2572, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_15_port, QN => n_1989);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n2571, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_14_port, QN => n_1990);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n2570, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_13_port, QN => n_1991);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n2569, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_12_port, QN => n_1992);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n2568, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_11_port, QN => n_1993);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n2567, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_10_port, QN => n_1994);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n2566, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_9_port, QN => n_1995);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n2565, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_8_port, QN => n_1996);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n2564, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_7_port, QN => n_1997);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n2563, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_6_port, QN => n_1998);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n2562, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_5_port, QN => n_1999);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n2561, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_4_port, QN => n_2000);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n2560, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_3_port, QN => n_2001);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n2559, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_2_port, QN => n_2002);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n2558, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_1_port, QN => n_2003);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n2557, CK => CLK, RN => 
                           RESET, Q => REGISTERS_26_0_port, QN => n_2004);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n2556, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_31_port, QN => n_2005);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n2555, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_30_port, QN => n_2006);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n2554, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_29_port, QN => n_2007);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n2553, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_28_port, QN => n_2008);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n2552, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_27_port, QN => n_2009);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n2551, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_26_port, QN => n_2010);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n2550, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_25_port, QN => n_2011);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n2549, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_24_port, QN => n_2012);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n2548, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_23_port, QN => n_2013);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n2547, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_22_port, QN => n_2014);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n2546, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_21_port, QN => n_2015);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n2545, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_20_port, QN => n_2016);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n2544, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_19_port, QN => n_2017);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n2543, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_18_port, QN => n_2018);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n2542, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_17_port, QN => n_2019);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n2541, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_16_port, QN => n_2020);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n2540, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_15_port, QN => n_2021);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n2539, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_14_port, QN => n_2022);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n2538, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_13_port, QN => n_2023);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n2537, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_12_port, QN => n_2024);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n2536, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_11_port, QN => n_2025);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n2535, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_10_port, QN => n_2026);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n2534, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_9_port, QN => n_2027);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n2533, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_8_port, QN => n_2028);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n2532, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_7_port, QN => n_2029);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n2531, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_6_port, QN => n_2030);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n2530, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_5_port, QN => n_2031);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n2529, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_4_port, QN => n_2032);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n2528, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_3_port, QN => n_2033);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n2527, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_2_port, QN => n_2034);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n2526, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_1_port, QN => n_2035);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n2525, CK => CLK, RN => 
                           RESET, Q => REGISTERS_27_0_port, QN => n_2036);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n2524, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_31_port, QN => n_2037);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n2523, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_30_port, QN => n_2038);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n2522, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_29_port, QN => n_2039);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n2521, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_28_port, QN => n_2040);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n2520, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_27_port, QN => n_2041);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n2519, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_26_port, QN => n_2042);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n2518, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_25_port, QN => n_2043);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n2517, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_24_port, QN => n_2044);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n2516, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_23_port, QN => n_2045);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n2515, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_22_port, QN => n_2046);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n2514, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_21_port, QN => n_2047);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n2513, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_20_port, QN => n_2048);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n2512, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_19_port, QN => n_2049);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n2511, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_18_port, QN => n_2050);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n2510, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_17_port, QN => n_2051);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n2509, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_16_port, QN => n_2052);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n2508, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_15_port, QN => n_2053);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n2507, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_14_port, QN => n_2054);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n2506, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_13_port, QN => n_2055);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n2505, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_12_port, QN => n_2056);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n2504, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_11_port, QN => n_2057);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n2503, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_10_port, QN => n_2058);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n2502, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_9_port, QN => n_2059);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n2501, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_8_port, QN => n_2060);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n2500, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_7_port, QN => n_2061);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n2499, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_6_port, QN => n_2062);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n2498, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_5_port, QN => n_2063);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n2497, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_4_port, QN => n_2064);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n2496, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_3_port, QN => n_2065);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n2495, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_2_port, QN => n_2066);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n2494, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_1_port, QN => n_2067);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n2493, CK => CLK, RN => 
                           RESET, Q => REGISTERS_28_0_port, QN => n_2068);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n2492, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_31_port, QN => n_2069);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n2491, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_30_port, QN => n_2070);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n2490, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_29_port, QN => n_2071);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n2489, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_28_port, QN => n_2072);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n2488, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_27_port, QN => n_2073);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n2487, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_26_port, QN => n_2074);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n2486, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_25_port, QN => n_2075);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n2485, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_24_port, QN => n_2076);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n2484, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_23_port, QN => n_2077);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n2483, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_22_port, QN => n_2078);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n2482, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_21_port, QN => n_2079);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n2481, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_20_port, QN => n_2080);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n2480, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_19_port, QN => n_2081);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n2479, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_18_port, QN => n_2082);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n2478, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_17_port, QN => n_2083);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n2477, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_16_port, QN => n_2084);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n2476, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_15_port, QN => n_2085);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n2475, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_14_port, QN => n_2086);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n2474, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_13_port, QN => n_2087);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n2473, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_12_port, QN => n_2088);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n2472, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_11_port, QN => n_2089);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n2471, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_10_port, QN => n_2090);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n2470, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_9_port, QN => n_2091);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n2469, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_8_port, QN => n_2092);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n2468, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_7_port, QN => n_2093);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n2467, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_6_port, QN => n_2094);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n2466, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_5_port, QN => n_2095);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n2465, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_4_port, QN => n_2096);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n2464, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_3_port, QN => n_2097);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n2463, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_2_port, QN => n_2098);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n2462, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_1_port, QN => n_2099);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n2461, CK => CLK, RN => 
                           RESET, Q => REGISTERS_29_0_port, QN => n_2100);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n2460, CK => CLK, RN => 
                           RESET, Q => n_2101, QN => n102);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n2459, CK => CLK, RN => 
                           RESET, Q => n_2102, QN => n101);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n2458, CK => CLK, RN => 
                           RESET, Q => n_2103, QN => n100);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n2457, CK => CLK, RN => 
                           RESET, Q => n_2104, QN => n99);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n2456, CK => CLK, RN => 
                           RESET, Q => n_2105, QN => n98);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n2455, CK => CLK, RN => 
                           RESET, Q => n_2106, QN => n97);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n2454, CK => CLK, RN => 
                           RESET, Q => n_2107, QN => n96);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n2453, CK => CLK, RN => 
                           RESET, Q => n_2108, QN => n95);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n2452, CK => CLK, RN => 
                           RESET, Q => n_2109, QN => n94);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n2451, CK => CLK, RN => 
                           RESET, Q => n_2110, QN => n93);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n2450, CK => CLK, RN => 
                           RESET, Q => n_2111, QN => n92);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n2449, CK => CLK, RN => 
                           RESET, Q => n_2112, QN => n91);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n2448, CK => CLK, RN => 
                           RESET, Q => n_2113, QN => n90);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n2447, CK => CLK, RN => 
                           RESET, Q => n_2114, QN => n89);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n2446, CK => CLK, RN => 
                           RESET, Q => n_2115, QN => n88);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n2445, CK => CLK, RN => 
                           RESET, Q => n_2116, QN => n87);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n2444, CK => CLK, RN => 
                           RESET, Q => n_2117, QN => n86);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n2443, CK => CLK, RN => 
                           RESET, Q => n_2118, QN => n85);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n2442, CK => CLK, RN => 
                           RESET, Q => n_2119, QN => n84);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n2441, CK => CLK, RN => 
                           RESET, Q => n_2120, QN => n83);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n2440, CK => CLK, RN => 
                           RESET, Q => n_2121, QN => n82);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n2439, CK => CLK, RN => 
                           RESET, Q => n_2122, QN => n81);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n2438, CK => CLK, RN => 
                           RESET, Q => n_2123, QN => n80);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n2437, CK => CLK, RN => 
                           RESET, Q => n_2124, QN => n79);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n2436, CK => CLK, RN => 
                           RESET, Q => n_2125, QN => n78);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n2435, CK => CLK, RN => 
                           RESET, Q => n_2126, QN => n77);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n2434, CK => CLK, RN => 
                           RESET, Q => n_2127, QN => n76);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n2433, CK => CLK, RN => 
                           RESET, Q => n_2128, QN => n75);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n2432, CK => CLK, RN => 
                           RESET, Q => n_2129, QN => n74);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n2431, CK => CLK, RN => 
                           RESET, Q => n_2130, QN => n73);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n2430, CK => CLK, RN => 
                           RESET, Q => n_2131, QN => n72);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n2429, CK => CLK, RN => 
                           RESET, Q => n_2132, QN => n71);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n2428, CK => CLK, RN => 
                           RESET, Q => n_2133, QN => n66);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n2427, CK => CLK, RN => 
                           RESET, Q => n_2134, QN => n64);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n2426, CK => CLK, RN => 
                           RESET, Q => n_2135, QN => n62);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n2425, CK => CLK, RN => 
                           RESET, Q => n_2136, QN => n60);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n2424, CK => CLK, RN => 
                           RESET, Q => n_2137, QN => n58);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n2423, CK => CLK, RN => 
                           RESET, Q => n_2138, QN => n56);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n2422, CK => CLK, RN => 
                           RESET, Q => n_2139, QN => n54);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n2421, CK => CLK, RN => 
                           RESET, Q => n_2140, QN => n52);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n2420, CK => CLK, RN => 
                           RESET, Q => n_2141, QN => n50);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n2419, CK => CLK, RN => 
                           RESET, Q => n_2142, QN => n48);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n2418, CK => CLK, RN => 
                           RESET, Q => n_2143, QN => n46);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n2417, CK => CLK, RN => 
                           RESET, Q => n_2144, QN => n44);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n2416, CK => CLK, RN => 
                           RESET, Q => n_2145, QN => n42);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n2415, CK => CLK, RN => 
                           RESET, Q => n_2146, QN => n40);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n2414, CK => CLK, RN => 
                           RESET, Q => n_2147, QN => n38);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n2413, CK => CLK, RN => 
                           RESET, Q => n_2148, QN => n36);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n2412, CK => CLK, RN => 
                           RESET, Q => n_2149, QN => n34);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n2411, CK => CLK, RN => 
                           RESET, Q => n_2150, QN => n32);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n2410, CK => CLK, RN => 
                           RESET, Q => n_2151, QN => n30);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n2409, CK => CLK, RN => 
                           RESET, Q => n_2152, QN => n28);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n2408, CK => CLK, RN => 
                           RESET, Q => n_2153, QN => n26);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n2407, CK => CLK, RN => 
                           RESET, Q => n_2154, QN => n24);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n2406, CK => CLK, RN => 
                           RESET, Q => n_2155, QN => n22);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n2405, CK => CLK, RN => 
                           RESET, Q => n_2156, QN => n20);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n2404, CK => CLK, RN => 
                           RESET, Q => n_2157, QN => n18);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n2403, CK => CLK, RN => 
                           RESET, Q => n_2158, QN => n16);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n2402, CK => CLK, RN => 
                           RESET, Q => n_2159, QN => n14);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n2401, CK => CLK, RN => 
                           RESET, Q => n_2160, QN => n12);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n2400, CK => CLK, RN => 
                           RESET, Q => n_2161, QN => n10);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n2399, CK => CLK, RN => 
                           RESET, Q => n_2162, QN => n8);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n2398, CK => CLK, RN => 
                           RESET, Q => n_2163, QN => n6);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n2397, CK => CLK, RN => 
                           RESET, Q => n_2164, QN => n4);
   OUT1_reg_31_inst : DLH_X1 port map( G => N286, D => N318, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => N286, D => N317, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => N286, D => N316, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => N286, D => N315, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => N286, D => N314, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => N286, D => N313, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => N286, D => N312, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => N286, D => N311, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => N286, D => N310, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => N286, D => N309, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => N286, D => N308, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => N286, D => N307, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => N286, D => N306, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => N286, D => N305, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => N286, D => N304, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => N286, D => N303, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => N286, D => N302, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => N286, D => N301, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => N286, D => N300, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => N286, D => N299, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => N286, D => N298, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => N286, D => N297, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => N286, D => N296, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => N286, D => N295, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => N286, D => N294, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => N286, D => N293, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => N286, D => N292, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => N286, D => N291, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => N286, D => N290, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => N286, D => N289, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => N286, D => N288, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => N286, D => N287, Q => OUT1(0));
   OUT2_reg_31_inst : DLH_X1 port map( G => N319, D => N351, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => N319, D => N350, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => N319, D => N349, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => N319, D => N348, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => N319, D => N347, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => N319, D => N346, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => N319, D => N345, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => N319, D => N344, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => N319, D => N343, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => N319, D => N342, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => N319, D => N341, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => N319, D => N340, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => N319, D => N339, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => N319, D => N338, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => N319, D => N337, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => N319, D => N336, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => N319, D => N335, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => N319, D => N334, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => N319, D => N333, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => N319, D => N332, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => N319, D => N331, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => N319, D => N330, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => N319, D => N329, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => N319, D => N328, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => N319, D => N327, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => N319, D => N326, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => N319, D => N325, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => N319, D => N324, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => N319, D => N323, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => N319, D => N322, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => N319, D => N321, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => N319, D => N320, Q => OUT2(0));
   U3 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => n2397)
                           ;
   U4 : OAI22_X1 port map( A1 => n1, A2 => n5, B1 => n3, B2 => n6, ZN => n2398)
                           ;
   U5 : OAI22_X1 port map( A1 => n1, A2 => n7, B1 => n3, B2 => n8, ZN => n2399)
                           ;
   U6 : OAI22_X1 port map( A1 => n1, A2 => n9, B1 => n3, B2 => n10, ZN => n2400
                           );
   U7 : OAI22_X1 port map( A1 => n1, A2 => n11, B1 => n3, B2 => n12, ZN => 
                           n2401);
   U8 : OAI22_X1 port map( A1 => n1, A2 => n13, B1 => n3, B2 => n14, ZN => 
                           n2402);
   U9 : OAI22_X1 port map( A1 => n1, A2 => n15, B1 => n3, B2 => n16, ZN => 
                           n2403);
   U10 : OAI22_X1 port map( A1 => n1, A2 => n17, B1 => n3, B2 => n18, ZN => 
                           n2404);
   U11 : OAI22_X1 port map( A1 => n1, A2 => n19, B1 => n3, B2 => n20, ZN => 
                           n2405);
   U12 : OAI22_X1 port map( A1 => n1, A2 => n21, B1 => n3, B2 => n22, ZN => 
                           n2406);
   U13 : OAI22_X1 port map( A1 => n1, A2 => n23, B1 => n3, B2 => n24, ZN => 
                           n2407);
   U14 : OAI22_X1 port map( A1 => n1, A2 => n25, B1 => n3, B2 => n26, ZN => 
                           n2408);
   U15 : OAI22_X1 port map( A1 => n1, A2 => n27, B1 => n3, B2 => n28, ZN => 
                           n2409);
   U16 : OAI22_X1 port map( A1 => n1, A2 => n29, B1 => n3, B2 => n30, ZN => 
                           n2410);
   U17 : OAI22_X1 port map( A1 => n1, A2 => n31, B1 => n3, B2 => n32, ZN => 
                           n2411);
   U18 : OAI22_X1 port map( A1 => n1, A2 => n33, B1 => n3, B2 => n34, ZN => 
                           n2412);
   U19 : OAI22_X1 port map( A1 => n1, A2 => n35, B1 => n3, B2 => n36, ZN => 
                           n2413);
   U20 : OAI22_X1 port map( A1 => n1, A2 => n37, B1 => n3, B2 => n38, ZN => 
                           n2414);
   U21 : OAI22_X1 port map( A1 => n1, A2 => n39, B1 => n3, B2 => n40, ZN => 
                           n2415);
   U22 : OAI22_X1 port map( A1 => n1, A2 => n41, B1 => n3, B2 => n42, ZN => 
                           n2416);
   U23 : OAI22_X1 port map( A1 => n1, A2 => n43, B1 => n3, B2 => n44, ZN => 
                           n2417);
   U24 : OAI22_X1 port map( A1 => n1, A2 => n45, B1 => n3, B2 => n46, ZN => 
                           n2418);
   U25 : OAI22_X1 port map( A1 => n1, A2 => n47, B1 => n3, B2 => n48, ZN => 
                           n2419);
   U26 : OAI22_X1 port map( A1 => n1, A2 => n49, B1 => n3, B2 => n50, ZN => 
                           n2420);
   U27 : OAI22_X1 port map( A1 => n1, A2 => n51, B1 => n3, B2 => n52, ZN => 
                           n2421);
   U28 : OAI22_X1 port map( A1 => n1, A2 => n53, B1 => n3, B2 => n54, ZN => 
                           n2422);
   U29 : OAI22_X1 port map( A1 => n1, A2 => n55, B1 => n3, B2 => n56, ZN => 
                           n2423);
   U30 : OAI22_X1 port map( A1 => n1, A2 => n57, B1 => n3, B2 => n58, ZN => 
                           n2424);
   U31 : OAI22_X1 port map( A1 => n1, A2 => n59, B1 => n3, B2 => n60, ZN => 
                           n2425);
   U32 : OAI22_X1 port map( A1 => n1, A2 => n61, B1 => n3, B2 => n62, ZN => 
                           n2426);
   U33 : OAI22_X1 port map( A1 => n1, A2 => n63, B1 => n3, B2 => n64, ZN => 
                           n2427);
   U34 : OAI22_X1 port map( A1 => n1, A2 => n65, B1 => n3, B2 => n66, ZN => 
                           n2428);
   U37 : OAI22_X1 port map( A1 => n2, A2 => n69, B1 => n70, B2 => n71, ZN => 
                           n2429);
   U38 : OAI22_X1 port map( A1 => n5, A2 => n69, B1 => n70, B2 => n72, ZN => 
                           n2430);
   U39 : OAI22_X1 port map( A1 => n7, A2 => n69, B1 => n70, B2 => n73, ZN => 
                           n2431);
   U40 : OAI22_X1 port map( A1 => n9, A2 => n69, B1 => n70, B2 => n74, ZN => 
                           n2432);
   U41 : OAI22_X1 port map( A1 => n11, A2 => n69, B1 => n70, B2 => n75, ZN => 
                           n2433);
   U42 : OAI22_X1 port map( A1 => n13, A2 => n69, B1 => n70, B2 => n76, ZN => 
                           n2434);
   U43 : OAI22_X1 port map( A1 => n15, A2 => n69, B1 => n70, B2 => n77, ZN => 
                           n2435);
   U44 : OAI22_X1 port map( A1 => n17, A2 => n69, B1 => n70, B2 => n78, ZN => 
                           n2436);
   U45 : OAI22_X1 port map( A1 => n19, A2 => n69, B1 => n70, B2 => n79, ZN => 
                           n2437);
   U46 : OAI22_X1 port map( A1 => n21, A2 => n69, B1 => n70, B2 => n80, ZN => 
                           n2438);
   U47 : OAI22_X1 port map( A1 => n23, A2 => n69, B1 => n70, B2 => n81, ZN => 
                           n2439);
   U48 : OAI22_X1 port map( A1 => n25, A2 => n69, B1 => n70, B2 => n82, ZN => 
                           n2440);
   U49 : OAI22_X1 port map( A1 => n27, A2 => n69, B1 => n70, B2 => n83, ZN => 
                           n2441);
   U50 : OAI22_X1 port map( A1 => n29, A2 => n69, B1 => n70, B2 => n84, ZN => 
                           n2442);
   U51 : OAI22_X1 port map( A1 => n31, A2 => n69, B1 => n70, B2 => n85, ZN => 
                           n2443);
   U52 : OAI22_X1 port map( A1 => n33, A2 => n69, B1 => n70, B2 => n86, ZN => 
                           n2444);
   U53 : OAI22_X1 port map( A1 => n35, A2 => n69, B1 => n70, B2 => n87, ZN => 
                           n2445);
   U54 : OAI22_X1 port map( A1 => n37, A2 => n69, B1 => n70, B2 => n88, ZN => 
                           n2446);
   U55 : OAI22_X1 port map( A1 => n39, A2 => n69, B1 => n70, B2 => n89, ZN => 
                           n2447);
   U56 : OAI22_X1 port map( A1 => n41, A2 => n69, B1 => n70, B2 => n90, ZN => 
                           n2448);
   U57 : OAI22_X1 port map( A1 => n43, A2 => n69, B1 => n70, B2 => n91, ZN => 
                           n2449);
   U58 : OAI22_X1 port map( A1 => n45, A2 => n69, B1 => n70, B2 => n92, ZN => 
                           n2450);
   U59 : OAI22_X1 port map( A1 => n47, A2 => n69, B1 => n70, B2 => n93, ZN => 
                           n2451);
   U60 : OAI22_X1 port map( A1 => n49, A2 => n69, B1 => n70, B2 => n94, ZN => 
                           n2452);
   U61 : OAI22_X1 port map( A1 => n51, A2 => n69, B1 => n70, B2 => n95, ZN => 
                           n2453);
   U62 : OAI22_X1 port map( A1 => n53, A2 => n69, B1 => n70, B2 => n96, ZN => 
                           n2454);
   U63 : OAI22_X1 port map( A1 => n55, A2 => n69, B1 => n70, B2 => n97, ZN => 
                           n2455);
   U64 : OAI22_X1 port map( A1 => n57, A2 => n69, B1 => n70, B2 => n98, ZN => 
                           n2456);
   U65 : OAI22_X1 port map( A1 => n59, A2 => n69, B1 => n70, B2 => n99, ZN => 
                           n2457);
   U66 : OAI22_X1 port map( A1 => n61, A2 => n69, B1 => n70, B2 => n100, ZN => 
                           n2458);
   U67 : OAI22_X1 port map( A1 => n63, A2 => n69, B1 => n70, B2 => n101, ZN => 
                           n2459);
   U68 : OAI22_X1 port map( A1 => n65, A2 => n69, B1 => n70, B2 => n102, ZN => 
                           n2460);
   U71 : INV_X1 port map( A => n104, ZN => n2461);
   U72 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_0_port, ZN => n104);
   U73 : INV_X1 port map( A => n107, ZN => n2462);
   U74 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_1_port, ZN => n107);
   U75 : INV_X1 port map( A => n108, ZN => n2463);
   U76 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_2_port, ZN => n108);
   U77 : INV_X1 port map( A => n109, ZN => n2464);
   U78 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_3_port, ZN => n109);
   U79 : INV_X1 port map( A => n110, ZN => n2465);
   U80 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_4_port, ZN => n110);
   U81 : INV_X1 port map( A => n111, ZN => n2466);
   U82 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_5_port, ZN => n111);
   U83 : INV_X1 port map( A => n112, ZN => n2467);
   U84 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_6_port, ZN => n112);
   U85 : INV_X1 port map( A => n113, ZN => n2468);
   U86 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_7_port, ZN => n113);
   U87 : INV_X1 port map( A => n114, ZN => n2469);
   U88 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_8_port, ZN => n114);
   U89 : INV_X1 port map( A => n115, ZN => n2470);
   U90 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_9_port, ZN => n115);
   U91 : INV_X1 port map( A => n116, ZN => n2471);
   U92 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_10_port, ZN => n116);
   U93 : INV_X1 port map( A => n117, ZN => n2472);
   U94 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_11_port, ZN => n117);
   U95 : INV_X1 port map( A => n118, ZN => n2473);
   U96 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_12_port, ZN => n118);
   U97 : INV_X1 port map( A => n119, ZN => n2474);
   U98 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_13_port, ZN => n119);
   U99 : INV_X1 port map( A => n120, ZN => n2475);
   U100 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_14_port, ZN => n120);
   U101 : INV_X1 port map( A => n121, ZN => n2476);
   U102 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_15_port, ZN => n121);
   U103 : INV_X1 port map( A => n122, ZN => n2477);
   U104 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_16_port, ZN => n122);
   U105 : INV_X1 port map( A => n123, ZN => n2478);
   U106 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_17_port, ZN => n123);
   U107 : INV_X1 port map( A => n124, ZN => n2479);
   U108 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_18_port, ZN => n124);
   U109 : INV_X1 port map( A => n125, ZN => n2480);
   U110 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_19_port, ZN => n125);
   U111 : INV_X1 port map( A => n126, ZN => n2481);
   U112 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_20_port, ZN => n126);
   U113 : INV_X1 port map( A => n127, ZN => n2482);
   U114 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_21_port, ZN => n127);
   U115 : INV_X1 port map( A => n128, ZN => n2483);
   U116 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_22_port, ZN => n128);
   U117 : INV_X1 port map( A => n129, ZN => n2484);
   U118 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_23_port, ZN => n129);
   U119 : INV_X1 port map( A => n130, ZN => n2485);
   U120 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_24_port, ZN => n130);
   U121 : INV_X1 port map( A => n131, ZN => n2486);
   U122 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_25_port, ZN => n131);
   U123 : INV_X1 port map( A => n132, ZN => n2487);
   U124 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_26_port, ZN => n132);
   U125 : INV_X1 port map( A => n133, ZN => n2488);
   U126 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_27_port, ZN => n133);
   U127 : INV_X1 port map( A => n134, ZN => n2489);
   U128 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_28_port, ZN => n134);
   U129 : INV_X1 port map( A => n135, ZN => n2490);
   U130 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_29_port, ZN => n135);
   U131 : INV_X1 port map( A => n136, ZN => n2491);
   U132 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_30_port, ZN => n136);
   U133 : INV_X1 port map( A => n137, ZN => n2492);
   U134 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n105, B1 => n106, B2 => 
                           REGISTERS_29_31_port, ZN => n137);
   U137 : INV_X1 port map( A => n139, ZN => n2493);
   U138 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_0_port, ZN => n139);
   U139 : INV_X1 port map( A => n142, ZN => n2494);
   U140 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_1_port, ZN => n142);
   U141 : INV_X1 port map( A => n143, ZN => n2495);
   U142 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_2_port, ZN => n143);
   U143 : INV_X1 port map( A => n144, ZN => n2496);
   U144 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_3_port, ZN => n144);
   U145 : INV_X1 port map( A => n145, ZN => n2497);
   U146 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_4_port, ZN => n145);
   U147 : INV_X1 port map( A => n146, ZN => n2498);
   U148 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_5_port, ZN => n146);
   U149 : INV_X1 port map( A => n147, ZN => n2499);
   U150 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_6_port, ZN => n147);
   U151 : INV_X1 port map( A => n148, ZN => n2500);
   U152 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_7_port, ZN => n148);
   U153 : INV_X1 port map( A => n149, ZN => n2501);
   U154 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_8_port, ZN => n149);
   U155 : INV_X1 port map( A => n150, ZN => n2502);
   U156 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_9_port, ZN => n150);
   U157 : INV_X1 port map( A => n151, ZN => n2503);
   U158 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_10_port, ZN => n151);
   U159 : INV_X1 port map( A => n152, ZN => n2504);
   U160 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_11_port, ZN => n152);
   U161 : INV_X1 port map( A => n153, ZN => n2505);
   U162 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_12_port, ZN => n153);
   U163 : INV_X1 port map( A => n154, ZN => n2506);
   U164 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_13_port, ZN => n154);
   U165 : INV_X1 port map( A => n155, ZN => n2507);
   U166 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_14_port, ZN => n155);
   U167 : INV_X1 port map( A => n156, ZN => n2508);
   U168 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_15_port, ZN => n156);
   U169 : INV_X1 port map( A => n157, ZN => n2509);
   U170 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_16_port, ZN => n157);
   U171 : INV_X1 port map( A => n158, ZN => n2510);
   U172 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_17_port, ZN => n158);
   U173 : INV_X1 port map( A => n159, ZN => n2511);
   U174 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_18_port, ZN => n159);
   U175 : INV_X1 port map( A => n160, ZN => n2512);
   U176 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_19_port, ZN => n160);
   U177 : INV_X1 port map( A => n161, ZN => n2513);
   U178 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_20_port, ZN => n161);
   U179 : INV_X1 port map( A => n162, ZN => n2514);
   U180 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_21_port, ZN => n162);
   U181 : INV_X1 port map( A => n163, ZN => n2515);
   U182 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_22_port, ZN => n163);
   U183 : INV_X1 port map( A => n164, ZN => n2516);
   U184 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_23_port, ZN => n164);
   U185 : INV_X1 port map( A => n165, ZN => n2517);
   U186 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_24_port, ZN => n165);
   U187 : INV_X1 port map( A => n166, ZN => n2518);
   U188 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_25_port, ZN => n166);
   U189 : INV_X1 port map( A => n167, ZN => n2519);
   U190 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_26_port, ZN => n167);
   U191 : INV_X1 port map( A => n168, ZN => n2520);
   U192 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_27_port, ZN => n168);
   U193 : INV_X1 port map( A => n169, ZN => n2521);
   U194 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_28_port, ZN => n169);
   U195 : INV_X1 port map( A => n170, ZN => n2522);
   U196 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_29_port, ZN => n170);
   U197 : INV_X1 port map( A => n171, ZN => n2523);
   U198 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_30_port, ZN => n171);
   U199 : INV_X1 port map( A => n172, ZN => n2524);
   U200 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n140, B1 => n141, B2 => 
                           REGISTERS_28_31_port, ZN => n172);
   U203 : INV_X1 port map( A => n174, ZN => n2525);
   U204 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_0_port, ZN => n174);
   U205 : INV_X1 port map( A => n177, ZN => n2526);
   U206 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_1_port, ZN => n177);
   U207 : INV_X1 port map( A => n178, ZN => n2527);
   U208 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_2_port, ZN => n178);
   U209 : INV_X1 port map( A => n179, ZN => n2528);
   U210 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_3_port, ZN => n179);
   U211 : INV_X1 port map( A => n180, ZN => n2529);
   U212 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_4_port, ZN => n180);
   U213 : INV_X1 port map( A => n181, ZN => n2530);
   U214 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_5_port, ZN => n181);
   U215 : INV_X1 port map( A => n182, ZN => n2531);
   U216 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_6_port, ZN => n182);
   U217 : INV_X1 port map( A => n183, ZN => n2532);
   U218 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_7_port, ZN => n183);
   U219 : INV_X1 port map( A => n184, ZN => n2533);
   U220 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_8_port, ZN => n184);
   U221 : INV_X1 port map( A => n185, ZN => n2534);
   U222 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_9_port, ZN => n185);
   U223 : INV_X1 port map( A => n186, ZN => n2535);
   U224 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_10_port, ZN => n186);
   U225 : INV_X1 port map( A => n187, ZN => n2536);
   U226 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_11_port, ZN => n187);
   U227 : INV_X1 port map( A => n188, ZN => n2537);
   U228 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_12_port, ZN => n188);
   U229 : INV_X1 port map( A => n189, ZN => n2538);
   U230 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_13_port, ZN => n189);
   U231 : INV_X1 port map( A => n190, ZN => n2539);
   U232 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_14_port, ZN => n190);
   U233 : INV_X1 port map( A => n191, ZN => n2540);
   U234 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_15_port, ZN => n191);
   U235 : INV_X1 port map( A => n192, ZN => n2541);
   U236 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_16_port, ZN => n192);
   U237 : INV_X1 port map( A => n193, ZN => n2542);
   U238 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_17_port, ZN => n193);
   U239 : INV_X1 port map( A => n194, ZN => n2543);
   U240 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_18_port, ZN => n194);
   U241 : INV_X1 port map( A => n195, ZN => n2544);
   U242 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_19_port, ZN => n195);
   U243 : INV_X1 port map( A => n196, ZN => n2545);
   U244 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_20_port, ZN => n196);
   U245 : INV_X1 port map( A => n197, ZN => n2546);
   U246 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_21_port, ZN => n197);
   U247 : INV_X1 port map( A => n198, ZN => n2547);
   U248 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_22_port, ZN => n198);
   U249 : INV_X1 port map( A => n199, ZN => n2548);
   U250 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_23_port, ZN => n199);
   U251 : INV_X1 port map( A => n200, ZN => n2549);
   U252 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_24_port, ZN => n200);
   U253 : INV_X1 port map( A => n201, ZN => n2550);
   U254 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_25_port, ZN => n201);
   U255 : INV_X1 port map( A => n202, ZN => n2551);
   U256 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_26_port, ZN => n202);
   U257 : INV_X1 port map( A => n203, ZN => n2552);
   U258 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_27_port, ZN => n203);
   U259 : INV_X1 port map( A => n204, ZN => n2553);
   U260 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_28_port, ZN => n204);
   U261 : INV_X1 port map( A => n205, ZN => n2554);
   U262 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_29_port, ZN => n205);
   U263 : INV_X1 port map( A => n206, ZN => n2555);
   U264 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_30_port, ZN => n206);
   U265 : INV_X1 port map( A => n207, ZN => n2556);
   U266 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n175, B1 => n176, B2 => 
                           REGISTERS_27_31_port, ZN => n207);
   U269 : INV_X1 port map( A => n209, ZN => n2557);
   U270 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_0_port, ZN => n209);
   U271 : INV_X1 port map( A => n212, ZN => n2558);
   U272 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_1_port, ZN => n212);
   U273 : INV_X1 port map( A => n213, ZN => n2559);
   U274 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_2_port, ZN => n213);
   U275 : INV_X1 port map( A => n214, ZN => n2560);
   U276 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_3_port, ZN => n214);
   U277 : INV_X1 port map( A => n215, ZN => n2561);
   U278 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_4_port, ZN => n215);
   U279 : INV_X1 port map( A => n216, ZN => n2562);
   U280 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_5_port, ZN => n216);
   U281 : INV_X1 port map( A => n217, ZN => n2563);
   U282 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_6_port, ZN => n217);
   U283 : INV_X1 port map( A => n218, ZN => n2564);
   U284 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_7_port, ZN => n218);
   U285 : INV_X1 port map( A => n219, ZN => n2565);
   U286 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_8_port, ZN => n219);
   U287 : INV_X1 port map( A => n220, ZN => n2566);
   U288 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_9_port, ZN => n220);
   U289 : INV_X1 port map( A => n221, ZN => n2567);
   U290 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_10_port, ZN => n221);
   U291 : INV_X1 port map( A => n222, ZN => n2568);
   U292 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_11_port, ZN => n222);
   U293 : INV_X1 port map( A => n223, ZN => n2569);
   U294 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_12_port, ZN => n223);
   U295 : INV_X1 port map( A => n224, ZN => n2570);
   U296 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_13_port, ZN => n224);
   U297 : INV_X1 port map( A => n225, ZN => n2571);
   U298 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_14_port, ZN => n225);
   U299 : INV_X1 port map( A => n226, ZN => n2572);
   U300 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_15_port, ZN => n226);
   U301 : INV_X1 port map( A => n227, ZN => n2573);
   U302 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_16_port, ZN => n227);
   U303 : INV_X1 port map( A => n228, ZN => n2574);
   U304 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_17_port, ZN => n228);
   U305 : INV_X1 port map( A => n229, ZN => n2575);
   U306 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_18_port, ZN => n229);
   U307 : INV_X1 port map( A => n230, ZN => n2576);
   U308 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_19_port, ZN => n230);
   U309 : INV_X1 port map( A => n231, ZN => n2577);
   U310 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_20_port, ZN => n231);
   U311 : INV_X1 port map( A => n232, ZN => n2578);
   U312 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_21_port, ZN => n232);
   U313 : INV_X1 port map( A => n233, ZN => n2579);
   U314 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_22_port, ZN => n233);
   U315 : INV_X1 port map( A => n234, ZN => n2580);
   U316 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_23_port, ZN => n234);
   U317 : INV_X1 port map( A => n235, ZN => n2581);
   U318 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_24_port, ZN => n235);
   U319 : INV_X1 port map( A => n236, ZN => n2582);
   U320 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_25_port, ZN => n236);
   U321 : INV_X1 port map( A => n237, ZN => n2583);
   U322 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_26_port, ZN => n237);
   U323 : INV_X1 port map( A => n238, ZN => n2584);
   U324 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_27_port, ZN => n238);
   U325 : INV_X1 port map( A => n239, ZN => n2585);
   U326 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_28_port, ZN => n239);
   U327 : INV_X1 port map( A => n240, ZN => n2586);
   U328 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_29_port, ZN => n240);
   U329 : INV_X1 port map( A => n241, ZN => n2587);
   U330 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_30_port, ZN => n241);
   U331 : INV_X1 port map( A => n242, ZN => n2588);
   U332 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n210, B1 => n211, B2 => 
                           REGISTERS_26_31_port, ZN => n242);
   U335 : OAI22_X1 port map( A1 => n2, A2 => n244, B1 => n245, B2 => n246, ZN 
                           => n2589);
   U336 : OAI22_X1 port map( A1 => n5, A2 => n244, B1 => n245, B2 => n247, ZN 
                           => n2590);
   U337 : OAI22_X1 port map( A1 => n7, A2 => n244, B1 => n245, B2 => n248, ZN 
                           => n2591);
   U338 : OAI22_X1 port map( A1 => n9, A2 => n244, B1 => n245, B2 => n249, ZN 
                           => n2592);
   U339 : OAI22_X1 port map( A1 => n11, A2 => n244, B1 => n245, B2 => n250, ZN 
                           => n2593);
   U340 : OAI22_X1 port map( A1 => n13, A2 => n244, B1 => n245, B2 => n251, ZN 
                           => n2594);
   U341 : OAI22_X1 port map( A1 => n15, A2 => n244, B1 => n245, B2 => n252, ZN 
                           => n2595);
   U342 : OAI22_X1 port map( A1 => n17, A2 => n244, B1 => n245, B2 => n253, ZN 
                           => n2596);
   U343 : OAI22_X1 port map( A1 => n19, A2 => n244, B1 => n245, B2 => n254, ZN 
                           => n2597);
   U344 : OAI22_X1 port map( A1 => n21, A2 => n244, B1 => n245, B2 => n255, ZN 
                           => n2598);
   U345 : OAI22_X1 port map( A1 => n23, A2 => n244, B1 => n245, B2 => n256, ZN 
                           => n2599);
   U346 : OAI22_X1 port map( A1 => n25, A2 => n244, B1 => n245, B2 => n257, ZN 
                           => n2600);
   U347 : OAI22_X1 port map( A1 => n27, A2 => n244, B1 => n245, B2 => n258, ZN 
                           => n2601);
   U348 : OAI22_X1 port map( A1 => n29, A2 => n244, B1 => n245, B2 => n259, ZN 
                           => n2602);
   U349 : OAI22_X1 port map( A1 => n31, A2 => n244, B1 => n245, B2 => n260, ZN 
                           => n2603);
   U350 : OAI22_X1 port map( A1 => n33, A2 => n244, B1 => n245, B2 => n261, ZN 
                           => n2604);
   U351 : OAI22_X1 port map( A1 => n35, A2 => n244, B1 => n245, B2 => n262, ZN 
                           => n2605);
   U352 : OAI22_X1 port map( A1 => n37, A2 => n244, B1 => n245, B2 => n263, ZN 
                           => n2606);
   U353 : OAI22_X1 port map( A1 => n39, A2 => n244, B1 => n245, B2 => n264, ZN 
                           => n2607);
   U354 : OAI22_X1 port map( A1 => n41, A2 => n244, B1 => n245, B2 => n265, ZN 
                           => n2608);
   U355 : OAI22_X1 port map( A1 => n43, A2 => n244, B1 => n245, B2 => n266, ZN 
                           => n2609);
   U356 : OAI22_X1 port map( A1 => n45, A2 => n244, B1 => n245, B2 => n267, ZN 
                           => n2610);
   U357 : OAI22_X1 port map( A1 => n47, A2 => n244, B1 => n245, B2 => n268, ZN 
                           => n2611);
   U358 : OAI22_X1 port map( A1 => n49, A2 => n244, B1 => n245, B2 => n269, ZN 
                           => n2612);
   U359 : OAI22_X1 port map( A1 => n51, A2 => n244, B1 => n245, B2 => n270, ZN 
                           => n2613);
   U360 : OAI22_X1 port map( A1 => n53, A2 => n244, B1 => n245, B2 => n271, ZN 
                           => n2614);
   U361 : OAI22_X1 port map( A1 => n55, A2 => n244, B1 => n245, B2 => n272, ZN 
                           => n2615);
   U362 : OAI22_X1 port map( A1 => n57, A2 => n244, B1 => n245, B2 => n273, ZN 
                           => n2616);
   U363 : OAI22_X1 port map( A1 => n59, A2 => n244, B1 => n245, B2 => n274, ZN 
                           => n2617);
   U364 : OAI22_X1 port map( A1 => n61, A2 => n244, B1 => n245, B2 => n275, ZN 
                           => n2618);
   U365 : OAI22_X1 port map( A1 => n63, A2 => n244, B1 => n245, B2 => n276, ZN 
                           => n2619);
   U366 : OAI22_X1 port map( A1 => n65, A2 => n244, B1 => n245, B2 => n277, ZN 
                           => n2620);
   U369 : OAI22_X1 port map( A1 => n2, A2 => n279, B1 => n280, B2 => n281, ZN 
                           => n2621);
   U370 : OAI22_X1 port map( A1 => n5, A2 => n279, B1 => n280, B2 => n282, ZN 
                           => n2622);
   U371 : OAI22_X1 port map( A1 => n7, A2 => n279, B1 => n280, B2 => n283, ZN 
                           => n2623);
   U372 : OAI22_X1 port map( A1 => n9, A2 => n279, B1 => n280, B2 => n284, ZN 
                           => n2624);
   U373 : OAI22_X1 port map( A1 => n11, A2 => n279, B1 => n280, B2 => n285, ZN 
                           => n2625);
   U374 : OAI22_X1 port map( A1 => n13, A2 => n279, B1 => n280, B2 => n286_port
                           , ZN => n2626);
   U375 : OAI22_X1 port map( A1 => n15, A2 => n279, B1 => n280, B2 => n287_port
                           , ZN => n2627);
   U376 : OAI22_X1 port map( A1 => n17, A2 => n279, B1 => n280, B2 => n288_port
                           , ZN => n2628);
   U377 : OAI22_X1 port map( A1 => n19, A2 => n279, B1 => n280, B2 => n289_port
                           , ZN => n2629);
   U378 : OAI22_X1 port map( A1 => n21, A2 => n279, B1 => n280, B2 => n290_port
                           , ZN => n2630);
   U379 : OAI22_X1 port map( A1 => n23, A2 => n279, B1 => n280, B2 => n291_port
                           , ZN => n2631);
   U380 : OAI22_X1 port map( A1 => n25, A2 => n279, B1 => n280, B2 => n292_port
                           , ZN => n2632);
   U381 : OAI22_X1 port map( A1 => n27, A2 => n279, B1 => n280, B2 => n293_port
                           , ZN => n2633);
   U382 : OAI22_X1 port map( A1 => n29, A2 => n279, B1 => n280, B2 => n294_port
                           , ZN => n2634);
   U383 : OAI22_X1 port map( A1 => n31, A2 => n279, B1 => n280, B2 => n295_port
                           , ZN => n2635);
   U384 : OAI22_X1 port map( A1 => n33, A2 => n279, B1 => n280, B2 => n296_port
                           , ZN => n2636);
   U385 : OAI22_X1 port map( A1 => n35, A2 => n279, B1 => n280, B2 => n297_port
                           , ZN => n2637);
   U386 : OAI22_X1 port map( A1 => n37, A2 => n279, B1 => n280, B2 => n298_port
                           , ZN => n2638);
   U387 : OAI22_X1 port map( A1 => n39, A2 => n279, B1 => n280, B2 => n299_port
                           , ZN => n2639);
   U388 : OAI22_X1 port map( A1 => n41, A2 => n279, B1 => n280, B2 => n300_port
                           , ZN => n2640);
   U389 : OAI22_X1 port map( A1 => n43, A2 => n279, B1 => n280, B2 => n301_port
                           , ZN => n2641);
   U390 : OAI22_X1 port map( A1 => n45, A2 => n279, B1 => n280, B2 => n302_port
                           , ZN => n2642);
   U391 : OAI22_X1 port map( A1 => n47, A2 => n279, B1 => n280, B2 => n303_port
                           , ZN => n2643);
   U392 : OAI22_X1 port map( A1 => n49, A2 => n279, B1 => n280, B2 => n304_port
                           , ZN => n2644);
   U393 : OAI22_X1 port map( A1 => n51, A2 => n279, B1 => n280, B2 => n305_port
                           , ZN => n2645);
   U394 : OAI22_X1 port map( A1 => n53, A2 => n279, B1 => n280, B2 => n306_port
                           , ZN => n2646);
   U395 : OAI22_X1 port map( A1 => n55, A2 => n279, B1 => n280, B2 => n307_port
                           , ZN => n2647);
   U396 : OAI22_X1 port map( A1 => n57, A2 => n279, B1 => n280, B2 => n308_port
                           , ZN => n2648);
   U397 : OAI22_X1 port map( A1 => n59, A2 => n279, B1 => n280, B2 => n309_port
                           , ZN => n2649);
   U398 : OAI22_X1 port map( A1 => n61, A2 => n279, B1 => n280, B2 => n310_port
                           , ZN => n2650);
   U399 : OAI22_X1 port map( A1 => n63, A2 => n279, B1 => n280, B2 => n311_port
                           , ZN => n2651);
   U400 : OAI22_X1 port map( A1 => n65, A2 => n279, B1 => n280, B2 => n312_port
                           , ZN => n2652);
   U403 : AND3_X1 port map( A1 => ADD_WR(3), A2 => n314_port, A3 => ADD_WR(4), 
                           ZN => n68);
   U404 : INV_X1 port map( A => n315_port, ZN => n2653);
   U405 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_0_port, ZN => n315_port);
   U406 : INV_X1 port map( A => n318_port, ZN => n2654);
   U407 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_1_port, ZN => n318_port);
   U408 : INV_X1 port map( A => n319_port, ZN => n2655);
   U409 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_2_port, ZN => n319_port);
   U410 : INV_X1 port map( A => n320_port, ZN => n2656);
   U411 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_3_port, ZN => n320_port);
   U412 : INV_X1 port map( A => n321_port, ZN => n2657);
   U413 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_4_port, ZN => n321_port);
   U414 : INV_X1 port map( A => n322_port, ZN => n2658);
   U415 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_5_port, ZN => n322_port);
   U416 : INV_X1 port map( A => n323_port, ZN => n2659);
   U417 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_6_port, ZN => n323_port);
   U418 : INV_X1 port map( A => n324_port, ZN => n2660);
   U419 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_7_port, ZN => n324_port);
   U420 : INV_X1 port map( A => n325_port, ZN => n2661);
   U421 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_8_port, ZN => n325_port);
   U422 : INV_X1 port map( A => n326_port, ZN => n2662);
   U423 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n316_port, B1 => n317_port,
                           B2 => REGISTERS_23_9_port, ZN => n326_port);
   U424 : INV_X1 port map( A => n327_port, ZN => n2663);
   U425 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_10_port, ZN => n327_port);
   U426 : INV_X1 port map( A => n328_port, ZN => n2664);
   U427 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_11_port, ZN => n328_port);
   U428 : INV_X1 port map( A => n329_port, ZN => n2665);
   U429 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_12_port, ZN => n329_port);
   U430 : INV_X1 port map( A => n330_port, ZN => n2666);
   U431 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_13_port, ZN => n330_port);
   U432 : INV_X1 port map( A => n331_port, ZN => n2667);
   U433 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_14_port, ZN => n331_port);
   U434 : INV_X1 port map( A => n332_port, ZN => n2668);
   U435 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_15_port, ZN => n332_port);
   U436 : INV_X1 port map( A => n333_port, ZN => n2669);
   U437 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_16_port, ZN => n333_port);
   U438 : INV_X1 port map( A => n334_port, ZN => n2670);
   U439 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_17_port, ZN => n334_port);
   U440 : INV_X1 port map( A => n335_port, ZN => n2671);
   U441 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_18_port, ZN => n335_port);
   U442 : INV_X1 port map( A => n336_port, ZN => n2672);
   U443 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_19_port, ZN => n336_port);
   U444 : INV_X1 port map( A => n337_port, ZN => n2673);
   U445 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_20_port, ZN => n337_port);
   U446 : INV_X1 port map( A => n338_port, ZN => n2674);
   U447 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_21_port, ZN => n338_port);
   U448 : INV_X1 port map( A => n339_port, ZN => n2675);
   U449 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_22_port, ZN => n339_port);
   U450 : INV_X1 port map( A => n340_port, ZN => n2676);
   U451 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_23_port, ZN => n340_port);
   U452 : INV_X1 port map( A => n341_port, ZN => n2677);
   U453 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_24_port, ZN => n341_port);
   U454 : INV_X1 port map( A => n342_port, ZN => n2678);
   U455 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_25_port, ZN => n342_port);
   U456 : INV_X1 port map( A => n343_port, ZN => n2679);
   U457 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_26_port, ZN => n343_port);
   U458 : INV_X1 port map( A => n344_port, ZN => n2680);
   U459 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_27_port, ZN => n344_port);
   U460 : INV_X1 port map( A => n345_port, ZN => n2681);
   U461 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_28_port, ZN => n345_port);
   U462 : INV_X1 port map( A => n346_port, ZN => n2682);
   U463 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_29_port, ZN => n346_port);
   U464 : INV_X1 port map( A => n347_port, ZN => n2683);
   U465 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_30_port, ZN => n347_port);
   U466 : INV_X1 port map( A => n348_port, ZN => n2684);
   U467 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n316_port, B1 => n317_port
                           , B2 => REGISTERS_23_31_port, ZN => n348_port);
   U470 : INV_X1 port map( A => n350_port, ZN => n2685);
   U471 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_0_port, ZN => n350_port);
   U472 : INV_X1 port map( A => n353, ZN => n2686);
   U473 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_1_port, ZN => n353);
   U474 : INV_X1 port map( A => n354, ZN => n2687);
   U475 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_2_port, ZN => n354);
   U476 : INV_X1 port map( A => n355, ZN => n2688);
   U477 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_3_port, ZN => n355);
   U478 : INV_X1 port map( A => n356, ZN => n2689);
   U479 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_4_port, ZN => n356);
   U480 : INV_X1 port map( A => n357, ZN => n2690);
   U481 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_5_port, ZN => n357);
   U482 : INV_X1 port map( A => n358, ZN => n2691);
   U483 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_6_port, ZN => n358);
   U484 : INV_X1 port map( A => n359, ZN => n2692);
   U485 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_7_port, ZN => n359);
   U486 : INV_X1 port map( A => n360, ZN => n2693);
   U487 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_8_port, ZN => n360);
   U488 : INV_X1 port map( A => n361, ZN => n2694);
   U489 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n351_port, B1 => n352_port,
                           B2 => REGISTERS_22_9_port, ZN => n361);
   U490 : INV_X1 port map( A => n362, ZN => n2695);
   U491 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_10_port, ZN => n362);
   U492 : INV_X1 port map( A => n363, ZN => n2696);
   U493 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_11_port, ZN => n363);
   U494 : INV_X1 port map( A => n364, ZN => n2697);
   U495 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_12_port, ZN => n364);
   U496 : INV_X1 port map( A => n365, ZN => n2698);
   U497 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_13_port, ZN => n365);
   U498 : INV_X1 port map( A => n366, ZN => n2699);
   U499 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_14_port, ZN => n366);
   U500 : INV_X1 port map( A => n367, ZN => n2700);
   U501 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_15_port, ZN => n367);
   U502 : INV_X1 port map( A => n368, ZN => n2701);
   U503 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_16_port, ZN => n368);
   U504 : INV_X1 port map( A => n369, ZN => n2702);
   U505 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_17_port, ZN => n369);
   U506 : INV_X1 port map( A => n370, ZN => n2703);
   U507 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_18_port, ZN => n370);
   U508 : INV_X1 port map( A => n371, ZN => n2704);
   U509 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_19_port, ZN => n371);
   U510 : INV_X1 port map( A => n372, ZN => n2705);
   U511 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_20_port, ZN => n372);
   U512 : INV_X1 port map( A => n373, ZN => n2706);
   U513 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_21_port, ZN => n373);
   U514 : INV_X1 port map( A => n374, ZN => n2707);
   U515 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_22_port, ZN => n374);
   U516 : INV_X1 port map( A => n375, ZN => n2708);
   U517 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_23_port, ZN => n375);
   U518 : INV_X1 port map( A => n376, ZN => n2709);
   U519 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_24_port, ZN => n376);
   U520 : INV_X1 port map( A => n377, ZN => n2710);
   U521 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_25_port, ZN => n377);
   U522 : INV_X1 port map( A => n378, ZN => n2711);
   U523 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_26_port, ZN => n378);
   U524 : INV_X1 port map( A => n379, ZN => n2712);
   U525 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_27_port, ZN => n379);
   U526 : INV_X1 port map( A => n380, ZN => n2713);
   U527 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_28_port, ZN => n380);
   U528 : INV_X1 port map( A => n381, ZN => n2714);
   U529 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_29_port, ZN => n381);
   U530 : INV_X1 port map( A => n382, ZN => n2715);
   U531 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_30_port, ZN => n382);
   U532 : INV_X1 port map( A => n383, ZN => n2716);
   U533 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n351_port, B1 => n352_port
                           , B2 => REGISTERS_22_31_port, ZN => n383);
   U536 : OAI22_X1 port map( A1 => n2, A2 => n384, B1 => n385, B2 => n386, ZN 
                           => n2717);
   U537 : OAI22_X1 port map( A1 => n5, A2 => n384, B1 => n385, B2 => n387, ZN 
                           => n2718);
   U538 : OAI22_X1 port map( A1 => n7, A2 => n384, B1 => n385, B2 => n388, ZN 
                           => n2719);
   U539 : OAI22_X1 port map( A1 => n9, A2 => n384, B1 => n385, B2 => n389, ZN 
                           => n2720);
   U540 : OAI22_X1 port map( A1 => n11, A2 => n384, B1 => n385, B2 => n390, ZN 
                           => n2721);
   U541 : OAI22_X1 port map( A1 => n13, A2 => n384, B1 => n385, B2 => n391, ZN 
                           => n2722);
   U542 : OAI22_X1 port map( A1 => n15, A2 => n384, B1 => n385, B2 => n392, ZN 
                           => n2723);
   U543 : OAI22_X1 port map( A1 => n17, A2 => n384, B1 => n385, B2 => n393, ZN 
                           => n2724);
   U544 : OAI22_X1 port map( A1 => n19, A2 => n384, B1 => n385, B2 => n394, ZN 
                           => n2725);
   U545 : OAI22_X1 port map( A1 => n21, A2 => n384, B1 => n385, B2 => n395, ZN 
                           => n2726);
   U546 : OAI22_X1 port map( A1 => n23, A2 => n384, B1 => n385, B2 => n396, ZN 
                           => n2727);
   U547 : OAI22_X1 port map( A1 => n25, A2 => n384, B1 => n385, B2 => n397, ZN 
                           => n2728);
   U548 : OAI22_X1 port map( A1 => n27, A2 => n384, B1 => n385, B2 => n398, ZN 
                           => n2729);
   U549 : OAI22_X1 port map( A1 => n29, A2 => n384, B1 => n385, B2 => n399, ZN 
                           => n2730);
   U550 : OAI22_X1 port map( A1 => n31, A2 => n384, B1 => n385, B2 => n400, ZN 
                           => n2731);
   U551 : OAI22_X1 port map( A1 => n33, A2 => n384, B1 => n385, B2 => n401, ZN 
                           => n2732);
   U552 : OAI22_X1 port map( A1 => n35, A2 => n384, B1 => n385, B2 => n402, ZN 
                           => n2733);
   U553 : OAI22_X1 port map( A1 => n37, A2 => n384, B1 => n385, B2 => n403, ZN 
                           => n2734);
   U554 : OAI22_X1 port map( A1 => n39, A2 => n384, B1 => n385, B2 => n404, ZN 
                           => n2735);
   U555 : OAI22_X1 port map( A1 => n41, A2 => n384, B1 => n385, B2 => n405, ZN 
                           => n2736);
   U556 : OAI22_X1 port map( A1 => n43, A2 => n384, B1 => n385, B2 => n406, ZN 
                           => n2737);
   U557 : OAI22_X1 port map( A1 => n45, A2 => n384, B1 => n385, B2 => n407, ZN 
                           => n2738);
   U558 : OAI22_X1 port map( A1 => n47, A2 => n384, B1 => n385, B2 => n408, ZN 
                           => n2739);
   U559 : OAI22_X1 port map( A1 => n49, A2 => n384, B1 => n385, B2 => n409, ZN 
                           => n2740);
   U560 : OAI22_X1 port map( A1 => n51, A2 => n384, B1 => n385, B2 => n410, ZN 
                           => n2741);
   U561 : OAI22_X1 port map( A1 => n53, A2 => n384, B1 => n385, B2 => n411, ZN 
                           => n2742);
   U562 : OAI22_X1 port map( A1 => n55, A2 => n384, B1 => n385, B2 => n412, ZN 
                           => n2743);
   U563 : OAI22_X1 port map( A1 => n57, A2 => n384, B1 => n385, B2 => n413, ZN 
                           => n2744);
   U564 : OAI22_X1 port map( A1 => n59, A2 => n384, B1 => n385, B2 => n414, ZN 
                           => n2745);
   U565 : OAI22_X1 port map( A1 => n61, A2 => n384, B1 => n385, B2 => n415, ZN 
                           => n2746);
   U566 : OAI22_X1 port map( A1 => n63, A2 => n384, B1 => n385, B2 => n416, ZN 
                           => n2747);
   U567 : OAI22_X1 port map( A1 => n65, A2 => n384, B1 => n385, B2 => n417, ZN 
                           => n2748);
   U570 : OAI22_X1 port map( A1 => n2, A2 => n418, B1 => n419, B2 => n420, ZN 
                           => n2749);
   U571 : OAI22_X1 port map( A1 => n5, A2 => n418, B1 => n419, B2 => n421, ZN 
                           => n2750);
   U572 : OAI22_X1 port map( A1 => n7, A2 => n418, B1 => n419, B2 => n422, ZN 
                           => n2751);
   U573 : OAI22_X1 port map( A1 => n9, A2 => n418, B1 => n419, B2 => n423, ZN 
                           => n2752);
   U574 : OAI22_X1 port map( A1 => n11, A2 => n418, B1 => n419, B2 => n424, ZN 
                           => n2753);
   U575 : OAI22_X1 port map( A1 => n13, A2 => n418, B1 => n419, B2 => n425, ZN 
                           => n2754);
   U576 : OAI22_X1 port map( A1 => n15, A2 => n418, B1 => n419, B2 => n426, ZN 
                           => n2755);
   U577 : OAI22_X1 port map( A1 => n17, A2 => n418, B1 => n419, B2 => n427, ZN 
                           => n2756);
   U578 : OAI22_X1 port map( A1 => n19, A2 => n418, B1 => n419, B2 => n428, ZN 
                           => n2757);
   U579 : OAI22_X1 port map( A1 => n21, A2 => n418, B1 => n419, B2 => n429, ZN 
                           => n2758);
   U580 : OAI22_X1 port map( A1 => n23, A2 => n418, B1 => n419, B2 => n430, ZN 
                           => n2759);
   U581 : OAI22_X1 port map( A1 => n25, A2 => n418, B1 => n419, B2 => n431, ZN 
                           => n2760);
   U582 : OAI22_X1 port map( A1 => n27, A2 => n418, B1 => n419, B2 => n432, ZN 
                           => n2761);
   U583 : OAI22_X1 port map( A1 => n29, A2 => n418, B1 => n419, B2 => n433, ZN 
                           => n2762);
   U584 : OAI22_X1 port map( A1 => n31, A2 => n418, B1 => n419, B2 => n434, ZN 
                           => n2763);
   U585 : OAI22_X1 port map( A1 => n33, A2 => n418, B1 => n419, B2 => n435, ZN 
                           => n2764);
   U586 : OAI22_X1 port map( A1 => n35, A2 => n418, B1 => n419, B2 => n436, ZN 
                           => n2765);
   U587 : OAI22_X1 port map( A1 => n37, A2 => n418, B1 => n419, B2 => n437, ZN 
                           => n2766);
   U588 : OAI22_X1 port map( A1 => n39, A2 => n418, B1 => n419, B2 => n438, ZN 
                           => n2767);
   U589 : OAI22_X1 port map( A1 => n41, A2 => n418, B1 => n419, B2 => n439, ZN 
                           => n2768);
   U590 : OAI22_X1 port map( A1 => n43, A2 => n418, B1 => n419, B2 => n440, ZN 
                           => n2769);
   U591 : OAI22_X1 port map( A1 => n45, A2 => n418, B1 => n419, B2 => n441, ZN 
                           => n2770);
   U592 : OAI22_X1 port map( A1 => n47, A2 => n418, B1 => n419, B2 => n442, ZN 
                           => n2771);
   U593 : OAI22_X1 port map( A1 => n49, A2 => n418, B1 => n419, B2 => n443, ZN 
                           => n2772);
   U594 : OAI22_X1 port map( A1 => n51, A2 => n418, B1 => n419, B2 => n444, ZN 
                           => n2773);
   U595 : OAI22_X1 port map( A1 => n53, A2 => n418, B1 => n419, B2 => n445, ZN 
                           => n2774);
   U596 : OAI22_X1 port map( A1 => n55, A2 => n418, B1 => n419, B2 => n446, ZN 
                           => n2775);
   U597 : OAI22_X1 port map( A1 => n57, A2 => n418, B1 => n419, B2 => n447, ZN 
                           => n2776);
   U598 : OAI22_X1 port map( A1 => n59, A2 => n418, B1 => n419, B2 => n448, ZN 
                           => n2777);
   U599 : OAI22_X1 port map( A1 => n61, A2 => n418, B1 => n419, B2 => n449, ZN 
                           => n2778);
   U600 : OAI22_X1 port map( A1 => n63, A2 => n418, B1 => n419, B2 => n450, ZN 
                           => n2779);
   U601 : OAI22_X1 port map( A1 => n65, A2 => n418, B1 => n419, B2 => n451, ZN 
                           => n2780);
   U604 : INV_X1 port map( A => n452, ZN => n2781);
   U605 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_0_port, ZN => n452);
   U606 : INV_X1 port map( A => n455, ZN => n2782);
   U607 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_1_port, ZN => n455);
   U608 : INV_X1 port map( A => n456, ZN => n2783);
   U609 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_2_port, ZN => n456);
   U610 : INV_X1 port map( A => n457, ZN => n2784);
   U611 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_3_port, ZN => n457);
   U612 : INV_X1 port map( A => n458, ZN => n2785);
   U613 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_4_port, ZN => n458);
   U614 : INV_X1 port map( A => n459, ZN => n2786);
   U615 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_5_port, ZN => n459);
   U616 : INV_X1 port map( A => n460, ZN => n2787);
   U617 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_6_port, ZN => n460);
   U618 : INV_X1 port map( A => n461, ZN => n2788);
   U619 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_7_port, ZN => n461);
   U620 : INV_X1 port map( A => n462, ZN => n2789);
   U621 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_8_port, ZN => n462);
   U622 : INV_X1 port map( A => n463, ZN => n2790);
   U623 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_9_port, ZN => n463);
   U624 : INV_X1 port map( A => n464, ZN => n2791);
   U625 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_10_port, ZN => n464);
   U626 : INV_X1 port map( A => n465, ZN => n2792);
   U627 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_11_port, ZN => n465);
   U628 : INV_X1 port map( A => n466, ZN => n2793);
   U629 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_12_port, ZN => n466);
   U630 : INV_X1 port map( A => n467, ZN => n2794);
   U631 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_13_port, ZN => n467);
   U632 : INV_X1 port map( A => n468, ZN => n2795);
   U633 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_14_port, ZN => n468);
   U634 : INV_X1 port map( A => n469, ZN => n2796);
   U635 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_15_port, ZN => n469);
   U636 : INV_X1 port map( A => n470, ZN => n2797);
   U637 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_16_port, ZN => n470);
   U638 : INV_X1 port map( A => n471, ZN => n2798);
   U639 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_17_port, ZN => n471);
   U640 : INV_X1 port map( A => n472, ZN => n2799);
   U641 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_18_port, ZN => n472);
   U642 : INV_X1 port map( A => n473, ZN => n2800);
   U643 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_19_port, ZN => n473);
   U644 : INV_X1 port map( A => n474, ZN => n2801);
   U645 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_20_port, ZN => n474);
   U646 : INV_X1 port map( A => n475, ZN => n2802);
   U647 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_21_port, ZN => n475);
   U648 : INV_X1 port map( A => n476, ZN => n2803);
   U649 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_22_port, ZN => n476);
   U650 : INV_X1 port map( A => n477, ZN => n2804);
   U651 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_23_port, ZN => n477);
   U652 : INV_X1 port map( A => n478, ZN => n2805);
   U653 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_24_port, ZN => n478);
   U654 : INV_X1 port map( A => n479, ZN => n2806);
   U655 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_25_port, ZN => n479);
   U656 : INV_X1 port map( A => n480, ZN => n2807);
   U657 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_26_port, ZN => n480);
   U658 : INV_X1 port map( A => n481, ZN => n2808);
   U659 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_27_port, ZN => n481);
   U660 : INV_X1 port map( A => n482, ZN => n2809);
   U661 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_28_port, ZN => n482);
   U662 : INV_X1 port map( A => n483, ZN => n2810);
   U663 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_29_port, ZN => n483);
   U664 : INV_X1 port map( A => n484, ZN => n2811);
   U665 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_30_port, ZN => n484);
   U666 : INV_X1 port map( A => n485, ZN => n2812);
   U667 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n453, B1 => n454, B2 => 
                           REGISTERS_19_31_port, ZN => n485);
   U670 : INV_X1 port map( A => n486, ZN => n2813);
   U671 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_0_port, ZN => n486);
   U672 : INV_X1 port map( A => n489, ZN => n2814);
   U673 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_1_port, ZN => n489);
   U674 : INV_X1 port map( A => n490, ZN => n2815);
   U675 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_2_port, ZN => n490);
   U676 : INV_X1 port map( A => n491, ZN => n2816);
   U677 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_3_port, ZN => n491);
   U678 : INV_X1 port map( A => n492, ZN => n2817);
   U679 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_4_port, ZN => n492);
   U680 : INV_X1 port map( A => n493, ZN => n2818);
   U681 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_5_port, ZN => n493);
   U682 : INV_X1 port map( A => n494, ZN => n2819);
   U683 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_6_port, ZN => n494);
   U684 : INV_X1 port map( A => n495, ZN => n2820);
   U685 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_7_port, ZN => n495);
   U686 : INV_X1 port map( A => n496, ZN => n2821);
   U687 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_8_port, ZN => n496);
   U688 : INV_X1 port map( A => n497, ZN => n2822);
   U689 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_9_port, ZN => n497);
   U690 : INV_X1 port map( A => n498, ZN => n2823);
   U691 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_10_port, ZN => n498);
   U692 : INV_X1 port map( A => n499, ZN => n2824);
   U693 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_11_port, ZN => n499);
   U694 : INV_X1 port map( A => n500, ZN => n2825);
   U695 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_12_port, ZN => n500);
   U696 : INV_X1 port map( A => n501, ZN => n2826);
   U697 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_13_port, ZN => n501);
   U698 : INV_X1 port map( A => n502, ZN => n2827);
   U699 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_14_port, ZN => n502);
   U700 : INV_X1 port map( A => n503, ZN => n2828);
   U701 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_15_port, ZN => n503);
   U702 : INV_X1 port map( A => n504, ZN => n2829);
   U703 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_16_port, ZN => n504);
   U704 : INV_X1 port map( A => n505, ZN => n2830);
   U705 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_17_port, ZN => n505);
   U706 : INV_X1 port map( A => n506, ZN => n2831);
   U707 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_18_port, ZN => n506);
   U708 : INV_X1 port map( A => n507, ZN => n2832);
   U709 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_19_port, ZN => n507);
   U710 : INV_X1 port map( A => n508, ZN => n2833);
   U711 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_20_port, ZN => n508);
   U712 : INV_X1 port map( A => n509, ZN => n2834);
   U713 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_21_port, ZN => n509);
   U714 : INV_X1 port map( A => n510, ZN => n2835);
   U715 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_22_port, ZN => n510);
   U716 : INV_X1 port map( A => n511, ZN => n2836);
   U717 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_23_port, ZN => n511);
   U718 : INV_X1 port map( A => n512, ZN => n2837);
   U719 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_24_port, ZN => n512);
   U720 : INV_X1 port map( A => n513, ZN => n2838);
   U721 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_25_port, ZN => n513);
   U722 : INV_X1 port map( A => n514, ZN => n2839);
   U723 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_26_port, ZN => n514);
   U724 : INV_X1 port map( A => n515, ZN => n2840);
   U725 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_27_port, ZN => n515);
   U726 : INV_X1 port map( A => n516, ZN => n2841);
   U727 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_28_port, ZN => n516);
   U728 : INV_X1 port map( A => n517, ZN => n2842);
   U729 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_29_port, ZN => n517);
   U730 : INV_X1 port map( A => n518, ZN => n2843);
   U731 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_30_port, ZN => n518);
   U732 : INV_X1 port map( A => n519, ZN => n2844);
   U733 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n487, B1 => n488, B2 => 
                           REGISTERS_18_31_port, ZN => n519);
   U736 : OAI22_X1 port map( A1 => n2, A2 => n520, B1 => n521, B2 => n522, ZN 
                           => n2845);
   U737 : OAI22_X1 port map( A1 => n5, A2 => n520, B1 => n521, B2 => n523, ZN 
                           => n2846);
   U738 : OAI22_X1 port map( A1 => n7, A2 => n520, B1 => n521, B2 => n524, ZN 
                           => n2847);
   U739 : OAI22_X1 port map( A1 => n9, A2 => n520, B1 => n521, B2 => n525, ZN 
                           => n2848);
   U740 : OAI22_X1 port map( A1 => n11, A2 => n520, B1 => n521, B2 => n526, ZN 
                           => n2849);
   U741 : OAI22_X1 port map( A1 => n13, A2 => n520, B1 => n521, B2 => n527, ZN 
                           => n2850);
   U742 : OAI22_X1 port map( A1 => n15, A2 => n520, B1 => n521, B2 => n528, ZN 
                           => n2851);
   U743 : OAI22_X1 port map( A1 => n17, A2 => n520, B1 => n521, B2 => n529, ZN 
                           => n2852);
   U744 : OAI22_X1 port map( A1 => n19, A2 => n520, B1 => n521, B2 => n530, ZN 
                           => n2853);
   U745 : OAI22_X1 port map( A1 => n21, A2 => n520, B1 => n521, B2 => n531, ZN 
                           => n2854);
   U746 : OAI22_X1 port map( A1 => n23, A2 => n520, B1 => n521, B2 => n532, ZN 
                           => n2855);
   U747 : OAI22_X1 port map( A1 => n25, A2 => n520, B1 => n521, B2 => n533, ZN 
                           => n2856);
   U748 : OAI22_X1 port map( A1 => n27, A2 => n520, B1 => n521, B2 => n534, ZN 
                           => n2857);
   U749 : OAI22_X1 port map( A1 => n29, A2 => n520, B1 => n521, B2 => n535, ZN 
                           => n2858);
   U750 : OAI22_X1 port map( A1 => n31, A2 => n520, B1 => n521, B2 => n536, ZN 
                           => n2859);
   U751 : OAI22_X1 port map( A1 => n33, A2 => n520, B1 => n521, B2 => n537, ZN 
                           => n2860);
   U752 : OAI22_X1 port map( A1 => n35, A2 => n520, B1 => n521, B2 => n538, ZN 
                           => n2861);
   U753 : OAI22_X1 port map( A1 => n37, A2 => n520, B1 => n521, B2 => n539, ZN 
                           => n2862);
   U754 : OAI22_X1 port map( A1 => n39, A2 => n520, B1 => n521, B2 => n540, ZN 
                           => n2863);
   U755 : OAI22_X1 port map( A1 => n41, A2 => n520, B1 => n521, B2 => n541, ZN 
                           => n2864);
   U756 : OAI22_X1 port map( A1 => n43, A2 => n520, B1 => n521, B2 => n542, ZN 
                           => n2865);
   U757 : OAI22_X1 port map( A1 => n45, A2 => n520, B1 => n521, B2 => n543, ZN 
                           => n2866);
   U758 : OAI22_X1 port map( A1 => n47, A2 => n520, B1 => n521, B2 => n544, ZN 
                           => n2867);
   U759 : OAI22_X1 port map( A1 => n49, A2 => n520, B1 => n521, B2 => n545, ZN 
                           => n2868);
   U760 : OAI22_X1 port map( A1 => n51, A2 => n520, B1 => n521, B2 => n546, ZN 
                           => n2869);
   U761 : OAI22_X1 port map( A1 => n53, A2 => n520, B1 => n521, B2 => n547, ZN 
                           => n2870);
   U762 : OAI22_X1 port map( A1 => n55, A2 => n520, B1 => n521, B2 => n548, ZN 
                           => n2871);
   U763 : OAI22_X1 port map( A1 => n57, A2 => n520, B1 => n521, B2 => n549, ZN 
                           => n2872);
   U764 : OAI22_X1 port map( A1 => n59, A2 => n520, B1 => n521, B2 => n550, ZN 
                           => n2873);
   U765 : OAI22_X1 port map( A1 => n61, A2 => n520, B1 => n521, B2 => n551, ZN 
                           => n2874);
   U766 : OAI22_X1 port map( A1 => n63, A2 => n520, B1 => n521, B2 => n552, ZN 
                           => n2875);
   U767 : OAI22_X1 port map( A1 => n65, A2 => n520, B1 => n521, B2 => n553, ZN 
                           => n2876);
   U770 : OAI22_X1 port map( A1 => n2, A2 => n554, B1 => n555, B2 => n556, ZN 
                           => n2877);
   U771 : OAI22_X1 port map( A1 => n5, A2 => n554, B1 => n555, B2 => n557, ZN 
                           => n2878);
   U772 : OAI22_X1 port map( A1 => n7, A2 => n554, B1 => n555, B2 => n558, ZN 
                           => n2879);
   U773 : OAI22_X1 port map( A1 => n9, A2 => n554, B1 => n555, B2 => n559, ZN 
                           => n2880);
   U774 : OAI22_X1 port map( A1 => n11, A2 => n554, B1 => n555, B2 => n560, ZN 
                           => n2881);
   U775 : OAI22_X1 port map( A1 => n13, A2 => n554, B1 => n555, B2 => n561, ZN 
                           => n2882);
   U776 : OAI22_X1 port map( A1 => n15, A2 => n554, B1 => n555, B2 => n562, ZN 
                           => n2883);
   U777 : OAI22_X1 port map( A1 => n17, A2 => n554, B1 => n555, B2 => n563, ZN 
                           => n2884);
   U778 : OAI22_X1 port map( A1 => n19, A2 => n554, B1 => n555, B2 => n564, ZN 
                           => n2885);
   U779 : OAI22_X1 port map( A1 => n21, A2 => n554, B1 => n555, B2 => n565, ZN 
                           => n2886);
   U780 : OAI22_X1 port map( A1 => n23, A2 => n554, B1 => n555, B2 => n566, ZN 
                           => n2887);
   U781 : OAI22_X1 port map( A1 => n25, A2 => n554, B1 => n555, B2 => n567, ZN 
                           => n2888);
   U782 : OAI22_X1 port map( A1 => n27, A2 => n554, B1 => n555, B2 => n568, ZN 
                           => n2889);
   U783 : OAI22_X1 port map( A1 => n29, A2 => n554, B1 => n555, B2 => n569, ZN 
                           => n2890);
   U784 : OAI22_X1 port map( A1 => n31, A2 => n554, B1 => n555, B2 => n570, ZN 
                           => n2891);
   U785 : OAI22_X1 port map( A1 => n33, A2 => n554, B1 => n555, B2 => n571, ZN 
                           => n2892);
   U786 : OAI22_X1 port map( A1 => n35, A2 => n554, B1 => n555, B2 => n572, ZN 
                           => n2893);
   U787 : OAI22_X1 port map( A1 => n37, A2 => n554, B1 => n555, B2 => n573, ZN 
                           => n2894);
   U788 : OAI22_X1 port map( A1 => n39, A2 => n554, B1 => n555, B2 => n574, ZN 
                           => n2895);
   U789 : OAI22_X1 port map( A1 => n41, A2 => n554, B1 => n555, B2 => n575, ZN 
                           => n2896);
   U790 : OAI22_X1 port map( A1 => n43, A2 => n554, B1 => n555, B2 => n576, ZN 
                           => n2897);
   U791 : OAI22_X1 port map( A1 => n45, A2 => n554, B1 => n555, B2 => n577, ZN 
                           => n2898);
   U792 : OAI22_X1 port map( A1 => n47, A2 => n554, B1 => n555, B2 => n578, ZN 
                           => n2899);
   U793 : OAI22_X1 port map( A1 => n49, A2 => n554, B1 => n555, B2 => n579, ZN 
                           => n2900);
   U794 : OAI22_X1 port map( A1 => n51, A2 => n554, B1 => n555, B2 => n580, ZN 
                           => n2901);
   U795 : OAI22_X1 port map( A1 => n53, A2 => n554, B1 => n555, B2 => n581, ZN 
                           => n2902);
   U796 : OAI22_X1 port map( A1 => n55, A2 => n554, B1 => n555, B2 => n582, ZN 
                           => n2903);
   U797 : OAI22_X1 port map( A1 => n57, A2 => n554, B1 => n555, B2 => n583, ZN 
                           => n2904);
   U798 : OAI22_X1 port map( A1 => n59, A2 => n554, B1 => n555, B2 => n584, ZN 
                           => n2905);
   U799 : OAI22_X1 port map( A1 => n61, A2 => n554, B1 => n555, B2 => n585, ZN 
                           => n2906);
   U800 : OAI22_X1 port map( A1 => n63, A2 => n554, B1 => n555, B2 => n586, ZN 
                           => n2907);
   U801 : OAI22_X1 port map( A1 => n65, A2 => n554, B1 => n555, B2 => n587, ZN 
                           => n2908);
   U804 : AND3_X1 port map( A1 => n314_port, A2 => n588, A3 => ADD_WR(4), ZN =>
                           n349_port);
   U805 : INV_X1 port map( A => n589, ZN => n2909);
   U806 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_0_port, ZN => n589);
   U807 : INV_X1 port map( A => n592, ZN => n2910);
   U808 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_1_port, ZN => n592);
   U809 : INV_X1 port map( A => n593, ZN => n2911);
   U810 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_2_port, ZN => n593);
   U811 : INV_X1 port map( A => n594, ZN => n2912);
   U812 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_3_port, ZN => n594);
   U813 : INV_X1 port map( A => n595, ZN => n2913);
   U814 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_4_port, ZN => n595);
   U815 : INV_X1 port map( A => n596, ZN => n2914);
   U816 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_5_port, ZN => n596);
   U817 : INV_X1 port map( A => n597, ZN => n2915);
   U818 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_6_port, ZN => n597);
   U819 : INV_X1 port map( A => n598, ZN => n2916);
   U820 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_7_port, ZN => n598);
   U821 : INV_X1 port map( A => n599, ZN => n2917);
   U822 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_8_port, ZN => n599);
   U823 : INV_X1 port map( A => n600, ZN => n2918);
   U824 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_9_port, ZN => n600);
   U825 : INV_X1 port map( A => n601, ZN => n2919);
   U826 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_10_port, ZN => n601);
   U827 : INV_X1 port map( A => n602, ZN => n2920);
   U828 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_11_port, ZN => n602);
   U829 : INV_X1 port map( A => n603, ZN => n2921);
   U830 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_12_port, ZN => n603);
   U831 : INV_X1 port map( A => n604, ZN => n2922);
   U832 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_13_port, ZN => n604);
   U833 : INV_X1 port map( A => n605, ZN => n2923);
   U834 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_14_port, ZN => n605);
   U835 : INV_X1 port map( A => n606, ZN => n2924);
   U836 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_15_port, ZN => n606);
   U837 : INV_X1 port map( A => n607, ZN => n2925);
   U838 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_16_port, ZN => n607);
   U839 : INV_X1 port map( A => n608, ZN => n2926);
   U840 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_17_port, ZN => n608);
   U841 : INV_X1 port map( A => n609, ZN => n2927);
   U842 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_18_port, ZN => n609);
   U843 : INV_X1 port map( A => n610, ZN => n2928);
   U844 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_19_port, ZN => n610);
   U845 : INV_X1 port map( A => n611, ZN => n2929);
   U846 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_20_port, ZN => n611);
   U847 : INV_X1 port map( A => n612, ZN => n2930);
   U848 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_21_port, ZN => n612);
   U849 : INV_X1 port map( A => n613, ZN => n2931);
   U850 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_22_port, ZN => n613);
   U851 : INV_X1 port map( A => n614, ZN => n2932);
   U852 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_23_port, ZN => n614);
   U853 : INV_X1 port map( A => n615, ZN => n2933);
   U854 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_24_port, ZN => n615);
   U855 : INV_X1 port map( A => n616, ZN => n2934);
   U856 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_25_port, ZN => n616);
   U857 : INV_X1 port map( A => n617, ZN => n2935);
   U858 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_26_port, ZN => n617);
   U859 : INV_X1 port map( A => n618, ZN => n2936);
   U860 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_27_port, ZN => n618);
   U861 : INV_X1 port map( A => n619, ZN => n2937);
   U862 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_28_port, ZN => n619);
   U863 : INV_X1 port map( A => n620, ZN => n2938);
   U864 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_29_port, ZN => n620);
   U865 : INV_X1 port map( A => n621, ZN => n2939);
   U866 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_30_port, ZN => n621);
   U867 : INV_X1 port map( A => n622, ZN => n2940);
   U868 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n590, B1 => n591, B2 => 
                           REGISTERS_15_31_port, ZN => n622);
   U871 : INV_X1 port map( A => n624, ZN => n2941);
   U872 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_0_port, ZN => n624);
   U873 : INV_X1 port map( A => n627, ZN => n2942);
   U874 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_1_port, ZN => n627);
   U875 : INV_X1 port map( A => n628, ZN => n2943);
   U876 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_2_port, ZN => n628);
   U877 : INV_X1 port map( A => n629, ZN => n2944);
   U878 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_3_port, ZN => n629);
   U879 : INV_X1 port map( A => n630, ZN => n2945);
   U880 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_4_port, ZN => n630);
   U881 : INV_X1 port map( A => n631, ZN => n2946);
   U882 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_5_port, ZN => n631);
   U883 : INV_X1 port map( A => n632, ZN => n2947);
   U884 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_6_port, ZN => n632);
   U885 : INV_X1 port map( A => n633, ZN => n2948);
   U886 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_7_port, ZN => n633);
   U887 : INV_X1 port map( A => n634, ZN => n2949);
   U888 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_8_port, ZN => n634);
   U889 : INV_X1 port map( A => n635, ZN => n2950);
   U890 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_9_port, ZN => n635);
   U891 : INV_X1 port map( A => n636, ZN => n2951);
   U892 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_10_port, ZN => n636);
   U893 : INV_X1 port map( A => n637, ZN => n2952);
   U894 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_11_port, ZN => n637);
   U895 : INV_X1 port map( A => n638, ZN => n2953);
   U896 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_12_port, ZN => n638);
   U897 : INV_X1 port map( A => n639, ZN => n2954);
   U898 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_13_port, ZN => n639);
   U899 : INV_X1 port map( A => n640, ZN => n2955);
   U900 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_14_port, ZN => n640);
   U901 : INV_X1 port map( A => n641, ZN => n2956);
   U902 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_15_port, ZN => n641);
   U903 : INV_X1 port map( A => n642, ZN => n2957);
   U904 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_16_port, ZN => n642);
   U905 : INV_X1 port map( A => n643, ZN => n2958);
   U906 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_17_port, ZN => n643);
   U907 : INV_X1 port map( A => n644, ZN => n2959);
   U908 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_18_port, ZN => n644);
   U909 : INV_X1 port map( A => n645, ZN => n2960);
   U910 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_19_port, ZN => n645);
   U911 : INV_X1 port map( A => n646, ZN => n2961);
   U912 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_20_port, ZN => n646);
   U913 : INV_X1 port map( A => n647, ZN => n2962);
   U914 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_21_port, ZN => n647);
   U915 : INV_X1 port map( A => n648, ZN => n2963);
   U916 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_22_port, ZN => n648);
   U917 : INV_X1 port map( A => n649, ZN => n2964);
   U918 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_23_port, ZN => n649);
   U919 : INV_X1 port map( A => n650, ZN => n2965);
   U920 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_24_port, ZN => n650);
   U921 : INV_X1 port map( A => n651, ZN => n2966);
   U922 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_25_port, ZN => n651);
   U923 : INV_X1 port map( A => n652, ZN => n2967);
   U924 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_26_port, ZN => n652);
   U925 : INV_X1 port map( A => n653, ZN => n2968);
   U926 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_27_port, ZN => n653);
   U927 : INV_X1 port map( A => n654, ZN => n2969);
   U928 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_28_port, ZN => n654);
   U929 : INV_X1 port map( A => n655, ZN => n2970);
   U930 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_29_port, ZN => n655);
   U931 : INV_X1 port map( A => n656, ZN => n2971);
   U932 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_30_port, ZN => n656);
   U933 : INV_X1 port map( A => n657, ZN => n2972);
   U934 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n625, B1 => n626, B2 => 
                           REGISTERS_14_31_port, ZN => n657);
   U937 : OAI22_X1 port map( A1 => n2, A2 => n658, B1 => n659, B2 => n660, ZN 
                           => n2973);
   U938 : OAI22_X1 port map( A1 => n5, A2 => n658, B1 => n659, B2 => n661, ZN 
                           => n2974);
   U939 : OAI22_X1 port map( A1 => n7, A2 => n658, B1 => n659, B2 => n662, ZN 
                           => n2975);
   U940 : OAI22_X1 port map( A1 => n9, A2 => n658, B1 => n659, B2 => n663, ZN 
                           => n2976);
   U941 : OAI22_X1 port map( A1 => n11, A2 => n658, B1 => n659, B2 => n664, ZN 
                           => n2977);
   U942 : OAI22_X1 port map( A1 => n13, A2 => n658, B1 => n659, B2 => n665, ZN 
                           => n2978);
   U943 : OAI22_X1 port map( A1 => n15, A2 => n658, B1 => n659, B2 => n666, ZN 
                           => n2979);
   U944 : OAI22_X1 port map( A1 => n17, A2 => n658, B1 => n659, B2 => n667, ZN 
                           => n2980);
   U945 : OAI22_X1 port map( A1 => n19, A2 => n658, B1 => n659, B2 => n668, ZN 
                           => n2981);
   U946 : OAI22_X1 port map( A1 => n21, A2 => n658, B1 => n659, B2 => n669, ZN 
                           => n2982);
   U947 : OAI22_X1 port map( A1 => n23, A2 => n658, B1 => n659, B2 => n670, ZN 
                           => n2983);
   U948 : OAI22_X1 port map( A1 => n25, A2 => n658, B1 => n659, B2 => n671, ZN 
                           => n2984);
   U949 : OAI22_X1 port map( A1 => n27, A2 => n658, B1 => n659, B2 => n672, ZN 
                           => n2985);
   U950 : OAI22_X1 port map( A1 => n29, A2 => n658, B1 => n659, B2 => n673, ZN 
                           => n2986);
   U951 : OAI22_X1 port map( A1 => n31, A2 => n658, B1 => n659, B2 => n674, ZN 
                           => n2987);
   U952 : OAI22_X1 port map( A1 => n33, A2 => n658, B1 => n659, B2 => n675, ZN 
                           => n2988);
   U953 : OAI22_X1 port map( A1 => n35, A2 => n658, B1 => n659, B2 => n676, ZN 
                           => n2989);
   U954 : OAI22_X1 port map( A1 => n37, A2 => n658, B1 => n659, B2 => n677, ZN 
                           => n2990);
   U955 : OAI22_X1 port map( A1 => n39, A2 => n658, B1 => n659, B2 => n678, ZN 
                           => n2991);
   U956 : OAI22_X1 port map( A1 => n41, A2 => n658, B1 => n659, B2 => n679, ZN 
                           => n2992);
   U957 : OAI22_X1 port map( A1 => n43, A2 => n658, B1 => n659, B2 => n680, ZN 
                           => n2993);
   U958 : OAI22_X1 port map( A1 => n45, A2 => n658, B1 => n659, B2 => n681, ZN 
                           => n2994);
   U959 : OAI22_X1 port map( A1 => n47, A2 => n658, B1 => n659, B2 => n682, ZN 
                           => n2995);
   U960 : OAI22_X1 port map( A1 => n49, A2 => n658, B1 => n659, B2 => n683, ZN 
                           => n2996);
   U961 : OAI22_X1 port map( A1 => n51, A2 => n658, B1 => n659, B2 => n684, ZN 
                           => n2997);
   U962 : OAI22_X1 port map( A1 => n53, A2 => n658, B1 => n659, B2 => n685, ZN 
                           => n2998);
   U963 : OAI22_X1 port map( A1 => n55, A2 => n658, B1 => n659, B2 => n686, ZN 
                           => n2999);
   U964 : OAI22_X1 port map( A1 => n57, A2 => n658, B1 => n659, B2 => n687, ZN 
                           => n3000);
   U965 : OAI22_X1 port map( A1 => n59, A2 => n658, B1 => n659, B2 => n688, ZN 
                           => n3001);
   U966 : OAI22_X1 port map( A1 => n61, A2 => n658, B1 => n659, B2 => n689, ZN 
                           => n3002);
   U967 : OAI22_X1 port map( A1 => n63, A2 => n658, B1 => n659, B2 => n690, ZN 
                           => n3003);
   U968 : OAI22_X1 port map( A1 => n65, A2 => n658, B1 => n659, B2 => n691, ZN 
                           => n3004);
   U971 : OAI22_X1 port map( A1 => n2, A2 => n692, B1 => n693, B2 => n694, ZN 
                           => n3005);
   U972 : OAI22_X1 port map( A1 => n5, A2 => n692, B1 => n693, B2 => n695, ZN 
                           => n3006);
   U973 : OAI22_X1 port map( A1 => n7, A2 => n692, B1 => n693, B2 => n696, ZN 
                           => n3007);
   U974 : OAI22_X1 port map( A1 => n9, A2 => n692, B1 => n693, B2 => n697, ZN 
                           => n3008);
   U975 : OAI22_X1 port map( A1 => n11, A2 => n692, B1 => n693, B2 => n698, ZN 
                           => n3009);
   U976 : OAI22_X1 port map( A1 => n13, A2 => n692, B1 => n693, B2 => n699, ZN 
                           => n3010);
   U977 : OAI22_X1 port map( A1 => n15, A2 => n692, B1 => n693, B2 => n700, ZN 
                           => n3011);
   U978 : OAI22_X1 port map( A1 => n17, A2 => n692, B1 => n693, B2 => n701, ZN 
                           => n3012);
   U979 : OAI22_X1 port map( A1 => n19, A2 => n692, B1 => n693, B2 => n702, ZN 
                           => n3013);
   U980 : OAI22_X1 port map( A1 => n21, A2 => n692, B1 => n693, B2 => n703, ZN 
                           => n3014);
   U981 : OAI22_X1 port map( A1 => n23, A2 => n692, B1 => n693, B2 => n704, ZN 
                           => n3015);
   U982 : OAI22_X1 port map( A1 => n25, A2 => n692, B1 => n693, B2 => n705, ZN 
                           => n3016);
   U983 : OAI22_X1 port map( A1 => n27, A2 => n692, B1 => n693, B2 => n706, ZN 
                           => n3017);
   U984 : OAI22_X1 port map( A1 => n29, A2 => n692, B1 => n693, B2 => n707, ZN 
                           => n3018);
   U985 : OAI22_X1 port map( A1 => n31, A2 => n692, B1 => n693, B2 => n708, ZN 
                           => n3019);
   U986 : OAI22_X1 port map( A1 => n33, A2 => n692, B1 => n693, B2 => n709, ZN 
                           => n3020);
   U987 : OAI22_X1 port map( A1 => n35, A2 => n692, B1 => n693, B2 => n710, ZN 
                           => n3021);
   U988 : OAI22_X1 port map( A1 => n37, A2 => n692, B1 => n693, B2 => n711, ZN 
                           => n3022);
   U989 : OAI22_X1 port map( A1 => n39, A2 => n692, B1 => n693, B2 => n712, ZN 
                           => n3023);
   U990 : OAI22_X1 port map( A1 => n41, A2 => n692, B1 => n693, B2 => n713, ZN 
                           => n3024);
   U991 : OAI22_X1 port map( A1 => n43, A2 => n692, B1 => n693, B2 => n714, ZN 
                           => n3025);
   U992 : OAI22_X1 port map( A1 => n45, A2 => n692, B1 => n693, B2 => n715, ZN 
                           => n3026);
   U993 : OAI22_X1 port map( A1 => n47, A2 => n692, B1 => n693, B2 => n716, ZN 
                           => n3027);
   U994 : OAI22_X1 port map( A1 => n49, A2 => n692, B1 => n693, B2 => n717, ZN 
                           => n3028);
   U995 : OAI22_X1 port map( A1 => n51, A2 => n692, B1 => n693, B2 => n718, ZN 
                           => n3029);
   U996 : OAI22_X1 port map( A1 => n53, A2 => n692, B1 => n693, B2 => n719, ZN 
                           => n3030);
   U997 : OAI22_X1 port map( A1 => n55, A2 => n692, B1 => n693, B2 => n720, ZN 
                           => n3031);
   U998 : OAI22_X1 port map( A1 => n57, A2 => n692, B1 => n693, B2 => n721, ZN 
                           => n3032);
   U999 : OAI22_X1 port map( A1 => n59, A2 => n692, B1 => n693, B2 => n722, ZN 
                           => n3033);
   U1000 : OAI22_X1 port map( A1 => n61, A2 => n692, B1 => n693, B2 => n723, ZN
                           => n3034);
   U1001 : OAI22_X1 port map( A1 => n63, A2 => n692, B1 => n693, B2 => n724, ZN
                           => n3035);
   U1002 : OAI22_X1 port map( A1 => n65, A2 => n692, B1 => n693, B2 => n725, ZN
                           => n3036);
   U1005 : INV_X1 port map( A => n726, ZN => n3037);
   U1006 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_0_port, ZN => n726);
   U1007 : INV_X1 port map( A => n729, ZN => n3038);
   U1008 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_1_port, ZN => n729);
   U1009 : INV_X1 port map( A => n730, ZN => n3039);
   U1010 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_2_port, ZN => n730);
   U1011 : INV_X1 port map( A => n731, ZN => n3040);
   U1012 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_3_port, ZN => n731);
   U1013 : INV_X1 port map( A => n732, ZN => n3041);
   U1014 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_4_port, ZN => n732);
   U1015 : INV_X1 port map( A => n733, ZN => n3042);
   U1016 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_5_port, ZN => n733);
   U1017 : INV_X1 port map( A => n734, ZN => n3043);
   U1018 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_6_port, ZN => n734);
   U1019 : INV_X1 port map( A => n735, ZN => n3044);
   U1020 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_7_port, ZN => n735);
   U1021 : INV_X1 port map( A => n736, ZN => n3045);
   U1022 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_8_port, ZN => n736);
   U1023 : INV_X1 port map( A => n737, ZN => n3046);
   U1024 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_9_port, ZN => n737);
   U1025 : INV_X1 port map( A => n738, ZN => n3047);
   U1026 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_10_port, ZN => n738);
   U1027 : INV_X1 port map( A => n739, ZN => n3048);
   U1028 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_11_port, ZN => n739);
   U1029 : INV_X1 port map( A => n740, ZN => n3049);
   U1030 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_12_port, ZN => n740);
   U1031 : INV_X1 port map( A => n741, ZN => n3050);
   U1032 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_13_port, ZN => n741);
   U1033 : INV_X1 port map( A => n742, ZN => n3051);
   U1034 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_14_port, ZN => n742);
   U1035 : INV_X1 port map( A => n743, ZN => n3052);
   U1036 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_15_port, ZN => n743);
   U1037 : INV_X1 port map( A => n744, ZN => n3053);
   U1038 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_16_port, ZN => n744);
   U1039 : INV_X1 port map( A => n745, ZN => n3054);
   U1040 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_17_port, ZN => n745);
   U1041 : INV_X1 port map( A => n746, ZN => n3055);
   U1042 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_18_port, ZN => n746);
   U1043 : INV_X1 port map( A => n747, ZN => n3056);
   U1044 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_19_port, ZN => n747);
   U1045 : INV_X1 port map( A => n748, ZN => n3057);
   U1046 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_20_port, ZN => n748);
   U1047 : INV_X1 port map( A => n749, ZN => n3058);
   U1048 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_21_port, ZN => n749);
   U1049 : INV_X1 port map( A => n750, ZN => n3059);
   U1050 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_22_port, ZN => n750);
   U1051 : INV_X1 port map( A => n751, ZN => n3060);
   U1052 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_23_port, ZN => n751);
   U1053 : INV_X1 port map( A => n752, ZN => n3061);
   U1054 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_24_port, ZN => n752);
   U1055 : INV_X1 port map( A => n753, ZN => n3062);
   U1056 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_25_port, ZN => n753);
   U1057 : INV_X1 port map( A => n754, ZN => n3063);
   U1058 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_26_port, ZN => n754);
   U1059 : INV_X1 port map( A => n755, ZN => n3064);
   U1060 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_27_port, ZN => n755);
   U1061 : INV_X1 port map( A => n756, ZN => n3065);
   U1062 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_28_port, ZN => n756);
   U1063 : INV_X1 port map( A => n757, ZN => n3066);
   U1064 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_29_port, ZN => n757);
   U1065 : INV_X1 port map( A => n758, ZN => n3067);
   U1066 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_30_port, ZN => n758);
   U1067 : INV_X1 port map( A => n759, ZN => n3068);
   U1068 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n727, B1 => n728, B2 => 
                           REGISTERS_11_31_port, ZN => n759);
   U1071 : INV_X1 port map( A => n760, ZN => n3069);
   U1072 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_0_port, ZN => n760);
   U1073 : INV_X1 port map( A => n763, ZN => n3070);
   U1074 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_1_port, ZN => n763);
   U1075 : INV_X1 port map( A => n764, ZN => n3071);
   U1076 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_2_port, ZN => n764);
   U1077 : INV_X1 port map( A => n765, ZN => n3072);
   U1078 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_3_port, ZN => n765);
   U1079 : INV_X1 port map( A => n766, ZN => n3073);
   U1080 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_4_port, ZN => n766);
   U1081 : INV_X1 port map( A => n767, ZN => n3074);
   U1082 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_5_port, ZN => n767);
   U1083 : INV_X1 port map( A => n768, ZN => n3075);
   U1084 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_6_port, ZN => n768);
   U1085 : INV_X1 port map( A => n769, ZN => n3076);
   U1086 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_7_port, ZN => n769);
   U1087 : INV_X1 port map( A => n770, ZN => n3077);
   U1088 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_8_port, ZN => n770);
   U1089 : INV_X1 port map( A => n771, ZN => n3078);
   U1090 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_9_port, ZN => n771);
   U1091 : INV_X1 port map( A => n772, ZN => n3079);
   U1092 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_10_port, ZN => n772);
   U1093 : INV_X1 port map( A => n773, ZN => n3080);
   U1094 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_11_port, ZN => n773);
   U1095 : INV_X1 port map( A => n774, ZN => n3081);
   U1096 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_12_port, ZN => n774);
   U1097 : INV_X1 port map( A => n775, ZN => n3082);
   U1098 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_13_port, ZN => n775);
   U1099 : INV_X1 port map( A => n776, ZN => n3083);
   U1100 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_14_port, ZN => n776);
   U1101 : INV_X1 port map( A => n777, ZN => n3084);
   U1102 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_15_port, ZN => n777);
   U1103 : INV_X1 port map( A => n778, ZN => n3085);
   U1104 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_16_port, ZN => n778);
   U1105 : INV_X1 port map( A => n779, ZN => n3086);
   U1106 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_17_port, ZN => n779);
   U1107 : INV_X1 port map( A => n780, ZN => n3087);
   U1108 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_18_port, ZN => n780);
   U1109 : INV_X1 port map( A => n781, ZN => n3088);
   U1110 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_19_port, ZN => n781);
   U1111 : INV_X1 port map( A => n782, ZN => n3089);
   U1112 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_20_port, ZN => n782);
   U1113 : INV_X1 port map( A => n783, ZN => n3090);
   U1114 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_21_port, ZN => n783);
   U1115 : INV_X1 port map( A => n784, ZN => n3091);
   U1116 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_22_port, ZN => n784);
   U1117 : INV_X1 port map( A => n785, ZN => n3092);
   U1118 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_23_port, ZN => n785);
   U1119 : INV_X1 port map( A => n786, ZN => n3093);
   U1120 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_24_port, ZN => n786);
   U1121 : INV_X1 port map( A => n787, ZN => n3094);
   U1122 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_25_port, ZN => n787);
   U1123 : INV_X1 port map( A => n788, ZN => n3095);
   U1124 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_26_port, ZN => n788);
   U1125 : INV_X1 port map( A => n789, ZN => n3096);
   U1126 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_27_port, ZN => n789);
   U1127 : INV_X1 port map( A => n790, ZN => n3097);
   U1128 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_28_port, ZN => n790);
   U1129 : INV_X1 port map( A => n791, ZN => n3098);
   U1130 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_29_port, ZN => n791);
   U1131 : INV_X1 port map( A => n792, ZN => n3099);
   U1132 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_30_port, ZN => n792);
   U1133 : INV_X1 port map( A => n793, ZN => n3100);
   U1134 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n761, B1 => n762, B2 => 
                           REGISTERS_10_31_port, ZN => n793);
   U1137 : OAI22_X1 port map( A1 => n2, A2 => n794, B1 => n795, B2 => n796, ZN 
                           => n3101);
   U1138 : OAI22_X1 port map( A1 => n5, A2 => n794, B1 => n795, B2 => n797, ZN 
                           => n3102);
   U1139 : OAI22_X1 port map( A1 => n7, A2 => n794, B1 => n795, B2 => n798, ZN 
                           => n3103);
   U1140 : OAI22_X1 port map( A1 => n9, A2 => n794, B1 => n795, B2 => n799, ZN 
                           => n3104);
   U1141 : OAI22_X1 port map( A1 => n11, A2 => n794, B1 => n795, B2 => n800, ZN
                           => n3105);
   U1142 : OAI22_X1 port map( A1 => n13, A2 => n794, B1 => n795, B2 => n801, ZN
                           => n3106);
   U1143 : OAI22_X1 port map( A1 => n15, A2 => n794, B1 => n795, B2 => n802, ZN
                           => n3107);
   U1144 : OAI22_X1 port map( A1 => n17, A2 => n794, B1 => n795, B2 => n803, ZN
                           => n3108);
   U1145 : OAI22_X1 port map( A1 => n19, A2 => n794, B1 => n795, B2 => n804, ZN
                           => n3109);
   U1146 : OAI22_X1 port map( A1 => n21, A2 => n794, B1 => n795, B2 => n805, ZN
                           => n3110);
   U1147 : OAI22_X1 port map( A1 => n23, A2 => n794, B1 => n795, B2 => n806, ZN
                           => n3111);
   U1148 : OAI22_X1 port map( A1 => n25, A2 => n794, B1 => n795, B2 => n807, ZN
                           => n3112);
   U1149 : OAI22_X1 port map( A1 => n27, A2 => n794, B1 => n795, B2 => n808, ZN
                           => n3113);
   U1150 : OAI22_X1 port map( A1 => n29, A2 => n794, B1 => n795, B2 => n809, ZN
                           => n3114);
   U1151 : OAI22_X1 port map( A1 => n31, A2 => n794, B1 => n795, B2 => n810, ZN
                           => n3115);
   U1152 : OAI22_X1 port map( A1 => n33, A2 => n794, B1 => n795, B2 => n811, ZN
                           => n3116);
   U1153 : OAI22_X1 port map( A1 => n35, A2 => n794, B1 => n795, B2 => n812, ZN
                           => n3117);
   U1154 : OAI22_X1 port map( A1 => n37, A2 => n794, B1 => n795, B2 => n813, ZN
                           => n3118);
   U1155 : OAI22_X1 port map( A1 => n39, A2 => n794, B1 => n795, B2 => n814, ZN
                           => n3119);
   U1156 : OAI22_X1 port map( A1 => n41, A2 => n794, B1 => n795, B2 => n815, ZN
                           => n3120);
   U1157 : OAI22_X1 port map( A1 => n43, A2 => n794, B1 => n795, B2 => n816, ZN
                           => n3121);
   U1158 : OAI22_X1 port map( A1 => n45, A2 => n794, B1 => n795, B2 => n817, ZN
                           => n3122);
   U1159 : OAI22_X1 port map( A1 => n47, A2 => n794, B1 => n795, B2 => n818, ZN
                           => n3123);
   U1160 : OAI22_X1 port map( A1 => n49, A2 => n794, B1 => n795, B2 => n819, ZN
                           => n3124);
   U1161 : OAI22_X1 port map( A1 => n51, A2 => n794, B1 => n795, B2 => n820, ZN
                           => n3125);
   U1162 : OAI22_X1 port map( A1 => n53, A2 => n794, B1 => n795, B2 => n821, ZN
                           => n3126);
   U1163 : OAI22_X1 port map( A1 => n55, A2 => n794, B1 => n795, B2 => n822, ZN
                           => n3127);
   U1164 : OAI22_X1 port map( A1 => n57, A2 => n794, B1 => n795, B2 => n823, ZN
                           => n3128);
   U1165 : OAI22_X1 port map( A1 => n59, A2 => n794, B1 => n795, B2 => n824, ZN
                           => n3129);
   U1166 : OAI22_X1 port map( A1 => n61, A2 => n794, B1 => n795, B2 => n825, ZN
                           => n3130);
   U1167 : OAI22_X1 port map( A1 => n63, A2 => n794, B1 => n795, B2 => n826, ZN
                           => n3131);
   U1168 : OAI22_X1 port map( A1 => n65, A2 => n794, B1 => n795, B2 => n827, ZN
                           => n3132);
   U1171 : OAI22_X1 port map( A1 => n2, A2 => n828, B1 => n829, B2 => n830, ZN 
                           => n3133);
   U1172 : OAI22_X1 port map( A1 => n5, A2 => n828, B1 => n829, B2 => n831, ZN 
                           => n3134);
   U1173 : OAI22_X1 port map( A1 => n7, A2 => n828, B1 => n829, B2 => n832, ZN 
                           => n3135);
   U1174 : OAI22_X1 port map( A1 => n9, A2 => n828, B1 => n829, B2 => n833, ZN 
                           => n3136);
   U1175 : OAI22_X1 port map( A1 => n11, A2 => n828, B1 => n829, B2 => n834, ZN
                           => n3137);
   U1176 : OAI22_X1 port map( A1 => n13, A2 => n828, B1 => n829, B2 => n835, ZN
                           => n3138);
   U1177 : OAI22_X1 port map( A1 => n15, A2 => n828, B1 => n829, B2 => n836, ZN
                           => n3139);
   U1178 : OAI22_X1 port map( A1 => n17, A2 => n828, B1 => n829, B2 => n837, ZN
                           => n3140);
   U1179 : OAI22_X1 port map( A1 => n19, A2 => n828, B1 => n829, B2 => n838, ZN
                           => n3141);
   U1180 : OAI22_X1 port map( A1 => n21, A2 => n828, B1 => n829, B2 => n839, ZN
                           => n3142);
   U1181 : OAI22_X1 port map( A1 => n23, A2 => n828, B1 => n829, B2 => n840, ZN
                           => n3143);
   U1182 : OAI22_X1 port map( A1 => n25, A2 => n828, B1 => n829, B2 => n841, ZN
                           => n3144);
   U1183 : OAI22_X1 port map( A1 => n27, A2 => n828, B1 => n829, B2 => n842, ZN
                           => n3145);
   U1184 : OAI22_X1 port map( A1 => n29, A2 => n828, B1 => n829, B2 => n843, ZN
                           => n3146);
   U1185 : OAI22_X1 port map( A1 => n31, A2 => n828, B1 => n829, B2 => n844, ZN
                           => n3147);
   U1186 : OAI22_X1 port map( A1 => n33, A2 => n828, B1 => n829, B2 => n845, ZN
                           => n3148);
   U1187 : OAI22_X1 port map( A1 => n35, A2 => n828, B1 => n829, B2 => n846, ZN
                           => n3149);
   U1188 : OAI22_X1 port map( A1 => n37, A2 => n828, B1 => n829, B2 => n847, ZN
                           => n3150);
   U1189 : OAI22_X1 port map( A1 => n39, A2 => n828, B1 => n829, B2 => n848, ZN
                           => n3151);
   U1190 : OAI22_X1 port map( A1 => n41, A2 => n828, B1 => n829, B2 => n849, ZN
                           => n3152);
   U1191 : OAI22_X1 port map( A1 => n43, A2 => n828, B1 => n829, B2 => n850, ZN
                           => n3153);
   U1192 : OAI22_X1 port map( A1 => n45, A2 => n828, B1 => n829, B2 => n851, ZN
                           => n3154);
   U1193 : OAI22_X1 port map( A1 => n47, A2 => n828, B1 => n829, B2 => n852, ZN
                           => n3155);
   U1194 : OAI22_X1 port map( A1 => n49, A2 => n828, B1 => n829, B2 => n853, ZN
                           => n3156);
   U1195 : OAI22_X1 port map( A1 => n51, A2 => n828, B1 => n829, B2 => n854, ZN
                           => n3157);
   U1196 : OAI22_X1 port map( A1 => n53, A2 => n828, B1 => n829, B2 => n855, ZN
                           => n3158);
   U1197 : OAI22_X1 port map( A1 => n55, A2 => n828, B1 => n829, B2 => n856, ZN
                           => n3159);
   U1198 : OAI22_X1 port map( A1 => n57, A2 => n828, B1 => n829, B2 => n857, ZN
                           => n3160);
   U1199 : OAI22_X1 port map( A1 => n59, A2 => n828, B1 => n829, B2 => n858, ZN
                           => n3161);
   U1200 : OAI22_X1 port map( A1 => n61, A2 => n828, B1 => n829, B2 => n859, ZN
                           => n3162);
   U1201 : OAI22_X1 port map( A1 => n63, A2 => n828, B1 => n829, B2 => n860, ZN
                           => n3163);
   U1202 : OAI22_X1 port map( A1 => n65, A2 => n828, B1 => n829, B2 => n861, ZN
                           => n3164);
   U1205 : AND3_X1 port map( A1 => n314_port, A2 => n862, A3 => ADD_WR(3), ZN 
                           => n623);
   U1206 : INV_X1 port map( A => n863, ZN => n3165);
   U1207 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_0_port, ZN => n863);
   U1208 : INV_X1 port map( A => n866, ZN => n3166);
   U1209 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_1_port, ZN => n866);
   U1210 : INV_X1 port map( A => n867, ZN => n3167);
   U1211 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_2_port, ZN => n867);
   U1212 : INV_X1 port map( A => n868, ZN => n3168);
   U1213 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_3_port, ZN => n868);
   U1214 : INV_X1 port map( A => n869, ZN => n3169);
   U1215 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_4_port, ZN => n869);
   U1216 : INV_X1 port map( A => n870, ZN => n3170);
   U1217 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_5_port, ZN => n870);
   U1218 : INV_X1 port map( A => n871, ZN => n3171);
   U1219 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_6_port, ZN => n871);
   U1220 : INV_X1 port map( A => n872, ZN => n3172);
   U1221 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_7_port, ZN => n872);
   U1222 : INV_X1 port map( A => n873, ZN => n3173);
   U1223 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_8_port, ZN => n873);
   U1224 : INV_X1 port map( A => n874, ZN => n3174);
   U1225 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_9_port, ZN => n874);
   U1226 : INV_X1 port map( A => n875, ZN => n3175);
   U1227 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_10_port, ZN => n875);
   U1228 : INV_X1 port map( A => n876, ZN => n3176);
   U1229 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_11_port, ZN => n876);
   U1230 : INV_X1 port map( A => n877, ZN => n3177);
   U1231 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_12_port, ZN => n877);
   U1232 : INV_X1 port map( A => n878, ZN => n3178);
   U1233 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_13_port, ZN => n878);
   U1234 : INV_X1 port map( A => n879, ZN => n3179);
   U1235 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_14_port, ZN => n879);
   U1236 : INV_X1 port map( A => n880, ZN => n3180);
   U1237 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_15_port, ZN => n880);
   U1238 : INV_X1 port map( A => n881, ZN => n3181);
   U1239 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_16_port, ZN => n881);
   U1240 : INV_X1 port map( A => n882, ZN => n3182);
   U1241 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_17_port, ZN => n882);
   U1242 : INV_X1 port map( A => n883, ZN => n3183);
   U1243 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_18_port, ZN => n883);
   U1244 : INV_X1 port map( A => n884, ZN => n3184);
   U1245 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_19_port, ZN => n884);
   U1246 : INV_X1 port map( A => n885, ZN => n3185);
   U1247 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_20_port, ZN => n885);
   U1248 : INV_X1 port map( A => n886, ZN => n3186);
   U1249 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_21_port, ZN => n886);
   U1250 : INV_X1 port map( A => n887, ZN => n3187);
   U1251 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_22_port, ZN => n887);
   U1252 : INV_X1 port map( A => n888, ZN => n3188);
   U1253 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_23_port, ZN => n888);
   U1254 : INV_X1 port map( A => n889, ZN => n3189);
   U1255 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_24_port, ZN => n889);
   U1256 : INV_X1 port map( A => n890, ZN => n3190);
   U1257 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_25_port, ZN => n890);
   U1258 : INV_X1 port map( A => n891, ZN => n3191);
   U1259 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_26_port, ZN => n891);
   U1260 : INV_X1 port map( A => n892, ZN => n3192);
   U1261 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_27_port, ZN => n892);
   U1262 : INV_X1 port map( A => n893, ZN => n3193);
   U1263 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_28_port, ZN => n893);
   U1264 : INV_X1 port map( A => n894, ZN => n3194);
   U1265 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_29_port, ZN => n894);
   U1266 : INV_X1 port map( A => n895, ZN => n3195);
   U1267 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_30_port, ZN => n895);
   U1268 : INV_X1 port map( A => n896, ZN => n3196);
   U1269 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n864, B1 => n865, B2 => 
                           REGISTERS_7_31_port, ZN => n896);
   U1272 : NOR3_X1 port map( A1 => n898, A2 => n899, A3 => n900, ZN => n67);
   U1273 : INV_X1 port map( A => n901, ZN => n3197);
   U1274 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_0_port, ZN => n901);
   U1275 : INV_X1 port map( A => n904, ZN => n3198);
   U1276 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_1_port, ZN => n904);
   U1277 : INV_X1 port map( A => n905, ZN => n3199);
   U1278 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_2_port, ZN => n905);
   U1279 : INV_X1 port map( A => n906, ZN => n3200);
   U1280 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_3_port, ZN => n906);
   U1281 : INV_X1 port map( A => n907, ZN => n3201);
   U1282 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_4_port, ZN => n907);
   U1283 : INV_X1 port map( A => n908, ZN => n3202);
   U1284 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_5_port, ZN => n908);
   U1285 : INV_X1 port map( A => n909, ZN => n3203);
   U1286 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_6_port, ZN => n909);
   U1287 : INV_X1 port map( A => n910, ZN => n3204);
   U1288 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_7_port, ZN => n910);
   U1289 : INV_X1 port map( A => n911, ZN => n3205);
   U1290 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_8_port, ZN => n911);
   U1291 : INV_X1 port map( A => n912, ZN => n3206);
   U1292 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_9_port, ZN => n912);
   U1293 : INV_X1 port map( A => n913, ZN => n3207);
   U1294 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_10_port, ZN => n913);
   U1295 : INV_X1 port map( A => n914, ZN => n3208);
   U1296 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_11_port, ZN => n914);
   U1297 : INV_X1 port map( A => n915, ZN => n3209);
   U1298 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_12_port, ZN => n915);
   U1299 : INV_X1 port map( A => n916, ZN => n3210);
   U1300 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_13_port, ZN => n916);
   U1301 : INV_X1 port map( A => n917, ZN => n3211);
   U1302 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_14_port, ZN => n917);
   U1303 : INV_X1 port map( A => n918, ZN => n3212);
   U1304 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_15_port, ZN => n918);
   U1305 : INV_X1 port map( A => n919, ZN => n3213);
   U1306 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_16_port, ZN => n919);
   U1307 : INV_X1 port map( A => n920, ZN => n3214);
   U1308 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_17_port, ZN => n920);
   U1309 : INV_X1 port map( A => n921, ZN => n3215);
   U1310 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_18_port, ZN => n921);
   U1311 : INV_X1 port map( A => n922, ZN => n3216);
   U1312 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_19_port, ZN => n922);
   U1313 : INV_X1 port map( A => n923, ZN => n3217);
   U1314 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_20_port, ZN => n923);
   U1315 : INV_X1 port map( A => n924, ZN => n3218);
   U1316 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_21_port, ZN => n924);
   U1317 : INV_X1 port map( A => n925, ZN => n3219);
   U1318 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_22_port, ZN => n925);
   U1319 : INV_X1 port map( A => n926, ZN => n3220);
   U1320 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_23_port, ZN => n926);
   U1321 : INV_X1 port map( A => n927, ZN => n3221);
   U1322 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_24_port, ZN => n927);
   U1323 : INV_X1 port map( A => n928, ZN => n3222);
   U1324 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_25_port, ZN => n928);
   U1325 : INV_X1 port map( A => n929, ZN => n3223);
   U1326 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_26_port, ZN => n929);
   U1327 : INV_X1 port map( A => n930, ZN => n3224);
   U1328 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_27_port, ZN => n930);
   U1329 : INV_X1 port map( A => n931, ZN => n3225);
   U1330 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_28_port, ZN => n931);
   U1331 : INV_X1 port map( A => n932, ZN => n3226);
   U1332 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_29_port, ZN => n932);
   U1333 : INV_X1 port map( A => n933, ZN => n3227);
   U1334 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_30_port, ZN => n933);
   U1335 : INV_X1 port map( A => n934, ZN => n3228);
   U1336 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n902, B1 => n903, B2 => 
                           REGISTERS_6_31_port, ZN => n934);
   U1339 : NOR3_X1 port map( A1 => n898, A2 => ADD_WR(0), A3 => n900, ZN => 
                           n103);
   U1340 : OAI22_X1 port map( A1 => n2, A2 => n935, B1 => n936, B2 => n937, ZN 
                           => n3229);
   U1341 : OAI22_X1 port map( A1 => n5, A2 => n935, B1 => n936, B2 => n938, ZN 
                           => n3230);
   U1342 : OAI22_X1 port map( A1 => n7, A2 => n935, B1 => n936, B2 => n939, ZN 
                           => n3231);
   U1343 : OAI22_X1 port map( A1 => n9, A2 => n935, B1 => n936, B2 => n940, ZN 
                           => n3232);
   U1344 : OAI22_X1 port map( A1 => n11, A2 => n935, B1 => n936, B2 => n941, ZN
                           => n3233);
   U1345 : OAI22_X1 port map( A1 => n13, A2 => n935, B1 => n936, B2 => n942, ZN
                           => n3234);
   U1346 : OAI22_X1 port map( A1 => n15, A2 => n935, B1 => n936, B2 => n943, ZN
                           => n3235);
   U1347 : OAI22_X1 port map( A1 => n17, A2 => n935, B1 => n936, B2 => n944, ZN
                           => n3236);
   U1348 : OAI22_X1 port map( A1 => n19, A2 => n935, B1 => n936, B2 => n945, ZN
                           => n3237);
   U1349 : OAI22_X1 port map( A1 => n21, A2 => n935, B1 => n936, B2 => n946, ZN
                           => n3238);
   U1350 : OAI22_X1 port map( A1 => n23, A2 => n935, B1 => n936, B2 => n947, ZN
                           => n3239);
   U1351 : OAI22_X1 port map( A1 => n25, A2 => n935, B1 => n936, B2 => n948, ZN
                           => n3240);
   U1352 : OAI22_X1 port map( A1 => n27, A2 => n935, B1 => n936, B2 => n949, ZN
                           => n3241);
   U1353 : OAI22_X1 port map( A1 => n29, A2 => n935, B1 => n936, B2 => n950, ZN
                           => n3242);
   U1354 : OAI22_X1 port map( A1 => n31, A2 => n935, B1 => n936, B2 => n951, ZN
                           => n3243);
   U1355 : OAI22_X1 port map( A1 => n33, A2 => n935, B1 => n936, B2 => n952, ZN
                           => n3244);
   U1356 : OAI22_X1 port map( A1 => n35, A2 => n935, B1 => n936, B2 => n953, ZN
                           => n3245);
   U1357 : OAI22_X1 port map( A1 => n37, A2 => n935, B1 => n936, B2 => n954, ZN
                           => n3246);
   U1358 : OAI22_X1 port map( A1 => n39, A2 => n935, B1 => n936, B2 => n955, ZN
                           => n3247);
   U1359 : OAI22_X1 port map( A1 => n41, A2 => n935, B1 => n936, B2 => n956, ZN
                           => n3248);
   U1360 : OAI22_X1 port map( A1 => n43, A2 => n935, B1 => n936, B2 => n957, ZN
                           => n3249);
   U1361 : OAI22_X1 port map( A1 => n45, A2 => n935, B1 => n936, B2 => n958, ZN
                           => n3250);
   U1362 : OAI22_X1 port map( A1 => n47, A2 => n935, B1 => n936, B2 => n959, ZN
                           => n3251);
   U1363 : OAI22_X1 port map( A1 => n49, A2 => n935, B1 => n936, B2 => n960, ZN
                           => n3252);
   U1364 : OAI22_X1 port map( A1 => n51, A2 => n935, B1 => n936, B2 => n961, ZN
                           => n3253);
   U1365 : OAI22_X1 port map( A1 => n53, A2 => n935, B1 => n936, B2 => n962, ZN
                           => n3254);
   U1366 : OAI22_X1 port map( A1 => n55, A2 => n935, B1 => n936, B2 => n963, ZN
                           => n3255);
   U1367 : OAI22_X1 port map( A1 => n57, A2 => n935, B1 => n936, B2 => n964, ZN
                           => n3256);
   U1368 : OAI22_X1 port map( A1 => n59, A2 => n935, B1 => n936, B2 => n965, ZN
                           => n3257);
   U1369 : OAI22_X1 port map( A1 => n61, A2 => n935, B1 => n936, B2 => n966, ZN
                           => n3258);
   U1370 : OAI22_X1 port map( A1 => n63, A2 => n935, B1 => n936, B2 => n967, ZN
                           => n3259);
   U1371 : OAI22_X1 port map( A1 => n65, A2 => n935, B1 => n936, B2 => n968, ZN
                           => n3260);
   U1374 : NOR3_X1 port map( A1 => n899, A2 => ADD_WR(1), A3 => n900, ZN => 
                           n138);
   U1375 : OAI22_X1 port map( A1 => n2, A2 => n969, B1 => n970, B2 => n971, ZN 
                           => n3261);
   U1376 : OAI22_X1 port map( A1 => n5, A2 => n969, B1 => n970, B2 => n972, ZN 
                           => n3262);
   U1377 : OAI22_X1 port map( A1 => n7, A2 => n969, B1 => n970, B2 => n973, ZN 
                           => n3263);
   U1378 : OAI22_X1 port map( A1 => n9, A2 => n969, B1 => n970, B2 => n974, ZN 
                           => n3264);
   U1379 : OAI22_X1 port map( A1 => n11, A2 => n969, B1 => n970, B2 => n975, ZN
                           => n3265);
   U1380 : OAI22_X1 port map( A1 => n13, A2 => n969, B1 => n970, B2 => n976, ZN
                           => n3266);
   U1381 : OAI22_X1 port map( A1 => n15, A2 => n969, B1 => n970, B2 => n977, ZN
                           => n3267);
   U1382 : OAI22_X1 port map( A1 => n17, A2 => n969, B1 => n970, B2 => n978, ZN
                           => n3268);
   U1383 : OAI22_X1 port map( A1 => n19, A2 => n969, B1 => n970, B2 => n979, ZN
                           => n3269);
   U1384 : OAI22_X1 port map( A1 => n21, A2 => n969, B1 => n970, B2 => n980, ZN
                           => n3270);
   U1385 : OAI22_X1 port map( A1 => n23, A2 => n969, B1 => n970, B2 => n981, ZN
                           => n3271);
   U1386 : OAI22_X1 port map( A1 => n25, A2 => n969, B1 => n970, B2 => n982, ZN
                           => n3272);
   U1387 : OAI22_X1 port map( A1 => n27, A2 => n969, B1 => n970, B2 => n983, ZN
                           => n3273);
   U1388 : OAI22_X1 port map( A1 => n29, A2 => n969, B1 => n970, B2 => n984, ZN
                           => n3274);
   U1389 : OAI22_X1 port map( A1 => n31, A2 => n969, B1 => n970, B2 => n985, ZN
                           => n3275);
   U1390 : OAI22_X1 port map( A1 => n33, A2 => n969, B1 => n970, B2 => n986, ZN
                           => n3276);
   U1391 : OAI22_X1 port map( A1 => n35, A2 => n969, B1 => n970, B2 => n987, ZN
                           => n3277);
   U1392 : OAI22_X1 port map( A1 => n37, A2 => n969, B1 => n970, B2 => n988, ZN
                           => n3278);
   U1393 : OAI22_X1 port map( A1 => n39, A2 => n969, B1 => n970, B2 => n989, ZN
                           => n3279);
   U1394 : OAI22_X1 port map( A1 => n41, A2 => n969, B1 => n970, B2 => n990, ZN
                           => n3280);
   U1395 : OAI22_X1 port map( A1 => n43, A2 => n969, B1 => n970, B2 => n991, ZN
                           => n3281);
   U1396 : OAI22_X1 port map( A1 => n45, A2 => n969, B1 => n970, B2 => n992, ZN
                           => n3282);
   U1397 : OAI22_X1 port map( A1 => n47, A2 => n969, B1 => n970, B2 => n993, ZN
                           => n3283);
   U1398 : OAI22_X1 port map( A1 => n49, A2 => n969, B1 => n970, B2 => n994, ZN
                           => n3284);
   U1399 : OAI22_X1 port map( A1 => n51, A2 => n969, B1 => n970, B2 => n995, ZN
                           => n3285);
   U1400 : OAI22_X1 port map( A1 => n53, A2 => n969, B1 => n970, B2 => n996, ZN
                           => n3286);
   U1401 : OAI22_X1 port map( A1 => n55, A2 => n969, B1 => n970, B2 => n997, ZN
                           => n3287);
   U1402 : OAI22_X1 port map( A1 => n57, A2 => n969, B1 => n970, B2 => n998, ZN
                           => n3288);
   U1403 : OAI22_X1 port map( A1 => n59, A2 => n969, B1 => n970, B2 => n999, ZN
                           => n3289);
   U1404 : OAI22_X1 port map( A1 => n61, A2 => n969, B1 => n970, B2 => n1000, 
                           ZN => n3290);
   U1405 : OAI22_X1 port map( A1 => n63, A2 => n969, B1 => n970, B2 => n1001, 
                           ZN => n3291);
   U1406 : OAI22_X1 port map( A1 => n65, A2 => n969, B1 => n970, B2 => n1002, 
                           ZN => n3292);
   U1409 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n900, ZN 
                           => n173);
   U1410 : INV_X1 port map( A => ADD_WR(2), ZN => n900);
   U1411 : INV_X1 port map( A => n1003, ZN => n3293);
   U1412 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_0_port, ZN => n1003);
   U1413 : INV_X1 port map( A => n1006, ZN => n3294);
   U1414 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_1_port, ZN => n1006);
   U1415 : INV_X1 port map( A => n1007, ZN => n3295);
   U1416 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_2_port, ZN => n1007);
   U1417 : INV_X1 port map( A => n1008, ZN => n3296);
   U1418 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_3_port, ZN => n1008);
   U1419 : INV_X1 port map( A => n1009, ZN => n3297);
   U1420 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_4_port, ZN => n1009);
   U1421 : INV_X1 port map( A => n1010, ZN => n3298);
   U1422 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_5_port, ZN => n1010);
   U1423 : INV_X1 port map( A => n1011, ZN => n3299);
   U1424 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_6_port, ZN => n1011);
   U1425 : INV_X1 port map( A => n1012, ZN => n3300);
   U1426 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_7_port, ZN => n1012);
   U1427 : INV_X1 port map( A => n1013, ZN => n3301);
   U1428 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_8_port, ZN => n1013);
   U1429 : INV_X1 port map( A => n1014, ZN => n3302);
   U1430 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n1004, B1 => n1005, B2 => 
                           REGISTERS_3_9_port, ZN => n1014);
   U1431 : INV_X1 port map( A => n1015, ZN => n3303);
   U1432 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_10_port, ZN => n1015);
   U1433 : INV_X1 port map( A => n1016, ZN => n3304);
   U1434 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_11_port, ZN => n1016);
   U1435 : INV_X1 port map( A => n1017, ZN => n3305);
   U1436 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_12_port, ZN => n1017);
   U1437 : INV_X1 port map( A => n1018, ZN => n3306);
   U1438 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_13_port, ZN => n1018);
   U1439 : INV_X1 port map( A => n1019, ZN => n3307);
   U1440 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_14_port, ZN => n1019);
   U1441 : INV_X1 port map( A => n1020, ZN => n3308);
   U1442 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_15_port, ZN => n1020);
   U1443 : INV_X1 port map( A => n1021, ZN => n3309);
   U1444 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_16_port, ZN => n1021);
   U1445 : INV_X1 port map( A => n1022, ZN => n3310);
   U1446 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_17_port, ZN => n1022);
   U1447 : INV_X1 port map( A => n1023, ZN => n3311);
   U1448 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_18_port, ZN => n1023);
   U1449 : INV_X1 port map( A => n1024, ZN => n3312);
   U1450 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_19_port, ZN => n1024);
   U1451 : INV_X1 port map( A => n1025, ZN => n3313);
   U1452 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_20_port, ZN => n1025);
   U1453 : INV_X1 port map( A => n1026, ZN => n3314);
   U1454 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_21_port, ZN => n1026);
   U1455 : INV_X1 port map( A => n1027, ZN => n3315);
   U1456 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_22_port, ZN => n1027);
   U1457 : INV_X1 port map( A => n1028, ZN => n3316);
   U1458 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_23_port, ZN => n1028);
   U1459 : INV_X1 port map( A => n1029, ZN => n3317);
   U1460 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_24_port, ZN => n1029);
   U1461 : INV_X1 port map( A => n1030, ZN => n3318);
   U1462 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_25_port, ZN => n1030);
   U1463 : INV_X1 port map( A => n1031, ZN => n3319);
   U1464 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_26_port, ZN => n1031);
   U1465 : INV_X1 port map( A => n1032, ZN => n3320);
   U1466 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_27_port, ZN => n1032);
   U1467 : INV_X1 port map( A => n1033, ZN => n3321);
   U1468 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_28_port, ZN => n1033);
   U1469 : INV_X1 port map( A => n1034, ZN => n3322);
   U1470 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_29_port, ZN => n1034);
   U1471 : INV_X1 port map( A => n1035, ZN => n3323);
   U1472 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_30_port, ZN => n1035);
   U1473 : INV_X1 port map( A => n1036, ZN => n3324);
   U1474 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n1004, B1 => n1005, B2 =>
                           REGISTERS_3_31_port, ZN => n1036);
   U1477 : NOR3_X1 port map( A1 => n899, A2 => ADD_WR(2), A3 => n898, ZN => 
                           n208);
   U1478 : INV_X1 port map( A => n1037, ZN => n3325);
   U1479 : AOI22_X1 port map( A1 => DATAIN(0), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_0_port, ZN => n1037);
   U1480 : INV_X1 port map( A => n1040, ZN => n3326);
   U1481 : AOI22_X1 port map( A1 => DATAIN(1), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_1_port, ZN => n1040);
   U1482 : INV_X1 port map( A => n1041, ZN => n3327);
   U1483 : AOI22_X1 port map( A1 => DATAIN(2), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_2_port, ZN => n1041);
   U1484 : INV_X1 port map( A => n1042, ZN => n3328);
   U1485 : AOI22_X1 port map( A1 => DATAIN(3), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_3_port, ZN => n1042);
   U1486 : INV_X1 port map( A => n1043, ZN => n3329);
   U1487 : AOI22_X1 port map( A1 => DATAIN(4), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_4_port, ZN => n1043);
   U1488 : INV_X1 port map( A => n1044, ZN => n3330);
   U1489 : AOI22_X1 port map( A1 => DATAIN(5), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_5_port, ZN => n1044);
   U1490 : INV_X1 port map( A => n1045, ZN => n3331);
   U1491 : AOI22_X1 port map( A1 => DATAIN(6), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_6_port, ZN => n1045);
   U1492 : INV_X1 port map( A => n1046, ZN => n3332);
   U1493 : AOI22_X1 port map( A1 => DATAIN(7), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_7_port, ZN => n1046);
   U1494 : INV_X1 port map( A => n1047, ZN => n3333);
   U1495 : AOI22_X1 port map( A1 => DATAIN(8), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_8_port, ZN => n1047);
   U1496 : INV_X1 port map( A => n1048, ZN => n3334);
   U1497 : AOI22_X1 port map( A1 => DATAIN(9), A2 => n1038, B1 => n1039, B2 => 
                           REGISTERS_2_9_port, ZN => n1048);
   U1498 : INV_X1 port map( A => n1049, ZN => n3335);
   U1499 : AOI22_X1 port map( A1 => DATAIN(10), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_10_port, ZN => n1049);
   U1500 : INV_X1 port map( A => n1050, ZN => n3336);
   U1501 : AOI22_X1 port map( A1 => DATAIN(11), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_11_port, ZN => n1050);
   U1502 : INV_X1 port map( A => n1051, ZN => n3337);
   U1503 : AOI22_X1 port map( A1 => DATAIN(12), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_12_port, ZN => n1051);
   U1504 : INV_X1 port map( A => n1052, ZN => n3338);
   U1505 : AOI22_X1 port map( A1 => DATAIN(13), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_13_port, ZN => n1052);
   U1506 : INV_X1 port map( A => n1053, ZN => n3339);
   U1507 : AOI22_X1 port map( A1 => DATAIN(14), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_14_port, ZN => n1053);
   U1508 : INV_X1 port map( A => n1054, ZN => n3340);
   U1509 : AOI22_X1 port map( A1 => DATAIN(15), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_15_port, ZN => n1054);
   U1510 : INV_X1 port map( A => n1055, ZN => n3341);
   U1511 : AOI22_X1 port map( A1 => DATAIN(16), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_16_port, ZN => n1055);
   U1512 : INV_X1 port map( A => n1056, ZN => n3342);
   U1513 : AOI22_X1 port map( A1 => DATAIN(17), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_17_port, ZN => n1056);
   U1514 : INV_X1 port map( A => n1057, ZN => n3343);
   U1515 : AOI22_X1 port map( A1 => DATAIN(18), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_18_port, ZN => n1057);
   U1516 : INV_X1 port map( A => n1058, ZN => n3344);
   U1517 : AOI22_X1 port map( A1 => DATAIN(19), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_19_port, ZN => n1058);
   U1518 : INV_X1 port map( A => n1059, ZN => n3345);
   U1519 : AOI22_X1 port map( A1 => DATAIN(20), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_20_port, ZN => n1059);
   U1520 : INV_X1 port map( A => n1060, ZN => n3346);
   U1521 : AOI22_X1 port map( A1 => DATAIN(21), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_21_port, ZN => n1060);
   U1522 : INV_X1 port map( A => n1061, ZN => n3347);
   U1523 : AOI22_X1 port map( A1 => DATAIN(22), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_22_port, ZN => n1061);
   U1524 : INV_X1 port map( A => n1062, ZN => n3348);
   U1525 : AOI22_X1 port map( A1 => DATAIN(23), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_23_port, ZN => n1062);
   U1526 : INV_X1 port map( A => n1063, ZN => n3349);
   U1527 : AOI22_X1 port map( A1 => DATAIN(24), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_24_port, ZN => n1063);
   U1528 : INV_X1 port map( A => n1064, ZN => n3350);
   U1529 : AOI22_X1 port map( A1 => DATAIN(25), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_25_port, ZN => n1064);
   U1530 : INV_X1 port map( A => n1065, ZN => n3351);
   U1531 : AOI22_X1 port map( A1 => DATAIN(26), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_26_port, ZN => n1065);
   U1532 : INV_X1 port map( A => n1066, ZN => n3352);
   U1533 : AOI22_X1 port map( A1 => DATAIN(27), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_27_port, ZN => n1066);
   U1534 : INV_X1 port map( A => n1067, ZN => n3353);
   U1535 : AOI22_X1 port map( A1 => DATAIN(28), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_28_port, ZN => n1067);
   U1536 : INV_X1 port map( A => n1068, ZN => n3354);
   U1537 : AOI22_X1 port map( A1 => DATAIN(29), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_29_port, ZN => n1068);
   U1538 : INV_X1 port map( A => n1069, ZN => n3355);
   U1539 : AOI22_X1 port map( A1 => DATAIN(30), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_30_port, ZN => n1069);
   U1540 : INV_X1 port map( A => n1070, ZN => n3356);
   U1541 : AOI22_X1 port map( A1 => DATAIN(31), A2 => n1038, B1 => n1039, B2 =>
                           REGISTERS_2_31_port, ZN => n1070);
   U1544 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n898, ZN 
                           => n243);
   U1545 : INV_X1 port map( A => ADD_WR(1), ZN => n898);
   U1546 : OAI22_X1 port map( A1 => n2, A2 => n1071, B1 => n1072, B2 => n1073, 
                           ZN => n3357);
   U1547 : OAI22_X1 port map( A1 => n5, A2 => n1071, B1 => n1072, B2 => n1074, 
                           ZN => n3358);
   U1548 : OAI22_X1 port map( A1 => n7, A2 => n1071, B1 => n1072, B2 => n1075, 
                           ZN => n3359);
   U1549 : OAI22_X1 port map( A1 => n9, A2 => n1071, B1 => n1072, B2 => n1076, 
                           ZN => n3360);
   U1550 : OAI22_X1 port map( A1 => n11, A2 => n1071, B1 => n1072, B2 => n1077,
                           ZN => n3361);
   U1551 : OAI22_X1 port map( A1 => n13, A2 => n1071, B1 => n1072, B2 => n1078,
                           ZN => n3362);
   U1552 : OAI22_X1 port map( A1 => n15, A2 => n1071, B1 => n1072, B2 => n1079,
                           ZN => n3363);
   U1553 : OAI22_X1 port map( A1 => n17, A2 => n1071, B1 => n1072, B2 => n1080,
                           ZN => n3364);
   U1554 : OAI22_X1 port map( A1 => n19, A2 => n1071, B1 => n1072, B2 => n1081,
                           ZN => n3365);
   U1555 : OAI22_X1 port map( A1 => n21, A2 => n1071, B1 => n1072, B2 => n1082,
                           ZN => n3366);
   U1556 : OAI22_X1 port map( A1 => n23, A2 => n1071, B1 => n1072, B2 => n1083,
                           ZN => n3367);
   U1557 : OAI22_X1 port map( A1 => n25, A2 => n1071, B1 => n1072, B2 => n1084,
                           ZN => n3368);
   U1558 : OAI22_X1 port map( A1 => n27, A2 => n1071, B1 => n1072, B2 => n1085,
                           ZN => n3369);
   U1559 : OAI22_X1 port map( A1 => n29, A2 => n1071, B1 => n1072, B2 => n1086,
                           ZN => n3370);
   U1560 : OAI22_X1 port map( A1 => n31, A2 => n1071, B1 => n1072, B2 => n1087,
                           ZN => n3371);
   U1561 : OAI22_X1 port map( A1 => n33, A2 => n1071, B1 => n1072, B2 => n1088,
                           ZN => n3372);
   U1562 : OAI22_X1 port map( A1 => n35, A2 => n1071, B1 => n1072, B2 => n1089,
                           ZN => n3373);
   U1563 : OAI22_X1 port map( A1 => n37, A2 => n1071, B1 => n1072, B2 => n1090,
                           ZN => n3374);
   U1564 : OAI22_X1 port map( A1 => n39, A2 => n1071, B1 => n1072, B2 => n1091,
                           ZN => n3375);
   U1565 : OAI22_X1 port map( A1 => n41, A2 => n1071, B1 => n1072, B2 => n1092,
                           ZN => n3376);
   U1566 : OAI22_X1 port map( A1 => n43, A2 => n1071, B1 => n1072, B2 => n1093,
                           ZN => n3377);
   U1567 : OAI22_X1 port map( A1 => n45, A2 => n1071, B1 => n1072, B2 => n1094,
                           ZN => n3378);
   U1568 : OAI22_X1 port map( A1 => n47, A2 => n1071, B1 => n1072, B2 => n1095,
                           ZN => n3379);
   U1569 : OAI22_X1 port map( A1 => n49, A2 => n1071, B1 => n1072, B2 => n1096,
                           ZN => n3380);
   U1570 : OAI22_X1 port map( A1 => n51, A2 => n1071, B1 => n1072, B2 => n1097,
                           ZN => n3381);
   U1571 : OAI22_X1 port map( A1 => n53, A2 => n1071, B1 => n1072, B2 => n1098,
                           ZN => n3382);
   U1572 : OAI22_X1 port map( A1 => n55, A2 => n1071, B1 => n1072, B2 => n1099,
                           ZN => n3383);
   U1573 : OAI22_X1 port map( A1 => n57, A2 => n1071, B1 => n1072, B2 => n1100,
                           ZN => n3384);
   U1574 : OAI22_X1 port map( A1 => n59, A2 => n1071, B1 => n1072, B2 => n1101,
                           ZN => n3385);
   U1575 : OAI22_X1 port map( A1 => n61, A2 => n1071, B1 => n1072, B2 => n1102,
                           ZN => n3386);
   U1576 : OAI22_X1 port map( A1 => n63, A2 => n1071, B1 => n1072, B2 => n1103,
                           ZN => n3387);
   U1577 : OAI22_X1 port map( A1 => n65, A2 => n1071, B1 => n1072, B2 => n1104,
                           ZN => n3388);
   U1580 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n899, ZN 
                           => n278);
   U1581 : INV_X1 port map( A => ADD_WR(0), ZN => n899);
   U1582 : OAI22_X1 port map( A1 => n2, A2 => n1105, B1 => n1106, B2 => n1107, 
                           ZN => n3389);
   U1583 : INV_X1 port map( A => DATAIN(0), ZN => n2);
   U1584 : OAI22_X1 port map( A1 => n5, A2 => n1105, B1 => n1106, B2 => n1108, 
                           ZN => n3390);
   U1585 : INV_X1 port map( A => DATAIN(1), ZN => n5);
   U1586 : OAI22_X1 port map( A1 => n7, A2 => n1105, B1 => n1106, B2 => n1109, 
                           ZN => n3391);
   U1587 : INV_X1 port map( A => DATAIN(2), ZN => n7);
   U1588 : OAI22_X1 port map( A1 => n9, A2 => n1105, B1 => n1106, B2 => n1110, 
                           ZN => n3392);
   U1589 : INV_X1 port map( A => DATAIN(3), ZN => n9);
   U1590 : OAI22_X1 port map( A1 => n11, A2 => n1105, B1 => n1106, B2 => n1111,
                           ZN => n3393);
   U1591 : INV_X1 port map( A => DATAIN(4), ZN => n11);
   U1592 : OAI22_X1 port map( A1 => n13, A2 => n1105, B1 => n1106, B2 => n1112,
                           ZN => n3394);
   U1593 : INV_X1 port map( A => DATAIN(5), ZN => n13);
   U1594 : OAI22_X1 port map( A1 => n15, A2 => n1105, B1 => n1106, B2 => n1113,
                           ZN => n3395);
   U1595 : INV_X1 port map( A => DATAIN(6), ZN => n15);
   U1596 : OAI22_X1 port map( A1 => n17, A2 => n1105, B1 => n1106, B2 => n1114,
                           ZN => n3396);
   U1597 : INV_X1 port map( A => DATAIN(7), ZN => n17);
   U1598 : OAI22_X1 port map( A1 => n19, A2 => n1105, B1 => n1106, B2 => n1115,
                           ZN => n3397);
   U1599 : INV_X1 port map( A => DATAIN(8), ZN => n19);
   U1600 : OAI22_X1 port map( A1 => n21, A2 => n1105, B1 => n1106, B2 => n1116,
                           ZN => n3398);
   U1601 : INV_X1 port map( A => DATAIN(9), ZN => n21);
   U1602 : OAI22_X1 port map( A1 => n23, A2 => n1105, B1 => n1106, B2 => n1117,
                           ZN => n3399);
   U1603 : INV_X1 port map( A => DATAIN(10), ZN => n23);
   U1604 : OAI22_X1 port map( A1 => n25, A2 => n1105, B1 => n1106, B2 => n1118,
                           ZN => n3400);
   U1605 : INV_X1 port map( A => DATAIN(11), ZN => n25);
   U1606 : OAI22_X1 port map( A1 => n27, A2 => n1105, B1 => n1106, B2 => n1119,
                           ZN => n3401);
   U1607 : INV_X1 port map( A => DATAIN(12), ZN => n27);
   U1608 : OAI22_X1 port map( A1 => n29, A2 => n1105, B1 => n1106, B2 => n1120,
                           ZN => n3402);
   U1609 : INV_X1 port map( A => DATAIN(13), ZN => n29);
   U1610 : OAI22_X1 port map( A1 => n31, A2 => n1105, B1 => n1106, B2 => n1121,
                           ZN => n3403);
   U1611 : INV_X1 port map( A => DATAIN(14), ZN => n31);
   U1612 : OAI22_X1 port map( A1 => n33, A2 => n1105, B1 => n1106, B2 => n1122,
                           ZN => n3404);
   U1613 : INV_X1 port map( A => DATAIN(15), ZN => n33);
   U1614 : OAI22_X1 port map( A1 => n35, A2 => n1105, B1 => n1106, B2 => n1123,
                           ZN => n3405);
   U1615 : INV_X1 port map( A => DATAIN(16), ZN => n35);
   U1616 : OAI22_X1 port map( A1 => n37, A2 => n1105, B1 => n1106, B2 => n1124,
                           ZN => n3406);
   U1617 : INV_X1 port map( A => DATAIN(17), ZN => n37);
   U1618 : OAI22_X1 port map( A1 => n39, A2 => n1105, B1 => n1106, B2 => n1125,
                           ZN => n3407);
   U1619 : INV_X1 port map( A => DATAIN(18), ZN => n39);
   U1620 : OAI22_X1 port map( A1 => n41, A2 => n1105, B1 => n1106, B2 => n1126,
                           ZN => n3408);
   U1621 : INV_X1 port map( A => DATAIN(19), ZN => n41);
   U1622 : OAI22_X1 port map( A1 => n43, A2 => n1105, B1 => n1106, B2 => n1127,
                           ZN => n3409);
   U1623 : INV_X1 port map( A => DATAIN(20), ZN => n43);
   U1624 : OAI22_X1 port map( A1 => n45, A2 => n1105, B1 => n1106, B2 => n1128,
                           ZN => n3410);
   U1625 : INV_X1 port map( A => DATAIN(21), ZN => n45);
   U1626 : OAI22_X1 port map( A1 => n47, A2 => n1105, B1 => n1106, B2 => n1129,
                           ZN => n3411);
   U1627 : INV_X1 port map( A => DATAIN(22), ZN => n47);
   U1628 : OAI22_X1 port map( A1 => n49, A2 => n1105, B1 => n1106, B2 => n1130,
                           ZN => n3412);
   U1629 : INV_X1 port map( A => DATAIN(23), ZN => n49);
   U1630 : OAI22_X1 port map( A1 => n51, A2 => n1105, B1 => n1106, B2 => n1131,
                           ZN => n3413);
   U1631 : INV_X1 port map( A => DATAIN(24), ZN => n51);
   U1632 : OAI22_X1 port map( A1 => n53, A2 => n1105, B1 => n1106, B2 => n1132,
                           ZN => n3414);
   U1633 : INV_X1 port map( A => DATAIN(25), ZN => n53);
   U1634 : OAI22_X1 port map( A1 => n55, A2 => n1105, B1 => n1106, B2 => n1133,
                           ZN => n3415);
   U1635 : INV_X1 port map( A => DATAIN(26), ZN => n55);
   U1636 : OAI22_X1 port map( A1 => n57, A2 => n1105, B1 => n1106, B2 => n1134,
                           ZN => n3416);
   U1637 : INV_X1 port map( A => DATAIN(27), ZN => n57);
   U1638 : OAI22_X1 port map( A1 => n59, A2 => n1105, B1 => n1106, B2 => n1135,
                           ZN => n3417);
   U1639 : INV_X1 port map( A => DATAIN(28), ZN => n59);
   U1640 : OAI22_X1 port map( A1 => n61, A2 => n1105, B1 => n1106, B2 => n1136,
                           ZN => n3418);
   U1641 : INV_X1 port map( A => DATAIN(29), ZN => n61);
   U1642 : OAI22_X1 port map( A1 => n63, A2 => n1105, B1 => n1106, B2 => n1137,
                           ZN => n3419);
   U1643 : INV_X1 port map( A => DATAIN(30), ZN => n63);
   U1644 : OAI22_X1 port map( A1 => n65, A2 => n1105, B1 => n1106, B2 => n1138,
                           ZN => n3420);
   U1647 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0),
                           ZN => n313_port);
   U1648 : AND3_X1 port map( A1 => n588, A2 => n862, A3 => n314_port, ZN => 
                           n897);
   U1649 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => wr_signal, ZN => 
                           n314_port);
   U1650 : INV_X1 port map( A => ADD_WR(4), ZN => n862);
   U1651 : INV_X1 port map( A => ADD_WR(3), ZN => n588);
   U1652 : INV_X1 port map( A => DATAIN(31), ZN => n65);
   U1653 : AOI21_X1 port map( B1 => n1139, B2 => n1140, A => N352, ZN => N351);
   U1654 : NOR4_X1 port map( A1 => n1141, A2 => n1142, A3 => n1143, A4 => n1144
                           , ZN => n1140);
   U1655 : OAI221_X1 port map( B1 => n553, B2 => n1145, C1 => n587, C2 => n1146
                           , A => n1147, ZN => n1144);
   U1656 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_31_port, B1 => 
                           n1149, B2 => REGISTERS_18_31_port, ZN => n1147);
   U1657 : OAI221_X1 port map( B1 => n417, B2 => n1150, C1 => n451, C2 => n1151
                           , A => n1152, ZN => n1143);
   U1658 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_31_port, B1 => 
                           n1154, B2 => REGISTERS_22_31_port, ZN => n1152);
   U1659 : OAI221_X1 port map( B1 => n277, B2 => n1155, C1 => n312_port, C2 => 
                           n1156, A => n1157, ZN => n1142);
   U1660 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_31_port, B1 => 
                           n1159, B2 => REGISTERS_26_31_port, ZN => n1157);
   U1661 : OAI221_X1 port map( B1 => n66, B2 => n1160, C1 => n102, C2 => n1161,
                           A => n1162, ZN => n1141);
   U1662 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_31_port, B1 => 
                           n1164, B2 => REGISTERS_28_31_port, ZN => n1162);
   U1663 : NOR4_X1 port map( A1 => n1165, A2 => n1166, A3 => n1167, A4 => n1168
                           , ZN => n1139);
   U1664 : OAI221_X1 port map( B1 => n1104, B2 => n1169, C1 => n1138, C2 => 
                           n1170, A => n1171, ZN => n1168);
   U1665 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_31_port, B1 => 
                           n1173, B2 => REGISTERS_2_31_port, ZN => n1171);
   U1666 : OAI221_X1 port map( B1 => n968, B2 => n1174, C1 => n1002, C2 => 
                           n1175, A => n1176, ZN => n1167);
   U1667 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_31_port, B1 => 
                           n1178, B2 => REGISTERS_6_31_port, ZN => n1176);
   U1668 : OAI221_X1 port map( B1 => n827, B2 => n1179, C1 => n861, C2 => n1180
                           , A => n1181, ZN => n1166);
   U1669 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_31_port, B1 => 
                           n1183, B2 => REGISTERS_10_31_port, ZN => n1181);
   U1670 : OAI221_X1 port map( B1 => n691, B2 => n1184, C1 => n725, C2 => n1185
                           , A => n1186, ZN => n1165);
   U1671 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_31_port, B1 => 
                           n1188, B2 => REGISTERS_14_31_port, ZN => n1186);
   U1672 : AOI21_X1 port map( B1 => n1189, B2 => n1190, A => N352, ZN => N350);
   U1673 : NOR4_X1 port map( A1 => n1191, A2 => n1192, A3 => n1193, A4 => n1194
                           , ZN => n1190);
   U1674 : OAI221_X1 port map( B1 => n552, B2 => n1145, C1 => n586, C2 => n1146
                           , A => n1195, ZN => n1194);
   U1675 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_30_port, B1 => 
                           n1149, B2 => REGISTERS_18_30_port, ZN => n1195);
   U1676 : OAI221_X1 port map( B1 => n416, B2 => n1150, C1 => n450, C2 => n1151
                           , A => n1196, ZN => n1193);
   U1677 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_30_port, B1 => 
                           n1154, B2 => REGISTERS_22_30_port, ZN => n1196);
   U1678 : OAI221_X1 port map( B1 => n276, B2 => n1155, C1 => n311_port, C2 => 
                           n1156, A => n1197, ZN => n1192);
   U1679 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_30_port, B1 => 
                           n1159, B2 => REGISTERS_26_30_port, ZN => n1197);
   U1680 : OAI221_X1 port map( B1 => n64, B2 => n1160, C1 => n101, C2 => n1161,
                           A => n1198, ZN => n1191);
   U1681 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_30_port, B1 => 
                           n1164, B2 => REGISTERS_28_30_port, ZN => n1198);
   U1682 : NOR4_X1 port map( A1 => n1199, A2 => n1200, A3 => n1201, A4 => n1202
                           , ZN => n1189);
   U1683 : OAI221_X1 port map( B1 => n1103, B2 => n1169, C1 => n1137, C2 => 
                           n1170, A => n1203, ZN => n1202);
   U1684 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_30_port, B1 => 
                           n1173, B2 => REGISTERS_2_30_port, ZN => n1203);
   U1685 : OAI221_X1 port map( B1 => n967, B2 => n1174, C1 => n1001, C2 => 
                           n1175, A => n1204, ZN => n1201);
   U1686 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_30_port, B1 => 
                           n1178, B2 => REGISTERS_6_30_port, ZN => n1204);
   U1687 : OAI221_X1 port map( B1 => n826, B2 => n1179, C1 => n860, C2 => n1180
                           , A => n1205, ZN => n1200);
   U1688 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_30_port, B1 => 
                           n1183, B2 => REGISTERS_10_30_port, ZN => n1205);
   U1689 : OAI221_X1 port map( B1 => n690, B2 => n1184, C1 => n724, C2 => n1185
                           , A => n1206, ZN => n1199);
   U1690 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_30_port, B1 => 
                           n1188, B2 => REGISTERS_14_30_port, ZN => n1206);
   U1691 : AOI21_X1 port map( B1 => n1207, B2 => n1208, A => N352, ZN => N349);
   U1692 : NOR4_X1 port map( A1 => n1209, A2 => n1210, A3 => n1211, A4 => n1212
                           , ZN => n1208);
   U1693 : OAI221_X1 port map( B1 => n551, B2 => n1145, C1 => n585, C2 => n1146
                           , A => n1213, ZN => n1212);
   U1694 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_29_port, B1 => 
                           n1149, B2 => REGISTERS_18_29_port, ZN => n1213);
   U1695 : OAI221_X1 port map( B1 => n415, B2 => n1150, C1 => n449, C2 => n1151
                           , A => n1214, ZN => n1211);
   U1696 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_29_port, B1 => 
                           n1154, B2 => REGISTERS_22_29_port, ZN => n1214);
   U1697 : OAI221_X1 port map( B1 => n275, B2 => n1155, C1 => n310_port, C2 => 
                           n1156, A => n1215, ZN => n1210);
   U1698 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_29_port, B1 => 
                           n1159, B2 => REGISTERS_26_29_port, ZN => n1215);
   U1699 : OAI221_X1 port map( B1 => n62, B2 => n1160, C1 => n100, C2 => n1161,
                           A => n1216, ZN => n1209);
   U1700 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_29_port, B1 => 
                           n1164, B2 => REGISTERS_28_29_port, ZN => n1216);
   U1701 : NOR4_X1 port map( A1 => n1217, A2 => n1218, A3 => n1219, A4 => n1220
                           , ZN => n1207);
   U1702 : OAI221_X1 port map( B1 => n1102, B2 => n1169, C1 => n1136, C2 => 
                           n1170, A => n1221, ZN => n1220);
   U1703 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_29_port, B1 => 
                           n1173, B2 => REGISTERS_2_29_port, ZN => n1221);
   U1704 : OAI221_X1 port map( B1 => n966, B2 => n1174, C1 => n1000, C2 => 
                           n1175, A => n1222, ZN => n1219);
   U1705 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_29_port, B1 => 
                           n1178, B2 => REGISTERS_6_29_port, ZN => n1222);
   U1706 : OAI221_X1 port map( B1 => n825, B2 => n1179, C1 => n859, C2 => n1180
                           , A => n1223, ZN => n1218);
   U1707 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_29_port, B1 => 
                           n1183, B2 => REGISTERS_10_29_port, ZN => n1223);
   U1708 : OAI221_X1 port map( B1 => n689, B2 => n1184, C1 => n723, C2 => n1185
                           , A => n1224, ZN => n1217);
   U1709 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_29_port, B1 => 
                           n1188, B2 => REGISTERS_14_29_port, ZN => n1224);
   U1710 : AOI21_X1 port map( B1 => n1225, B2 => n1226, A => N352, ZN => N348);
   U1711 : NOR4_X1 port map( A1 => n1227, A2 => n1228, A3 => n1229, A4 => n1230
                           , ZN => n1226);
   U1712 : OAI221_X1 port map( B1 => n550, B2 => n1145, C1 => n584, C2 => n1146
                           , A => n1231, ZN => n1230);
   U1713 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_28_port, B1 => 
                           n1149, B2 => REGISTERS_18_28_port, ZN => n1231);
   U1714 : OAI221_X1 port map( B1 => n414, B2 => n1150, C1 => n448, C2 => n1151
                           , A => n1232, ZN => n1229);
   U1715 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_28_port, B1 => 
                           n1154, B2 => REGISTERS_22_28_port, ZN => n1232);
   U1716 : OAI221_X1 port map( B1 => n274, B2 => n1155, C1 => n309_port, C2 => 
                           n1156, A => n1233, ZN => n1228);
   U1717 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_28_port, B1 => 
                           n1159, B2 => REGISTERS_26_28_port, ZN => n1233);
   U1718 : OAI221_X1 port map( B1 => n60, B2 => n1160, C1 => n99, C2 => n1161, 
                           A => n1234, ZN => n1227);
   U1719 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_28_port, B1 => 
                           n1164, B2 => REGISTERS_28_28_port, ZN => n1234);
   U1720 : NOR4_X1 port map( A1 => n1235, A2 => n1236, A3 => n1237, A4 => n1238
                           , ZN => n1225);
   U1721 : OAI221_X1 port map( B1 => n1101, B2 => n1169, C1 => n1135, C2 => 
                           n1170, A => n1239, ZN => n1238);
   U1722 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_28_port, B1 => 
                           n1173, B2 => REGISTERS_2_28_port, ZN => n1239);
   U1723 : OAI221_X1 port map( B1 => n965, B2 => n1174, C1 => n999, C2 => n1175
                           , A => n1240, ZN => n1237);
   U1724 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_28_port, B1 => 
                           n1178, B2 => REGISTERS_6_28_port, ZN => n1240);
   U1725 : OAI221_X1 port map( B1 => n824, B2 => n1179, C1 => n858, C2 => n1180
                           , A => n1241, ZN => n1236);
   U1726 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_28_port, B1 => 
                           n1183, B2 => REGISTERS_10_28_port, ZN => n1241);
   U1727 : OAI221_X1 port map( B1 => n688, B2 => n1184, C1 => n722, C2 => n1185
                           , A => n1242, ZN => n1235);
   U1728 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_28_port, B1 => 
                           n1188, B2 => REGISTERS_14_28_port, ZN => n1242);
   U1729 : AOI21_X1 port map( B1 => n1243, B2 => n1244, A => N352, ZN => N347);
   U1730 : NOR4_X1 port map( A1 => n1245, A2 => n1246, A3 => n1247, A4 => n1248
                           , ZN => n1244);
   U1731 : OAI221_X1 port map( B1 => n549, B2 => n1145, C1 => n583, C2 => n1146
                           , A => n1249, ZN => n1248);
   U1732 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_27_port, B1 => 
                           n1149, B2 => REGISTERS_18_27_port, ZN => n1249);
   U1733 : OAI221_X1 port map( B1 => n413, B2 => n1150, C1 => n447, C2 => n1151
                           , A => n1250, ZN => n1247);
   U1734 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_27_port, B1 => 
                           n1154, B2 => REGISTERS_22_27_port, ZN => n1250);
   U1735 : OAI221_X1 port map( B1 => n273, B2 => n1155, C1 => n308_port, C2 => 
                           n1156, A => n1251, ZN => n1246);
   U1736 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_27_port, B1 => 
                           n1159, B2 => REGISTERS_26_27_port, ZN => n1251);
   U1737 : OAI221_X1 port map( B1 => n58, B2 => n1160, C1 => n98, C2 => n1161, 
                           A => n1252, ZN => n1245);
   U1738 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_27_port, B1 => 
                           n1164, B2 => REGISTERS_28_27_port, ZN => n1252);
   U1739 : NOR4_X1 port map( A1 => n1253, A2 => n1254, A3 => n1255, A4 => n1256
                           , ZN => n1243);
   U1740 : OAI221_X1 port map( B1 => n1100, B2 => n1169, C1 => n1134, C2 => 
                           n1170, A => n1257, ZN => n1256);
   U1741 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_27_port, B1 => 
                           n1173, B2 => REGISTERS_2_27_port, ZN => n1257);
   U1742 : OAI221_X1 port map( B1 => n964, B2 => n1174, C1 => n998, C2 => n1175
                           , A => n1258, ZN => n1255);
   U1743 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_27_port, B1 => 
                           n1178, B2 => REGISTERS_6_27_port, ZN => n1258);
   U1744 : OAI221_X1 port map( B1 => n823, B2 => n1179, C1 => n857, C2 => n1180
                           , A => n1259, ZN => n1254);
   U1745 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_27_port, B1 => 
                           n1183, B2 => REGISTERS_10_27_port, ZN => n1259);
   U1746 : OAI221_X1 port map( B1 => n687, B2 => n1184, C1 => n721, C2 => n1185
                           , A => n1260, ZN => n1253);
   U1747 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_27_port, B1 => 
                           n1188, B2 => REGISTERS_14_27_port, ZN => n1260);
   U1748 : AOI21_X1 port map( B1 => n1261, B2 => n1262, A => N352, ZN => N346);
   U1749 : NOR4_X1 port map( A1 => n1263, A2 => n1264, A3 => n1265, A4 => n1266
                           , ZN => n1262);
   U1750 : OAI221_X1 port map( B1 => n548, B2 => n1145, C1 => n582, C2 => n1146
                           , A => n1267, ZN => n1266);
   U1751 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_26_port, B1 => 
                           n1149, B2 => REGISTERS_18_26_port, ZN => n1267);
   U1752 : OAI221_X1 port map( B1 => n412, B2 => n1150, C1 => n446, C2 => n1151
                           , A => n1268, ZN => n1265);
   U1753 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_26_port, B1 => 
                           n1154, B2 => REGISTERS_22_26_port, ZN => n1268);
   U1754 : OAI221_X1 port map( B1 => n272, B2 => n1155, C1 => n307_port, C2 => 
                           n1156, A => n1269, ZN => n1264);
   U1755 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_26_port, B1 => 
                           n1159, B2 => REGISTERS_26_26_port, ZN => n1269);
   U1756 : OAI221_X1 port map( B1 => n56, B2 => n1160, C1 => n97, C2 => n1161, 
                           A => n1270, ZN => n1263);
   U1757 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_26_port, B1 => 
                           n1164, B2 => REGISTERS_28_26_port, ZN => n1270);
   U1758 : NOR4_X1 port map( A1 => n1271, A2 => n1272, A3 => n1273, A4 => n1274
                           , ZN => n1261);
   U1759 : OAI221_X1 port map( B1 => n1099, B2 => n1169, C1 => n1133, C2 => 
                           n1170, A => n1275, ZN => n1274);
   U1760 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_26_port, B1 => 
                           n1173, B2 => REGISTERS_2_26_port, ZN => n1275);
   U1761 : OAI221_X1 port map( B1 => n963, B2 => n1174, C1 => n997, C2 => n1175
                           , A => n1276, ZN => n1273);
   U1762 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_26_port, B1 => 
                           n1178, B2 => REGISTERS_6_26_port, ZN => n1276);
   U1763 : OAI221_X1 port map( B1 => n822, B2 => n1179, C1 => n856, C2 => n1180
                           , A => n1277, ZN => n1272);
   U1764 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_26_port, B1 => 
                           n1183, B2 => REGISTERS_10_26_port, ZN => n1277);
   U1765 : OAI221_X1 port map( B1 => n686, B2 => n1184, C1 => n720, C2 => n1185
                           , A => n1278, ZN => n1271);
   U1766 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_26_port, B1 => 
                           n1188, B2 => REGISTERS_14_26_port, ZN => n1278);
   U1767 : AOI21_X1 port map( B1 => n1279, B2 => n1280, A => N352, ZN => N345);
   U1768 : NOR4_X1 port map( A1 => n1281, A2 => n1282, A3 => n1283, A4 => n1284
                           , ZN => n1280);
   U1769 : OAI221_X1 port map( B1 => n547, B2 => n1145, C1 => n581, C2 => n1146
                           , A => n1285, ZN => n1284);
   U1770 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_25_port, B1 => 
                           n1149, B2 => REGISTERS_18_25_port, ZN => n1285);
   U1771 : OAI221_X1 port map( B1 => n411, B2 => n1150, C1 => n445, C2 => n1151
                           , A => n1286, ZN => n1283);
   U1772 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_25_port, B1 => 
                           n1154, B2 => REGISTERS_22_25_port, ZN => n1286);
   U1773 : OAI221_X1 port map( B1 => n271, B2 => n1155, C1 => n306_port, C2 => 
                           n1156, A => n1287, ZN => n1282);
   U1774 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_25_port, B1 => 
                           n1159, B2 => REGISTERS_26_25_port, ZN => n1287);
   U1775 : OAI221_X1 port map( B1 => n54, B2 => n1160, C1 => n96, C2 => n1161, 
                           A => n1288, ZN => n1281);
   U1776 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_25_port, B1 => 
                           n1164, B2 => REGISTERS_28_25_port, ZN => n1288);
   U1777 : NOR4_X1 port map( A1 => n1289, A2 => n1290, A3 => n1291, A4 => n1292
                           , ZN => n1279);
   U1778 : OAI221_X1 port map( B1 => n1098, B2 => n1169, C1 => n1132, C2 => 
                           n1170, A => n1293, ZN => n1292);
   U1779 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_25_port, B1 => 
                           n1173, B2 => REGISTERS_2_25_port, ZN => n1293);
   U1780 : OAI221_X1 port map( B1 => n962, B2 => n1174, C1 => n996, C2 => n1175
                           , A => n1294, ZN => n1291);
   U1781 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_25_port, B1 => 
                           n1178, B2 => REGISTERS_6_25_port, ZN => n1294);
   U1782 : OAI221_X1 port map( B1 => n821, B2 => n1179, C1 => n855, C2 => n1180
                           , A => n1295, ZN => n1290);
   U1783 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_25_port, B1 => 
                           n1183, B2 => REGISTERS_10_25_port, ZN => n1295);
   U1784 : OAI221_X1 port map( B1 => n685, B2 => n1184, C1 => n719, C2 => n1185
                           , A => n1296, ZN => n1289);
   U1785 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_25_port, B1 => 
                           n1188, B2 => REGISTERS_14_25_port, ZN => n1296);
   U1786 : AOI21_X1 port map( B1 => n1297, B2 => n1298, A => N352, ZN => N344);
   U1787 : NOR4_X1 port map( A1 => n1299, A2 => n1300, A3 => n1301, A4 => n1302
                           , ZN => n1298);
   U1788 : OAI221_X1 port map( B1 => n546, B2 => n1145, C1 => n580, C2 => n1146
                           , A => n1303, ZN => n1302);
   U1789 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_24_port, B1 => 
                           n1149, B2 => REGISTERS_18_24_port, ZN => n1303);
   U1790 : OAI221_X1 port map( B1 => n410, B2 => n1150, C1 => n444, C2 => n1151
                           , A => n1304, ZN => n1301);
   U1791 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_24_port, B1 => 
                           n1154, B2 => REGISTERS_22_24_port, ZN => n1304);
   U1792 : OAI221_X1 port map( B1 => n270, B2 => n1155, C1 => n305_port, C2 => 
                           n1156, A => n1305, ZN => n1300);
   U1793 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_24_port, B1 => 
                           n1159, B2 => REGISTERS_26_24_port, ZN => n1305);
   U1794 : OAI221_X1 port map( B1 => n52, B2 => n1160, C1 => n95, C2 => n1161, 
                           A => n1306, ZN => n1299);
   U1795 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_24_port, B1 => 
                           n1164, B2 => REGISTERS_28_24_port, ZN => n1306);
   U1796 : NOR4_X1 port map( A1 => n1307, A2 => n1308, A3 => n1309, A4 => n1310
                           , ZN => n1297);
   U1797 : OAI221_X1 port map( B1 => n1097, B2 => n1169, C1 => n1131, C2 => 
                           n1170, A => n1311, ZN => n1310);
   U1798 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_24_port, B1 => 
                           n1173, B2 => REGISTERS_2_24_port, ZN => n1311);
   U1799 : OAI221_X1 port map( B1 => n961, B2 => n1174, C1 => n995, C2 => n1175
                           , A => n1312, ZN => n1309);
   U1800 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_24_port, B1 => 
                           n1178, B2 => REGISTERS_6_24_port, ZN => n1312);
   U1801 : OAI221_X1 port map( B1 => n820, B2 => n1179, C1 => n854, C2 => n1180
                           , A => n1313, ZN => n1308);
   U1802 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_24_port, B1 => 
                           n1183, B2 => REGISTERS_10_24_port, ZN => n1313);
   U1803 : OAI221_X1 port map( B1 => n684, B2 => n1184, C1 => n718, C2 => n1185
                           , A => n1314, ZN => n1307);
   U1804 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_24_port, B1 => 
                           n1188, B2 => REGISTERS_14_24_port, ZN => n1314);
   U1805 : AOI21_X1 port map( B1 => n1315, B2 => n1316, A => N352, ZN => N343);
   U1806 : NOR4_X1 port map( A1 => n1317, A2 => n1318, A3 => n1319, A4 => n1320
                           , ZN => n1316);
   U1807 : OAI221_X1 port map( B1 => n545, B2 => n1145, C1 => n579, C2 => n1146
                           , A => n1321, ZN => n1320);
   U1808 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_23_port, B1 => 
                           n1149, B2 => REGISTERS_18_23_port, ZN => n1321);
   U1809 : OAI221_X1 port map( B1 => n409, B2 => n1150, C1 => n443, C2 => n1151
                           , A => n1322, ZN => n1319);
   U1810 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_23_port, B1 => 
                           n1154, B2 => REGISTERS_22_23_port, ZN => n1322);
   U1811 : OAI221_X1 port map( B1 => n269, B2 => n1155, C1 => n304_port, C2 => 
                           n1156, A => n1323, ZN => n1318);
   U1812 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_23_port, B1 => 
                           n1159, B2 => REGISTERS_26_23_port, ZN => n1323);
   U1813 : OAI221_X1 port map( B1 => n50, B2 => n1160, C1 => n94, C2 => n1161, 
                           A => n1324, ZN => n1317);
   U1814 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_23_port, B1 => 
                           n1164, B2 => REGISTERS_28_23_port, ZN => n1324);
   U1815 : NOR4_X1 port map( A1 => n1325, A2 => n1326, A3 => n1327, A4 => n1328
                           , ZN => n1315);
   U1816 : OAI221_X1 port map( B1 => n1096, B2 => n1169, C1 => n1130, C2 => 
                           n1170, A => n1329, ZN => n1328);
   U1817 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_23_port, B1 => 
                           n1173, B2 => REGISTERS_2_23_port, ZN => n1329);
   U1818 : OAI221_X1 port map( B1 => n960, B2 => n1174, C1 => n994, C2 => n1175
                           , A => n1330, ZN => n1327);
   U1819 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_23_port, B1 => 
                           n1178, B2 => REGISTERS_6_23_port, ZN => n1330);
   U1820 : OAI221_X1 port map( B1 => n819, B2 => n1179, C1 => n853, C2 => n1180
                           , A => n1331, ZN => n1326);
   U1821 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_23_port, B1 => 
                           n1183, B2 => REGISTERS_10_23_port, ZN => n1331);
   U1822 : OAI221_X1 port map( B1 => n683, B2 => n1184, C1 => n717, C2 => n1185
                           , A => n1332, ZN => n1325);
   U1823 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_23_port, B1 => 
                           n1188, B2 => REGISTERS_14_23_port, ZN => n1332);
   U1824 : AOI21_X1 port map( B1 => n1333, B2 => n1334, A => N352, ZN => N342);
   U1825 : NOR4_X1 port map( A1 => n1335, A2 => n1336, A3 => n1337, A4 => n1338
                           , ZN => n1334);
   U1826 : OAI221_X1 port map( B1 => n544, B2 => n1145, C1 => n578, C2 => n1146
                           , A => n1339, ZN => n1338);
   U1827 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_22_port, B1 => 
                           n1149, B2 => REGISTERS_18_22_port, ZN => n1339);
   U1828 : OAI221_X1 port map( B1 => n408, B2 => n1150, C1 => n442, C2 => n1151
                           , A => n1340, ZN => n1337);
   U1829 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_22_port, B1 => 
                           n1154, B2 => REGISTERS_22_22_port, ZN => n1340);
   U1830 : OAI221_X1 port map( B1 => n268, B2 => n1155, C1 => n303_port, C2 => 
                           n1156, A => n1341, ZN => n1336);
   U1831 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_22_port, B1 => 
                           n1159, B2 => REGISTERS_26_22_port, ZN => n1341);
   U1832 : OAI221_X1 port map( B1 => n48, B2 => n1160, C1 => n93, C2 => n1161, 
                           A => n1342, ZN => n1335);
   U1833 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_22_port, B1 => 
                           n1164, B2 => REGISTERS_28_22_port, ZN => n1342);
   U1834 : NOR4_X1 port map( A1 => n1343, A2 => n1344, A3 => n1345, A4 => n1346
                           , ZN => n1333);
   U1835 : OAI221_X1 port map( B1 => n1095, B2 => n1169, C1 => n1129, C2 => 
                           n1170, A => n1347, ZN => n1346);
   U1836 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_22_port, B1 => 
                           n1173, B2 => REGISTERS_2_22_port, ZN => n1347);
   U1837 : OAI221_X1 port map( B1 => n959, B2 => n1174, C1 => n993, C2 => n1175
                           , A => n1348, ZN => n1345);
   U1838 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_22_port, B1 => 
                           n1178, B2 => REGISTERS_6_22_port, ZN => n1348);
   U1839 : OAI221_X1 port map( B1 => n818, B2 => n1179, C1 => n852, C2 => n1180
                           , A => n1349, ZN => n1344);
   U1840 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_22_port, B1 => 
                           n1183, B2 => REGISTERS_10_22_port, ZN => n1349);
   U1841 : OAI221_X1 port map( B1 => n682, B2 => n1184, C1 => n716, C2 => n1185
                           , A => n1350, ZN => n1343);
   U1842 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_22_port, B1 => 
                           n1188, B2 => REGISTERS_14_22_port, ZN => n1350);
   U1843 : AOI21_X1 port map( B1 => n1351, B2 => n1352, A => N352, ZN => N341);
   U1844 : NOR4_X1 port map( A1 => n1353, A2 => n1354, A3 => n1355, A4 => n1356
                           , ZN => n1352);
   U1845 : OAI221_X1 port map( B1 => n543, B2 => n1145, C1 => n577, C2 => n1146
                           , A => n1357, ZN => n1356);
   U1846 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_21_port, B1 => 
                           n1149, B2 => REGISTERS_18_21_port, ZN => n1357);
   U1847 : OAI221_X1 port map( B1 => n407, B2 => n1150, C1 => n441, C2 => n1151
                           , A => n1358, ZN => n1355);
   U1848 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_21_port, B1 => 
                           n1154, B2 => REGISTERS_22_21_port, ZN => n1358);
   U1849 : OAI221_X1 port map( B1 => n267, B2 => n1155, C1 => n302_port, C2 => 
                           n1156, A => n1359, ZN => n1354);
   U1850 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_21_port, B1 => 
                           n1159, B2 => REGISTERS_26_21_port, ZN => n1359);
   U1851 : OAI221_X1 port map( B1 => n46, B2 => n1160, C1 => n92, C2 => n1161, 
                           A => n1360, ZN => n1353);
   U1852 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_21_port, B1 => 
                           n1164, B2 => REGISTERS_28_21_port, ZN => n1360);
   U1853 : NOR4_X1 port map( A1 => n1361, A2 => n1362, A3 => n1363, A4 => n1364
                           , ZN => n1351);
   U1854 : OAI221_X1 port map( B1 => n1094, B2 => n1169, C1 => n1128, C2 => 
                           n1170, A => n1365, ZN => n1364);
   U1855 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_21_port, B1 => 
                           n1173, B2 => REGISTERS_2_21_port, ZN => n1365);
   U1856 : OAI221_X1 port map( B1 => n958, B2 => n1174, C1 => n992, C2 => n1175
                           , A => n1366, ZN => n1363);
   U1857 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_21_port, B1 => 
                           n1178, B2 => REGISTERS_6_21_port, ZN => n1366);
   U1858 : OAI221_X1 port map( B1 => n817, B2 => n1179, C1 => n851, C2 => n1180
                           , A => n1367, ZN => n1362);
   U1859 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_21_port, B1 => 
                           n1183, B2 => REGISTERS_10_21_port, ZN => n1367);
   U1860 : OAI221_X1 port map( B1 => n681, B2 => n1184, C1 => n715, C2 => n1185
                           , A => n1368, ZN => n1361);
   U1861 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_21_port, B1 => 
                           n1188, B2 => REGISTERS_14_21_port, ZN => n1368);
   U1862 : AOI21_X1 port map( B1 => n1369, B2 => n1370, A => N352, ZN => N340);
   U1863 : NOR4_X1 port map( A1 => n1371, A2 => n1372, A3 => n1373, A4 => n1374
                           , ZN => n1370);
   U1864 : OAI221_X1 port map( B1 => n542, B2 => n1145, C1 => n576, C2 => n1146
                           , A => n1375, ZN => n1374);
   U1865 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_20_port, B1 => 
                           n1149, B2 => REGISTERS_18_20_port, ZN => n1375);
   U1866 : OAI221_X1 port map( B1 => n406, B2 => n1150, C1 => n440, C2 => n1151
                           , A => n1376, ZN => n1373);
   U1867 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_20_port, B1 => 
                           n1154, B2 => REGISTERS_22_20_port, ZN => n1376);
   U1868 : OAI221_X1 port map( B1 => n266, B2 => n1155, C1 => n301_port, C2 => 
                           n1156, A => n1377, ZN => n1372);
   U1869 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_20_port, B1 => 
                           n1159, B2 => REGISTERS_26_20_port, ZN => n1377);
   U1870 : OAI221_X1 port map( B1 => n44, B2 => n1160, C1 => n91, C2 => n1161, 
                           A => n1378, ZN => n1371);
   U1871 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_20_port, B1 => 
                           n1164, B2 => REGISTERS_28_20_port, ZN => n1378);
   U1872 : NOR4_X1 port map( A1 => n1379, A2 => n1380, A3 => n1381, A4 => n1382
                           , ZN => n1369);
   U1873 : OAI221_X1 port map( B1 => n1093, B2 => n1169, C1 => n1127, C2 => 
                           n1170, A => n1383, ZN => n1382);
   U1874 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_20_port, B1 => 
                           n1173, B2 => REGISTERS_2_20_port, ZN => n1383);
   U1875 : OAI221_X1 port map( B1 => n957, B2 => n1174, C1 => n991, C2 => n1175
                           , A => n1384, ZN => n1381);
   U1876 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_20_port, B1 => 
                           n1178, B2 => REGISTERS_6_20_port, ZN => n1384);
   U1877 : OAI221_X1 port map( B1 => n816, B2 => n1179, C1 => n850, C2 => n1180
                           , A => n1385, ZN => n1380);
   U1878 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_20_port, B1 => 
                           n1183, B2 => REGISTERS_10_20_port, ZN => n1385);
   U1879 : OAI221_X1 port map( B1 => n680, B2 => n1184, C1 => n714, C2 => n1185
                           , A => n1386, ZN => n1379);
   U1880 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_20_port, B1 => 
                           n1188, B2 => REGISTERS_14_20_port, ZN => n1386);
   U1881 : AOI21_X1 port map( B1 => n1387, B2 => n1388, A => N352, ZN => N339);
   U1882 : NOR4_X1 port map( A1 => n1389, A2 => n1390, A3 => n1391, A4 => n1392
                           , ZN => n1388);
   U1883 : OAI221_X1 port map( B1 => n541, B2 => n1145, C1 => n575, C2 => n1146
                           , A => n1393, ZN => n1392);
   U1884 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_19_port, B1 => 
                           n1149, B2 => REGISTERS_18_19_port, ZN => n1393);
   U1885 : OAI221_X1 port map( B1 => n405, B2 => n1150, C1 => n439, C2 => n1151
                           , A => n1394, ZN => n1391);
   U1886 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_19_port, B1 => 
                           n1154, B2 => REGISTERS_22_19_port, ZN => n1394);
   U1887 : OAI221_X1 port map( B1 => n265, B2 => n1155, C1 => n300_port, C2 => 
                           n1156, A => n1395, ZN => n1390);
   U1888 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_19_port, B1 => 
                           n1159, B2 => REGISTERS_26_19_port, ZN => n1395);
   U1889 : OAI221_X1 port map( B1 => n42, B2 => n1160, C1 => n90, C2 => n1161, 
                           A => n1396, ZN => n1389);
   U1890 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_19_port, B1 => 
                           n1164, B2 => REGISTERS_28_19_port, ZN => n1396);
   U1891 : NOR4_X1 port map( A1 => n1397, A2 => n1398, A3 => n1399, A4 => n1400
                           , ZN => n1387);
   U1892 : OAI221_X1 port map( B1 => n1092, B2 => n1169, C1 => n1126, C2 => 
                           n1170, A => n1401, ZN => n1400);
   U1893 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_19_port, B1 => 
                           n1173, B2 => REGISTERS_2_19_port, ZN => n1401);
   U1894 : OAI221_X1 port map( B1 => n956, B2 => n1174, C1 => n990, C2 => n1175
                           , A => n1402, ZN => n1399);
   U1895 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_19_port, B1 => 
                           n1178, B2 => REGISTERS_6_19_port, ZN => n1402);
   U1896 : OAI221_X1 port map( B1 => n815, B2 => n1179, C1 => n849, C2 => n1180
                           , A => n1403, ZN => n1398);
   U1897 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_19_port, B1 => 
                           n1183, B2 => REGISTERS_10_19_port, ZN => n1403);
   U1898 : OAI221_X1 port map( B1 => n679, B2 => n1184, C1 => n713, C2 => n1185
                           , A => n1404, ZN => n1397);
   U1899 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_19_port, B1 => 
                           n1188, B2 => REGISTERS_14_19_port, ZN => n1404);
   U1900 : AOI21_X1 port map( B1 => n1405, B2 => n1406, A => N352, ZN => N338);
   U1901 : NOR4_X1 port map( A1 => n1407, A2 => n1408, A3 => n1409, A4 => n1410
                           , ZN => n1406);
   U1902 : OAI221_X1 port map( B1 => n540, B2 => n1145, C1 => n574, C2 => n1146
                           , A => n1411, ZN => n1410);
   U1903 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_18_port, B1 => 
                           n1149, B2 => REGISTERS_18_18_port, ZN => n1411);
   U1904 : OAI221_X1 port map( B1 => n404, B2 => n1150, C1 => n438, C2 => n1151
                           , A => n1412, ZN => n1409);
   U1905 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_18_port, B1 => 
                           n1154, B2 => REGISTERS_22_18_port, ZN => n1412);
   U1906 : OAI221_X1 port map( B1 => n264, B2 => n1155, C1 => n299_port, C2 => 
                           n1156, A => n1413, ZN => n1408);
   U1907 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_18_port, B1 => 
                           n1159, B2 => REGISTERS_26_18_port, ZN => n1413);
   U1908 : OAI221_X1 port map( B1 => n40, B2 => n1160, C1 => n89, C2 => n1161, 
                           A => n1414, ZN => n1407);
   U1909 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_18_port, B1 => 
                           n1164, B2 => REGISTERS_28_18_port, ZN => n1414);
   U1910 : NOR4_X1 port map( A1 => n1415, A2 => n1416, A3 => n1417, A4 => n1418
                           , ZN => n1405);
   U1911 : OAI221_X1 port map( B1 => n1091, B2 => n1169, C1 => n1125, C2 => 
                           n1170, A => n1419, ZN => n1418);
   U1912 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_18_port, B1 => 
                           n1173, B2 => REGISTERS_2_18_port, ZN => n1419);
   U1913 : OAI221_X1 port map( B1 => n955, B2 => n1174, C1 => n989, C2 => n1175
                           , A => n1420, ZN => n1417);
   U1914 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_18_port, B1 => 
                           n1178, B2 => REGISTERS_6_18_port, ZN => n1420);
   U1915 : OAI221_X1 port map( B1 => n814, B2 => n1179, C1 => n848, C2 => n1180
                           , A => n1421, ZN => n1416);
   U1916 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_18_port, B1 => 
                           n1183, B2 => REGISTERS_10_18_port, ZN => n1421);
   U1917 : OAI221_X1 port map( B1 => n678, B2 => n1184, C1 => n712, C2 => n1185
                           , A => n1422, ZN => n1415);
   U1918 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_18_port, B1 => 
                           n1188, B2 => REGISTERS_14_18_port, ZN => n1422);
   U1919 : AOI21_X1 port map( B1 => n1423, B2 => n1424, A => N352, ZN => N337);
   U1920 : NOR4_X1 port map( A1 => n1425, A2 => n1426, A3 => n1427, A4 => n1428
                           , ZN => n1424);
   U1921 : OAI221_X1 port map( B1 => n539, B2 => n1145, C1 => n573, C2 => n1146
                           , A => n1429, ZN => n1428);
   U1922 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_17_port, B1 => 
                           n1149, B2 => REGISTERS_18_17_port, ZN => n1429);
   U1923 : OAI221_X1 port map( B1 => n403, B2 => n1150, C1 => n437, C2 => n1151
                           , A => n1430, ZN => n1427);
   U1924 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_17_port, B1 => 
                           n1154, B2 => REGISTERS_22_17_port, ZN => n1430);
   U1925 : OAI221_X1 port map( B1 => n263, B2 => n1155, C1 => n298_port, C2 => 
                           n1156, A => n1431, ZN => n1426);
   U1926 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_17_port, B1 => 
                           n1159, B2 => REGISTERS_26_17_port, ZN => n1431);
   U1927 : OAI221_X1 port map( B1 => n38, B2 => n1160, C1 => n88, C2 => n1161, 
                           A => n1432, ZN => n1425);
   U1928 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_17_port, B1 => 
                           n1164, B2 => REGISTERS_28_17_port, ZN => n1432);
   U1929 : NOR4_X1 port map( A1 => n1433, A2 => n1434, A3 => n1435, A4 => n1436
                           , ZN => n1423);
   U1930 : OAI221_X1 port map( B1 => n1090, B2 => n1169, C1 => n1124, C2 => 
                           n1170, A => n1437, ZN => n1436);
   U1931 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_17_port, B1 => 
                           n1173, B2 => REGISTERS_2_17_port, ZN => n1437);
   U1932 : OAI221_X1 port map( B1 => n954, B2 => n1174, C1 => n988, C2 => n1175
                           , A => n1438, ZN => n1435);
   U1933 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_17_port, B1 => 
                           n1178, B2 => REGISTERS_6_17_port, ZN => n1438);
   U1934 : OAI221_X1 port map( B1 => n813, B2 => n1179, C1 => n847, C2 => n1180
                           , A => n1439, ZN => n1434);
   U1935 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_17_port, B1 => 
                           n1183, B2 => REGISTERS_10_17_port, ZN => n1439);
   U1936 : OAI221_X1 port map( B1 => n677, B2 => n1184, C1 => n711, C2 => n1185
                           , A => n1440, ZN => n1433);
   U1937 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_17_port, B1 => 
                           n1188, B2 => REGISTERS_14_17_port, ZN => n1440);
   U1938 : AOI21_X1 port map( B1 => n1441, B2 => n1442, A => N352, ZN => N336);
   U1939 : NOR4_X1 port map( A1 => n1443, A2 => n1444, A3 => n1445, A4 => n1446
                           , ZN => n1442);
   U1940 : OAI221_X1 port map( B1 => n538, B2 => n1145, C1 => n572, C2 => n1146
                           , A => n1447, ZN => n1446);
   U1941 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_16_port, B1 => 
                           n1149, B2 => REGISTERS_18_16_port, ZN => n1447);
   U1942 : OAI221_X1 port map( B1 => n402, B2 => n1150, C1 => n436, C2 => n1151
                           , A => n1448, ZN => n1445);
   U1943 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_16_port, B1 => 
                           n1154, B2 => REGISTERS_22_16_port, ZN => n1448);
   U1944 : OAI221_X1 port map( B1 => n262, B2 => n1155, C1 => n297_port, C2 => 
                           n1156, A => n1449, ZN => n1444);
   U1945 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_16_port, B1 => 
                           n1159, B2 => REGISTERS_26_16_port, ZN => n1449);
   U1946 : OAI221_X1 port map( B1 => n36, B2 => n1160, C1 => n87, C2 => n1161, 
                           A => n1450, ZN => n1443);
   U1947 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_16_port, B1 => 
                           n1164, B2 => REGISTERS_28_16_port, ZN => n1450);
   U1948 : NOR4_X1 port map( A1 => n1451, A2 => n1452, A3 => n1453, A4 => n1454
                           , ZN => n1441);
   U1949 : OAI221_X1 port map( B1 => n1089, B2 => n1169, C1 => n1123, C2 => 
                           n1170, A => n1455, ZN => n1454);
   U1950 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_16_port, B1 => 
                           n1173, B2 => REGISTERS_2_16_port, ZN => n1455);
   U1951 : OAI221_X1 port map( B1 => n953, B2 => n1174, C1 => n987, C2 => n1175
                           , A => n1456, ZN => n1453);
   U1952 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_16_port, B1 => 
                           n1178, B2 => REGISTERS_6_16_port, ZN => n1456);
   U1953 : OAI221_X1 port map( B1 => n812, B2 => n1179, C1 => n846, C2 => n1180
                           , A => n1457, ZN => n1452);
   U1954 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_16_port, B1 => 
                           n1183, B2 => REGISTERS_10_16_port, ZN => n1457);
   U1955 : OAI221_X1 port map( B1 => n676, B2 => n1184, C1 => n710, C2 => n1185
                           , A => n1458, ZN => n1451);
   U1956 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_16_port, B1 => 
                           n1188, B2 => REGISTERS_14_16_port, ZN => n1458);
   U1957 : AOI21_X1 port map( B1 => n1459, B2 => n1460, A => N352, ZN => N335);
   U1958 : NOR4_X1 port map( A1 => n1461, A2 => n1462, A3 => n1463, A4 => n1464
                           , ZN => n1460);
   U1959 : OAI221_X1 port map( B1 => n537, B2 => n1145, C1 => n571, C2 => n1146
                           , A => n1465, ZN => n1464);
   U1960 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_15_port, B1 => 
                           n1149, B2 => REGISTERS_18_15_port, ZN => n1465);
   U1961 : OAI221_X1 port map( B1 => n401, B2 => n1150, C1 => n435, C2 => n1151
                           , A => n1466, ZN => n1463);
   U1962 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_15_port, B1 => 
                           n1154, B2 => REGISTERS_22_15_port, ZN => n1466);
   U1963 : OAI221_X1 port map( B1 => n261, B2 => n1155, C1 => n296_port, C2 => 
                           n1156, A => n1467, ZN => n1462);
   U1964 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_15_port, B1 => 
                           n1159, B2 => REGISTERS_26_15_port, ZN => n1467);
   U1965 : OAI221_X1 port map( B1 => n34, B2 => n1160, C1 => n86, C2 => n1161, 
                           A => n1468, ZN => n1461);
   U1966 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_15_port, B1 => 
                           n1164, B2 => REGISTERS_28_15_port, ZN => n1468);
   U1967 : NOR4_X1 port map( A1 => n1469, A2 => n1470, A3 => n1471, A4 => n1472
                           , ZN => n1459);
   U1968 : OAI221_X1 port map( B1 => n1088, B2 => n1169, C1 => n1122, C2 => 
                           n1170, A => n1473, ZN => n1472);
   U1969 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_15_port, B1 => 
                           n1173, B2 => REGISTERS_2_15_port, ZN => n1473);
   U1970 : OAI221_X1 port map( B1 => n952, B2 => n1174, C1 => n986, C2 => n1175
                           , A => n1474, ZN => n1471);
   U1971 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_15_port, B1 => 
                           n1178, B2 => REGISTERS_6_15_port, ZN => n1474);
   U1972 : OAI221_X1 port map( B1 => n811, B2 => n1179, C1 => n845, C2 => n1180
                           , A => n1475, ZN => n1470);
   U1973 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_15_port, B1 => 
                           n1183, B2 => REGISTERS_10_15_port, ZN => n1475);
   U1974 : OAI221_X1 port map( B1 => n675, B2 => n1184, C1 => n709, C2 => n1185
                           , A => n1476, ZN => n1469);
   U1975 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_15_port, B1 => 
                           n1188, B2 => REGISTERS_14_15_port, ZN => n1476);
   U1976 : AOI21_X1 port map( B1 => n1477, B2 => n1478, A => N352, ZN => N334);
   U1977 : NOR4_X1 port map( A1 => n1479, A2 => n1480, A3 => n1481, A4 => n1482
                           , ZN => n1478);
   U1978 : OAI221_X1 port map( B1 => n536, B2 => n1145, C1 => n570, C2 => n1146
                           , A => n1483, ZN => n1482);
   U1979 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_14_port, B1 => 
                           n1149, B2 => REGISTERS_18_14_port, ZN => n1483);
   U1980 : OAI221_X1 port map( B1 => n400, B2 => n1150, C1 => n434, C2 => n1151
                           , A => n1484, ZN => n1481);
   U1981 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_14_port, B1 => 
                           n1154, B2 => REGISTERS_22_14_port, ZN => n1484);
   U1982 : OAI221_X1 port map( B1 => n260, B2 => n1155, C1 => n295_port, C2 => 
                           n1156, A => n1485, ZN => n1480);
   U1983 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_14_port, B1 => 
                           n1159, B2 => REGISTERS_26_14_port, ZN => n1485);
   U1984 : OAI221_X1 port map( B1 => n32, B2 => n1160, C1 => n85, C2 => n1161, 
                           A => n1486, ZN => n1479);
   U1985 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_14_port, B1 => 
                           n1164, B2 => REGISTERS_28_14_port, ZN => n1486);
   U1986 : NOR4_X1 port map( A1 => n1487, A2 => n1488, A3 => n1489, A4 => n1490
                           , ZN => n1477);
   U1987 : OAI221_X1 port map( B1 => n1087, B2 => n1169, C1 => n1121, C2 => 
                           n1170, A => n1491, ZN => n1490);
   U1988 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_14_port, B1 => 
                           n1173, B2 => REGISTERS_2_14_port, ZN => n1491);
   U1989 : OAI221_X1 port map( B1 => n951, B2 => n1174, C1 => n985, C2 => n1175
                           , A => n1492, ZN => n1489);
   U1990 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_14_port, B1 => 
                           n1178, B2 => REGISTERS_6_14_port, ZN => n1492);
   U1991 : OAI221_X1 port map( B1 => n810, B2 => n1179, C1 => n844, C2 => n1180
                           , A => n1493, ZN => n1488);
   U1992 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_14_port, B1 => 
                           n1183, B2 => REGISTERS_10_14_port, ZN => n1493);
   U1993 : OAI221_X1 port map( B1 => n674, B2 => n1184, C1 => n708, C2 => n1185
                           , A => n1494, ZN => n1487);
   U1994 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_14_port, B1 => 
                           n1188, B2 => REGISTERS_14_14_port, ZN => n1494);
   U1995 : AOI21_X1 port map( B1 => n1495, B2 => n1496, A => N352, ZN => N333);
   U1996 : NOR4_X1 port map( A1 => n1497, A2 => n1498, A3 => n1499, A4 => n1500
                           , ZN => n1496);
   U1997 : OAI221_X1 port map( B1 => n535, B2 => n1145, C1 => n569, C2 => n1146
                           , A => n1501, ZN => n1500);
   U1998 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_13_port, B1 => 
                           n1149, B2 => REGISTERS_18_13_port, ZN => n1501);
   U1999 : OAI221_X1 port map( B1 => n399, B2 => n1150, C1 => n433, C2 => n1151
                           , A => n1502, ZN => n1499);
   U2000 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_13_port, B1 => 
                           n1154, B2 => REGISTERS_22_13_port, ZN => n1502);
   U2001 : OAI221_X1 port map( B1 => n259, B2 => n1155, C1 => n294_port, C2 => 
                           n1156, A => n1503, ZN => n1498);
   U2002 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_13_port, B1 => 
                           n1159, B2 => REGISTERS_26_13_port, ZN => n1503);
   U2003 : OAI221_X1 port map( B1 => n30, B2 => n1160, C1 => n84, C2 => n1161, 
                           A => n1504, ZN => n1497);
   U2004 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_13_port, B1 => 
                           n1164, B2 => REGISTERS_28_13_port, ZN => n1504);
   U2005 : NOR4_X1 port map( A1 => n1505, A2 => n1506, A3 => n1507, A4 => n1508
                           , ZN => n1495);
   U2006 : OAI221_X1 port map( B1 => n1086, B2 => n1169, C1 => n1120, C2 => 
                           n1170, A => n1509, ZN => n1508);
   U2007 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_13_port, B1 => 
                           n1173, B2 => REGISTERS_2_13_port, ZN => n1509);
   U2008 : OAI221_X1 port map( B1 => n950, B2 => n1174, C1 => n984, C2 => n1175
                           , A => n1510, ZN => n1507);
   U2009 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_13_port, B1 => 
                           n1178, B2 => REGISTERS_6_13_port, ZN => n1510);
   U2010 : OAI221_X1 port map( B1 => n809, B2 => n1179, C1 => n843, C2 => n1180
                           , A => n1511, ZN => n1506);
   U2011 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_13_port, B1 => 
                           n1183, B2 => REGISTERS_10_13_port, ZN => n1511);
   U2012 : OAI221_X1 port map( B1 => n673, B2 => n1184, C1 => n707, C2 => n1185
                           , A => n1512, ZN => n1505);
   U2013 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_13_port, B1 => 
                           n1188, B2 => REGISTERS_14_13_port, ZN => n1512);
   U2014 : AOI21_X1 port map( B1 => n1513, B2 => n1514, A => N352, ZN => N332);
   U2015 : NOR4_X1 port map( A1 => n1515, A2 => n1516, A3 => n1517, A4 => n1518
                           , ZN => n1514);
   U2016 : OAI221_X1 port map( B1 => n534, B2 => n1145, C1 => n568, C2 => n1146
                           , A => n1519, ZN => n1518);
   U2017 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_12_port, B1 => 
                           n1149, B2 => REGISTERS_18_12_port, ZN => n1519);
   U2018 : OAI221_X1 port map( B1 => n398, B2 => n1150, C1 => n432, C2 => n1151
                           , A => n1520, ZN => n1517);
   U2019 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_12_port, B1 => 
                           n1154, B2 => REGISTERS_22_12_port, ZN => n1520);
   U2020 : OAI221_X1 port map( B1 => n258, B2 => n1155, C1 => n293_port, C2 => 
                           n1156, A => n1521, ZN => n1516);
   U2021 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_12_port, B1 => 
                           n1159, B2 => REGISTERS_26_12_port, ZN => n1521);
   U2022 : OAI221_X1 port map( B1 => n28, B2 => n1160, C1 => n83, C2 => n1161, 
                           A => n1522, ZN => n1515);
   U2023 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_12_port, B1 => 
                           n1164, B2 => REGISTERS_28_12_port, ZN => n1522);
   U2024 : NOR4_X1 port map( A1 => n1523, A2 => n1524, A3 => n1525, A4 => n1526
                           , ZN => n1513);
   U2025 : OAI221_X1 port map( B1 => n1085, B2 => n1169, C1 => n1119, C2 => 
                           n1170, A => n1527, ZN => n1526);
   U2026 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_12_port, B1 => 
                           n1173, B2 => REGISTERS_2_12_port, ZN => n1527);
   U2027 : OAI221_X1 port map( B1 => n949, B2 => n1174, C1 => n983, C2 => n1175
                           , A => n1528, ZN => n1525);
   U2028 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_12_port, B1 => 
                           n1178, B2 => REGISTERS_6_12_port, ZN => n1528);
   U2029 : OAI221_X1 port map( B1 => n808, B2 => n1179, C1 => n842, C2 => n1180
                           , A => n1529, ZN => n1524);
   U2030 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_12_port, B1 => 
                           n1183, B2 => REGISTERS_10_12_port, ZN => n1529);
   U2031 : OAI221_X1 port map( B1 => n672, B2 => n1184, C1 => n706, C2 => n1185
                           , A => n1530, ZN => n1523);
   U2032 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_12_port, B1 => 
                           n1188, B2 => REGISTERS_14_12_port, ZN => n1530);
   U2033 : AOI21_X1 port map( B1 => n1531, B2 => n1532, A => N352, ZN => N331);
   U2034 : NOR4_X1 port map( A1 => n1533, A2 => n1534, A3 => n1535, A4 => n1536
                           , ZN => n1532);
   U2035 : OAI221_X1 port map( B1 => n533, B2 => n1145, C1 => n567, C2 => n1146
                           , A => n1537, ZN => n1536);
   U2036 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_11_port, B1 => 
                           n1149, B2 => REGISTERS_18_11_port, ZN => n1537);
   U2037 : OAI221_X1 port map( B1 => n397, B2 => n1150, C1 => n431, C2 => n1151
                           , A => n1538, ZN => n1535);
   U2038 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_11_port, B1 => 
                           n1154, B2 => REGISTERS_22_11_port, ZN => n1538);
   U2039 : OAI221_X1 port map( B1 => n257, B2 => n1155, C1 => n292_port, C2 => 
                           n1156, A => n1539, ZN => n1534);
   U2040 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_11_port, B1 => 
                           n1159, B2 => REGISTERS_26_11_port, ZN => n1539);
   U2041 : OAI221_X1 port map( B1 => n26, B2 => n1160, C1 => n82, C2 => n1161, 
                           A => n1540, ZN => n1533);
   U2042 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_11_port, B1 => 
                           n1164, B2 => REGISTERS_28_11_port, ZN => n1540);
   U2043 : NOR4_X1 port map( A1 => n1541, A2 => n1542, A3 => n1543, A4 => n1544
                           , ZN => n1531);
   U2044 : OAI221_X1 port map( B1 => n1084, B2 => n1169, C1 => n1118, C2 => 
                           n1170, A => n1545, ZN => n1544);
   U2045 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_11_port, B1 => 
                           n1173, B2 => REGISTERS_2_11_port, ZN => n1545);
   U2046 : OAI221_X1 port map( B1 => n948, B2 => n1174, C1 => n982, C2 => n1175
                           , A => n1546, ZN => n1543);
   U2047 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_11_port, B1 => 
                           n1178, B2 => REGISTERS_6_11_port, ZN => n1546);
   U2048 : OAI221_X1 port map( B1 => n807, B2 => n1179, C1 => n841, C2 => n1180
                           , A => n1547, ZN => n1542);
   U2049 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_11_port, B1 => 
                           n1183, B2 => REGISTERS_10_11_port, ZN => n1547);
   U2050 : OAI221_X1 port map( B1 => n671, B2 => n1184, C1 => n705, C2 => n1185
                           , A => n1548, ZN => n1541);
   U2051 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_11_port, B1 => 
                           n1188, B2 => REGISTERS_14_11_port, ZN => n1548);
   U2052 : AOI21_X1 port map( B1 => n1549, B2 => n1550, A => N352, ZN => N330);
   U2053 : NOR4_X1 port map( A1 => n1551, A2 => n1552, A3 => n1553, A4 => n1554
                           , ZN => n1550);
   U2054 : OAI221_X1 port map( B1 => n532, B2 => n1145, C1 => n566, C2 => n1146
                           , A => n1555, ZN => n1554);
   U2055 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_10_port, B1 => 
                           n1149, B2 => REGISTERS_18_10_port, ZN => n1555);
   U2056 : OAI221_X1 port map( B1 => n396, B2 => n1150, C1 => n430, C2 => n1151
                           , A => n1556, ZN => n1553);
   U2057 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_10_port, B1 => 
                           n1154, B2 => REGISTERS_22_10_port, ZN => n1556);
   U2058 : OAI221_X1 port map( B1 => n256, B2 => n1155, C1 => n291_port, C2 => 
                           n1156, A => n1557, ZN => n1552);
   U2059 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_10_port, B1 => 
                           n1159, B2 => REGISTERS_26_10_port, ZN => n1557);
   U2060 : OAI221_X1 port map( B1 => n24, B2 => n1160, C1 => n81, C2 => n1161, 
                           A => n1558, ZN => n1551);
   U2061 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_10_port, B1 => 
                           n1164, B2 => REGISTERS_28_10_port, ZN => n1558);
   U2062 : NOR4_X1 port map( A1 => n1559, A2 => n1560, A3 => n1561, A4 => n1562
                           , ZN => n1549);
   U2063 : OAI221_X1 port map( B1 => n1083, B2 => n1169, C1 => n1117, C2 => 
                           n1170, A => n1563, ZN => n1562);
   U2064 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_10_port, B1 => 
                           n1173, B2 => REGISTERS_2_10_port, ZN => n1563);
   U2065 : OAI221_X1 port map( B1 => n947, B2 => n1174, C1 => n981, C2 => n1175
                           , A => n1564, ZN => n1561);
   U2066 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_10_port, B1 => 
                           n1178, B2 => REGISTERS_6_10_port, ZN => n1564);
   U2067 : OAI221_X1 port map( B1 => n806, B2 => n1179, C1 => n840, C2 => n1180
                           , A => n1565, ZN => n1560);
   U2068 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_10_port, B1 => 
                           n1183, B2 => REGISTERS_10_10_port, ZN => n1565);
   U2069 : OAI221_X1 port map( B1 => n670, B2 => n1184, C1 => n704, C2 => n1185
                           , A => n1566, ZN => n1559);
   U2070 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_10_port, B1 => 
                           n1188, B2 => REGISTERS_14_10_port, ZN => n1566);
   U2071 : AOI21_X1 port map( B1 => n1567, B2 => n1568, A => N352, ZN => N329);
   U2072 : NOR4_X1 port map( A1 => n1569, A2 => n1570, A3 => n1571, A4 => n1572
                           , ZN => n1568);
   U2073 : OAI221_X1 port map( B1 => n531, B2 => n1145, C1 => n565, C2 => n1146
                           , A => n1573, ZN => n1572);
   U2074 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_9_port, B1 => 
                           n1149, B2 => REGISTERS_18_9_port, ZN => n1573);
   U2075 : OAI221_X1 port map( B1 => n395, B2 => n1150, C1 => n429, C2 => n1151
                           , A => n1574, ZN => n1571);
   U2076 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_9_port, B1 => 
                           n1154, B2 => REGISTERS_22_9_port, ZN => n1574);
   U2077 : OAI221_X1 port map( B1 => n255, B2 => n1155, C1 => n290_port, C2 => 
                           n1156, A => n1575, ZN => n1570);
   U2078 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_9_port, B1 => 
                           n1159, B2 => REGISTERS_26_9_port, ZN => n1575);
   U2079 : OAI221_X1 port map( B1 => n22, B2 => n1160, C1 => n80, C2 => n1161, 
                           A => n1576, ZN => n1569);
   U2080 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_9_port, B1 => 
                           n1164, B2 => REGISTERS_28_9_port, ZN => n1576);
   U2081 : NOR4_X1 port map( A1 => n1577, A2 => n1578, A3 => n1579, A4 => n1580
                           , ZN => n1567);
   U2082 : OAI221_X1 port map( B1 => n1082, B2 => n1169, C1 => n1116, C2 => 
                           n1170, A => n1581, ZN => n1580);
   U2083 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_9_port, B1 => 
                           n1173, B2 => REGISTERS_2_9_port, ZN => n1581);
   U2084 : OAI221_X1 port map( B1 => n946, B2 => n1174, C1 => n980, C2 => n1175
                           , A => n1582, ZN => n1579);
   U2085 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_9_port, B1 => 
                           n1178, B2 => REGISTERS_6_9_port, ZN => n1582);
   U2086 : OAI221_X1 port map( B1 => n805, B2 => n1179, C1 => n839, C2 => n1180
                           , A => n1583, ZN => n1578);
   U2087 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_9_port, B1 => 
                           n1183, B2 => REGISTERS_10_9_port, ZN => n1583);
   U2088 : OAI221_X1 port map( B1 => n669, B2 => n1184, C1 => n703, C2 => n1185
                           , A => n1584, ZN => n1577);
   U2089 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_9_port, B1 => 
                           n1188, B2 => REGISTERS_14_9_port, ZN => n1584);
   U2090 : AOI21_X1 port map( B1 => n1585, B2 => n1586, A => N352, ZN => N328);
   U2091 : NOR4_X1 port map( A1 => n1587, A2 => n1588, A3 => n1589, A4 => n1590
                           , ZN => n1586);
   U2092 : OAI221_X1 port map( B1 => n530, B2 => n1145, C1 => n564, C2 => n1146
                           , A => n1591, ZN => n1590);
   U2093 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_8_port, B1 => 
                           n1149, B2 => REGISTERS_18_8_port, ZN => n1591);
   U2094 : OAI221_X1 port map( B1 => n394, B2 => n1150, C1 => n428, C2 => n1151
                           , A => n1592, ZN => n1589);
   U2095 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_8_port, B1 => 
                           n1154, B2 => REGISTERS_22_8_port, ZN => n1592);
   U2096 : OAI221_X1 port map( B1 => n254, B2 => n1155, C1 => n289_port, C2 => 
                           n1156, A => n1593, ZN => n1588);
   U2097 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_8_port, B1 => 
                           n1159, B2 => REGISTERS_26_8_port, ZN => n1593);
   U2098 : OAI221_X1 port map( B1 => n20, B2 => n1160, C1 => n79, C2 => n1161, 
                           A => n1594, ZN => n1587);
   U2099 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_8_port, B1 => 
                           n1164, B2 => REGISTERS_28_8_port, ZN => n1594);
   U2100 : NOR4_X1 port map( A1 => n1595, A2 => n1596, A3 => n1597, A4 => n1598
                           , ZN => n1585);
   U2101 : OAI221_X1 port map( B1 => n1081, B2 => n1169, C1 => n1115, C2 => 
                           n1170, A => n1599, ZN => n1598);
   U2102 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_8_port, B1 => 
                           n1173, B2 => REGISTERS_2_8_port, ZN => n1599);
   U2103 : OAI221_X1 port map( B1 => n945, B2 => n1174, C1 => n979, C2 => n1175
                           , A => n1600, ZN => n1597);
   U2104 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_8_port, B1 => 
                           n1178, B2 => REGISTERS_6_8_port, ZN => n1600);
   U2105 : OAI221_X1 port map( B1 => n804, B2 => n1179, C1 => n838, C2 => n1180
                           , A => n1601, ZN => n1596);
   U2106 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_8_port, B1 => 
                           n1183, B2 => REGISTERS_10_8_port, ZN => n1601);
   U2107 : OAI221_X1 port map( B1 => n668, B2 => n1184, C1 => n702, C2 => n1185
                           , A => n1602, ZN => n1595);
   U2108 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_8_port, B1 => 
                           n1188, B2 => REGISTERS_14_8_port, ZN => n1602);
   U2109 : AOI21_X1 port map( B1 => n1603, B2 => n1604, A => N352, ZN => N327);
   U2110 : NOR4_X1 port map( A1 => n1605, A2 => n1606, A3 => n1607, A4 => n1608
                           , ZN => n1604);
   U2111 : OAI221_X1 port map( B1 => n529, B2 => n1145, C1 => n563, C2 => n1146
                           , A => n1609, ZN => n1608);
   U2112 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_7_port, B1 => 
                           n1149, B2 => REGISTERS_18_7_port, ZN => n1609);
   U2113 : OAI221_X1 port map( B1 => n393, B2 => n1150, C1 => n427, C2 => n1151
                           , A => n1610, ZN => n1607);
   U2114 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_7_port, B1 => 
                           n1154, B2 => REGISTERS_22_7_port, ZN => n1610);
   U2115 : OAI221_X1 port map( B1 => n253, B2 => n1155, C1 => n288_port, C2 => 
                           n1156, A => n1611, ZN => n1606);
   U2116 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_7_port, B1 => 
                           n1159, B2 => REGISTERS_26_7_port, ZN => n1611);
   U2117 : OAI221_X1 port map( B1 => n18, B2 => n1160, C1 => n78, C2 => n1161, 
                           A => n1612, ZN => n1605);
   U2118 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_7_port, B1 => 
                           n1164, B2 => REGISTERS_28_7_port, ZN => n1612);
   U2119 : NOR4_X1 port map( A1 => n1613, A2 => n1614, A3 => n1615, A4 => n1616
                           , ZN => n1603);
   U2120 : OAI221_X1 port map( B1 => n1080, B2 => n1169, C1 => n1114, C2 => 
                           n1170, A => n1617, ZN => n1616);
   U2121 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_7_port, B1 => 
                           n1173, B2 => REGISTERS_2_7_port, ZN => n1617);
   U2122 : OAI221_X1 port map( B1 => n944, B2 => n1174, C1 => n978, C2 => n1175
                           , A => n1618, ZN => n1615);
   U2123 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_7_port, B1 => 
                           n1178, B2 => REGISTERS_6_7_port, ZN => n1618);
   U2124 : OAI221_X1 port map( B1 => n803, B2 => n1179, C1 => n837, C2 => n1180
                           , A => n1619, ZN => n1614);
   U2125 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_7_port, B1 => 
                           n1183, B2 => REGISTERS_10_7_port, ZN => n1619);
   U2126 : OAI221_X1 port map( B1 => n667, B2 => n1184, C1 => n701, C2 => n1185
                           , A => n1620, ZN => n1613);
   U2127 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_7_port, B1 => 
                           n1188, B2 => REGISTERS_14_7_port, ZN => n1620);
   U2128 : AOI21_X1 port map( B1 => n1621, B2 => n1622, A => N352, ZN => N326);
   U2129 : NOR4_X1 port map( A1 => n1623, A2 => n1624, A3 => n1625, A4 => n1626
                           , ZN => n1622);
   U2130 : OAI221_X1 port map( B1 => n528, B2 => n1145, C1 => n562, C2 => n1146
                           , A => n1627, ZN => n1626);
   U2131 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_6_port, B1 => 
                           n1149, B2 => REGISTERS_18_6_port, ZN => n1627);
   U2132 : OAI221_X1 port map( B1 => n392, B2 => n1150, C1 => n426, C2 => n1151
                           , A => n1628, ZN => n1625);
   U2133 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_6_port, B1 => 
                           n1154, B2 => REGISTERS_22_6_port, ZN => n1628);
   U2134 : OAI221_X1 port map( B1 => n252, B2 => n1155, C1 => n287_port, C2 => 
                           n1156, A => n1629, ZN => n1624);
   U2135 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_6_port, B1 => 
                           n1159, B2 => REGISTERS_26_6_port, ZN => n1629);
   U2136 : OAI221_X1 port map( B1 => n16, B2 => n1160, C1 => n77, C2 => n1161, 
                           A => n1630, ZN => n1623);
   U2137 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_6_port, B1 => 
                           n1164, B2 => REGISTERS_28_6_port, ZN => n1630);
   U2138 : NOR4_X1 port map( A1 => n1631, A2 => n1632, A3 => n1633, A4 => n1634
                           , ZN => n1621);
   U2139 : OAI221_X1 port map( B1 => n1079, B2 => n1169, C1 => n1113, C2 => 
                           n1170, A => n1635, ZN => n1634);
   U2140 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_6_port, B1 => 
                           n1173, B2 => REGISTERS_2_6_port, ZN => n1635);
   U2141 : OAI221_X1 port map( B1 => n943, B2 => n1174, C1 => n977, C2 => n1175
                           , A => n1636, ZN => n1633);
   U2142 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_6_port, B1 => 
                           n1178, B2 => REGISTERS_6_6_port, ZN => n1636);
   U2143 : OAI221_X1 port map( B1 => n802, B2 => n1179, C1 => n836, C2 => n1180
                           , A => n1637, ZN => n1632);
   U2144 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_6_port, B1 => 
                           n1183, B2 => REGISTERS_10_6_port, ZN => n1637);
   U2145 : OAI221_X1 port map( B1 => n666, B2 => n1184, C1 => n700, C2 => n1185
                           , A => n1638, ZN => n1631);
   U2146 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_6_port, B1 => 
                           n1188, B2 => REGISTERS_14_6_port, ZN => n1638);
   U2147 : AOI21_X1 port map( B1 => n1639, B2 => n1640, A => N352, ZN => N325);
   U2148 : NOR4_X1 port map( A1 => n1641, A2 => n1642, A3 => n1643, A4 => n1644
                           , ZN => n1640);
   U2149 : OAI221_X1 port map( B1 => n527, B2 => n1145, C1 => n561, C2 => n1146
                           , A => n1645, ZN => n1644);
   U2150 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_5_port, B1 => 
                           n1149, B2 => REGISTERS_18_5_port, ZN => n1645);
   U2151 : OAI221_X1 port map( B1 => n391, B2 => n1150, C1 => n425, C2 => n1151
                           , A => n1646, ZN => n1643);
   U2152 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_5_port, B1 => 
                           n1154, B2 => REGISTERS_22_5_port, ZN => n1646);
   U2153 : OAI221_X1 port map( B1 => n251, B2 => n1155, C1 => n286_port, C2 => 
                           n1156, A => n1647, ZN => n1642);
   U2154 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_5_port, B1 => 
                           n1159, B2 => REGISTERS_26_5_port, ZN => n1647);
   U2155 : OAI221_X1 port map( B1 => n14, B2 => n1160, C1 => n76, C2 => n1161, 
                           A => n1648, ZN => n1641);
   U2156 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_5_port, B1 => 
                           n1164, B2 => REGISTERS_28_5_port, ZN => n1648);
   U2157 : NOR4_X1 port map( A1 => n1649, A2 => n1650, A3 => n1651, A4 => n1652
                           , ZN => n1639);
   U2158 : OAI221_X1 port map( B1 => n1078, B2 => n1169, C1 => n1112, C2 => 
                           n1170, A => n1653, ZN => n1652);
   U2159 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_5_port, B1 => 
                           n1173, B2 => REGISTERS_2_5_port, ZN => n1653);
   U2160 : OAI221_X1 port map( B1 => n942, B2 => n1174, C1 => n976, C2 => n1175
                           , A => n1654, ZN => n1651);
   U2161 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_5_port, B1 => 
                           n1178, B2 => REGISTERS_6_5_port, ZN => n1654);
   U2162 : OAI221_X1 port map( B1 => n801, B2 => n1179, C1 => n835, C2 => n1180
                           , A => n1655, ZN => n1650);
   U2163 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_5_port, B1 => 
                           n1183, B2 => REGISTERS_10_5_port, ZN => n1655);
   U2164 : OAI221_X1 port map( B1 => n665, B2 => n1184, C1 => n699, C2 => n1185
                           , A => n1656, ZN => n1649);
   U2165 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_5_port, B1 => 
                           n1188, B2 => REGISTERS_14_5_port, ZN => n1656);
   U2166 : AOI21_X1 port map( B1 => n1657, B2 => n1658, A => N352, ZN => N324);
   U2167 : NOR4_X1 port map( A1 => n1659, A2 => n1660, A3 => n1661, A4 => n1662
                           , ZN => n1658);
   U2168 : OAI221_X1 port map( B1 => n526, B2 => n1145, C1 => n560, C2 => n1146
                           , A => n1663, ZN => n1662);
   U2169 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_4_port, B1 => 
                           n1149, B2 => REGISTERS_18_4_port, ZN => n1663);
   U2170 : OAI221_X1 port map( B1 => n390, B2 => n1150, C1 => n424, C2 => n1151
                           , A => n1664, ZN => n1661);
   U2171 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_4_port, B1 => 
                           n1154, B2 => REGISTERS_22_4_port, ZN => n1664);
   U2172 : OAI221_X1 port map( B1 => n250, B2 => n1155, C1 => n285, C2 => n1156
                           , A => n1665, ZN => n1660);
   U2173 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_4_port, B1 => 
                           n1159, B2 => REGISTERS_26_4_port, ZN => n1665);
   U2174 : OAI221_X1 port map( B1 => n12, B2 => n1160, C1 => n75, C2 => n1161, 
                           A => n1666, ZN => n1659);
   U2175 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_4_port, B1 => 
                           n1164, B2 => REGISTERS_28_4_port, ZN => n1666);
   U2176 : NOR4_X1 port map( A1 => n1667, A2 => n1668, A3 => n1669, A4 => n1670
                           , ZN => n1657);
   U2177 : OAI221_X1 port map( B1 => n1077, B2 => n1169, C1 => n1111, C2 => 
                           n1170, A => n1671, ZN => n1670);
   U2178 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_4_port, B1 => 
                           n1173, B2 => REGISTERS_2_4_port, ZN => n1671);
   U2179 : OAI221_X1 port map( B1 => n941, B2 => n1174, C1 => n975, C2 => n1175
                           , A => n1672, ZN => n1669);
   U2180 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_4_port, B1 => 
                           n1178, B2 => REGISTERS_6_4_port, ZN => n1672);
   U2181 : OAI221_X1 port map( B1 => n800, B2 => n1179, C1 => n834, C2 => n1180
                           , A => n1673, ZN => n1668);
   U2182 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_4_port, B1 => 
                           n1183, B2 => REGISTERS_10_4_port, ZN => n1673);
   U2183 : OAI221_X1 port map( B1 => n664, B2 => n1184, C1 => n698, C2 => n1185
                           , A => n1674, ZN => n1667);
   U2184 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_4_port, B1 => 
                           n1188, B2 => REGISTERS_14_4_port, ZN => n1674);
   U2185 : AOI21_X1 port map( B1 => n1675, B2 => n1676, A => N352, ZN => N323);
   U2186 : NOR4_X1 port map( A1 => n1677, A2 => n1678, A3 => n1679, A4 => n1680
                           , ZN => n1676);
   U2187 : OAI221_X1 port map( B1 => n525, B2 => n1145, C1 => n559, C2 => n1146
                           , A => n1681, ZN => n1680);
   U2188 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_3_port, B1 => 
                           n1149, B2 => REGISTERS_18_3_port, ZN => n1681);
   U2189 : OAI221_X1 port map( B1 => n389, B2 => n1150, C1 => n423, C2 => n1151
                           , A => n1682, ZN => n1679);
   U2190 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_3_port, B1 => 
                           n1154, B2 => REGISTERS_22_3_port, ZN => n1682);
   U2191 : OAI221_X1 port map( B1 => n249, B2 => n1155, C1 => n284, C2 => n1156
                           , A => n1683, ZN => n1678);
   U2192 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_3_port, B1 => 
                           n1159, B2 => REGISTERS_26_3_port, ZN => n1683);
   U2193 : OAI221_X1 port map( B1 => n10, B2 => n1160, C1 => n74, C2 => n1161, 
                           A => n1684, ZN => n1677);
   U2194 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_3_port, B1 => 
                           n1164, B2 => REGISTERS_28_3_port, ZN => n1684);
   U2195 : NOR4_X1 port map( A1 => n1685, A2 => n1686, A3 => n1687, A4 => n1688
                           , ZN => n1675);
   U2196 : OAI221_X1 port map( B1 => n1076, B2 => n1169, C1 => n1110, C2 => 
                           n1170, A => n1689, ZN => n1688);
   U2197 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_3_port, B1 => 
                           n1173, B2 => REGISTERS_2_3_port, ZN => n1689);
   U2198 : OAI221_X1 port map( B1 => n940, B2 => n1174, C1 => n974, C2 => n1175
                           , A => n1690, ZN => n1687);
   U2199 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_3_port, B1 => 
                           n1178, B2 => REGISTERS_6_3_port, ZN => n1690);
   U2200 : OAI221_X1 port map( B1 => n799, B2 => n1179, C1 => n833, C2 => n1180
                           , A => n1691, ZN => n1686);
   U2201 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_3_port, B1 => 
                           n1183, B2 => REGISTERS_10_3_port, ZN => n1691);
   U2202 : OAI221_X1 port map( B1 => n663, B2 => n1184, C1 => n697, C2 => n1185
                           , A => n1692, ZN => n1685);
   U2203 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_3_port, B1 => 
                           n1188, B2 => REGISTERS_14_3_port, ZN => n1692);
   U2204 : AOI21_X1 port map( B1 => n1693, B2 => n1694, A => N352, ZN => N322);
   U2205 : NOR4_X1 port map( A1 => n1695, A2 => n1696, A3 => n1697, A4 => n1698
                           , ZN => n1694);
   U2206 : OAI221_X1 port map( B1 => n524, B2 => n1145, C1 => n558, C2 => n1146
                           , A => n1699, ZN => n1698);
   U2207 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_2_port, B1 => 
                           n1149, B2 => REGISTERS_18_2_port, ZN => n1699);
   U2208 : OAI221_X1 port map( B1 => n388, B2 => n1150, C1 => n422, C2 => n1151
                           , A => n1700, ZN => n1697);
   U2209 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_2_port, B1 => 
                           n1154, B2 => REGISTERS_22_2_port, ZN => n1700);
   U2210 : OAI221_X1 port map( B1 => n248, B2 => n1155, C1 => n283, C2 => n1156
                           , A => n1701, ZN => n1696);
   U2211 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_2_port, B1 => 
                           n1159, B2 => REGISTERS_26_2_port, ZN => n1701);
   U2212 : OAI221_X1 port map( B1 => n8, B2 => n1160, C1 => n73, C2 => n1161, A
                           => n1702, ZN => n1695);
   U2213 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_2_port, B1 => 
                           n1164, B2 => REGISTERS_28_2_port, ZN => n1702);
   U2214 : NOR4_X1 port map( A1 => n1703, A2 => n1704, A3 => n1705, A4 => n1706
                           , ZN => n1693);
   U2215 : OAI221_X1 port map( B1 => n1075, B2 => n1169, C1 => n1109, C2 => 
                           n1170, A => n1707, ZN => n1706);
   U2216 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_2_port, B1 => 
                           n1173, B2 => REGISTERS_2_2_port, ZN => n1707);
   U2217 : OAI221_X1 port map( B1 => n939, B2 => n1174, C1 => n973, C2 => n1175
                           , A => n1708, ZN => n1705);
   U2218 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_2_port, B1 => 
                           n1178, B2 => REGISTERS_6_2_port, ZN => n1708);
   U2219 : OAI221_X1 port map( B1 => n798, B2 => n1179, C1 => n832, C2 => n1180
                           , A => n1709, ZN => n1704);
   U2220 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_2_port, B1 => 
                           n1183, B2 => REGISTERS_10_2_port, ZN => n1709);
   U2221 : OAI221_X1 port map( B1 => n662, B2 => n1184, C1 => n696, C2 => n1185
                           , A => n1710, ZN => n1703);
   U2222 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_2_port, B1 => 
                           n1188, B2 => REGISTERS_14_2_port, ZN => n1710);
   U2223 : AOI21_X1 port map( B1 => n1711, B2 => n1712, A => N352, ZN => N321);
   U2224 : NOR4_X1 port map( A1 => n1713, A2 => n1714, A3 => n1715, A4 => n1716
                           , ZN => n1712);
   U2225 : OAI221_X1 port map( B1 => n523, B2 => n1145, C1 => n557, C2 => n1146
                           , A => n1717, ZN => n1716);
   U2226 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_1_port, B1 => 
                           n1149, B2 => REGISTERS_18_1_port, ZN => n1717);
   U2227 : OAI221_X1 port map( B1 => n387, B2 => n1150, C1 => n421, C2 => n1151
                           , A => n1718, ZN => n1715);
   U2228 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_1_port, B1 => 
                           n1154, B2 => REGISTERS_22_1_port, ZN => n1718);
   U2229 : OAI221_X1 port map( B1 => n247, B2 => n1155, C1 => n282, C2 => n1156
                           , A => n1719, ZN => n1714);
   U2230 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_1_port, B1 => 
                           n1159, B2 => REGISTERS_26_1_port, ZN => n1719);
   U2231 : OAI221_X1 port map( B1 => n6, B2 => n1160, C1 => n72, C2 => n1161, A
                           => n1720, ZN => n1713);
   U2232 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_1_port, B1 => 
                           n1164, B2 => REGISTERS_28_1_port, ZN => n1720);
   U2233 : NOR4_X1 port map( A1 => n1721, A2 => n1722, A3 => n1723, A4 => n1724
                           , ZN => n1711);
   U2234 : OAI221_X1 port map( B1 => n1074, B2 => n1169, C1 => n1108, C2 => 
                           n1170, A => n1725, ZN => n1724);
   U2235 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_1_port, B1 => 
                           n1173, B2 => REGISTERS_2_1_port, ZN => n1725);
   U2236 : OAI221_X1 port map( B1 => n938, B2 => n1174, C1 => n972, C2 => n1175
                           , A => n1726, ZN => n1723);
   U2237 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_1_port, B1 => 
                           n1178, B2 => REGISTERS_6_1_port, ZN => n1726);
   U2238 : OAI221_X1 port map( B1 => n797, B2 => n1179, C1 => n831, C2 => n1180
                           , A => n1727, ZN => n1722);
   U2239 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_1_port, B1 => 
                           n1183, B2 => REGISTERS_10_1_port, ZN => n1727);
   U2240 : OAI221_X1 port map( B1 => n661, B2 => n1184, C1 => n695, C2 => n1185
                           , A => n1728, ZN => n1721);
   U2241 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_1_port, B1 => 
                           n1188, B2 => REGISTERS_14_1_port, ZN => n1728);
   U2242 : AOI21_X1 port map( B1 => n1729, B2 => n1730, A => N352, ZN => N320);
   U2243 : NOR4_X1 port map( A1 => n1731, A2 => n1732, A3 => n1733, A4 => n1734
                           , ZN => n1730);
   U2244 : OAI221_X1 port map( B1 => n522, B2 => n1145, C1 => n556, C2 => n1146
                           , A => n1735, ZN => n1734);
   U2245 : AOI22_X1 port map( A1 => n1148, A2 => REGISTERS_19_0_port, B1 => 
                           n1149, B2 => REGISTERS_18_0_port, ZN => n1735);
   U2250 : OAI221_X1 port map( B1 => n386, B2 => n1150, C1 => n420, C2 => n1151
                           , A => n1740, ZN => n1733);
   U2251 : AOI22_X1 port map( A1 => n1153, A2 => REGISTERS_23_0_port, B1 => 
                           n1154, B2 => REGISTERS_22_0_port, ZN => n1740);
   U2255 : AND2_X1 port map( A1 => n1743, A2 => n1744, ZN => n1736);
   U2257 : AND2_X1 port map( A1 => n1743, A2 => ADD_RD2(0), ZN => n1738);
   U2258 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => n1745, ZN => n1743);
   U2259 : OAI221_X1 port map( B1 => n246, B2 => n1155, C1 => n281, C2 => n1156
                           , A => n1746, ZN => n1732);
   U2260 : AOI22_X1 port map( A1 => n1158, A2 => REGISTERS_27_0_port, B1 => 
                           n1159, B2 => REGISTERS_26_0_port, ZN => n1746);
   U2265 : OAI221_X1 port map( B1 => n4, B2 => n1160, C1 => n71, C2 => n1161, A
                           => n1749, ZN => n1731);
   U2266 : AOI22_X1 port map( A1 => n1163, A2 => REGISTERS_29_0_port, B1 => 
                           n1164, B2 => REGISTERS_28_0_port, ZN => n1749);
   U2270 : AND2_X1 port map( A1 => n1750, A2 => n1744, ZN => n1747);
   U2272 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n1750, ZN => n1748);
   U2273 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1750);
   U2274 : NOR4_X1 port map( A1 => n1751, A2 => n1752, A3 => n1753, A4 => n1754
                           , ZN => n1729);
   U2275 : OAI221_X1 port map( B1 => n1073, B2 => n1169, C1 => n1107, C2 => 
                           n1170, A => n1755, ZN => n1754);
   U2276 : AOI22_X1 port map( A1 => n1172, A2 => REGISTERS_3_0_port, B1 => 
                           n1173, B2 => REGISTERS_2_0_port, ZN => n1755);
   U2281 : OAI221_X1 port map( B1 => n937, B2 => n1174, C1 => n971, C2 => n1175
                           , A => n1758, ZN => n1753);
   U2282 : AOI22_X1 port map( A1 => n1177, A2 => REGISTERS_7_0_port, B1 => 
                           n1178, B2 => REGISTERS_6_0_port, ZN => n1758);
   U2286 : AND2_X1 port map( A1 => n1759, A2 => n1744, ZN => n1756);
   U2288 : AND2_X1 port map( A1 => n1759, A2 => ADD_RD2(0), ZN => n1757);
   U2289 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n1759);
   U2290 : OAI221_X1 port map( B1 => n796, B2 => n1179, C1 => n830, C2 => n1180
                           , A => n1760, ZN => n1752);
   U2291 : AOI22_X1 port map( A1 => n1182, A2 => REGISTERS_11_0_port, B1 => 
                           n1183, B2 => REGISTERS_10_0_port, ZN => n1760);
   U2294 : NOR2_X1 port map( A1 => n1763, A2 => ADD_RD2(2), ZN => n1737);
   U2298 : OAI221_X1 port map( B1 => n660, B2 => n1184, C1 => n694, C2 => n1185
                           , A => n1764, ZN => n1751);
   U2299 : AOI22_X1 port map( A1 => n1187, A2 => REGISTERS_15_0_port, B1 => 
                           n1188, B2 => REGISTERS_14_0_port, ZN => n1764);
   U2302 : NOR2_X1 port map( A1 => n1765, A2 => n1763, ZN => n1741);
   U2303 : INV_X1 port map( A => ADD_RD2(1), ZN => n1763);
   U2305 : AND2_X1 port map( A1 => n1766, A2 => n1744, ZN => n1761);
   U2306 : INV_X1 port map( A => ADD_RD2(0), ZN => n1744);
   U2309 : INV_X1 port map( A => ADD_RD2(2), ZN => n1765);
   U2310 : AND2_X1 port map( A1 => n1766, A2 => ADD_RD2(0), ZN => n1762);
   U2311 : NOR2_X1 port map( A1 => n1745, A2 => ADD_RD2(4), ZN => n1766);
   U2312 : INV_X1 port map( A => ADD_RD2(3), ZN => n1745);
   U2313 : NAND2_X1 port map( A1 => n1767, A2 => RESET, ZN => N319);
   U2314 : NAND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n1767);
   U2315 : AOI21_X1 port map( B1 => n1768, B2 => n1769, A => N352, ZN => N318);
   U2316 : NOR4_X1 port map( A1 => n1770, A2 => n1771, A3 => n1772, A4 => n1773
                           , ZN => n1769);
   U2317 : OAI221_X1 port map( B1 => n553, B2 => n1774, C1 => n587, C2 => n1775
                           , A => n1776, ZN => n1773);
   U2318 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_31_port, B1 => 
                           n1778, B2 => REGISTERS_18_31_port, ZN => n1776);
   U2319 : OAI221_X1 port map( B1 => n417, B2 => n1779, C1 => n451, C2 => n1780
                           , A => n1781, ZN => n1772);
   U2320 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_31_port, B1 => 
                           n1783, B2 => REGISTERS_22_31_port, ZN => n1781);
   U2321 : OAI221_X1 port map( B1 => n277, B2 => n1784, C1 => n312_port, C2 => 
                           n1785, A => n1786, ZN => n1771);
   U2322 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_31_port, B1 => 
                           n1788, B2 => REGISTERS_26_31_port, ZN => n1786);
   U2323 : OAI221_X1 port map( B1 => n66, B2 => n1789, C1 => n102, C2 => n1790,
                           A => n1791, ZN => n1770);
   U2324 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_31_port, B1 => 
                           n1793, B2 => REGISTERS_28_31_port, ZN => n1791);
   U2325 : NOR4_X1 port map( A1 => n1794, A2 => n1795, A3 => n1796, A4 => n1797
                           , ZN => n1768);
   U2326 : OAI221_X1 port map( B1 => n1104, B2 => n1798, C1 => n1138, C2 => 
                           n1799, A => n1800, ZN => n1797);
   U2327 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_31_port, B1 => 
                           n1802, B2 => REGISTERS_2_31_port, ZN => n1800);
   U2328 : OAI221_X1 port map( B1 => n968, B2 => n1803, C1 => n1002, C2 => 
                           n1804, A => n1805, ZN => n1796);
   U2329 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_31_port, B1 => 
                           n1807, B2 => REGISTERS_6_31_port, ZN => n1805);
   U2330 : OAI221_X1 port map( B1 => n827, B2 => n1808, C1 => n861, C2 => n1809
                           , A => n1810, ZN => n1795);
   U2331 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_31_port, B1 => 
                           n1812, B2 => REGISTERS_10_31_port, ZN => n1810);
   U2332 : OAI221_X1 port map( B1 => n691, B2 => n1813, C1 => n725, C2 => n1814
                           , A => n1815, ZN => n1794);
   U2333 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_31_port, B1 => 
                           n1817, B2 => REGISTERS_14_31_port, ZN => n1815);
   U2334 : AOI21_X1 port map( B1 => n1818, B2 => n1819, A => N352, ZN => N317);
   U2335 : NOR4_X1 port map( A1 => n1820, A2 => n1821, A3 => n1822, A4 => n1823
                           , ZN => n1819);
   U2336 : OAI221_X1 port map( B1 => n552, B2 => n1774, C1 => n586, C2 => n1775
                           , A => n1824, ZN => n1823);
   U2337 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_30_port, B1 => 
                           n1778, B2 => REGISTERS_18_30_port, ZN => n1824);
   U2338 : OAI221_X1 port map( B1 => n416, B2 => n1779, C1 => n450, C2 => n1780
                           , A => n1825, ZN => n1822);
   U2339 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_30_port, B1 => 
                           n1783, B2 => REGISTERS_22_30_port, ZN => n1825);
   U2340 : OAI221_X1 port map( B1 => n276, B2 => n1784, C1 => n311_port, C2 => 
                           n1785, A => n1826, ZN => n1821);
   U2341 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_30_port, B1 => 
                           n1788, B2 => REGISTERS_26_30_port, ZN => n1826);
   U2342 : OAI221_X1 port map( B1 => n64, B2 => n1789, C1 => n101, C2 => n1790,
                           A => n1827, ZN => n1820);
   U2343 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_30_port, B1 => 
                           n1793, B2 => REGISTERS_28_30_port, ZN => n1827);
   U2344 : NOR4_X1 port map( A1 => n1828, A2 => n1829, A3 => n1830, A4 => n1831
                           , ZN => n1818);
   U2345 : OAI221_X1 port map( B1 => n1103, B2 => n1798, C1 => n1137, C2 => 
                           n1799, A => n1832, ZN => n1831);
   U2346 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_30_port, B1 => 
                           n1802, B2 => REGISTERS_2_30_port, ZN => n1832);
   U2347 : OAI221_X1 port map( B1 => n967, B2 => n1803, C1 => n1001, C2 => 
                           n1804, A => n1833, ZN => n1830);
   U2348 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_30_port, B1 => 
                           n1807, B2 => REGISTERS_6_30_port, ZN => n1833);
   U2349 : OAI221_X1 port map( B1 => n826, B2 => n1808, C1 => n860, C2 => n1809
                           , A => n1834, ZN => n1829);
   U2350 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_30_port, B1 => 
                           n1812, B2 => REGISTERS_10_30_port, ZN => n1834);
   U2351 : OAI221_X1 port map( B1 => n690, B2 => n1813, C1 => n724, C2 => n1814
                           , A => n1835, ZN => n1828);
   U2352 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_30_port, B1 => 
                           n1817, B2 => REGISTERS_14_30_port, ZN => n1835);
   U2353 : AOI21_X1 port map( B1 => n1836, B2 => n1837, A => N352, ZN => N316);
   U2354 : NOR4_X1 port map( A1 => n1838, A2 => n1839, A3 => n1840, A4 => n1841
                           , ZN => n1837);
   U2355 : OAI221_X1 port map( B1 => n551, B2 => n1774, C1 => n585, C2 => n1775
                           , A => n1842, ZN => n1841);
   U2356 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_29_port, B1 => 
                           n1778, B2 => REGISTERS_18_29_port, ZN => n1842);
   U2357 : OAI221_X1 port map( B1 => n415, B2 => n1779, C1 => n449, C2 => n1780
                           , A => n1843, ZN => n1840);
   U2358 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_29_port, B1 => 
                           n1783, B2 => REGISTERS_22_29_port, ZN => n1843);
   U2359 : OAI221_X1 port map( B1 => n275, B2 => n1784, C1 => n310_port, C2 => 
                           n1785, A => n1844, ZN => n1839);
   U2360 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_29_port, B1 => 
                           n1788, B2 => REGISTERS_26_29_port, ZN => n1844);
   U2361 : OAI221_X1 port map( B1 => n62, B2 => n1789, C1 => n100, C2 => n1790,
                           A => n1845, ZN => n1838);
   U2362 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_29_port, B1 => 
                           n1793, B2 => REGISTERS_28_29_port, ZN => n1845);
   U2363 : NOR4_X1 port map( A1 => n1846, A2 => n1847, A3 => n1848, A4 => n1849
                           , ZN => n1836);
   U2364 : OAI221_X1 port map( B1 => n1102, B2 => n1798, C1 => n1136, C2 => 
                           n1799, A => n1850, ZN => n1849);
   U2365 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_29_port, B1 => 
                           n1802, B2 => REGISTERS_2_29_port, ZN => n1850);
   U2366 : OAI221_X1 port map( B1 => n966, B2 => n1803, C1 => n1000, C2 => 
                           n1804, A => n1851, ZN => n1848);
   U2367 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_29_port, B1 => 
                           n1807, B2 => REGISTERS_6_29_port, ZN => n1851);
   U2368 : OAI221_X1 port map( B1 => n825, B2 => n1808, C1 => n859, C2 => n1809
                           , A => n1852, ZN => n1847);
   U2369 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_29_port, B1 => 
                           n1812, B2 => REGISTERS_10_29_port, ZN => n1852);
   U2370 : OAI221_X1 port map( B1 => n689, B2 => n1813, C1 => n723, C2 => n1814
                           , A => n1853, ZN => n1846);
   U2371 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_29_port, B1 => 
                           n1817, B2 => REGISTERS_14_29_port, ZN => n1853);
   U2372 : AOI21_X1 port map( B1 => n1854, B2 => n1855, A => N352, ZN => N315);
   U2373 : NOR4_X1 port map( A1 => n1856, A2 => n1857, A3 => n1858, A4 => n1859
                           , ZN => n1855);
   U2374 : OAI221_X1 port map( B1 => n550, B2 => n1774, C1 => n584, C2 => n1775
                           , A => n1860, ZN => n1859);
   U2375 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_28_port, B1 => 
                           n1778, B2 => REGISTERS_18_28_port, ZN => n1860);
   U2376 : OAI221_X1 port map( B1 => n414, B2 => n1779, C1 => n448, C2 => n1780
                           , A => n1861, ZN => n1858);
   U2377 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_28_port, B1 => 
                           n1783, B2 => REGISTERS_22_28_port, ZN => n1861);
   U2378 : OAI221_X1 port map( B1 => n274, B2 => n1784, C1 => n309_port, C2 => 
                           n1785, A => n1862, ZN => n1857);
   U2379 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_28_port, B1 => 
                           n1788, B2 => REGISTERS_26_28_port, ZN => n1862);
   U2380 : OAI221_X1 port map( B1 => n60, B2 => n1789, C1 => n99, C2 => n1790, 
                           A => n1863, ZN => n1856);
   U2381 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_28_port, B1 => 
                           n1793, B2 => REGISTERS_28_28_port, ZN => n1863);
   U2382 : NOR4_X1 port map( A1 => n1864, A2 => n1865, A3 => n1866, A4 => n1867
                           , ZN => n1854);
   U2383 : OAI221_X1 port map( B1 => n1101, B2 => n1798, C1 => n1135, C2 => 
                           n1799, A => n1868, ZN => n1867);
   U2384 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_28_port, B1 => 
                           n1802, B2 => REGISTERS_2_28_port, ZN => n1868);
   U2385 : OAI221_X1 port map( B1 => n965, B2 => n1803, C1 => n999, C2 => n1804
                           , A => n1869, ZN => n1866);
   U2386 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_28_port, B1 => 
                           n1807, B2 => REGISTERS_6_28_port, ZN => n1869);
   U2387 : OAI221_X1 port map( B1 => n824, B2 => n1808, C1 => n858, C2 => n1809
                           , A => n1870, ZN => n1865);
   U2388 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_28_port, B1 => 
                           n1812, B2 => REGISTERS_10_28_port, ZN => n1870);
   U2389 : OAI221_X1 port map( B1 => n688, B2 => n1813, C1 => n722, C2 => n1814
                           , A => n1871, ZN => n1864);
   U2390 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_28_port, B1 => 
                           n1817, B2 => REGISTERS_14_28_port, ZN => n1871);
   U2391 : AOI21_X1 port map( B1 => n1872, B2 => n1873, A => N352, ZN => N314);
   U2392 : NOR4_X1 port map( A1 => n1874, A2 => n1875, A3 => n1876, A4 => n1877
                           , ZN => n1873);
   U2393 : OAI221_X1 port map( B1 => n549, B2 => n1774, C1 => n583, C2 => n1775
                           , A => n1878, ZN => n1877);
   U2394 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_27_port, B1 => 
                           n1778, B2 => REGISTERS_18_27_port, ZN => n1878);
   U2395 : OAI221_X1 port map( B1 => n413, B2 => n1779, C1 => n447, C2 => n1780
                           , A => n1879, ZN => n1876);
   U2396 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_27_port, B1 => 
                           n1783, B2 => REGISTERS_22_27_port, ZN => n1879);
   U2397 : OAI221_X1 port map( B1 => n273, B2 => n1784, C1 => n308_port, C2 => 
                           n1785, A => n1880, ZN => n1875);
   U2398 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_27_port, B1 => 
                           n1788, B2 => REGISTERS_26_27_port, ZN => n1880);
   U2399 : OAI221_X1 port map( B1 => n58, B2 => n1789, C1 => n98, C2 => n1790, 
                           A => n1881, ZN => n1874);
   U2400 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_27_port, B1 => 
                           n1793, B2 => REGISTERS_28_27_port, ZN => n1881);
   U2401 : NOR4_X1 port map( A1 => n1882, A2 => n1883, A3 => n1884, A4 => n1885
                           , ZN => n1872);
   U2402 : OAI221_X1 port map( B1 => n1100, B2 => n1798, C1 => n1134, C2 => 
                           n1799, A => n1886, ZN => n1885);
   U2403 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_27_port, B1 => 
                           n1802, B2 => REGISTERS_2_27_port, ZN => n1886);
   U2404 : OAI221_X1 port map( B1 => n964, B2 => n1803, C1 => n998, C2 => n1804
                           , A => n1887, ZN => n1884);
   U2405 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_27_port, B1 => 
                           n1807, B2 => REGISTERS_6_27_port, ZN => n1887);
   U2406 : OAI221_X1 port map( B1 => n823, B2 => n1808, C1 => n857, C2 => n1809
                           , A => n1888, ZN => n1883);
   U2407 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_27_port, B1 => 
                           n1812, B2 => REGISTERS_10_27_port, ZN => n1888);
   U2408 : OAI221_X1 port map( B1 => n687, B2 => n1813, C1 => n721, C2 => n1814
                           , A => n1889, ZN => n1882);
   U2409 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_27_port, B1 => 
                           n1817, B2 => REGISTERS_14_27_port, ZN => n1889);
   U2410 : AOI21_X1 port map( B1 => n1890, B2 => n1891, A => N352, ZN => N313);
   U2411 : NOR4_X1 port map( A1 => n1892, A2 => n1893, A3 => n1894, A4 => n1895
                           , ZN => n1891);
   U2412 : OAI221_X1 port map( B1 => n548, B2 => n1774, C1 => n582, C2 => n1775
                           , A => n1896, ZN => n1895);
   U2413 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_26_port, B1 => 
                           n1778, B2 => REGISTERS_18_26_port, ZN => n1896);
   U2414 : OAI221_X1 port map( B1 => n412, B2 => n1779, C1 => n446, C2 => n1780
                           , A => n1897, ZN => n1894);
   U2415 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_26_port, B1 => 
                           n1783, B2 => REGISTERS_22_26_port, ZN => n1897);
   U2416 : OAI221_X1 port map( B1 => n272, B2 => n1784, C1 => n307_port, C2 => 
                           n1785, A => n1898, ZN => n1893);
   U2417 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_26_port, B1 => 
                           n1788, B2 => REGISTERS_26_26_port, ZN => n1898);
   U2418 : OAI221_X1 port map( B1 => n56, B2 => n1789, C1 => n97, C2 => n1790, 
                           A => n1899, ZN => n1892);
   U2419 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_26_port, B1 => 
                           n1793, B2 => REGISTERS_28_26_port, ZN => n1899);
   U2420 : NOR4_X1 port map( A1 => n1900, A2 => n1901, A3 => n1902, A4 => n1903
                           , ZN => n1890);
   U2421 : OAI221_X1 port map( B1 => n1099, B2 => n1798, C1 => n1133, C2 => 
                           n1799, A => n1904, ZN => n1903);
   U2422 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_26_port, B1 => 
                           n1802, B2 => REGISTERS_2_26_port, ZN => n1904);
   U2423 : OAI221_X1 port map( B1 => n963, B2 => n1803, C1 => n997, C2 => n1804
                           , A => n1905, ZN => n1902);
   U2424 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_26_port, B1 => 
                           n1807, B2 => REGISTERS_6_26_port, ZN => n1905);
   U2425 : OAI221_X1 port map( B1 => n822, B2 => n1808, C1 => n856, C2 => n1809
                           , A => n1906, ZN => n1901);
   U2426 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_26_port, B1 => 
                           n1812, B2 => REGISTERS_10_26_port, ZN => n1906);
   U2427 : OAI221_X1 port map( B1 => n686, B2 => n1813, C1 => n720, C2 => n1814
                           , A => n1907, ZN => n1900);
   U2428 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_26_port, B1 => 
                           n1817, B2 => REGISTERS_14_26_port, ZN => n1907);
   U2429 : AOI21_X1 port map( B1 => n1908, B2 => n1909, A => N352, ZN => N312);
   U2430 : NOR4_X1 port map( A1 => n1910, A2 => n1911, A3 => n1912, A4 => n1913
                           , ZN => n1909);
   U2431 : OAI221_X1 port map( B1 => n547, B2 => n1774, C1 => n581, C2 => n1775
                           , A => n1914, ZN => n1913);
   U2432 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_25_port, B1 => 
                           n1778, B2 => REGISTERS_18_25_port, ZN => n1914);
   U2433 : OAI221_X1 port map( B1 => n411, B2 => n1779, C1 => n445, C2 => n1780
                           , A => n1915, ZN => n1912);
   U2434 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_25_port, B1 => 
                           n1783, B2 => REGISTERS_22_25_port, ZN => n1915);
   U2435 : OAI221_X1 port map( B1 => n271, B2 => n1784, C1 => n306_port, C2 => 
                           n1785, A => n1916, ZN => n1911);
   U2436 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_25_port, B1 => 
                           n1788, B2 => REGISTERS_26_25_port, ZN => n1916);
   U2437 : OAI221_X1 port map( B1 => n54, B2 => n1789, C1 => n96, C2 => n1790, 
                           A => n1917, ZN => n1910);
   U2438 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_25_port, B1 => 
                           n1793, B2 => REGISTERS_28_25_port, ZN => n1917);
   U2439 : NOR4_X1 port map( A1 => n1918, A2 => n1919, A3 => n1920, A4 => n1921
                           , ZN => n1908);
   U2440 : OAI221_X1 port map( B1 => n1098, B2 => n1798, C1 => n1132, C2 => 
                           n1799, A => n1922, ZN => n1921);
   U2441 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_25_port, B1 => 
                           n1802, B2 => REGISTERS_2_25_port, ZN => n1922);
   U2442 : OAI221_X1 port map( B1 => n962, B2 => n1803, C1 => n996, C2 => n1804
                           , A => n1923, ZN => n1920);
   U2443 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_25_port, B1 => 
                           n1807, B2 => REGISTERS_6_25_port, ZN => n1923);
   U2444 : OAI221_X1 port map( B1 => n821, B2 => n1808, C1 => n855, C2 => n1809
                           , A => n1924, ZN => n1919);
   U2445 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_25_port, B1 => 
                           n1812, B2 => REGISTERS_10_25_port, ZN => n1924);
   U2446 : OAI221_X1 port map( B1 => n685, B2 => n1813, C1 => n719, C2 => n1814
                           , A => n1925, ZN => n1918);
   U2447 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_25_port, B1 => 
                           n1817, B2 => REGISTERS_14_25_port, ZN => n1925);
   U2448 : AOI21_X1 port map( B1 => n1926, B2 => n1927, A => N352, ZN => N311);
   U2449 : NOR4_X1 port map( A1 => n1928, A2 => n1929, A3 => n1930, A4 => n1931
                           , ZN => n1927);
   U2450 : OAI221_X1 port map( B1 => n546, B2 => n1774, C1 => n580, C2 => n1775
                           , A => n1932, ZN => n1931);
   U2451 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_24_port, B1 => 
                           n1778, B2 => REGISTERS_18_24_port, ZN => n1932);
   U2452 : OAI221_X1 port map( B1 => n410, B2 => n1779, C1 => n444, C2 => n1780
                           , A => n1933, ZN => n1930);
   U2453 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_24_port, B1 => 
                           n1783, B2 => REGISTERS_22_24_port, ZN => n1933);
   U2454 : OAI221_X1 port map( B1 => n270, B2 => n1784, C1 => n305_port, C2 => 
                           n1785, A => n1934, ZN => n1929);
   U2455 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_24_port, B1 => 
                           n1788, B2 => REGISTERS_26_24_port, ZN => n1934);
   U2456 : OAI221_X1 port map( B1 => n52, B2 => n1789, C1 => n95, C2 => n1790, 
                           A => n1935, ZN => n1928);
   U2457 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_24_port, B1 => 
                           n1793, B2 => REGISTERS_28_24_port, ZN => n1935);
   U2458 : NOR4_X1 port map( A1 => n1936, A2 => n1937, A3 => n1938, A4 => n1939
                           , ZN => n1926);
   U2459 : OAI221_X1 port map( B1 => n1097, B2 => n1798, C1 => n1131, C2 => 
                           n1799, A => n1940, ZN => n1939);
   U2460 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_24_port, B1 => 
                           n1802, B2 => REGISTERS_2_24_port, ZN => n1940);
   U2461 : OAI221_X1 port map( B1 => n961, B2 => n1803, C1 => n995, C2 => n1804
                           , A => n1941, ZN => n1938);
   U2462 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_24_port, B1 => 
                           n1807, B2 => REGISTERS_6_24_port, ZN => n1941);
   U2463 : OAI221_X1 port map( B1 => n820, B2 => n1808, C1 => n854, C2 => n1809
                           , A => n1942, ZN => n1937);
   U2464 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_24_port, B1 => 
                           n1812, B2 => REGISTERS_10_24_port, ZN => n1942);
   U2465 : OAI221_X1 port map( B1 => n684, B2 => n1813, C1 => n718, C2 => n1814
                           , A => n1943, ZN => n1936);
   U2466 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_24_port, B1 => 
                           n1817, B2 => REGISTERS_14_24_port, ZN => n1943);
   U2467 : AOI21_X1 port map( B1 => n1944, B2 => n1945, A => N352, ZN => N310);
   U2468 : NOR4_X1 port map( A1 => n1946, A2 => n1947, A3 => n1948, A4 => n1949
                           , ZN => n1945);
   U2469 : OAI221_X1 port map( B1 => n545, B2 => n1774, C1 => n579, C2 => n1775
                           , A => n1950, ZN => n1949);
   U2470 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_23_port, B1 => 
                           n1778, B2 => REGISTERS_18_23_port, ZN => n1950);
   U2471 : OAI221_X1 port map( B1 => n409, B2 => n1779, C1 => n443, C2 => n1780
                           , A => n1951, ZN => n1948);
   U2472 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_23_port, B1 => 
                           n1783, B2 => REGISTERS_22_23_port, ZN => n1951);
   U2473 : OAI221_X1 port map( B1 => n269, B2 => n1784, C1 => n304_port, C2 => 
                           n1785, A => n1952, ZN => n1947);
   U2474 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_23_port, B1 => 
                           n1788, B2 => REGISTERS_26_23_port, ZN => n1952);
   U2475 : OAI221_X1 port map( B1 => n50, B2 => n1789, C1 => n94, C2 => n1790, 
                           A => n1953, ZN => n1946);
   U2476 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_23_port, B1 => 
                           n1793, B2 => REGISTERS_28_23_port, ZN => n1953);
   U2477 : NOR4_X1 port map( A1 => n1954, A2 => n1955, A3 => n1956, A4 => n1957
                           , ZN => n1944);
   U2478 : OAI221_X1 port map( B1 => n1096, B2 => n1798, C1 => n1130, C2 => 
                           n1799, A => n1958, ZN => n1957);
   U2479 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_23_port, B1 => 
                           n1802, B2 => REGISTERS_2_23_port, ZN => n1958);
   U2480 : OAI221_X1 port map( B1 => n960, B2 => n1803, C1 => n994, C2 => n1804
                           , A => n1959, ZN => n1956);
   U2481 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_23_port, B1 => 
                           n1807, B2 => REGISTERS_6_23_port, ZN => n1959);
   U2482 : OAI221_X1 port map( B1 => n819, B2 => n1808, C1 => n853, C2 => n1809
                           , A => n1960, ZN => n1955);
   U2483 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_23_port, B1 => 
                           n1812, B2 => REGISTERS_10_23_port, ZN => n1960);
   U2484 : OAI221_X1 port map( B1 => n683, B2 => n1813, C1 => n717, C2 => n1814
                           , A => n1961, ZN => n1954);
   U2485 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_23_port, B1 => 
                           n1817, B2 => REGISTERS_14_23_port, ZN => n1961);
   U2486 : AOI21_X1 port map( B1 => n1962, B2 => n1963, A => N352, ZN => N309);
   U2487 : NOR4_X1 port map( A1 => n1964, A2 => n1965, A3 => n1966, A4 => n1967
                           , ZN => n1963);
   U2488 : OAI221_X1 port map( B1 => n544, B2 => n1774, C1 => n578, C2 => n1775
                           , A => n1968, ZN => n1967);
   U2489 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_22_port, B1 => 
                           n1778, B2 => REGISTERS_18_22_port, ZN => n1968);
   U2490 : OAI221_X1 port map( B1 => n408, B2 => n1779, C1 => n442, C2 => n1780
                           , A => n1969, ZN => n1966);
   U2491 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_22_port, B1 => 
                           n1783, B2 => REGISTERS_22_22_port, ZN => n1969);
   U2492 : OAI221_X1 port map( B1 => n268, B2 => n1784, C1 => n303_port, C2 => 
                           n1785, A => n1970, ZN => n1965);
   U2493 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_22_port, B1 => 
                           n1788, B2 => REGISTERS_26_22_port, ZN => n1970);
   U2494 : OAI221_X1 port map( B1 => n48, B2 => n1789, C1 => n93, C2 => n1790, 
                           A => n1971, ZN => n1964);
   U2495 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_22_port, B1 => 
                           n1793, B2 => REGISTERS_28_22_port, ZN => n1971);
   U2496 : NOR4_X1 port map( A1 => n1972, A2 => n1973, A3 => n1974, A4 => n1975
                           , ZN => n1962);
   U2497 : OAI221_X1 port map( B1 => n1095, B2 => n1798, C1 => n1129, C2 => 
                           n1799, A => n1976, ZN => n1975);
   U2498 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_22_port, B1 => 
                           n1802, B2 => REGISTERS_2_22_port, ZN => n1976);
   U2499 : OAI221_X1 port map( B1 => n959, B2 => n1803, C1 => n993, C2 => n1804
                           , A => n1977, ZN => n1974);
   U2500 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_22_port, B1 => 
                           n1807, B2 => REGISTERS_6_22_port, ZN => n1977);
   U2501 : OAI221_X1 port map( B1 => n818, B2 => n1808, C1 => n852, C2 => n1809
                           , A => n1978, ZN => n1973);
   U2502 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_22_port, B1 => 
                           n1812, B2 => REGISTERS_10_22_port, ZN => n1978);
   U2503 : OAI221_X1 port map( B1 => n682, B2 => n1813, C1 => n716, C2 => n1814
                           , A => n1979, ZN => n1972);
   U2504 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_22_port, B1 => 
                           n1817, B2 => REGISTERS_14_22_port, ZN => n1979);
   U2505 : AOI21_X1 port map( B1 => n1980, B2 => n1981, A => N352, ZN => N308);
   U2506 : NOR4_X1 port map( A1 => n1982, A2 => n1983, A3 => n1984, A4 => n1985
                           , ZN => n1981);
   U2507 : OAI221_X1 port map( B1 => n543, B2 => n1774, C1 => n577, C2 => n1775
                           , A => n1986, ZN => n1985);
   U2508 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_21_port, B1 => 
                           n1778, B2 => REGISTERS_18_21_port, ZN => n1986);
   U2509 : OAI221_X1 port map( B1 => n407, B2 => n1779, C1 => n441, C2 => n1780
                           , A => n1987, ZN => n1984);
   U2510 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_21_port, B1 => 
                           n1783, B2 => REGISTERS_22_21_port, ZN => n1987);
   U2511 : OAI221_X1 port map( B1 => n267, B2 => n1784, C1 => n302_port, C2 => 
                           n1785, A => n1988, ZN => n1983);
   U2512 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_21_port, B1 => 
                           n1788, B2 => REGISTERS_26_21_port, ZN => n1988);
   U2513 : OAI221_X1 port map( B1 => n46, B2 => n1789, C1 => n92, C2 => n1790, 
                           A => n1989, ZN => n1982);
   U2514 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_21_port, B1 => 
                           n1793, B2 => REGISTERS_28_21_port, ZN => n1989);
   U2515 : NOR4_X1 port map( A1 => n1990, A2 => n1991, A3 => n1992, A4 => n1993
                           , ZN => n1980);
   U2516 : OAI221_X1 port map( B1 => n1094, B2 => n1798, C1 => n1128, C2 => 
                           n1799, A => n1994, ZN => n1993);
   U2517 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_21_port, B1 => 
                           n1802, B2 => REGISTERS_2_21_port, ZN => n1994);
   U2518 : OAI221_X1 port map( B1 => n958, B2 => n1803, C1 => n992, C2 => n1804
                           , A => n1995, ZN => n1992);
   U2519 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_21_port, B1 => 
                           n1807, B2 => REGISTERS_6_21_port, ZN => n1995);
   U2520 : OAI221_X1 port map( B1 => n817, B2 => n1808, C1 => n851, C2 => n1809
                           , A => n1996, ZN => n1991);
   U2521 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_21_port, B1 => 
                           n1812, B2 => REGISTERS_10_21_port, ZN => n1996);
   U2522 : OAI221_X1 port map( B1 => n681, B2 => n1813, C1 => n715, C2 => n1814
                           , A => n1997, ZN => n1990);
   U2523 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_21_port, B1 => 
                           n1817, B2 => REGISTERS_14_21_port, ZN => n1997);
   U2524 : AOI21_X1 port map( B1 => n1998, B2 => n1999, A => N352, ZN => N307);
   U2525 : NOR4_X1 port map( A1 => n2000, A2 => n2001, A3 => n2002, A4 => n2003
                           , ZN => n1999);
   U2526 : OAI221_X1 port map( B1 => n542, B2 => n1774, C1 => n576, C2 => n1775
                           , A => n2004, ZN => n2003);
   U2527 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_20_port, B1 => 
                           n1778, B2 => REGISTERS_18_20_port, ZN => n2004);
   U2528 : OAI221_X1 port map( B1 => n406, B2 => n1779, C1 => n440, C2 => n1780
                           , A => n2005, ZN => n2002);
   U2529 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_20_port, B1 => 
                           n1783, B2 => REGISTERS_22_20_port, ZN => n2005);
   U2530 : OAI221_X1 port map( B1 => n266, B2 => n1784, C1 => n301_port, C2 => 
                           n1785, A => n2006, ZN => n2001);
   U2531 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_20_port, B1 => 
                           n1788, B2 => REGISTERS_26_20_port, ZN => n2006);
   U2532 : OAI221_X1 port map( B1 => n44, B2 => n1789, C1 => n91, C2 => n1790, 
                           A => n2007, ZN => n2000);
   U2533 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_20_port, B1 => 
                           n1793, B2 => REGISTERS_28_20_port, ZN => n2007);
   U2534 : NOR4_X1 port map( A1 => n2008, A2 => n2009, A3 => n2010, A4 => n2011
                           , ZN => n1998);
   U2535 : OAI221_X1 port map( B1 => n1093, B2 => n1798, C1 => n1127, C2 => 
                           n1799, A => n2012, ZN => n2011);
   U2536 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_20_port, B1 => 
                           n1802, B2 => REGISTERS_2_20_port, ZN => n2012);
   U2537 : OAI221_X1 port map( B1 => n957, B2 => n1803, C1 => n991, C2 => n1804
                           , A => n2013, ZN => n2010);
   U2538 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_20_port, B1 => 
                           n1807, B2 => REGISTERS_6_20_port, ZN => n2013);
   U2539 : OAI221_X1 port map( B1 => n816, B2 => n1808, C1 => n850, C2 => n1809
                           , A => n2014, ZN => n2009);
   U2540 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_20_port, B1 => 
                           n1812, B2 => REGISTERS_10_20_port, ZN => n2014);
   U2541 : OAI221_X1 port map( B1 => n680, B2 => n1813, C1 => n714, C2 => n1814
                           , A => n2015, ZN => n2008);
   U2542 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_20_port, B1 => 
                           n1817, B2 => REGISTERS_14_20_port, ZN => n2015);
   U2543 : AOI21_X1 port map( B1 => n2016, B2 => n2017, A => N352, ZN => N306);
   U2544 : NOR4_X1 port map( A1 => n2018, A2 => n2019, A3 => n2020, A4 => n2021
                           , ZN => n2017);
   U2545 : OAI221_X1 port map( B1 => n541, B2 => n1774, C1 => n575, C2 => n1775
                           , A => n2022, ZN => n2021);
   U2546 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_19_port, B1 => 
                           n1778, B2 => REGISTERS_18_19_port, ZN => n2022);
   U2547 : OAI221_X1 port map( B1 => n405, B2 => n1779, C1 => n439, C2 => n1780
                           , A => n2023, ZN => n2020);
   U2548 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_19_port, B1 => 
                           n1783, B2 => REGISTERS_22_19_port, ZN => n2023);
   U2549 : OAI221_X1 port map( B1 => n265, B2 => n1784, C1 => n300_port, C2 => 
                           n1785, A => n2024, ZN => n2019);
   U2550 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_19_port, B1 => 
                           n1788, B2 => REGISTERS_26_19_port, ZN => n2024);
   U2551 : OAI221_X1 port map( B1 => n42, B2 => n1789, C1 => n90, C2 => n1790, 
                           A => n2025, ZN => n2018);
   U2552 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_19_port, B1 => 
                           n1793, B2 => REGISTERS_28_19_port, ZN => n2025);
   U2553 : NOR4_X1 port map( A1 => n2026, A2 => n2027, A3 => n2028, A4 => n2029
                           , ZN => n2016);
   U2554 : OAI221_X1 port map( B1 => n1092, B2 => n1798, C1 => n1126, C2 => 
                           n1799, A => n2030, ZN => n2029);
   U2555 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_19_port, B1 => 
                           n1802, B2 => REGISTERS_2_19_port, ZN => n2030);
   U2556 : OAI221_X1 port map( B1 => n956, B2 => n1803, C1 => n990, C2 => n1804
                           , A => n2031, ZN => n2028);
   U2557 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_19_port, B1 => 
                           n1807, B2 => REGISTERS_6_19_port, ZN => n2031);
   U2558 : OAI221_X1 port map( B1 => n815, B2 => n1808, C1 => n849, C2 => n1809
                           , A => n2032, ZN => n2027);
   U2559 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_19_port, B1 => 
                           n1812, B2 => REGISTERS_10_19_port, ZN => n2032);
   U2560 : OAI221_X1 port map( B1 => n679, B2 => n1813, C1 => n713, C2 => n1814
                           , A => n2033, ZN => n2026);
   U2561 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_19_port, B1 => 
                           n1817, B2 => REGISTERS_14_19_port, ZN => n2033);
   U2562 : AOI21_X1 port map( B1 => n2034, B2 => n2035, A => N352, ZN => N305);
   U2563 : NOR4_X1 port map( A1 => n2036, A2 => n2037, A3 => n2038, A4 => n2039
                           , ZN => n2035);
   U2564 : OAI221_X1 port map( B1 => n540, B2 => n1774, C1 => n574, C2 => n1775
                           , A => n2040, ZN => n2039);
   U2565 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_18_port, B1 => 
                           n1778, B2 => REGISTERS_18_18_port, ZN => n2040);
   U2566 : OAI221_X1 port map( B1 => n404, B2 => n1779, C1 => n438, C2 => n1780
                           , A => n2041, ZN => n2038);
   U2567 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_18_port, B1 => 
                           n1783, B2 => REGISTERS_22_18_port, ZN => n2041);
   U2568 : OAI221_X1 port map( B1 => n264, B2 => n1784, C1 => n299_port, C2 => 
                           n1785, A => n2042, ZN => n2037);
   U2569 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_18_port, B1 => 
                           n1788, B2 => REGISTERS_26_18_port, ZN => n2042);
   U2570 : OAI221_X1 port map( B1 => n40, B2 => n1789, C1 => n89, C2 => n1790, 
                           A => n2043, ZN => n2036);
   U2571 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_18_port, B1 => 
                           n1793, B2 => REGISTERS_28_18_port, ZN => n2043);
   U2572 : NOR4_X1 port map( A1 => n2044, A2 => n2045, A3 => n2046, A4 => n2047
                           , ZN => n2034);
   U2573 : OAI221_X1 port map( B1 => n1091, B2 => n1798, C1 => n1125, C2 => 
                           n1799, A => n2048, ZN => n2047);
   U2574 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_18_port, B1 => 
                           n1802, B2 => REGISTERS_2_18_port, ZN => n2048);
   U2575 : OAI221_X1 port map( B1 => n955, B2 => n1803, C1 => n989, C2 => n1804
                           , A => n2049, ZN => n2046);
   U2576 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_18_port, B1 => 
                           n1807, B2 => REGISTERS_6_18_port, ZN => n2049);
   U2577 : OAI221_X1 port map( B1 => n814, B2 => n1808, C1 => n848, C2 => n1809
                           , A => n2050, ZN => n2045);
   U2578 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_18_port, B1 => 
                           n1812, B2 => REGISTERS_10_18_port, ZN => n2050);
   U2579 : OAI221_X1 port map( B1 => n678, B2 => n1813, C1 => n712, C2 => n1814
                           , A => n2051, ZN => n2044);
   U2580 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_18_port, B1 => 
                           n1817, B2 => REGISTERS_14_18_port, ZN => n2051);
   U2581 : AOI21_X1 port map( B1 => n2052, B2 => n2053, A => N352, ZN => N304);
   U2582 : NOR4_X1 port map( A1 => n2054, A2 => n2055, A3 => n2056, A4 => n2057
                           , ZN => n2053);
   U2583 : OAI221_X1 port map( B1 => n539, B2 => n1774, C1 => n573, C2 => n1775
                           , A => n2058, ZN => n2057);
   U2584 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_17_port, B1 => 
                           n1778, B2 => REGISTERS_18_17_port, ZN => n2058);
   U2585 : OAI221_X1 port map( B1 => n403, B2 => n1779, C1 => n437, C2 => n1780
                           , A => n2059, ZN => n2056);
   U2586 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_17_port, B1 => 
                           n1783, B2 => REGISTERS_22_17_port, ZN => n2059);
   U2587 : OAI221_X1 port map( B1 => n263, B2 => n1784, C1 => n298_port, C2 => 
                           n1785, A => n2060, ZN => n2055);
   U2588 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_17_port, B1 => 
                           n1788, B2 => REGISTERS_26_17_port, ZN => n2060);
   U2589 : OAI221_X1 port map( B1 => n38, B2 => n1789, C1 => n88, C2 => n1790, 
                           A => n2061, ZN => n2054);
   U2590 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_17_port, B1 => 
                           n1793, B2 => REGISTERS_28_17_port, ZN => n2061);
   U2591 : NOR4_X1 port map( A1 => n2062, A2 => n2063, A3 => n2064, A4 => n2065
                           , ZN => n2052);
   U2592 : OAI221_X1 port map( B1 => n1090, B2 => n1798, C1 => n1124, C2 => 
                           n1799, A => n2066, ZN => n2065);
   U2593 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_17_port, B1 => 
                           n1802, B2 => REGISTERS_2_17_port, ZN => n2066);
   U2594 : OAI221_X1 port map( B1 => n954, B2 => n1803, C1 => n988, C2 => n1804
                           , A => n2067, ZN => n2064);
   U2595 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_17_port, B1 => 
                           n1807, B2 => REGISTERS_6_17_port, ZN => n2067);
   U2596 : OAI221_X1 port map( B1 => n813, B2 => n1808, C1 => n847, C2 => n1809
                           , A => n2068, ZN => n2063);
   U2597 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_17_port, B1 => 
                           n1812, B2 => REGISTERS_10_17_port, ZN => n2068);
   U2598 : OAI221_X1 port map( B1 => n677, B2 => n1813, C1 => n711, C2 => n1814
                           , A => n2069, ZN => n2062);
   U2599 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_17_port, B1 => 
                           n1817, B2 => REGISTERS_14_17_port, ZN => n2069);
   U2600 : AOI21_X1 port map( B1 => n2070, B2 => n2071, A => N352, ZN => N303);
   U2601 : NOR4_X1 port map( A1 => n2072, A2 => n2073, A3 => n2074, A4 => n2075
                           , ZN => n2071);
   U2602 : OAI221_X1 port map( B1 => n538, B2 => n1774, C1 => n572, C2 => n1775
                           , A => n2076, ZN => n2075);
   U2603 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_16_port, B1 => 
                           n1778, B2 => REGISTERS_18_16_port, ZN => n2076);
   U2604 : OAI221_X1 port map( B1 => n402, B2 => n1779, C1 => n436, C2 => n1780
                           , A => n2077, ZN => n2074);
   U2605 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_16_port, B1 => 
                           n1783, B2 => REGISTERS_22_16_port, ZN => n2077);
   U2606 : OAI221_X1 port map( B1 => n262, B2 => n1784, C1 => n297_port, C2 => 
                           n1785, A => n2078, ZN => n2073);
   U2607 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_16_port, B1 => 
                           n1788, B2 => REGISTERS_26_16_port, ZN => n2078);
   U2608 : OAI221_X1 port map( B1 => n36, B2 => n1789, C1 => n87, C2 => n1790, 
                           A => n2079, ZN => n2072);
   U2609 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_16_port, B1 => 
                           n1793, B2 => REGISTERS_28_16_port, ZN => n2079);
   U2610 : NOR4_X1 port map( A1 => n2080, A2 => n2081, A3 => n2082, A4 => n2083
                           , ZN => n2070);
   U2611 : OAI221_X1 port map( B1 => n1089, B2 => n1798, C1 => n1123, C2 => 
                           n1799, A => n2084, ZN => n2083);
   U2612 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_16_port, B1 => 
                           n1802, B2 => REGISTERS_2_16_port, ZN => n2084);
   U2613 : OAI221_X1 port map( B1 => n953, B2 => n1803, C1 => n987, C2 => n1804
                           , A => n2085, ZN => n2082);
   U2614 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_16_port, B1 => 
                           n1807, B2 => REGISTERS_6_16_port, ZN => n2085);
   U2615 : OAI221_X1 port map( B1 => n812, B2 => n1808, C1 => n846, C2 => n1809
                           , A => n2086, ZN => n2081);
   U2616 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_16_port, B1 => 
                           n1812, B2 => REGISTERS_10_16_port, ZN => n2086);
   U2617 : OAI221_X1 port map( B1 => n676, B2 => n1813, C1 => n710, C2 => n1814
                           , A => n2087, ZN => n2080);
   U2618 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_16_port, B1 => 
                           n1817, B2 => REGISTERS_14_16_port, ZN => n2087);
   U2619 : AOI21_X1 port map( B1 => n2088, B2 => n2089, A => N352, ZN => N302);
   U2620 : NOR4_X1 port map( A1 => n2090, A2 => n2091, A3 => n2092, A4 => n2093
                           , ZN => n2089);
   U2621 : OAI221_X1 port map( B1 => n537, B2 => n1774, C1 => n571, C2 => n1775
                           , A => n2094, ZN => n2093);
   U2622 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_15_port, B1 => 
                           n1778, B2 => REGISTERS_18_15_port, ZN => n2094);
   U2623 : OAI221_X1 port map( B1 => n401, B2 => n1779, C1 => n435, C2 => n1780
                           , A => n2095, ZN => n2092);
   U2624 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_15_port, B1 => 
                           n1783, B2 => REGISTERS_22_15_port, ZN => n2095);
   U2625 : OAI221_X1 port map( B1 => n261, B2 => n1784, C1 => n296_port, C2 => 
                           n1785, A => n2096, ZN => n2091);
   U2626 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_15_port, B1 => 
                           n1788, B2 => REGISTERS_26_15_port, ZN => n2096);
   U2627 : OAI221_X1 port map( B1 => n34, B2 => n1789, C1 => n86, C2 => n1790, 
                           A => n2097, ZN => n2090);
   U2628 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_15_port, B1 => 
                           n1793, B2 => REGISTERS_28_15_port, ZN => n2097);
   U2629 : NOR4_X1 port map( A1 => n2098, A2 => n2099, A3 => n2100, A4 => n2101
                           , ZN => n2088);
   U2630 : OAI221_X1 port map( B1 => n1088, B2 => n1798, C1 => n1122, C2 => 
                           n1799, A => n2102, ZN => n2101);
   U2631 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_15_port, B1 => 
                           n1802, B2 => REGISTERS_2_15_port, ZN => n2102);
   U2632 : OAI221_X1 port map( B1 => n952, B2 => n1803, C1 => n986, C2 => n1804
                           , A => n2103, ZN => n2100);
   U2633 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_15_port, B1 => 
                           n1807, B2 => REGISTERS_6_15_port, ZN => n2103);
   U2634 : OAI221_X1 port map( B1 => n811, B2 => n1808, C1 => n845, C2 => n1809
                           , A => n2104, ZN => n2099);
   U2635 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_15_port, B1 => 
                           n1812, B2 => REGISTERS_10_15_port, ZN => n2104);
   U2636 : OAI221_X1 port map( B1 => n675, B2 => n1813, C1 => n709, C2 => n1814
                           , A => n2105, ZN => n2098);
   U2637 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_15_port, B1 => 
                           n1817, B2 => REGISTERS_14_15_port, ZN => n2105);
   U2638 : AOI21_X1 port map( B1 => n2106, B2 => n2107, A => N352, ZN => N301);
   U2639 : NOR4_X1 port map( A1 => n2108, A2 => n2109, A3 => n2110, A4 => n2111
                           , ZN => n2107);
   U2640 : OAI221_X1 port map( B1 => n536, B2 => n1774, C1 => n570, C2 => n1775
                           , A => n2112, ZN => n2111);
   U2641 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_14_port, B1 => 
                           n1778, B2 => REGISTERS_18_14_port, ZN => n2112);
   U2642 : OAI221_X1 port map( B1 => n400, B2 => n1779, C1 => n434, C2 => n1780
                           , A => n2113, ZN => n2110);
   U2643 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_14_port, B1 => 
                           n1783, B2 => REGISTERS_22_14_port, ZN => n2113);
   U2644 : OAI221_X1 port map( B1 => n260, B2 => n1784, C1 => n295_port, C2 => 
                           n1785, A => n2114, ZN => n2109);
   U2645 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_14_port, B1 => 
                           n1788, B2 => REGISTERS_26_14_port, ZN => n2114);
   U2646 : OAI221_X1 port map( B1 => n32, B2 => n1789, C1 => n85, C2 => n1790, 
                           A => n2115, ZN => n2108);
   U2647 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_14_port, B1 => 
                           n1793, B2 => REGISTERS_28_14_port, ZN => n2115);
   U2648 : NOR4_X1 port map( A1 => n2116, A2 => n2117, A3 => n2118, A4 => n2119
                           , ZN => n2106);
   U2649 : OAI221_X1 port map( B1 => n1087, B2 => n1798, C1 => n1121, C2 => 
                           n1799, A => n2120, ZN => n2119);
   U2650 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_14_port, B1 => 
                           n1802, B2 => REGISTERS_2_14_port, ZN => n2120);
   U2651 : OAI221_X1 port map( B1 => n951, B2 => n1803, C1 => n985, C2 => n1804
                           , A => n2121, ZN => n2118);
   U2652 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_14_port, B1 => 
                           n1807, B2 => REGISTERS_6_14_port, ZN => n2121);
   U2653 : OAI221_X1 port map( B1 => n810, B2 => n1808, C1 => n844, C2 => n1809
                           , A => n2122, ZN => n2117);
   U2654 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_14_port, B1 => 
                           n1812, B2 => REGISTERS_10_14_port, ZN => n2122);
   U2655 : OAI221_X1 port map( B1 => n674, B2 => n1813, C1 => n708, C2 => n1814
                           , A => n2123, ZN => n2116);
   U2656 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_14_port, B1 => 
                           n1817, B2 => REGISTERS_14_14_port, ZN => n2123);
   U2657 : AOI21_X1 port map( B1 => n2124, B2 => n2125, A => N352, ZN => N300);
   U2658 : NOR4_X1 port map( A1 => n2126, A2 => n2127, A3 => n2128, A4 => n2129
                           , ZN => n2125);
   U2659 : OAI221_X1 port map( B1 => n535, B2 => n1774, C1 => n569, C2 => n1775
                           , A => n2130, ZN => n2129);
   U2660 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_13_port, B1 => 
                           n1778, B2 => REGISTERS_18_13_port, ZN => n2130);
   U2661 : OAI221_X1 port map( B1 => n399, B2 => n1779, C1 => n433, C2 => n1780
                           , A => n2131, ZN => n2128);
   U2662 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_13_port, B1 => 
                           n1783, B2 => REGISTERS_22_13_port, ZN => n2131);
   U2663 : OAI221_X1 port map( B1 => n259, B2 => n1784, C1 => n294_port, C2 => 
                           n1785, A => n2132, ZN => n2127);
   U2664 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_13_port, B1 => 
                           n1788, B2 => REGISTERS_26_13_port, ZN => n2132);
   U2665 : OAI221_X1 port map( B1 => n30, B2 => n1789, C1 => n84, C2 => n1790, 
                           A => n2133, ZN => n2126);
   U2666 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_13_port, B1 => 
                           n1793, B2 => REGISTERS_28_13_port, ZN => n2133);
   U2667 : NOR4_X1 port map( A1 => n2134, A2 => n2135, A3 => n2136, A4 => n2137
                           , ZN => n2124);
   U2668 : OAI221_X1 port map( B1 => n1086, B2 => n1798, C1 => n1120, C2 => 
                           n1799, A => n2138, ZN => n2137);
   U2669 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_13_port, B1 => 
                           n1802, B2 => REGISTERS_2_13_port, ZN => n2138);
   U2670 : OAI221_X1 port map( B1 => n950, B2 => n1803, C1 => n984, C2 => n1804
                           , A => n2139, ZN => n2136);
   U2671 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_13_port, B1 => 
                           n1807, B2 => REGISTERS_6_13_port, ZN => n2139);
   U2672 : OAI221_X1 port map( B1 => n809, B2 => n1808, C1 => n843, C2 => n1809
                           , A => n2140, ZN => n2135);
   U2673 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_13_port, B1 => 
                           n1812, B2 => REGISTERS_10_13_port, ZN => n2140);
   U2674 : OAI221_X1 port map( B1 => n673, B2 => n1813, C1 => n707, C2 => n1814
                           , A => n2141, ZN => n2134);
   U2675 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_13_port, B1 => 
                           n1817, B2 => REGISTERS_14_13_port, ZN => n2141);
   U2676 : AOI21_X1 port map( B1 => n2142, B2 => n2143, A => N352, ZN => N299);
   U2677 : NOR4_X1 port map( A1 => n2144, A2 => n2145, A3 => n2146, A4 => n2147
                           , ZN => n2143);
   U2678 : OAI221_X1 port map( B1 => n534, B2 => n1774, C1 => n568, C2 => n1775
                           , A => n2148, ZN => n2147);
   U2679 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_12_port, B1 => 
                           n1778, B2 => REGISTERS_18_12_port, ZN => n2148);
   U2680 : OAI221_X1 port map( B1 => n398, B2 => n1779, C1 => n432, C2 => n1780
                           , A => n2149, ZN => n2146);
   U2681 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_12_port, B1 => 
                           n1783, B2 => REGISTERS_22_12_port, ZN => n2149);
   U2682 : OAI221_X1 port map( B1 => n258, B2 => n1784, C1 => n293_port, C2 => 
                           n1785, A => n2150, ZN => n2145);
   U2683 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_12_port, B1 => 
                           n1788, B2 => REGISTERS_26_12_port, ZN => n2150);
   U2684 : OAI221_X1 port map( B1 => n28, B2 => n1789, C1 => n83, C2 => n1790, 
                           A => n2151, ZN => n2144);
   U2685 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_12_port, B1 => 
                           n1793, B2 => REGISTERS_28_12_port, ZN => n2151);
   U2686 : NOR4_X1 port map( A1 => n2152, A2 => n2153, A3 => n2154, A4 => n2155
                           , ZN => n2142);
   U2687 : OAI221_X1 port map( B1 => n1085, B2 => n1798, C1 => n1119, C2 => 
                           n1799, A => n2156, ZN => n2155);
   U2688 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_12_port, B1 => 
                           n1802, B2 => REGISTERS_2_12_port, ZN => n2156);
   U2689 : OAI221_X1 port map( B1 => n949, B2 => n1803, C1 => n983, C2 => n1804
                           , A => n2157, ZN => n2154);
   U2690 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_12_port, B1 => 
                           n1807, B2 => REGISTERS_6_12_port, ZN => n2157);
   U2691 : OAI221_X1 port map( B1 => n808, B2 => n1808, C1 => n842, C2 => n1809
                           , A => n2158, ZN => n2153);
   U2692 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_12_port, B1 => 
                           n1812, B2 => REGISTERS_10_12_port, ZN => n2158);
   U2693 : OAI221_X1 port map( B1 => n672, B2 => n1813, C1 => n706, C2 => n1814
                           , A => n2159, ZN => n2152);
   U2694 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_12_port, B1 => 
                           n1817, B2 => REGISTERS_14_12_port, ZN => n2159);
   U2695 : AOI21_X1 port map( B1 => n2160, B2 => n2161, A => N352, ZN => N298);
   U2696 : NOR4_X1 port map( A1 => n2162, A2 => n2163, A3 => n2164, A4 => n2165
                           , ZN => n2161);
   U2697 : OAI221_X1 port map( B1 => n533, B2 => n1774, C1 => n567, C2 => n1775
                           , A => n2166, ZN => n2165);
   U2698 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_11_port, B1 => 
                           n1778, B2 => REGISTERS_18_11_port, ZN => n2166);
   U2699 : OAI221_X1 port map( B1 => n397, B2 => n1779, C1 => n431, C2 => n1780
                           , A => n2167, ZN => n2164);
   U2700 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_11_port, B1 => 
                           n1783, B2 => REGISTERS_22_11_port, ZN => n2167);
   U2701 : OAI221_X1 port map( B1 => n257, B2 => n1784, C1 => n292_port, C2 => 
                           n1785, A => n2168, ZN => n2163);
   U2702 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_11_port, B1 => 
                           n1788, B2 => REGISTERS_26_11_port, ZN => n2168);
   U2703 : OAI221_X1 port map( B1 => n26, B2 => n1789, C1 => n82, C2 => n1790, 
                           A => n2169, ZN => n2162);
   U2704 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_11_port, B1 => 
                           n1793, B2 => REGISTERS_28_11_port, ZN => n2169);
   U2705 : NOR4_X1 port map( A1 => n2170, A2 => n2171, A3 => n2172, A4 => n2173
                           , ZN => n2160);
   U2706 : OAI221_X1 port map( B1 => n1084, B2 => n1798, C1 => n1118, C2 => 
                           n1799, A => n2174, ZN => n2173);
   U2707 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_11_port, B1 => 
                           n1802, B2 => REGISTERS_2_11_port, ZN => n2174);
   U2708 : OAI221_X1 port map( B1 => n948, B2 => n1803, C1 => n982, C2 => n1804
                           , A => n2175, ZN => n2172);
   U2709 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_11_port, B1 => 
                           n1807, B2 => REGISTERS_6_11_port, ZN => n2175);
   U2710 : OAI221_X1 port map( B1 => n807, B2 => n1808, C1 => n841, C2 => n1809
                           , A => n2176, ZN => n2171);
   U2711 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_11_port, B1 => 
                           n1812, B2 => REGISTERS_10_11_port, ZN => n2176);
   U2712 : OAI221_X1 port map( B1 => n671, B2 => n1813, C1 => n705, C2 => n1814
                           , A => n2177, ZN => n2170);
   U2713 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_11_port, B1 => 
                           n1817, B2 => REGISTERS_14_11_port, ZN => n2177);
   U2714 : AOI21_X1 port map( B1 => n2178, B2 => n2179, A => N352, ZN => N297);
   U2715 : NOR4_X1 port map( A1 => n2180, A2 => n2181, A3 => n2182, A4 => n2183
                           , ZN => n2179);
   U2716 : OAI221_X1 port map( B1 => n532, B2 => n1774, C1 => n566, C2 => n1775
                           , A => n2184, ZN => n2183);
   U2717 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_10_port, B1 => 
                           n1778, B2 => REGISTERS_18_10_port, ZN => n2184);
   U2718 : OAI221_X1 port map( B1 => n396, B2 => n1779, C1 => n430, C2 => n1780
                           , A => n2185, ZN => n2182);
   U2719 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_10_port, B1 => 
                           n1783, B2 => REGISTERS_22_10_port, ZN => n2185);
   U2720 : OAI221_X1 port map( B1 => n256, B2 => n1784, C1 => n291_port, C2 => 
                           n1785, A => n2186, ZN => n2181);
   U2721 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_10_port, B1 => 
                           n1788, B2 => REGISTERS_26_10_port, ZN => n2186);
   U2722 : OAI221_X1 port map( B1 => n24, B2 => n1789, C1 => n81, C2 => n1790, 
                           A => n2187, ZN => n2180);
   U2723 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_10_port, B1 => 
                           n1793, B2 => REGISTERS_28_10_port, ZN => n2187);
   U2724 : NOR4_X1 port map( A1 => n2188, A2 => n2189, A3 => n2190, A4 => n2191
                           , ZN => n2178);
   U2725 : OAI221_X1 port map( B1 => n1083, B2 => n1798, C1 => n1117, C2 => 
                           n1799, A => n2192, ZN => n2191);
   U2726 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_10_port, B1 => 
                           n1802, B2 => REGISTERS_2_10_port, ZN => n2192);
   U2727 : OAI221_X1 port map( B1 => n947, B2 => n1803, C1 => n981, C2 => n1804
                           , A => n2193, ZN => n2190);
   U2728 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_10_port, B1 => 
                           n1807, B2 => REGISTERS_6_10_port, ZN => n2193);
   U2729 : OAI221_X1 port map( B1 => n806, B2 => n1808, C1 => n840, C2 => n1809
                           , A => n2194, ZN => n2189);
   U2730 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_10_port, B1 => 
                           n1812, B2 => REGISTERS_10_10_port, ZN => n2194);
   U2731 : OAI221_X1 port map( B1 => n670, B2 => n1813, C1 => n704, C2 => n1814
                           , A => n2195, ZN => n2188);
   U2732 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_10_port, B1 => 
                           n1817, B2 => REGISTERS_14_10_port, ZN => n2195);
   U2733 : AOI21_X1 port map( B1 => n2196, B2 => n2197, A => N352, ZN => N296);
   U2734 : NOR4_X1 port map( A1 => n2198, A2 => n2199, A3 => n2200, A4 => n2201
                           , ZN => n2197);
   U2735 : OAI221_X1 port map( B1 => n531, B2 => n1774, C1 => n565, C2 => n1775
                           , A => n2202, ZN => n2201);
   U2736 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_9_port, B1 => 
                           n1778, B2 => REGISTERS_18_9_port, ZN => n2202);
   U2737 : OAI221_X1 port map( B1 => n395, B2 => n1779, C1 => n429, C2 => n1780
                           , A => n2203, ZN => n2200);
   U2738 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_9_port, B1 => 
                           n1783, B2 => REGISTERS_22_9_port, ZN => n2203);
   U2739 : OAI221_X1 port map( B1 => n255, B2 => n1784, C1 => n290_port, C2 => 
                           n1785, A => n2204, ZN => n2199);
   U2740 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_9_port, B1 => 
                           n1788, B2 => REGISTERS_26_9_port, ZN => n2204);
   U2741 : OAI221_X1 port map( B1 => n22, B2 => n1789, C1 => n80, C2 => n1790, 
                           A => n2205, ZN => n2198);
   U2742 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_9_port, B1 => 
                           n1793, B2 => REGISTERS_28_9_port, ZN => n2205);
   U2743 : NOR4_X1 port map( A1 => n2206, A2 => n2207, A3 => n2208, A4 => n2209
                           , ZN => n2196);
   U2744 : OAI221_X1 port map( B1 => n1082, B2 => n1798, C1 => n1116, C2 => 
                           n1799, A => n2210, ZN => n2209);
   U2745 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_9_port, B1 => 
                           n1802, B2 => REGISTERS_2_9_port, ZN => n2210);
   U2746 : OAI221_X1 port map( B1 => n946, B2 => n1803, C1 => n980, C2 => n1804
                           , A => n2211, ZN => n2208);
   U2747 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_9_port, B1 => 
                           n1807, B2 => REGISTERS_6_9_port, ZN => n2211);
   U2748 : OAI221_X1 port map( B1 => n805, B2 => n1808, C1 => n839, C2 => n1809
                           , A => n2212, ZN => n2207);
   U2749 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_9_port, B1 => 
                           n1812, B2 => REGISTERS_10_9_port, ZN => n2212);
   U2750 : OAI221_X1 port map( B1 => n669, B2 => n1813, C1 => n703, C2 => n1814
                           , A => n2213, ZN => n2206);
   U2751 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_9_port, B1 => 
                           n1817, B2 => REGISTERS_14_9_port, ZN => n2213);
   U2752 : AOI21_X1 port map( B1 => n2214, B2 => n2215, A => N352, ZN => N295);
   U2753 : NOR4_X1 port map( A1 => n2216, A2 => n2217, A3 => n2218, A4 => n2219
                           , ZN => n2215);
   U2754 : OAI221_X1 port map( B1 => n530, B2 => n1774, C1 => n564, C2 => n1775
                           , A => n2220, ZN => n2219);
   U2755 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_8_port, B1 => 
                           n1778, B2 => REGISTERS_18_8_port, ZN => n2220);
   U2756 : OAI221_X1 port map( B1 => n394, B2 => n1779, C1 => n428, C2 => n1780
                           , A => n2221, ZN => n2218);
   U2757 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_8_port, B1 => 
                           n1783, B2 => REGISTERS_22_8_port, ZN => n2221);
   U2758 : OAI221_X1 port map( B1 => n254, B2 => n1784, C1 => n289_port, C2 => 
                           n1785, A => n2222, ZN => n2217);
   U2759 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_8_port, B1 => 
                           n1788, B2 => REGISTERS_26_8_port, ZN => n2222);
   U2760 : OAI221_X1 port map( B1 => n20, B2 => n1789, C1 => n79, C2 => n1790, 
                           A => n2223, ZN => n2216);
   U2761 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_8_port, B1 => 
                           n1793, B2 => REGISTERS_28_8_port, ZN => n2223);
   U2762 : NOR4_X1 port map( A1 => n2224, A2 => n2225, A3 => n2226, A4 => n2227
                           , ZN => n2214);
   U2763 : OAI221_X1 port map( B1 => n1081, B2 => n1798, C1 => n1115, C2 => 
                           n1799, A => n2228, ZN => n2227);
   U2764 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_8_port, B1 => 
                           n1802, B2 => REGISTERS_2_8_port, ZN => n2228);
   U2765 : OAI221_X1 port map( B1 => n945, B2 => n1803, C1 => n979, C2 => n1804
                           , A => n2229, ZN => n2226);
   U2766 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_8_port, B1 => 
                           n1807, B2 => REGISTERS_6_8_port, ZN => n2229);
   U2767 : OAI221_X1 port map( B1 => n804, B2 => n1808, C1 => n838, C2 => n1809
                           , A => n2230, ZN => n2225);
   U2768 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_8_port, B1 => 
                           n1812, B2 => REGISTERS_10_8_port, ZN => n2230);
   U2769 : OAI221_X1 port map( B1 => n668, B2 => n1813, C1 => n702, C2 => n1814
                           , A => n2231, ZN => n2224);
   U2770 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_8_port, B1 => 
                           n1817, B2 => REGISTERS_14_8_port, ZN => n2231);
   U2771 : AOI21_X1 port map( B1 => n2232, B2 => n2233, A => N352, ZN => N294);
   U2772 : NOR4_X1 port map( A1 => n2234, A2 => n2235, A3 => n2236, A4 => n2237
                           , ZN => n2233);
   U2773 : OAI221_X1 port map( B1 => n529, B2 => n1774, C1 => n563, C2 => n1775
                           , A => n2238, ZN => n2237);
   U2774 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_7_port, B1 => 
                           n1778, B2 => REGISTERS_18_7_port, ZN => n2238);
   U2775 : OAI221_X1 port map( B1 => n393, B2 => n1779, C1 => n427, C2 => n1780
                           , A => n2239, ZN => n2236);
   U2776 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_7_port, B1 => 
                           n1783, B2 => REGISTERS_22_7_port, ZN => n2239);
   U2777 : OAI221_X1 port map( B1 => n253, B2 => n1784, C1 => n288_port, C2 => 
                           n1785, A => n2240, ZN => n2235);
   U2778 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_7_port, B1 => 
                           n1788, B2 => REGISTERS_26_7_port, ZN => n2240);
   U2779 : OAI221_X1 port map( B1 => n18, B2 => n1789, C1 => n78, C2 => n1790, 
                           A => n2241, ZN => n2234);
   U2780 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_7_port, B1 => 
                           n1793, B2 => REGISTERS_28_7_port, ZN => n2241);
   U2781 : NOR4_X1 port map( A1 => n2242, A2 => n2243, A3 => n2244, A4 => n2245
                           , ZN => n2232);
   U2782 : OAI221_X1 port map( B1 => n1080, B2 => n1798, C1 => n1114, C2 => 
                           n1799, A => n2246, ZN => n2245);
   U2783 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_7_port, B1 => 
                           n1802, B2 => REGISTERS_2_7_port, ZN => n2246);
   U2784 : OAI221_X1 port map( B1 => n944, B2 => n1803, C1 => n978, C2 => n1804
                           , A => n2247, ZN => n2244);
   U2785 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_7_port, B1 => 
                           n1807, B2 => REGISTERS_6_7_port, ZN => n2247);
   U2786 : OAI221_X1 port map( B1 => n803, B2 => n1808, C1 => n837, C2 => n1809
                           , A => n2248, ZN => n2243);
   U2787 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_7_port, B1 => 
                           n1812, B2 => REGISTERS_10_7_port, ZN => n2248);
   U2788 : OAI221_X1 port map( B1 => n667, B2 => n1813, C1 => n701, C2 => n1814
                           , A => n2249, ZN => n2242);
   U2789 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_7_port, B1 => 
                           n1817, B2 => REGISTERS_14_7_port, ZN => n2249);
   U2790 : AOI21_X1 port map( B1 => n2250, B2 => n2251, A => N352, ZN => N293);
   U2791 : NOR4_X1 port map( A1 => n2252, A2 => n2253, A3 => n2254, A4 => n2255
                           , ZN => n2251);
   U2792 : OAI221_X1 port map( B1 => n528, B2 => n1774, C1 => n562, C2 => n1775
                           , A => n2256, ZN => n2255);
   U2793 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_6_port, B1 => 
                           n1778, B2 => REGISTERS_18_6_port, ZN => n2256);
   U2794 : OAI221_X1 port map( B1 => n392, B2 => n1779, C1 => n426, C2 => n1780
                           , A => n2257, ZN => n2254);
   U2795 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_6_port, B1 => 
                           n1783, B2 => REGISTERS_22_6_port, ZN => n2257);
   U2796 : OAI221_X1 port map( B1 => n252, B2 => n1784, C1 => n287_port, C2 => 
                           n1785, A => n2258, ZN => n2253);
   U2797 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_6_port, B1 => 
                           n1788, B2 => REGISTERS_26_6_port, ZN => n2258);
   U2798 : OAI221_X1 port map( B1 => n16, B2 => n1789, C1 => n77, C2 => n1790, 
                           A => n2259, ZN => n2252);
   U2799 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_6_port, B1 => 
                           n1793, B2 => REGISTERS_28_6_port, ZN => n2259);
   U2800 : NOR4_X1 port map( A1 => n2260, A2 => n2261, A3 => n2262, A4 => n2263
                           , ZN => n2250);
   U2801 : OAI221_X1 port map( B1 => n1079, B2 => n1798, C1 => n1113, C2 => 
                           n1799, A => n2264, ZN => n2263);
   U2802 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_6_port, B1 => 
                           n1802, B2 => REGISTERS_2_6_port, ZN => n2264);
   U2803 : OAI221_X1 port map( B1 => n943, B2 => n1803, C1 => n977, C2 => n1804
                           , A => n2265, ZN => n2262);
   U2804 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_6_port, B1 => 
                           n1807, B2 => REGISTERS_6_6_port, ZN => n2265);
   U2805 : OAI221_X1 port map( B1 => n802, B2 => n1808, C1 => n836, C2 => n1809
                           , A => n2266, ZN => n2261);
   U2806 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_6_port, B1 => 
                           n1812, B2 => REGISTERS_10_6_port, ZN => n2266);
   U2807 : OAI221_X1 port map( B1 => n666, B2 => n1813, C1 => n700, C2 => n1814
                           , A => n2267, ZN => n2260);
   U2808 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_6_port, B1 => 
                           n1817, B2 => REGISTERS_14_6_port, ZN => n2267);
   U2809 : AOI21_X1 port map( B1 => n2268, B2 => n2269, A => N352, ZN => N292);
   U2810 : NOR4_X1 port map( A1 => n2270, A2 => n2271, A3 => n2272, A4 => n2273
                           , ZN => n2269);
   U2811 : OAI221_X1 port map( B1 => n527, B2 => n1774, C1 => n561, C2 => n1775
                           , A => n2274, ZN => n2273);
   U2812 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_5_port, B1 => 
                           n1778, B2 => REGISTERS_18_5_port, ZN => n2274);
   U2813 : OAI221_X1 port map( B1 => n391, B2 => n1779, C1 => n425, C2 => n1780
                           , A => n2275, ZN => n2272);
   U2814 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_5_port, B1 => 
                           n1783, B2 => REGISTERS_22_5_port, ZN => n2275);
   U2815 : OAI221_X1 port map( B1 => n251, B2 => n1784, C1 => n286_port, C2 => 
                           n1785, A => n2276, ZN => n2271);
   U2816 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_5_port, B1 => 
                           n1788, B2 => REGISTERS_26_5_port, ZN => n2276);
   U2817 : OAI221_X1 port map( B1 => n14, B2 => n1789, C1 => n76, C2 => n1790, 
                           A => n2277, ZN => n2270);
   U2818 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_5_port, B1 => 
                           n1793, B2 => REGISTERS_28_5_port, ZN => n2277);
   U2819 : NOR4_X1 port map( A1 => n2278, A2 => n2279, A3 => n2280, A4 => n2281
                           , ZN => n2268);
   U2820 : OAI221_X1 port map( B1 => n1078, B2 => n1798, C1 => n1112, C2 => 
                           n1799, A => n2282, ZN => n2281);
   U2821 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_5_port, B1 => 
                           n1802, B2 => REGISTERS_2_5_port, ZN => n2282);
   U2822 : OAI221_X1 port map( B1 => n942, B2 => n1803, C1 => n976, C2 => n1804
                           , A => n2283, ZN => n2280);
   U2823 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_5_port, B1 => 
                           n1807, B2 => REGISTERS_6_5_port, ZN => n2283);
   U2824 : OAI221_X1 port map( B1 => n801, B2 => n1808, C1 => n835, C2 => n1809
                           , A => n2284, ZN => n2279);
   U2825 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_5_port, B1 => 
                           n1812, B2 => REGISTERS_10_5_port, ZN => n2284);
   U2826 : OAI221_X1 port map( B1 => n665, B2 => n1813, C1 => n699, C2 => n1814
                           , A => n2285, ZN => n2278);
   U2827 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_5_port, B1 => 
                           n1817, B2 => REGISTERS_14_5_port, ZN => n2285);
   U2828 : AOI21_X1 port map( B1 => n2286, B2 => n2287, A => N352, ZN => N291);
   U2829 : NOR4_X1 port map( A1 => n2288, A2 => n2289, A3 => n2290, A4 => n2291
                           , ZN => n2287);
   U2830 : OAI221_X1 port map( B1 => n526, B2 => n1774, C1 => n560, C2 => n1775
                           , A => n2292, ZN => n2291);
   U2831 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_4_port, B1 => 
                           n1778, B2 => REGISTERS_18_4_port, ZN => n2292);
   U2832 : OAI221_X1 port map( B1 => n390, B2 => n1779, C1 => n424, C2 => n1780
                           , A => n2293, ZN => n2290);
   U2833 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_4_port, B1 => 
                           n1783, B2 => REGISTERS_22_4_port, ZN => n2293);
   U2834 : OAI221_X1 port map( B1 => n250, B2 => n1784, C1 => n285, C2 => n1785
                           , A => n2294, ZN => n2289);
   U2835 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_4_port, B1 => 
                           n1788, B2 => REGISTERS_26_4_port, ZN => n2294);
   U2836 : OAI221_X1 port map( B1 => n12, B2 => n1789, C1 => n75, C2 => n1790, 
                           A => n2295, ZN => n2288);
   U2837 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_4_port, B1 => 
                           n1793, B2 => REGISTERS_28_4_port, ZN => n2295);
   U2838 : NOR4_X1 port map( A1 => n2296, A2 => n2297, A3 => n2298, A4 => n2299
                           , ZN => n2286);
   U2839 : OAI221_X1 port map( B1 => n1077, B2 => n1798, C1 => n1111, C2 => 
                           n1799, A => n2300, ZN => n2299);
   U2840 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_4_port, B1 => 
                           n1802, B2 => REGISTERS_2_4_port, ZN => n2300);
   U2841 : OAI221_X1 port map( B1 => n941, B2 => n1803, C1 => n975, C2 => n1804
                           , A => n2301, ZN => n2298);
   U2842 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_4_port, B1 => 
                           n1807, B2 => REGISTERS_6_4_port, ZN => n2301);
   U2843 : OAI221_X1 port map( B1 => n800, B2 => n1808, C1 => n834, C2 => n1809
                           , A => n2302, ZN => n2297);
   U2844 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_4_port, B1 => 
                           n1812, B2 => REGISTERS_10_4_port, ZN => n2302);
   U2845 : OAI221_X1 port map( B1 => n664, B2 => n1813, C1 => n698, C2 => n1814
                           , A => n2303, ZN => n2296);
   U2846 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_4_port, B1 => 
                           n1817, B2 => REGISTERS_14_4_port, ZN => n2303);
   U2847 : AOI21_X1 port map( B1 => n2304, B2 => n2305, A => N352, ZN => N290);
   U2848 : NOR4_X1 port map( A1 => n2306, A2 => n2307, A3 => n2308, A4 => n2309
                           , ZN => n2305);
   U2849 : OAI221_X1 port map( B1 => n525, B2 => n1774, C1 => n559, C2 => n1775
                           , A => n2310, ZN => n2309);
   U2850 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_3_port, B1 => 
                           n1778, B2 => REGISTERS_18_3_port, ZN => n2310);
   U2851 : OAI221_X1 port map( B1 => n389, B2 => n1779, C1 => n423, C2 => n1780
                           , A => n2311, ZN => n2308);
   U2852 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_3_port, B1 => 
                           n1783, B2 => REGISTERS_22_3_port, ZN => n2311);
   U2853 : OAI221_X1 port map( B1 => n249, B2 => n1784, C1 => n284, C2 => n1785
                           , A => n2312, ZN => n2307);
   U2854 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_3_port, B1 => 
                           n1788, B2 => REGISTERS_26_3_port, ZN => n2312);
   U2855 : OAI221_X1 port map( B1 => n10, B2 => n1789, C1 => n74, C2 => n1790, 
                           A => n2313, ZN => n2306);
   U2856 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_3_port, B1 => 
                           n1793, B2 => REGISTERS_28_3_port, ZN => n2313);
   U2857 : NOR4_X1 port map( A1 => n2314, A2 => n2315, A3 => n2316, A4 => n2317
                           , ZN => n2304);
   U2858 : OAI221_X1 port map( B1 => n1076, B2 => n1798, C1 => n1110, C2 => 
                           n1799, A => n2318, ZN => n2317);
   U2859 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_3_port, B1 => 
                           n1802, B2 => REGISTERS_2_3_port, ZN => n2318);
   U2860 : OAI221_X1 port map( B1 => n940, B2 => n1803, C1 => n974, C2 => n1804
                           , A => n2319, ZN => n2316);
   U2861 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_3_port, B1 => 
                           n1807, B2 => REGISTERS_6_3_port, ZN => n2319);
   U2862 : OAI221_X1 port map( B1 => n799, B2 => n1808, C1 => n833, C2 => n1809
                           , A => n2320, ZN => n2315);
   U2863 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_3_port, B1 => 
                           n1812, B2 => REGISTERS_10_3_port, ZN => n2320);
   U2864 : OAI221_X1 port map( B1 => n663, B2 => n1813, C1 => n697, C2 => n1814
                           , A => n2321, ZN => n2314);
   U2865 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_3_port, B1 => 
                           n1817, B2 => REGISTERS_14_3_port, ZN => n2321);
   U2866 : AOI21_X1 port map( B1 => n2322, B2 => n2323, A => N352, ZN => N289);
   U2867 : NOR4_X1 port map( A1 => n2324, A2 => n2325, A3 => n2326, A4 => n2327
                           , ZN => n2323);
   U2868 : OAI221_X1 port map( B1 => n524, B2 => n1774, C1 => n558, C2 => n1775
                           , A => n2328, ZN => n2327);
   U2869 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_2_port, B1 => 
                           n1778, B2 => REGISTERS_18_2_port, ZN => n2328);
   U2870 : OAI221_X1 port map( B1 => n388, B2 => n1779, C1 => n422, C2 => n1780
                           , A => n2329, ZN => n2326);
   U2871 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_2_port, B1 => 
                           n1783, B2 => REGISTERS_22_2_port, ZN => n2329);
   U2872 : OAI221_X1 port map( B1 => n248, B2 => n1784, C1 => n283, C2 => n1785
                           , A => n2330, ZN => n2325);
   U2873 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_2_port, B1 => 
                           n1788, B2 => REGISTERS_26_2_port, ZN => n2330);
   U2874 : OAI221_X1 port map( B1 => n8, B2 => n1789, C1 => n73, C2 => n1790, A
                           => n2331, ZN => n2324);
   U2875 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_2_port, B1 => 
                           n1793, B2 => REGISTERS_28_2_port, ZN => n2331);
   U2876 : NOR4_X1 port map( A1 => n2332, A2 => n2333, A3 => n2334, A4 => n2335
                           , ZN => n2322);
   U2877 : OAI221_X1 port map( B1 => n1075, B2 => n1798, C1 => n1109, C2 => 
                           n1799, A => n2336, ZN => n2335);
   U2878 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_2_port, B1 => 
                           n1802, B2 => REGISTERS_2_2_port, ZN => n2336);
   U2879 : OAI221_X1 port map( B1 => n939, B2 => n1803, C1 => n973, C2 => n1804
                           , A => n2337, ZN => n2334);
   U2880 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_2_port, B1 => 
                           n1807, B2 => REGISTERS_6_2_port, ZN => n2337);
   U2881 : OAI221_X1 port map( B1 => n798, B2 => n1808, C1 => n832, C2 => n1809
                           , A => n2338, ZN => n2333);
   U2882 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_2_port, B1 => 
                           n1812, B2 => REGISTERS_10_2_port, ZN => n2338);
   U2883 : OAI221_X1 port map( B1 => n662, B2 => n1813, C1 => n696, C2 => n1814
                           , A => n2339, ZN => n2332);
   U2884 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_2_port, B1 => 
                           n1817, B2 => REGISTERS_14_2_port, ZN => n2339);
   U2885 : AOI21_X1 port map( B1 => n2340, B2 => n2341, A => N352, ZN => N288);
   U2886 : NOR4_X1 port map( A1 => n2342, A2 => n2343, A3 => n2344, A4 => n2345
                           , ZN => n2341);
   U2887 : OAI221_X1 port map( B1 => n523, B2 => n1774, C1 => n557, C2 => n1775
                           , A => n2346, ZN => n2345);
   U2888 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_1_port, B1 => 
                           n1778, B2 => REGISTERS_18_1_port, ZN => n2346);
   U2889 : OAI221_X1 port map( B1 => n387, B2 => n1779, C1 => n421, C2 => n1780
                           , A => n2347, ZN => n2344);
   U2890 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_1_port, B1 => 
                           n1783, B2 => REGISTERS_22_1_port, ZN => n2347);
   U2891 : OAI221_X1 port map( B1 => n247, B2 => n1784, C1 => n282, C2 => n1785
                           , A => n2348, ZN => n2343);
   U2892 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_1_port, B1 => 
                           n1788, B2 => REGISTERS_26_1_port, ZN => n2348);
   U2893 : OAI221_X1 port map( B1 => n6, B2 => n1789, C1 => n72, C2 => n1790, A
                           => n2349, ZN => n2342);
   U2894 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_1_port, B1 => 
                           n1793, B2 => REGISTERS_28_1_port, ZN => n2349);
   U2895 : NOR4_X1 port map( A1 => n2350, A2 => n2351, A3 => n2352, A4 => n2353
                           , ZN => n2340);
   U2896 : OAI221_X1 port map( B1 => n1074, B2 => n1798, C1 => n1108, C2 => 
                           n1799, A => n2354, ZN => n2353);
   U2897 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_1_port, B1 => 
                           n1802, B2 => REGISTERS_2_1_port, ZN => n2354);
   U2898 : OAI221_X1 port map( B1 => n938, B2 => n1803, C1 => n972, C2 => n1804
                           , A => n2355, ZN => n2352);
   U2899 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_1_port, B1 => 
                           n1807, B2 => REGISTERS_6_1_port, ZN => n2355);
   U2900 : OAI221_X1 port map( B1 => n797, B2 => n1808, C1 => n831, C2 => n1809
                           , A => n2356, ZN => n2351);
   U2901 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_1_port, B1 => 
                           n1812, B2 => REGISTERS_10_1_port, ZN => n2356);
   U2902 : OAI221_X1 port map( B1 => n661, B2 => n1813, C1 => n695, C2 => n1814
                           , A => n2357, ZN => n2350);
   U2903 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_1_port, B1 => 
                           n1817, B2 => REGISTERS_14_1_port, ZN => n2357);
   U2904 : AOI21_X1 port map( B1 => n2358, B2 => n2359, A => N352, ZN => N287);
   U2906 : NOR4_X1 port map( A1 => n2360, A2 => n2361, A3 => n2362, A4 => n2363
                           , ZN => n2359);
   U2907 : OAI221_X1 port map( B1 => n522, B2 => n1774, C1 => n556, C2 => n1775
                           , A => n2364, ZN => n2363);
   U2908 : AOI22_X1 port map( A1 => n1777, A2 => REGISTERS_19_0_port, B1 => 
                           n1778, B2 => REGISTERS_18_0_port, ZN => n2364);
   U2913 : OAI221_X1 port map( B1 => n386, B2 => n1779, C1 => n420, C2 => n1780
                           , A => n2369, ZN => n2362);
   U2914 : AOI22_X1 port map( A1 => n1782, A2 => REGISTERS_23_0_port, B1 => 
                           n1783, B2 => REGISTERS_22_0_port, ZN => n2369);
   U2918 : AND2_X1 port map( A1 => n2372, A2 => n2373, ZN => n2365);
   U2920 : AND2_X1 port map( A1 => n2372, A2 => ADD_RD1(0), ZN => n2367);
   U2921 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => n2374, ZN => n2372);
   U2922 : OAI221_X1 port map( B1 => n246, B2 => n1784, C1 => n281, C2 => n1785
                           , A => n2375, ZN => n2361);
   U2923 : AOI22_X1 port map( A1 => n1787, A2 => REGISTERS_27_0_port, B1 => 
                           n1788, B2 => REGISTERS_26_0_port, ZN => n2375);
   U2928 : OAI221_X1 port map( B1 => n4, B2 => n1789, C1 => n71, C2 => n1790, A
                           => n2378, ZN => n2360);
   U2929 : AOI22_X1 port map( A1 => n1792, A2 => REGISTERS_29_0_port, B1 => 
                           n1793, B2 => REGISTERS_28_0_port, ZN => n2378);
   U2933 : AND2_X1 port map( A1 => n2379, A2 => n2373, ZN => n2376);
   U2935 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n2379, ZN => n2377);
   U2936 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n2379);
   U2937 : NOR4_X1 port map( A1 => n2380, A2 => n2381, A3 => n2382, A4 => n2383
                           , ZN => n2358);
   U2938 : OAI221_X1 port map( B1 => n1073, B2 => n1798, C1 => n1107, C2 => 
                           n1799, A => n2384, ZN => n2383);
   U2939 : AOI22_X1 port map( A1 => n1801, A2 => REGISTERS_3_0_port, B1 => 
                           n1802, B2 => REGISTERS_2_0_port, ZN => n2384);
   U2944 : OAI221_X1 port map( B1 => n937, B2 => n1803, C1 => n971, C2 => n1804
                           , A => n2387, ZN => n2382);
   U2945 : AOI22_X1 port map( A1 => n1806, A2 => REGISTERS_7_0_port, B1 => 
                           n1807, B2 => REGISTERS_6_0_port, ZN => n2387);
   U2949 : AND2_X1 port map( A1 => n2388, A2 => n2373, ZN => n2385);
   U2951 : AND2_X1 port map( A1 => n2388, A2 => ADD_RD1(0), ZN => n2386);
   U2952 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n2388);
   U2953 : OAI221_X1 port map( B1 => n796, B2 => n1808, C1 => n830, C2 => n1809
                           , A => n2389, ZN => n2381);
   U2954 : AOI22_X1 port map( A1 => n1811, A2 => REGISTERS_11_0_port, B1 => 
                           n1812, B2 => REGISTERS_10_0_port, ZN => n2389);
   U2957 : NOR2_X1 port map( A1 => n2392, A2 => ADD_RD1(2), ZN => n2366);
   U2961 : OAI221_X1 port map( B1 => n660, B2 => n1813, C1 => n694, C2 => n1814
                           , A => n2393, ZN => n2380);
   U2962 : AOI22_X1 port map( A1 => n1816, A2 => REGISTERS_15_0_port, B1 => 
                           n1817, B2 => REGISTERS_14_0_port, ZN => n2393);
   U2965 : NOR2_X1 port map( A1 => n2394, A2 => n2392, ZN => n2370);
   U2966 : INV_X1 port map( A => ADD_RD1(1), ZN => n2392);
   U2968 : AND2_X1 port map( A1 => n2395, A2 => n2373, ZN => n2390);
   U2969 : INV_X1 port map( A => ADD_RD1(0), ZN => n2373);
   U2972 : INV_X1 port map( A => ADD_RD1(2), ZN => n2394);
   U2973 : AND2_X1 port map( A1 => n2395, A2 => ADD_RD1(0), ZN => n2391);
   U2974 : NOR2_X1 port map( A1 => n2374, A2 => ADD_RD1(4), ZN => n2395);
   U2975 : INV_X1 port map( A => ADD_RD1(3), ZN => n2374);
   U2976 : NAND2_X1 port map( A1 => n2396, A2 => RESET, ZN => N286);
   U2977 : NAND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n2396);
   U35 : AND2_X2 port map( A1 => n2390, A2 => n2370, ZN => n1817);
   U36 : AND2_X2 port map( A1 => n2390, A2 => n2366, ZN => n1812);
   U69 : AND2_X2 port map( A1 => n2385, A2 => n2370, ZN => n1807);
   U70 : AND2_X2 port map( A1 => n2385, A2 => n2366, ZN => n1802);
   U135 : AND2_X2 port map( A1 => n2371, A2 => n2376, ZN => n1793);
   U136 : AND2_X2 port map( A1 => n2366, A2 => n2376, ZN => n1788);
   U201 : AND2_X2 port map( A1 => n2365, A2 => n2370, ZN => n1783);
   U202 : AND2_X2 port map( A1 => n2365, A2 => n2366, ZN => n1778);
   U267 : AND2_X2 port map( A1 => n1761, A2 => n1741, ZN => n1188);
   U268 : AND2_X2 port map( A1 => n1761, A2 => n1737, ZN => n1183);
   U333 : AND2_X2 port map( A1 => n1756, A2 => n1741, ZN => n1178);
   U334 : AND2_X2 port map( A1 => n1756, A2 => n1737, ZN => n1173);
   U367 : AND2_X2 port map( A1 => n1742, A2 => n1747, ZN => n1164);
   U368 : AND2_X2 port map( A1 => n1737, A2 => n1747, ZN => n1159);
   U401 : AND2_X2 port map( A1 => n1736, A2 => n1741, ZN => n1154);
   U402 : AND2_X2 port map( A1 => n1736, A2 => n1737, ZN => n1149);
   U468 : NAND2_X2 port map( A1 => n2385, A2 => n2368, ZN => n1799);
   U469 : NAND2_X2 port map( A1 => n2376, A2 => n2370, ZN => n1790);
   U534 : NAND2_X2 port map( A1 => n2368, A2 => n2376, ZN => n1785);
   U535 : NAND2_X2 port map( A1 => n2365, A2 => n2371, ZN => n1780);
   U568 : NOR2_X2 port map( A1 => n2394, A2 => ADD_RD1(1), ZN => n2371);
   U569 : NAND2_X2 port map( A1 => n2365, A2 => n2368, ZN => n1775);
   U602 : NOR2_X2 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n2368);
   U603 : NAND2_X2 port map( A1 => n1761, A2 => n1742, ZN => n1185);
   U668 : NOR2_X2 port map( A1 => n1765, A2 => ADD_RD2(1), ZN => n1742);
   U669 : NAND2_X2 port map( A1 => n1761, A2 => n1739, ZN => n1180);
   U734 : NAND2_X2 port map( A1 => n1756, A2 => n1742, ZN => n1175);
   U735 : NAND2_X2 port map( A1 => n1756, A2 => n1739, ZN => n1170);
   U768 : NAND2_X2 port map( A1 => n1747, A2 => n1741, ZN => n1161);
   U769 : NAND2_X2 port map( A1 => n1739, A2 => n1747, ZN => n1156);
   U802 : NOR2_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1739);
   U803 : NAND2_X2 port map( A1 => n1736, A2 => n1742, ZN => n1151);
   U869 : NAND2_X2 port map( A1 => n1736, A2 => n1739, ZN => n1146);
   U870 : NAND2_X2 port map( A1 => n2390, A2 => n2368, ZN => n1809);
   U935 : NAND2_X2 port map( A1 => n2385, A2 => n2371, ZN => n1804);
   U936 : NAND2_X2 port map( A1 => n2390, A2 => n2371, ZN => n1814);
   U969 : NAND2_X2 port map( A1 => n1738, A2 => n1739, ZN => n1145);
   U970 : NAND2_X2 port map( A1 => n1739, A2 => n1748, ZN => n1155);
   U1003 : NAND2_X2 port map( A1 => n1738, A2 => n1742, ZN => n1150);
   U1004 : NAND2_X2 port map( A1 => n1757, A2 => n1739, ZN => n1169);
   U1069 : NAND2_X2 port map( A1 => n1741, A2 => n1748, ZN => n1160);
   U1070 : NAND2_X2 port map( A1 => n1762, A2 => n1739, ZN => n1179);
   U1135 : NAND2_X2 port map( A1 => n1757, A2 => n1742, ZN => n1174);
   U1136 : NAND2_X2 port map( A1 => n2367, A2 => n2368, ZN => n1774);
   U1169 : NAND2_X2 port map( A1 => n1762, A2 => n1742, ZN => n1184);
   U1170 : NAND2_X2 port map( A1 => n2368, A2 => n2377, ZN => n1784);
   U1203 : NAND2_X2 port map( A1 => n2367, A2 => n2371, ZN => n1779);
   U1204 : NAND2_X2 port map( A1 => n2386, A2 => n2368, ZN => n1798);
   U1270 : NAND2_X2 port map( A1 => n2370, A2 => n2377, ZN => n1789);
   U1271 : NAND2_X2 port map( A1 => n2391, A2 => n2368, ZN => n1808);
   U1337 : NAND2_X2 port map( A1 => n2386, A2 => n2371, ZN => n1803);
   U1338 : NAND2_X2 port map( A1 => n2391, A2 => n2371, ZN => n1813);
   U1372 : AND2_X2 port map( A1 => n1738, A2 => n1741, ZN => n1153);
   U1373 : AND2_X2 port map( A1 => n1738, A2 => n1737, ZN => n1148);
   U1407 : AND2_X2 port map( A1 => n1742, A2 => n1748, ZN => n1163);
   U1408 : AND2_X2 port map( A1 => n1737, A2 => n1748, ZN => n1158);
   U1475 : AND2_X2 port map( A1 => n1757, A2 => n1741, ZN => n1177);
   U1476 : AND2_X2 port map( A1 => n1757, A2 => n1737, ZN => n1172);
   U1542 : AND2_X2 port map( A1 => n1762, A2 => n1741, ZN => n1187);
   U1543 : AND2_X2 port map( A1 => n1762, A2 => n1737, ZN => n1182);
   U1578 : AND2_X2 port map( A1 => n2367, A2 => n2370, ZN => n1782);
   U1579 : AND2_X2 port map( A1 => n2367, A2 => n2366, ZN => n1777);
   U1645 : AND2_X2 port map( A1 => n2371, A2 => n2377, ZN => n1792);
   U1646 : AND2_X2 port map( A1 => n2366, A2 => n2377, ZN => n1787);
   U2246 : AND2_X2 port map( A1 => n2386, A2 => n2370, ZN => n1806);
   U2247 : AND2_X2 port map( A1 => n2386, A2 => n2366, ZN => n1801);
   U2248 : AND2_X2 port map( A1 => n2391, A2 => n2370, ZN => n1816);
   U2249 : AND2_X2 port map( A1 => n2391, A2 => n2366, ZN => n1811);
   U2252 : INV_X2 port map( A => n106, ZN => n105);
   U2253 : NAND2_X2 port map( A1 => n138, A2 => n68, ZN => n106);
   U2254 : INV_X2 port map( A => n176, ZN => n175);
   U2256 : NAND2_X2 port map( A1 => n208, A2 => n68, ZN => n176);
   U2261 : INV_X2 port map( A => n141, ZN => n140);
   U2262 : NAND2_X2 port map( A1 => n173, A2 => n68, ZN => n141);
   U2263 : INV_X2 port map( A => n317_port, ZN => n316_port);
   U2264 : NAND2_X2 port map( A1 => n349_port, A2 => n67, ZN => n317_port);
   U2267 : INV_X2 port map( A => n211, ZN => n210);
   U2268 : NAND2_X2 port map( A1 => n243, A2 => n68, ZN => n211);
   U2269 : INV_X2 port map( A => n454, ZN => n453);
   U2271 : NAND2_X2 port map( A1 => n349_port, A2 => n208, ZN => n454);
   U2277 : INV_X2 port map( A => n352_port, ZN => n351_port);
   U2278 : NAND2_X2 port map( A1 => n349_port, A2 => n103, ZN => n352_port);
   U2279 : INV_X2 port map( A => n591, ZN => n590);
   U2280 : NAND2_X2 port map( A1 => n623, A2 => n67, ZN => n591);
   U2283 : INV_X2 port map( A => n488, ZN => n487);
   U2284 : NAND2_X2 port map( A1 => n349_port, A2 => n243, ZN => n488);
   U2285 : INV_X2 port map( A => n728, ZN => n727);
   U2287 : NAND2_X2 port map( A1 => n623, A2 => n208, ZN => n728);
   U2292 : INV_X2 port map( A => n626, ZN => n625);
   U2293 : NAND2_X2 port map( A1 => n623, A2 => n103, ZN => n626);
   U2295 : INV_X2 port map( A => n865, ZN => n864);
   U2296 : NAND2_X2 port map( A1 => n897, A2 => n67, ZN => n865);
   U2297 : INV_X2 port map( A => n762, ZN => n761);
   U2300 : NAND2_X2 port map( A1 => n623, A2 => n243, ZN => n762);
   U2301 : INV_X2 port map( A => n1005, ZN => n1004);
   U2304 : NAND2_X2 port map( A1 => n897, A2 => n208, ZN => n1005);
   U2307 : INV_X2 port map( A => n903, ZN => n902);
   U2308 : NAND2_X2 port map( A1 => n897, A2 => n103, ZN => n903);
   U2905 : INV_X2 port map( A => n69, ZN => n70);
   U2909 : NAND2_X2 port map( A1 => n103, A2 => n68, ZN => n69);
   U2910 : INV_X2 port map( A => n1039, ZN => n1038);
   U2911 : NAND2_X2 port map( A1 => n897, A2 => n243, ZN => n1039);
   U2912 : INV_X2 port map( A => n279, ZN => n280);
   U2915 : NAND2_X2 port map( A1 => n313_port, A2 => n68, ZN => n279);
   U2916 : INV_X2 port map( A => n244, ZN => n245);
   U2917 : NAND2_X2 port map( A1 => n278, A2 => n68, ZN => n244);
   U2919 : INV_X2 port map( A => n418, ZN => n419);
   U2924 : NAND2_X2 port map( A1 => n349_port, A2 => n173, ZN => n418);
   U2925 : INV_X2 port map( A => n384, ZN => n385);
   U2926 : NAND2_X2 port map( A1 => n349_port, A2 => n138, ZN => n384);
   U2927 : INV_X2 port map( A => n554, ZN => n555);
   U2930 : NAND2_X2 port map( A1 => n349_port, A2 => n313_port, ZN => n554);
   U2931 : INV_X2 port map( A => n520, ZN => n521);
   U2932 : NAND2_X2 port map( A1 => n349_port, A2 => n278, ZN => n520);
   U2934 : INV_X2 port map( A => n692, ZN => n693);
   U2940 : NAND2_X2 port map( A1 => n623, A2 => n173, ZN => n692);
   U2941 : INV_X2 port map( A => n658, ZN => n659);
   U2942 : NAND2_X2 port map( A1 => n623, A2 => n138, ZN => n658);
   U2943 : INV_X2 port map( A => n828, ZN => n829);
   U2946 : NAND2_X2 port map( A1 => n623, A2 => n313_port, ZN => n828);
   U2947 : INV_X2 port map( A => n794, ZN => n795);
   U2948 : NAND2_X2 port map( A1 => n623, A2 => n278, ZN => n794);
   U2950 : INV_X2 port map( A => n969, ZN => n970);
   U2955 : NAND2_X2 port map( A1 => n897, A2 => n173, ZN => n969);
   U2956 : INV_X2 port map( A => n935, ZN => n936);
   U2958 : NAND2_X2 port map( A1 => n897, A2 => n138, ZN => n935);
   U2959 : INV_X2 port map( A => n1105, ZN => n1106);
   U2960 : NAND2_X2 port map( A1 => n897, A2 => n313_port, ZN => n1105);
   U2963 : INV_X2 port map( A => n1071, ZN => n1072);
   U2964 : NAND2_X2 port map( A1 => n897, A2 => n278, ZN => n1071);
   U2967 : INV_X2 port map( A => n1, ZN => n3);
   U2970 : NAND2_X2 port map( A1 => n67, A2 => n68, ZN => n1);
   U2971 : INV_X4 port map( A => RESET, ZN => N352);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IR_DECODE_NBIT32_opBIT6_regBIT5 is

   port( CLK : in std_logic;  IR_26 : in std_logic_vector (25 downto 0);  
         OPCODE : in std_logic_vector (5 downto 0);  is_signed : in std_logic; 
         RS1, RS2, RD : out std_logic_vector (4 downto 0);  IMMEDIATE : out 
         std_logic_vector (31 downto 0));

end IR_DECODE_NBIT32_opBIT6_regBIT5;

architecture SYN_BEHAV of IR_DECODE_NBIT32_opBIT6_regBIT5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component sign_eval_N_in26_N_out32
      port( IR_out : in std_logic_vector (25 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_eval_N_in16_N_out32
      port( IR_out : in std_logic_vector (15 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_eval_N_in5_N_out32
      port( IR_out : in std_logic_vector (4 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic0_port, IMMEDIATE_16_31_port, IMMEDIATE_16_15_port, 
      IMMEDIATE_16_14_port, IMMEDIATE_16_13_port, IMMEDIATE_16_12_port, 
      IMMEDIATE_16_11_port, IMMEDIATE_16_10_port, IMMEDIATE_16_9_port, 
      IMMEDIATE_16_8_port, IMMEDIATE_16_7_port, IMMEDIATE_16_6_port, 
      IMMEDIATE_16_5_port, IMMEDIATE_16_4_port, IMMEDIATE_16_3_port, 
      IMMEDIATE_16_2_port, IMMEDIATE_16_1_port, IMMEDIATE_16_0_port, N143, N144
      , N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
      N157, N158, N159, N160, N161, N162, N163, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173,
      n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, 
      n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, 
      n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, 
      n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, 
      n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, 
      n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, 
      n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, 
      n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243 : std_logic;

begin
   
   X_Logic0_port <= '0';
   RD_reg_4_inst : DLH_X1 port map( G => CLK, D => N147, Q => RD(4));
   RD_reg_3_inst : DLH_X1 port map( G => CLK, D => N146, Q => RD(3));
   RD_reg_2_inst : DLH_X1 port map( G => CLK, D => N145, Q => RD(2));
   RD_reg_1_inst : DLH_X1 port map( G => CLK, D => N144, Q => RD(1));
   RD_reg_0_inst : DLH_X1 port map( G => CLK, D => N143, Q => RD(0));
   IMMEDIATE_reg_31_inst : DLH_X1 port map( G => CLK, D => n36, Q => 
                           IMMEDIATE(31));
   IMMEDIATE_reg_30_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(30));
   IMMEDIATE_reg_29_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(29));
   IMMEDIATE_reg_28_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(28));
   IMMEDIATE_reg_27_inst : DLH_X1 port map( G => CLK, D => n36, Q => 
                           IMMEDIATE(27));
   IMMEDIATE_reg_26_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(26));
   IMMEDIATE_reg_25_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(25));
   IMMEDIATE_reg_24_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(24));
   IMMEDIATE_reg_23_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(23));
   IMMEDIATE_reg_22_inst : DLH_X1 port map( G => CLK, D => n36, Q => 
                           IMMEDIATE(22));
   IMMEDIATE_reg_21_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(21));
   IMMEDIATE_reg_20_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(20));
   IMMEDIATE_reg_19_inst : DLH_X1 port map( G => CLK, D => n36, Q => 
                           IMMEDIATE(19));
   IMMEDIATE_reg_18_inst : DLH_X1 port map( G => CLK, D => n36, Q => 
                           IMMEDIATE(18));
   IMMEDIATE_reg_17_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(17));
   IMMEDIATE_reg_16_inst : DLH_X1 port map( G => CLK, D => n32, Q => 
                           IMMEDIATE(16));
   IMMEDIATE_reg_15_inst : DLH_X1 port map( G => CLK, D => N163, Q => 
                           IMMEDIATE(15));
   IMMEDIATE_reg_14_inst : DLH_X1 port map( G => CLK, D => N162, Q => 
                           IMMEDIATE(14));
   IMMEDIATE_reg_13_inst : DLH_X1 port map( G => CLK, D => N161, Q => 
                           IMMEDIATE(13));
   IMMEDIATE_reg_12_inst : DLH_X1 port map( G => CLK, D => N160, Q => 
                           IMMEDIATE(12));
   IMMEDIATE_reg_11_inst : DLH_X1 port map( G => CLK, D => N159, Q => 
                           IMMEDIATE(11));
   IMMEDIATE_reg_10_inst : DLH_X1 port map( G => CLK, D => N158, Q => 
                           IMMEDIATE(10));
   IMMEDIATE_reg_9_inst : DLH_X1 port map( G => CLK, D => N157, Q => 
                           IMMEDIATE(9));
   IMMEDIATE_reg_8_inst : DLH_X1 port map( G => CLK, D => N156, Q => 
                           IMMEDIATE(8));
   IMMEDIATE_reg_7_inst : DLH_X1 port map( G => CLK, D => N155, Q => 
                           IMMEDIATE(7));
   IMMEDIATE_reg_6_inst : DLH_X1 port map( G => CLK, D => N154, Q => 
                           IMMEDIATE(6));
   IMMEDIATE_reg_5_inst : DLH_X1 port map( G => CLK, D => N153, Q => 
                           IMMEDIATE(5));
   IMMEDIATE_reg_4_inst : DLH_X1 port map( G => CLK, D => N152, Q => 
                           IMMEDIATE(4));
   IMMEDIATE_reg_3_inst : DLH_X1 port map( G => CLK, D => N151, Q => 
                           IMMEDIATE(3));
   IMMEDIATE_reg_2_inst : DLH_X1 port map( G => CLK, D => N150, Q => 
                           IMMEDIATE(2));
   IMMEDIATE_reg_1_inst : DLH_X1 port map( G => CLK, D => N149, Q => 
                           IMMEDIATE(1));
   IMMEDIATE_reg_0_inst : DLH_X1 port map( G => CLK, D => N148, Q => 
                           IMMEDIATE(0));
   RS1_reg_4_inst : DLH_X1 port map( G => CLK, D => IR_26(25), Q => RS1(4));
   RS1_reg_3_inst : DLH_X1 port map( G => CLK, D => IR_26(24), Q => RS1(3));
   RS1_reg_2_inst : DLH_X1 port map( G => CLK, D => IR_26(23), Q => RS1(2));
   RS1_reg_1_inst : DLH_X1 port map( G => CLK, D => IR_26(22), Q => RS1(1));
   RS1_reg_0_inst : DLH_X1 port map( G => CLK, D => IR_26(21), Q => RS1(0));
   RS2_reg_4_inst : DLH_X1 port map( G => CLK, D => IR_26(20), Q => RS2(4));
   RS2_reg_3_inst : DLH_X1 port map( G => CLK, D => IR_26(19), Q => RS2(3));
   RS2_reg_2_inst : DLH_X1 port map( G => CLK, D => IR_26(18), Q => RS2(2));
   RS2_reg_1_inst : DLH_X1 port map( G => CLK, D => IR_26(17), Q => RS2(1));
   RS2_reg_0_inst : DLH_X1 port map( G => CLK, D => IR_26(16), Q => RS2(0));
   SIGN_EXTENSION_imm5 : sign_eval_N_in5_N_out32 port map( IR_out(4) => 
                           IR_26(15), IR_out(3) => IR_26(14), IR_out(2) => 
                           IR_26(13), IR_out(1) => IR_26(12), IR_out(0) => 
                           IR_26(11), signed_val => is_signed, Immediate(31) =>
                           n_2165, Immediate(30) => n_2166, Immediate(29) => 
                           n_2167, Immediate(28) => n_2168, Immediate(27) => 
                           n_2169, Immediate(26) => n_2170, Immediate(25) => 
                           n_2171, Immediate(24) => n_2172, Immediate(23) => 
                           n_2173, Immediate(22) => n_2174, Immediate(21) => 
                           n_2175, Immediate(20) => n_2176, Immediate(19) => 
                           n_2177, Immediate(18) => n_2178, Immediate(17) => 
                           n_2179, Immediate(16) => n_2180, Immediate(15) => 
                           n_2181, Immediate(14) => n_2182, Immediate(13) => 
                           n_2183, Immediate(12) => n_2184, Immediate(11) => 
                           n_2185, Immediate(10) => n_2186, Immediate(9) => 
                           n_2187, Immediate(8) => n_2188, Immediate(7) => 
                           n_2189, Immediate(6) => n_2190, Immediate(5) => 
                           n_2191, Immediate(4) => n_2192, Immediate(3) => 
                           n_2193, Immediate(2) => n_2194, Immediate(1) => 
                           n_2195, Immediate(0) => n_2196);
   SIGN_EXTENSION_imm16 : sign_eval_N_in16_N_out32 port map( IR_out(15) => 
                           IR_26(15), IR_out(14) => IR_26(14), IR_out(13) => 
                           IR_26(13), IR_out(12) => IR_26(12), IR_out(11) => 
                           IR_26(11), IR_out(10) => IR_26(10), IR_out(9) => 
                           IR_26(9), IR_out(8) => IR_26(8), IR_out(7) => 
                           IR_26(7), IR_out(6) => IR_26(6), IR_out(5) => 
                           IR_26(5), IR_out(4) => IR_26(4), IR_out(3) => 
                           IR_26(3), IR_out(2) => IR_26(2), IR_out(1) => 
                           IR_26(1), IR_out(0) => IR_26(0), signed_val => 
                           is_signed, Immediate(31) => IMMEDIATE_16_31_port, 
                           Immediate(30) => n_2197, Immediate(29) => n_2198, 
                           Immediate(28) => n_2199, Immediate(27) => n_2200, 
                           Immediate(26) => n_2201, Immediate(25) => n_2202, 
                           Immediate(24) => n_2203, Immediate(23) => n_2204, 
                           Immediate(22) => n_2205, Immediate(21) => n_2206, 
                           Immediate(20) => n_2207, Immediate(19) => n_2208, 
                           Immediate(18) => n_2209, Immediate(17) => n_2210, 
                           Immediate(16) => n_2211, Immediate(15) => 
                           IMMEDIATE_16_15_port, Immediate(14) => 
                           IMMEDIATE_16_14_port, Immediate(13) => 
                           IMMEDIATE_16_13_port, Immediate(12) => 
                           IMMEDIATE_16_12_port, Immediate(11) => 
                           IMMEDIATE_16_11_port, Immediate(10) => 
                           IMMEDIATE_16_10_port, Immediate(9) => 
                           IMMEDIATE_16_9_port, Immediate(8) => 
                           IMMEDIATE_16_8_port, Immediate(7) => 
                           IMMEDIATE_16_7_port, Immediate(6) => 
                           IMMEDIATE_16_6_port, Immediate(5) => 
                           IMMEDIATE_16_5_port, Immediate(4) => 
                           IMMEDIATE_16_4_port, Immediate(3) => 
                           IMMEDIATE_16_3_port, Immediate(2) => 
                           IMMEDIATE_16_2_port, Immediate(1) => 
                           IMMEDIATE_16_1_port, Immediate(0) => 
                           IMMEDIATE_16_0_port);
   SIGN_EXTENSION_imm26 : sign_eval_N_in26_N_out32 port map( IR_out(25) => 
                           IR_26(25), IR_out(24) => IR_26(24), IR_out(23) => 
                           IR_26(23), IR_out(22) => IR_26(22), IR_out(21) => 
                           IR_26(21), IR_out(20) => IR_26(20), IR_out(19) => 
                           IR_26(19), IR_out(18) => IR_26(18), IR_out(17) => 
                           IR_26(17), IR_out(16) => IR_26(16), IR_out(15) => 
                           IR_26(15), IR_out(14) => IR_26(14), IR_out(13) => 
                           IR_26(13), IR_out(12) => IR_26(12), IR_out(11) => 
                           IR_26(11), IR_out(10) => IR_26(10), IR_out(9) => 
                           IR_26(9), IR_out(8) => IR_26(8), IR_out(7) => 
                           IR_26(7), IR_out(6) => IR_26(6), IR_out(5) => 
                           IR_26(5), IR_out(4) => IR_26(4), IR_out(3) => 
                           IR_26(3), IR_out(2) => IR_26(2), IR_out(1) => 
                           IR_26(1), IR_out(0) => IR_26(0), signed_val => 
                           X_Logic0_port, Immediate(31) => n_2212, 
                           Immediate(30) => n_2213, Immediate(29) => n_2214, 
                           Immediate(28) => n_2215, Immediate(27) => n_2216, 
                           Immediate(26) => n_2217, Immediate(25) => n_2218, 
                           Immediate(24) => n_2219, Immediate(23) => n_2220, 
                           Immediate(22) => n_2221, Immediate(21) => n_2222, 
                           Immediate(20) => n_2223, Immediate(19) => n_2224, 
                           Immediate(18) => n_2225, Immediate(17) => n_2226, 
                           Immediate(16) => n_2227, Immediate(15) => n_2228, 
                           Immediate(14) => n_2229, Immediate(13) => n_2230, 
                           Immediate(12) => n_2231, Immediate(11) => n_2232, 
                           Immediate(10) => n_2233, Immediate(9) => n_2234, 
                           Immediate(8) => n_2235, Immediate(7) => n_2236, 
                           Immediate(6) => n_2237, Immediate(5) => n_2238, 
                           Immediate(4) => n_2239, Immediate(3) => n_2240, 
                           Immediate(2) => n_2241, Immediate(1) => n_2242, 
                           Immediate(0) => n_2243);
   U3 : NAND4_X1 port map( A1 => n8, A2 => n21, A3 => n22, A4 => n23, ZN => n1)
                           ;
   U4 : NAND4_X1 port map( A1 => n8, A2 => n21, A3 => n22, A4 => n23, ZN => n38
                           );
   U5 : NAND4_X1 port map( A1 => n7, A2 => n24, A3 => n25, A4 => n26, ZN => n2)
                           ;
   U6 : INV_X1 port map( A => OPCODE(3), ZN => n3);
   U7 : AND3_X2 port map( A1 => n3, A2 => n28, A3 => n27, ZN => n8);
   U8 : MUX2_X1 port map( A => IR_26(15), B => IR_26(20), S => n4, Z => N147);
   U9 : NAND4_X1 port map( A1 => n8, A2 => n19, A3 => n20, A4 => n23, ZN => n4)
                           ;
   U10 : AND3_X1 port map( A1 => n11, A2 => n12, A3 => n29, ZN => n5);
   U11 : AND3_X1 port map( A1 => n11, A2 => n12, A3 => n3, ZN => n7);
   U12 : MUX2_X1 port map( A => IR_26(14), B => IR_26(19), S => n35, Z => N146)
                           ;
   U13 : AND3_X2 port map( A1 => n11, A2 => n29, A3 => n12, ZN => n6);
   U14 : AND2_X2 port map( A1 => n34, A2 => IMMEDIATE_16_31_port, ZN => n32);
   U15 : NAND3_X1 port map( A1 => n28, A2 => n13, A3 => n27, ZN => n9);
   U16 : NAND4_X1 port map( A1 => n6, A2 => n24, A3 => n25, A4 => n15, ZN => 
                           n33);
   U17 : NAND4_X1 port map( A1 => n6, A2 => n16, A3 => n14, A4 => n15, ZN => 
                           n10);
   U18 : INV_X1 port map( A => OPCODE(5), ZN => n11);
   U19 : INV_X1 port map( A => OPCODE(4), ZN => n12);
   U20 : INV_X1 port map( A => OPCODE(3), ZN => n13);
   U21 : NAND4_X1 port map( A1 => n6, A2 => n21, A3 => n14, A4 => n15, ZN => 
                           n34);
   U22 : INV_X1 port map( A => OPCODE(0), ZN => n14);
   U23 : INV_X1 port map( A => OPCODE(2), ZN => n15);
   U24 : NAND4_X1 port map( A1 => n5, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n35);
   U25 : INV_X1 port map( A => OPCODE(1), ZN => n16);
   U26 : INV_X1 port map( A => OPCODE(2), ZN => n17);
   U27 : INV_X1 port map( A => OPCODE(0), ZN => n18);
   U28 : NAND4_X1 port map( A1 => n17, A2 => n19, A3 => n20, A4 => n6, ZN => 
                           n30);
   U29 : INV_X1 port map( A => OPCODE(1), ZN => n19);
   U30 : INV_X1 port map( A => OPCODE(0), ZN => n20);
   U31 : INV_X1 port map( A => OPCODE(1), ZN => n21);
   U32 : INV_X1 port map( A => OPCODE(0), ZN => n22);
   U33 : INV_X1 port map( A => OPCODE(2), ZN => n23);
   U34 : NAND4_X1 port map( A1 => n7, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           n37);
   U35 : INV_X1 port map( A => OPCODE(1), ZN => n24);
   U36 : INV_X1 port map( A => OPCODE(0), ZN => n25);
   U37 : INV_X1 port map( A => OPCODE(2), ZN => n26);
   U38 : INV_X1 port map( A => OPCODE(5), ZN => n27);
   U39 : INV_X1 port map( A => OPCODE(4), ZN => n28);
   U40 : INV_X1 port map( A => OPCODE(3), ZN => n29);
   U41 : MUX2_X1 port map( A => IR_26(18), B => IR_26(13), S => n31, Z => N145)
                           ;
   U42 : NOR4_X1 port map( A1 => n9, A2 => OPCODE(1), A3 => OPCODE(0), A4 => 
                           OPCODE(2), ZN => n31);
   U43 : AND2_X1 port map( A1 => n33, A2 => IMMEDIATE_16_31_port, ZN => n36);
   U44 : AND2_X1 port map( A1 => n1, A2 => IMMEDIATE_16_15_port, ZN => N163);
   U45 : AND2_X1 port map( A1 => n10, A2 => IMMEDIATE_16_14_port, ZN => N162);
   U46 : AND2_X1 port map( A1 => n33, A2 => IMMEDIATE_16_13_port, ZN => N161);
   U47 : AND2_X1 port map( A1 => n1, A2 => IMMEDIATE_16_12_port, ZN => N160);
   U48 : AND2_X1 port map( A1 => n38, A2 => IMMEDIATE_16_11_port, ZN => N159);
   U49 : AND2_X1 port map( A1 => n1, A2 => IMMEDIATE_16_10_port, ZN => N158);
   U50 : AND2_X1 port map( A1 => n10, A2 => IMMEDIATE_16_9_port, ZN => N157);
   U51 : AND2_X1 port map( A1 => n1, A2 => IMMEDIATE_16_8_port, ZN => N156);
   U52 : AND2_X1 port map( A1 => n38, A2 => IMMEDIATE_16_7_port, ZN => N155);
   U53 : AND2_X1 port map( A1 => n30, A2 => IMMEDIATE_16_6_port, ZN => N154);
   U54 : AND2_X1 port map( A1 => n30, A2 => IMMEDIATE_16_5_port, ZN => N153);
   U55 : AND2_X1 port map( A1 => n38, A2 => IMMEDIATE_16_4_port, ZN => N152);
   U56 : AND2_X1 port map( A1 => n38, A2 => IMMEDIATE_16_3_port, ZN => N151);
   U57 : AND2_X1 port map( A1 => n10, A2 => IMMEDIATE_16_2_port, ZN => N150);
   U58 : AND2_X1 port map( A1 => n10, A2 => IMMEDIATE_16_1_port, ZN => N149);
   U59 : AND2_X1 port map( A1 => n30, A2 => IMMEDIATE_16_0_port, ZN => N148);
   U60 : MUX2_X1 port map( A => IR_26(12), B => IR_26(17), S => n2, Z => N144);
   U61 : MUX2_X1 port map( A => IR_26(11), B => IR_26(16), S => n37, Z => N143)
                           ;

end SYN_BEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_0;

architecture SYN_struct of MUX21_GENERIC_NBIT32_0 is

   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_225
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_226
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_227
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_228
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_229
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_230
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_231
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_232
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_233
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_234
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_235
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_236
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_237
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_238
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_239
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_240
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_241
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_242
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_243
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_244
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_245
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_246
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_247
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_248
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_249
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_250
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_251
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_252
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_253
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_254
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_255
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   gen1_0 : MUX21_0 port map( A => A(0), B => B(0), S => n3, Y => Y(0));
   gen1_1 : MUX21_255 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   gen1_2 : MUX21_254 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   gen1_3 : MUX21_253 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   gen1_4 : MUX21_252 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   gen1_5 : MUX21_251 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   gen1_6 : MUX21_250 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   gen1_7 : MUX21_249 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   gen1_8 : MUX21_248 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   gen1_9 : MUX21_247 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   gen1_10 : MUX21_246 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   gen1_11 : MUX21_245 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   gen1_12 : MUX21_244 port map( A => A(12), B => B(12), S => n1, Y => Y(12));
   gen1_13 : MUX21_243 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   gen1_14 : MUX21_242 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   gen1_15 : MUX21_241 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   gen1_16 : MUX21_240 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   gen1_17 : MUX21_239 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   gen1_18 : MUX21_238 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   gen1_19 : MUX21_237 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   gen1_20 : MUX21_236 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   gen1_21 : MUX21_235 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   gen1_22 : MUX21_234 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   gen1_23 : MUX21_233 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   gen1_24 : MUX21_232 port map( A => A(24), B => B(24), S => n2, Y => Y(24));
   gen1_25 : MUX21_231 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   gen1_26 : MUX21_230 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   gen1_27 : MUX21_229 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   gen1_28 : MUX21_228 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   gen1_29 : MUX21_227 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   gen1_30 : MUX21_226 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   gen1_31 : MUX21_225 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : CLKBUF_X3 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X3 port map( A => SEL, Z => n2);
   U3 : CLKBUF_X3 port map( A => SEL, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n96, CK => CK, RN => RESET, Q => 
                           Q(31), QN => n64);
   Q_reg_30_inst : DFFR_X1 port map( D => n95, CK => CK, RN => RESET, Q => 
                           Q(30), QN => n63);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => CK, RN => RESET, Q => 
                           Q(29), QN => n62);
   Q_reg_28_inst : DFFR_X1 port map( D => n93, CK => CK, RN => RESET, Q => 
                           Q(28), QN => n61);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => CK, RN => RESET, Q => 
                           Q(27), QN => n60);
   Q_reg_26_inst : DFFR_X1 port map( D => n91, CK => CK, RN => RESET, Q => 
                           Q(26), QN => n59);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => CK, RN => RESET, Q => 
                           Q(25), QN => n58);
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => CK, RN => RESET, Q => 
                           Q(24), QN => n57);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => CK, RN => RESET, Q => 
                           Q(23), QN => n56);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => CK, RN => RESET, Q => 
                           Q(22), QN => n55);
   Q_reg_21_inst : DFFR_X1 port map( D => n86, CK => CK, RN => RESET, Q => 
                           Q(21), QN => n54);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => CK, RN => RESET, Q => 
                           Q(20), QN => n53);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => CK, RN => RESET, Q => 
                           Q(19), QN => n52);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => CK, RN => RESET, Q => 
                           Q(18), QN => n51);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => CK, RN => RESET, Q => 
                           Q(17), QN => n50);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => CK, RN => RESET, Q => 
                           Q(16), QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => CK, RN => RESET, Q => 
                           Q(15), QN => n48);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => CK, RN => RESET, Q => 
                           Q(14), QN => n47);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => CK, RN => RESET, Q => 
                           Q(13), QN => n46);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => CK, RN => RESET, Q => 
                           Q(12), QN => n45);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => CK, RN => RESET, Q => 
                           Q(11), QN => n44);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => CK, RN => RESET, Q => 
                           Q(10), QN => n43);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => CK, RN => RESET, Q => Q(9),
                           QN => n42);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => CK, RN => RESET, Q => Q(8),
                           QN => n41);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => CK, RN => RESET, Q => Q(7),
                           QN => n40);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => CK, RN => RESET, Q => Q(6),
                           QN => n39);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => CK, RN => RESET, Q => Q(5),
                           QN => n38);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => CK, RN => RESET, Q => Q(4),
                           QN => n37);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => CK, RN => RESET, Q => Q(3),
                           QN => n36);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => CK, RN => RESET, Q => Q(2),
                           QN => n35);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => CK, RN => RESET, Q => Q(1),
                           QN => n34);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => CK, RN => RESET, Q => Q(0),
                           QN => n33);
   U2 : OAI21_X1 port map( B1 => n33, B2 => ENABLE, A => n1, ZN => n65);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => n34, B2 => ENABLE, A => n2, ZN => n66);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n35, B2 => ENABLE, A => n3, ZN => n67);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n36, B2 => ENABLE, A => n4, ZN => n68);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n4);
   U10 : OAI21_X1 port map( B1 => n37, B2 => ENABLE, A => n5, ZN => n69);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n5);
   U12 : OAI21_X1 port map( B1 => n38, B2 => ENABLE, A => n6, ZN => n70);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n6);
   U14 : OAI21_X1 port map( B1 => n39, B2 => ENABLE, A => n7, ZN => n71);
   U15 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n7);
   U16 : OAI21_X1 port map( B1 => n40, B2 => ENABLE, A => n8, ZN => n72);
   U17 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n8);
   U18 : OAI21_X1 port map( B1 => n41, B2 => ENABLE, A => n9, ZN => n73);
   U19 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n9);
   U20 : OAI21_X1 port map( B1 => n42, B2 => ENABLE, A => n10, ZN => n74);
   U21 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n10);
   U22 : OAI21_X1 port map( B1 => n43, B2 => ENABLE, A => n11, ZN => n75);
   U23 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n11);
   U24 : OAI21_X1 port map( B1 => n44, B2 => ENABLE, A => n12, ZN => n76);
   U25 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n12);
   U26 : OAI21_X1 port map( B1 => n45, B2 => ENABLE, A => n13, ZN => n77);
   U27 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n13);
   U28 : OAI21_X1 port map( B1 => n46, B2 => ENABLE, A => n14, ZN => n78);
   U29 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n14);
   U30 : OAI21_X1 port map( B1 => n47, B2 => ENABLE, A => n15, ZN => n79);
   U31 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n15);
   U32 : OAI21_X1 port map( B1 => n48, B2 => ENABLE, A => n16, ZN => n80);
   U33 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n16);
   U34 : OAI21_X1 port map( B1 => n49, B2 => ENABLE, A => n17, ZN => n81);
   U35 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n17);
   U36 : OAI21_X1 port map( B1 => n50, B2 => ENABLE, A => n18, ZN => n82);
   U37 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n18);
   U38 : OAI21_X1 port map( B1 => n51, B2 => ENABLE, A => n19, ZN => n83);
   U39 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n19);
   U40 : OAI21_X1 port map( B1 => n52, B2 => ENABLE, A => n20, ZN => n84);
   U41 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n20);
   U42 : OAI21_X1 port map( B1 => n53, B2 => ENABLE, A => n21, ZN => n85);
   U43 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n21);
   U44 : OAI21_X1 port map( B1 => n54, B2 => ENABLE, A => n22, ZN => n86);
   U45 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n22);
   U46 : OAI21_X1 port map( B1 => n55, B2 => ENABLE, A => n23, ZN => n87);
   U47 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n23);
   U48 : OAI21_X1 port map( B1 => n56, B2 => ENABLE, A => n24, ZN => n88);
   U49 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n24);
   U50 : OAI21_X1 port map( B1 => n57, B2 => ENABLE, A => n25, ZN => n89);
   U51 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n25);
   U52 : OAI21_X1 port map( B1 => n58, B2 => ENABLE, A => n26, ZN => n90);
   U53 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n26);
   U54 : OAI21_X1 port map( B1 => n59, B2 => ENABLE, A => n27, ZN => n91);
   U55 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n27);
   U56 : OAI21_X1 port map( B1 => n60, B2 => ENABLE, A => n28, ZN => n92);
   U57 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n28);
   U58 : OAI21_X1 port map( B1 => n61, B2 => ENABLE, A => n29, ZN => n93);
   U59 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n29);
   U60 : OAI21_X1 port map( B1 => n62, B2 => ENABLE, A => n30, ZN => n94);
   U61 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n30);
   U62 : OAI21_X1 port map( B1 => n63, B2 => ENABLE, A => n31, ZN => n95);
   U63 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n31);
   U64 : OAI21_X1 port map( B1 => n64, B2 => ENABLE, A => n32, ZN => n96);
   U65 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n32);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DATAPTH_NBIT32_REG_BIT5 is

   port( CLK, RST : in std_logic;  PC, IR : in std_logic_vector (31 downto 0); 
         PC_OUT : out std_logic_vector (31 downto 0);  NPC_LATCH_EN, 
         ir_LATCH_EN, signed_op, RF1, RF2, WF1, regImm_LATCH_EN, S1, S2, EN2, 
         lhi_sel, jump_en, branch_cond, sb_op, RM, WM, EN3, S3 : in std_logic; 
         instruction_alu : in std_logic_vector (0 to 5);  DATA_MEM_ADDR, 
         DATA_MEM_IN : out std_logic_vector (31 downto 0);  DATA_MEM_OUT : in 
         std_logic_vector (31 downto 0);  DATA_MEM_ENABLE, DATA_MEM_RM, 
         DATA_MEM_WM : out std_logic);

end DATAPTH_NBIT32_REG_BIT5;

architecture SYN_STRUCTURAL of DATAPTH_NBIT32_REG_BIT5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DATAPTH_NBIT32_REG_BIT5_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_1
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FF_2
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FF_3
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_2
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_3
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component load_data
      port( data_in : in std_logic_vector (31 downto 0);  signed_val, load_op :
            in std_logic;  load_type : in std_logic_vector (1 downto 0);  
            data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT6_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 
            downto 0);  Q : out std_logic_vector (5 downto 0));
   end component;
   
   component FF_4
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_2
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_4
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_5
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT32_5
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_6
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component COND_BT_NBIT32
      port( ZERO_BIT, OPCODE_0, branch_op : in std_logic;  con_sign : out 
            std_logic);
   end component;
   
   component zero_eval_NBIT32
      port( input : in std_logic_vector (31 downto 0);  res : out std_logic);
   end component;
   
   component ALU_N32
      port( CLK : in std_logic;  FUNC : in std_logic_vector (0 to 5);  DATA1, 
            DATA2 : in std_logic_vector (31 downto 0);  OUT_ALU : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_6
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT6_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 
            downto 0);  Q : out std_logic_vector (5 downto 0));
   end component;
   
   component FF_7
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_7
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_8
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_9
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_10
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_0
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component register_file
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0);  wr_signal : in std_logic);
   end component;
   
   component IR_DECODE_NBIT32_opBIT6_regBIT5
      port( CLK : in std_logic;  IR_26 : in std_logic_vector (25 downto 0);  
            OPCODE : in std_logic_vector (5 downto 0);  is_signed : in 
            std_logic;  RS1, RS2, RD : out std_logic_vector (4 downto 0);  
            IMMEDIATE : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_11
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_12
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_13
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_14
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_15
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_16
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_17
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_18
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, PC_fetch0_31_port, PC_fetch0_30_port, 
      PC_fetch0_29_port, PC_fetch0_28_port, PC_fetch0_27_port, 
      PC_fetch0_26_port, PC_fetch0_25_port, PC_fetch0_24_port, 
      PC_fetch0_23_port, PC_fetch0_22_port, PC_fetch0_21_port, 
      PC_fetch0_20_port, PC_fetch0_19_port, PC_fetch0_18_port, 
      PC_fetch0_17_port, PC_fetch0_16_port, PC_fetch0_15_port, 
      PC_fetch0_14_port, PC_fetch0_13_port, PC_fetch0_12_port, 
      PC_fetch0_11_port, PC_fetch0_10_port, PC_fetch0_9_port, PC_fetch0_8_port,
      PC_fetch0_7_port, PC_fetch0_6_port, PC_fetch0_5_port, PC_fetch0_4_port, 
      PC_fetch0_3_port, PC_fetch0_2_port, PC_fetch0_1_port, PC_fetch0_0_port, 
      NPC_31_port, NPC_30_port, NPC_29_port, NPC_28_port, NPC_27_port, 
      NPC_26_port, NPC_25_port, NPC_24_port, NPC_23_port, NPC_22_port, 
      NPC_21_port, NPC_20_port, NPC_19_port, NPC_18_port, NPC_17_port, 
      NPC_16_port, NPC_15_port, NPC_14_port, NPC_13_port, NPC_12_port, 
      NPC_11_port, NPC_10_port, NPC_9_port, NPC_8_port, NPC_7_port, NPC_6_port,
      NPC_5_port, NPC_4_port, NPC_3_port, NPC_2_port, NPC_1_port, NPC_0_port, 
      NPC_fetch1_31_port, NPC_fetch1_30_port, NPC_fetch1_29_port, 
      NPC_fetch1_28_port, NPC_fetch1_27_port, NPC_fetch1_26_port, 
      NPC_fetch1_25_port, NPC_fetch1_24_port, NPC_fetch1_23_port, 
      NPC_fetch1_22_port, NPC_fetch1_21_port, NPC_fetch1_20_port, 
      NPC_fetch1_19_port, NPC_fetch1_18_port, NPC_fetch1_17_port, 
      NPC_fetch1_16_port, NPC_fetch1_15_port, NPC_fetch1_14_port, 
      NPC_fetch1_13_port, NPC_fetch1_12_port, NPC_fetch1_11_port, 
      NPC_fetch1_10_port, NPC_fetch1_9_port, NPC_fetch1_8_port, 
      NPC_fetch1_7_port, NPC_fetch1_6_port, NPC_fetch1_5_port, 
      NPC_fetch1_4_port, NPC_fetch1_3_port, NPC_fetch1_2_port, 
      NPC_fetch1_1_port, NPC_fetch1_0_port, PC_fetch1_31_port, 
      PC_fetch1_30_port, PC_fetch1_29_port, PC_fetch1_28_port, 
      PC_fetch1_27_port, PC_fetch1_26_port, PC_fetch1_25_port, 
      PC_fetch1_24_port, PC_fetch1_23_port, PC_fetch1_22_port, 
      PC_fetch1_21_port, PC_fetch1_20_port, PC_fetch1_19_port, 
      PC_fetch1_18_port, PC_fetch1_17_port, PC_fetch1_16_port, 
      PC_fetch1_15_port, PC_fetch1_14_port, PC_fetch1_13_port, 
      PC_fetch1_12_port, PC_fetch1_11_port, PC_fetch1_10_port, PC_fetch1_9_port
      , PC_fetch1_8_port, PC_fetch1_7_port, PC_fetch1_6_port, PC_fetch1_5_port,
      PC_fetch1_4_port, PC_fetch1_3_port, PC_fetch1_2_port, PC_fetch1_1_port, 
      PC_fetch1_0_port, PC_OUT_i_31_port, PC_OUT_i_30_port, PC_OUT_i_29_port, 
      PC_OUT_i_28_port, PC_OUT_i_27_port, PC_OUT_i_26_port, PC_OUT_i_25_port, 
      PC_OUT_i_24_port, PC_OUT_i_23_port, PC_OUT_i_22_port, PC_OUT_i_21_port, 
      PC_OUT_i_20_port, PC_OUT_i_19_port, PC_OUT_i_18_port, PC_OUT_i_17_port, 
      PC_OUT_i_16_port, PC_OUT_i_15_port, PC_OUT_i_14_port, PC_OUT_i_13_port, 
      PC_OUT_i_12_port, PC_OUT_i_11_port, PC_OUT_i_10_port, PC_OUT_i_9_port, 
      PC_OUT_i_8_port, PC_OUT_i_7_port, PC_OUT_i_6_port, PC_OUT_i_5_port, 
      PC_OUT_i_4_port, PC_OUT_i_3_port, PC_OUT_i_2_port, PC_OUT_i_1_port, 
      PC_OUT_i_0_port, sel_npc, NPC_fetch_31_port, NPC_fetch_30_port, 
      NPC_fetch_29_port, NPC_fetch_28_port, NPC_fetch_27_port, 
      NPC_fetch_26_port, NPC_fetch_25_port, NPC_fetch_24_port, 
      NPC_fetch_23_port, NPC_fetch_22_port, NPC_fetch_21_port, 
      NPC_fetch_20_port, NPC_fetch_19_port, NPC_fetch_18_port, 
      NPC_fetch_17_port, NPC_fetch_16_port, NPC_fetch_15_port, 
      NPC_fetch_14_port, NPC_fetch_13_port, NPC_fetch_12_port, 
      NPC_fetch_11_port, NPC_fetch_10_port, NPC_fetch_9_port, NPC_fetch_8_port,
      NPC_fetch_7_port, NPC_fetch_6_port, NPC_fetch_5_port, NPC_fetch_4_port, 
      NPC_fetch_3_port, NPC_fetch_2_port, NPC_fetch_1_port, NPC_fetch_0_port, 
      PC_fetch_31_port, PC_fetch_30_port, PC_fetch_29_port, PC_fetch_28_port, 
      PC_fetch_27_port, PC_fetch_26_port, PC_fetch_25_port, PC_fetch_24_port, 
      PC_fetch_23_port, PC_fetch_22_port, PC_fetch_21_port, PC_fetch_20_port, 
      PC_fetch_19_port, PC_fetch_18_port, PC_fetch_17_port, PC_fetch_16_port, 
      PC_fetch_15_port, PC_fetch_14_port, PC_fetch_13_port, PC_fetch_12_port, 
      PC_fetch_11_port, PC_fetch_10_port, PC_fetch_9_port, PC_fetch_8_port, 
      PC_fetch_7_port, PC_fetch_6_port, PC_fetch_5_port, PC_fetch_4_port, 
      PC_fetch_3_port, PC_fetch_2_port, PC_fetch_1_port, PC_fetch_0_port, 
      ir_fetch_31_port, ir_fetch_30_port, ir_fetch_29_port, ir_fetch_28_port, 
      ir_fetch_27_port, ir_fetch_26_port, ir_fetch_25_port, ir_fetch_24_port, 
      ir_fetch_23_port, ir_fetch_22_port, ir_fetch_21_port, ir_fetch_20_port, 
      ir_fetch_19_port, ir_fetch_18_port, ir_fetch_17_port, ir_fetch_16_port, 
      ir_fetch_15_port, ir_fetch_14_port, ir_fetch_13_port, ir_fetch_12_port, 
      ir_fetch_11_port, ir_fetch_10_port, ir_fetch_9_port, ir_fetch_8_port, 
      ir_fetch_7_port, ir_fetch_6_port, ir_fetch_5_port, ir_fetch_4_port, 
      ir_fetch_3_port, ir_fetch_2_port, ir_fetch_1_port, ir_fetch_0_port, 
      NPC_Dec_31_port, NPC_Dec_30_port, NPC_Dec_29_port, NPC_Dec_28_port, 
      NPC_Dec_27_port, NPC_Dec_26_port, NPC_Dec_25_port, NPC_Dec_24_port, 
      NPC_Dec_23_port, NPC_Dec_22_port, NPC_Dec_21_port, NPC_Dec_20_port, 
      NPC_Dec_19_port, NPC_Dec_18_port, NPC_Dec_17_port, NPC_Dec_16_port, 
      NPC_Dec_15_port, NPC_Dec_14_port, NPC_Dec_13_port, NPC_Dec_12_port, 
      NPC_Dec_11_port, NPC_Dec_10_port, NPC_Dec_9_port, NPC_Dec_8_port, 
      NPC_Dec_7_port, NPC_Dec_6_port, NPC_Dec_5_port, NPC_Dec_4_port, 
      NPC_Dec_3_port, NPC_Dec_2_port, NPC_Dec_1_port, NPC_Dec_0_port, 
      IR_Dec_31_port, IR_Dec_30_port, IR_Dec_29_port, IR_Dec_28_port, 
      IR_Dec_27_port, IR_Dec_26_port, IR_Dec_25_port, IR_Dec_24_port, 
      IR_Dec_23_port, IR_Dec_22_port, IR_Dec_21_port, IR_Dec_20_port, 
      IR_Dec_19_port, IR_Dec_18_port, IR_Dec_17_port, IR_Dec_16_port, 
      IR_Dec_15_port, IR_Dec_14_port, IR_Dec_13_port, IR_Dec_12_port, 
      IR_Dec_11_port, IR_Dec_10_port, IR_Dec_9_port, IR_Dec_8_port, 
      IR_Dec_7_port, IR_Dec_6_port, IR_Dec_5_port, IR_Dec_4_port, IR_Dec_3_port
      , IR_Dec_2_port, IR_Dec_1_port, IR_Dec_0_port, RS1_4_port, RS1_3_port, 
      RS1_2_port, RS1_1_port, RS1_0_port, RS2_4_port, RS2_3_port, RS2_2_port, 
      RS2_1_port, RS2_0_port, RD_4_port, RD_3_port, RD_2_port, RD_1_port, 
      RD_0_port, Imm_31_port, Imm_30_port, Imm_29_port, Imm_28_port, 
      Imm_27_port, Imm_26_port, Imm_25_port, Imm_24_port, Imm_23_port, 
      Imm_22_port, Imm_21_port, Imm_20_port, Imm_19_port, Imm_18_port, 
      Imm_17_port, Imm_16_port, Imm_15_port, Imm_14_port, Imm_13_port, 
      Imm_12_port, Imm_11_port, Imm_10_port, Imm_9_port, Imm_8_port, Imm_7_port
      , Imm_6_port, Imm_5_port, Imm_4_port, Imm_3_port, Imm_2_port, Imm_1_port,
      Imm_0_port, wr_signal, RD_wb_4_port, RD_wb_3_port, RD_wb_2_port, 
      RD_wb_1_port, RD_wb_0_port, OUT_data_31_port, OUT_data_30_port, 
      OUT_data_29_port, OUT_data_28_port, OUT_data_27_port, OUT_data_26_port, 
      OUT_data_25_port, OUT_data_24_port, OUT_data_23_port, OUT_data_22_port, 
      OUT_data_21_port, OUT_data_20_port, OUT_data_19_port, OUT_data_18_port, 
      OUT_data_17_port, OUT_data_16_port, OUT_data_15_port, OUT_data_14_port, 
      OUT_data_13_port, OUT_data_12_port, OUT_data_11_port, OUT_data_10_port, 
      OUT_data_9_port, OUT_data_8_port, OUT_data_7_port, OUT_data_6_port, 
      OUT_data_5_port, OUT_data_4_port, OUT_data_3_port, OUT_data_2_port, 
      OUT_data_1_port, OUT_data_0_port, regA_31_port, regA_30_port, 
      regA_29_port, regA_28_port, regA_27_port, regA_26_port, regA_25_port, 
      regA_24_port, regA_23_port, regA_22_port, regA_21_port, regA_20_port, 
      regA_19_port, regA_18_port, regA_17_port, regA_16_port, regA_15_port, 
      regA_14_port, regA_13_port, regA_12_port, regA_11_port, regA_10_port, 
      regA_9_port, regA_8_port, regA_7_port, regA_6_port, regA_5_port, 
      regA_4_port, regA_3_port, regA_2_port, regA_1_port, regA_0_port, 
      regB_31_port, regB_30_port, regB_29_port, regB_28_port, regB_27_port, 
      regB_26_port, regB_25_port, regB_24_port, regB_23_port, regB_22_port, 
      regB_21_port, regB_20_port, regB_19_port, regB_18_port, regB_17_port, 
      regB_16_port, regB_15_port, regB_14_port, regB_13_port, regB_12_port, 
      regB_11_port, regB_10_port, regB_9_port, regB_8_port, regB_7_port, 
      regB_6_port, regB_5_port, regB_4_port, regB_3_port, regB_2_port, 
      regB_1_port, regB_0_port, wr_signal_wb, signed_op_ex, NPC_ex_31_port, 
      NPC_ex_30_port, NPC_ex_29_port, NPC_ex_28_port, NPC_ex_27_port, 
      NPC_ex_26_port, NPC_ex_25_port, NPC_ex_24_port, NPC_ex_23_port, 
      NPC_ex_22_port, NPC_ex_21_port, NPC_ex_20_port, NPC_ex_19_port, 
      NPC_ex_18_port, NPC_ex_17_port, NPC_ex_16_port, NPC_ex_15_port, 
      NPC_ex_14_port, NPC_ex_13_port, NPC_ex_12_port, NPC_ex_11_port, 
      NPC_ex_10_port, NPC_ex_9_port, NPC_ex_8_port, NPC_ex_7_port, 
      NPC_ex_6_port, NPC_ex_5_port, NPC_ex_4_port, NPC_ex_3_port, NPC_ex_2_port
      , NPC_ex_1_port, NPC_ex_0_port, regA_ex_31_port, regA_ex_30_port, 
      regA_ex_29_port, regA_ex_28_port, regA_ex_27_port, regA_ex_26_port, 
      regA_ex_25_port, regA_ex_24_port, regA_ex_23_port, regA_ex_22_port, 
      regA_ex_21_port, regA_ex_20_port, regA_ex_19_port, regA_ex_18_port, 
      regA_ex_17_port, regA_ex_16_port, regA_ex_15_port, regA_ex_14_port, 
      regA_ex_13_port, regA_ex_12_port, regA_ex_11_port, regA_ex_10_port, 
      regA_ex_9_port, regA_ex_8_port, regA_ex_7_port, regA_ex_6_port, 
      regA_ex_5_port, regA_ex_4_port, regA_ex_3_port, regA_ex_2_port, 
      regA_ex_1_port, regA_ex_0_port, regB_ex_31_port, regB_ex_30_port, 
      regB_ex_29_port, regB_ex_28_port, regB_ex_27_port, regB_ex_26_port, 
      regB_ex_25_port, regB_ex_24_port, regB_ex_23_port, regB_ex_22_port, 
      regB_ex_21_port, regB_ex_20_port, regB_ex_19_port, regB_ex_18_port, 
      regB_ex_17_port, regB_ex_16_port, regB_ex_15_port, regB_ex_14_port, 
      regB_ex_13_port, regB_ex_12_port, regB_ex_11_port, regB_ex_10_port, 
      regB_ex_9_port, regB_ex_8_port, regB_ex_7_port, regB_ex_6_port, 
      regB_ex_5_port, regB_ex_4_port, regB_ex_3_port, regB_ex_2_port, 
      regB_ex_1_port, regB_ex_0_port, Imm_ex_31_port, Imm_ex_30_port, 
      Imm_ex_29_port, Imm_ex_28_port, Imm_ex_27_port, Imm_ex_26_port, 
      Imm_ex_25_port, Imm_ex_24_port, Imm_ex_23_port, Imm_ex_22_port, 
      Imm_ex_21_port, Imm_ex_20_port, Imm_ex_19_port, Imm_ex_18_port, 
      Imm_ex_17_port, Imm_ex_16_port, Imm_ex_15_port, Imm_ex_14_port, 
      Imm_ex_13_port, Imm_ex_12_port, Imm_ex_11_port, Imm_ex_10_port, 
      Imm_ex_9_port, Imm_ex_8_port, Imm_ex_7_port, Imm_ex_6_port, Imm_ex_5_port
      , Imm_ex_4_port, Imm_ex_3_port, Imm_ex_2_port, Imm_ex_1_port, 
      Imm_ex_0_port, RD_ex_4_port, RD_ex_3_port, RD_ex_2_port, RD_ex_1_port, 
      RD_ex_0_port, wr_signal_exe, IR_26_ex_5_port, IR_26_ex_4_port, 
      IR_26_ex_3_port, IR_26_ex_2_port, IR_26_ex_1_port, IR_26_ex_0_port, 
      LHI_ex_31_port, LHI_ex_30_port, LHI_ex_29_port, LHI_ex_28_port, 
      LHI_ex_27_port, LHI_ex_26_port, LHI_ex_25_port, LHI_ex_24_port, 
      LHI_ex_23_port, LHI_ex_22_port, LHI_ex_21_port, LHI_ex_20_port, 
      LHI_ex_19_port, LHI_ex_18_port, LHI_ex_17_port, LHI_ex_16_port, 
      LHI_ex_15_port, LHI_ex_14_port, LHI_ex_13_port, LHI_ex_12_port, 
      LHI_ex_11_port, LHI_ex_10_port, LHI_ex_9_port, LHI_ex_8_port, 
      LHI_ex_7_port, LHI_ex_6_port, LHI_ex_5_port, LHI_ex_4_port, LHI_ex_3_port
      , LHI_ex_2_port, LHI_ex_1_port, LHI_ex_0_port, input1_ALU_31_port, 
      input1_ALU_30_port, input1_ALU_29_port, input1_ALU_28_port, 
      input1_ALU_27_port, input1_ALU_26_port, input1_ALU_25_port, 
      input1_ALU_24_port, input1_ALU_23_port, input1_ALU_22_port, 
      input1_ALU_21_port, input1_ALU_20_port, input1_ALU_19_port, 
      input1_ALU_18_port, input1_ALU_17_port, input1_ALU_16_port, 
      input1_ALU_15_port, input1_ALU_14_port, input1_ALU_13_port, 
      input1_ALU_12_port, input1_ALU_11_port, input1_ALU_10_port, 
      input1_ALU_9_port, input1_ALU_8_port, input1_ALU_7_port, 
      input1_ALU_6_port, input1_ALU_5_port, input1_ALU_4_port, 
      input1_ALU_3_port, input1_ALU_2_port, input1_ALU_1_port, 
      input1_ALU_0_port, input2_ALU_31_port, input2_ALU_30_port, 
      input2_ALU_29_port, input2_ALU_28_port, input2_ALU_27_port, 
      input2_ALU_26_port, input2_ALU_25_port, input2_ALU_24_port, 
      input2_ALU_23_port, input2_ALU_22_port, input2_ALU_21_port, 
      input2_ALU_20_port, input2_ALU_19_port, input2_ALU_18_port, 
      input2_ALU_17_port, input2_ALU_16_port, input2_ALU_15_port, 
      input2_ALU_14_port, input2_ALU_13_port, input2_ALU_12_port, 
      input2_ALU_11_port, input2_ALU_10_port, input2_ALU_9_port, 
      input2_ALU_8_port, input2_ALU_7_port, input2_ALU_6_port, 
      input2_ALU_5_port, input2_ALU_4_port, input2_ALU_3_port, 
      input2_ALU_2_port, input2_ALU_1_port, input2_ALU_0_port, ALU_out_31_port,
      ALU_out_30_port, ALU_out_29_port, ALU_out_28_port, ALU_out_27_port, 
      ALU_out_26_port, ALU_out_25_port, ALU_out_24_port, ALU_out_23_port, 
      ALU_out_22_port, ALU_out_21_port, ALU_out_20_port, ALU_out_19_port, 
      ALU_out_18_port, ALU_out_17_port, ALU_out_16_port, ALU_out_15_port, 
      ALU_out_14_port, ALU_out_13_port, ALU_out_12_port, ALU_out_11_port, 
      ALU_out_10_port, ALU_out_9_port, ALU_out_8_port, ALU_out_7_port, 
      ALU_out_6_port, ALU_out_5_port, ALU_out_4_port, ALU_out_3_port, 
      ALU_out_2_port, ALU_out_1_port, ALU_out_0_port, is_zero, cond, 
      ALU_ex_31_port, ALU_ex_30_port, ALU_ex_29_port, ALU_ex_28_port, 
      ALU_ex_27_port, ALU_ex_26_port, ALU_ex_25_port, ALU_ex_24_port, 
      ALU_ex_23_port, ALU_ex_22_port, ALU_ex_21_port, ALU_ex_20_port, 
      ALU_ex_19_port, ALU_ex_18_port, ALU_ex_17_port, ALU_ex_16_port, 
      ALU_ex_15_port, ALU_ex_14_port, ALU_ex_13_port, ALU_ex_12_port, 
      ALU_ex_11_port, ALU_ex_10_port, ALU_ex_9_port, ALU_ex_8_port, 
      ALU_ex_7_port, ALU_ex_6_port, ALU_ex_5_port, ALU_ex_4_port, ALU_ex_3_port
      , ALU_ex_2_port, ALU_ex_1_port, ALU_ex_0_port, signed_op_mem, 
      NPC_mem_31_port, NPC_mem_30_port, NPC_mem_29_port, NPC_mem_28_port, 
      NPC_mem_27_port, NPC_mem_26_port, NPC_mem_25_port, NPC_mem_24_port, 
      NPC_mem_23_port, NPC_mem_22_port, NPC_mem_21_port, NPC_mem_20_port, 
      NPC_mem_19_port, NPC_mem_18_port, NPC_mem_17_port, NPC_mem_16_port, 
      NPC_mem_15_port, NPC_mem_14_port, NPC_mem_13_port, NPC_mem_12_port, 
      NPC_mem_11_port, NPC_mem_10_port, NPC_mem_9_port, NPC_mem_8_port, 
      NPC_mem_7_port, NPC_mem_6_port, NPC_mem_5_port, NPC_mem_4_port, 
      NPC_mem_3_port, NPC_mem_2_port, NPC_mem_1_port, NPC_mem_0_port, cond_mem,
      regB_mem_31_port, regB_mem_30_port, regB_mem_29_port, regB_mem_28_port, 
      regB_mem_27_port, regB_mem_26_port, regB_mem_25_port, regB_mem_24_port, 
      regB_mem_23_port, regB_mem_22_port, regB_mem_21_port, regB_mem_20_port, 
      regB_mem_19_port, regB_mem_18_port, regB_mem_17_port, regB_mem_16_port, 
      regB_mem_15_port, regB_mem_14_port, regB_mem_13_port, regB_mem_12_port, 
      regB_mem_11_port, regB_mem_10_port, regB_mem_9_port, regB_mem_8_port, 
      regB_mem_7_port, regB_mem_6_port, regB_mem_5_port, regB_mem_4_port, 
      regB_mem_3_port, regB_mem_2_port, regB_mem_1_port, regB_mem_0_port, 
      RD_mem_4_port, RD_mem_3_port, RD_mem_2_port, RD_mem_1_port, RD_mem_0_port
      , wr_signal_mem, IR_26_mem_5_port, IR_26_mem_4_port, IR_26_mem_3_port, 
      IR_26_mem_2_port, IR_26_mem_1_port, IR_26_mem_0_port, sel_saved_reg, N14,
      wr_signal_mem1, LMD_out_31_port, LMD_out_30_port, LMD_out_29_port, 
      LMD_out_28_port, LMD_out_27_port, LMD_out_26_port, LMD_out_25_port, 
      LMD_out_24_port, LMD_out_23_port, LMD_out_22_port, LMD_out_21_port, 
      LMD_out_20_port, LMD_out_19_port, LMD_out_18_port, LMD_out_17_port, 
      LMD_out_16_port, LMD_out_15_port, LMD_out_14_port, LMD_out_13_port, 
      LMD_out_12_port, LMD_out_11_port, LMD_out_10_port, LMD_out_9_port, 
      LMD_out_8_port, LMD_out_7_port, LMD_out_6_port, LMD_out_5_port, 
      LMD_out_4_port, LMD_out_3_port, LMD_out_2_port, LMD_out_1_port, 
      LMD_out_0_port, ALU_wb_31_port, ALU_wb_30_port, ALU_wb_29_port, 
      ALU_wb_28_port, ALU_wb_27_port, ALU_wb_26_port, ALU_wb_25_port, 
      ALU_wb_24_port, ALU_wb_23_port, ALU_wb_22_port, ALU_wb_21_port, 
      ALU_wb_20_port, ALU_wb_19_port, ALU_wb_18_port, ALU_wb_17_port, 
      ALU_wb_16_port, ALU_wb_15_port, ALU_wb_14_port, ALU_wb_13_port, 
      ALU_wb_12_port, ALU_wb_11_port, ALU_wb_10_port, ALU_wb_9_port, 
      ALU_wb_8_port, ALU_wb_7_port, ALU_wb_6_port, ALU_wb_5_port, ALU_wb_4_port
      , ALU_wb_3_port, ALU_wb_2_port, ALU_wb_1_port, ALU_wb_0_port, 
      LMD_wb_31_port, LMD_wb_30_port, LMD_wb_29_port, LMD_wb_28_port, 
      LMD_wb_27_port, LMD_wb_26_port, LMD_wb_25_port, LMD_wb_24_port, 
      LMD_wb_23_port, LMD_wb_22_port, LMD_wb_21_port, LMD_wb_20_port, 
      LMD_wb_19_port, LMD_wb_18_port, LMD_wb_17_port, LMD_wb_16_port, 
      LMD_wb_15_port, LMD_wb_14_port, LMD_wb_13_port, LMD_wb_12_port, 
      LMD_wb_11_port, LMD_wb_10_port, LMD_wb_9_port, LMD_wb_8_port, 
      LMD_wb_7_port, LMD_wb_6_port, LMD_wb_5_port, LMD_wb_4_port, LMD_wb_3_port
      , LMD_wb_2_port, LMD_wb_1_port, LMD_wb_0_port, sel_saved_reg_wb, 
      NPC_wb_31_port, NPC_wb_30_port, NPC_wb_29_port, NPC_wb_28_port, 
      NPC_wb_27_port, NPC_wb_26_port, NPC_wb_25_port, NPC_wb_24_port, 
      NPC_wb_23_port, NPC_wb_22_port, NPC_wb_21_port, NPC_wb_20_port, 
      NPC_wb_19_port, NPC_wb_18_port, NPC_wb_17_port, NPC_wb_16_port, 
      NPC_wb_15_port, NPC_wb_14_port, NPC_wb_13_port, NPC_wb_12_port, 
      NPC_wb_11_port, NPC_wb_10_port, NPC_wb_9_port, NPC_wb_8_port, 
      NPC_wb_7_port, NPC_wb_6_port, NPC_wb_5_port, NPC_wb_4_port, NPC_wb_3_port
      , NPC_wb_2_port, NPC_wb_1_port, NPC_wb_0_port, n1, n2, n3, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14_port, n15, n16, n17, n18, n19, n20, n21
      , n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n_2244, n_2245, n_2246,
      n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, 
      n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, 
      n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, 
      n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, 
      n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, 
      n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, 
      n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308 : 
      std_logic;

begin
   DATA_MEM_RM <= RM;
   DATA_MEM_WM <= WM;
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   DATA_MEM_ADDR_reg_31_inst : DLH_X1 port map( G => N14, D => ALU_ex_31_port, 
                           Q => DATA_MEM_ADDR(31));
   DATA_MEM_ADDR_reg_30_inst : DLH_X1 port map( G => N14, D => ALU_ex_30_port, 
                           Q => DATA_MEM_ADDR(30));
   DATA_MEM_ADDR_reg_29_inst : DLH_X1 port map( G => N14, D => ALU_ex_29_port, 
                           Q => DATA_MEM_ADDR(29));
   DATA_MEM_ADDR_reg_28_inst : DLH_X1 port map( G => N14, D => ALU_ex_28_port, 
                           Q => DATA_MEM_ADDR(28));
   DATA_MEM_ADDR_reg_27_inst : DLH_X1 port map( G => N14, D => ALU_ex_27_port, 
                           Q => DATA_MEM_ADDR(27));
   DATA_MEM_ADDR_reg_26_inst : DLH_X1 port map( G => N14, D => ALU_ex_26_port, 
                           Q => DATA_MEM_ADDR(26));
   DATA_MEM_ADDR_reg_25_inst : DLH_X1 port map( G => N14, D => ALU_ex_25_port, 
                           Q => DATA_MEM_ADDR(25));
   DATA_MEM_ADDR_reg_24_inst : DLH_X1 port map( G => N14, D => ALU_ex_24_port, 
                           Q => DATA_MEM_ADDR(24));
   DATA_MEM_ADDR_reg_23_inst : DLH_X1 port map( G => N14, D => ALU_ex_23_port, 
                           Q => DATA_MEM_ADDR(23));
   DATA_MEM_ADDR_reg_22_inst : DLH_X1 port map( G => N14, D => ALU_ex_22_port, 
                           Q => DATA_MEM_ADDR(22));
   DATA_MEM_ADDR_reg_21_inst : DLH_X1 port map( G => N14, D => ALU_ex_21_port, 
                           Q => DATA_MEM_ADDR(21));
   DATA_MEM_ADDR_reg_20_inst : DLH_X1 port map( G => N14, D => ALU_ex_20_port, 
                           Q => DATA_MEM_ADDR(20));
   DATA_MEM_ADDR_reg_19_inst : DLH_X1 port map( G => N14, D => ALU_ex_19_port, 
                           Q => DATA_MEM_ADDR(19));
   DATA_MEM_ADDR_reg_18_inst : DLH_X1 port map( G => N14, D => ALU_ex_18_port, 
                           Q => DATA_MEM_ADDR(18));
   DATA_MEM_ADDR_reg_17_inst : DLH_X1 port map( G => N14, D => ALU_ex_17_port, 
                           Q => DATA_MEM_ADDR(17));
   DATA_MEM_ADDR_reg_16_inst : DLH_X1 port map( G => N14, D => ALU_ex_16_port, 
                           Q => DATA_MEM_ADDR(16));
   DATA_MEM_ADDR_reg_15_inst : DLH_X1 port map( G => N14, D => ALU_ex_15_port, 
                           Q => DATA_MEM_ADDR(15));
   DATA_MEM_ADDR_reg_14_inst : DLH_X1 port map( G => N14, D => ALU_ex_14_port, 
                           Q => DATA_MEM_ADDR(14));
   DATA_MEM_ADDR_reg_13_inst : DLH_X1 port map( G => N14, D => ALU_ex_13_port, 
                           Q => DATA_MEM_ADDR(13));
   DATA_MEM_ADDR_reg_12_inst : DLH_X1 port map( G => N14, D => ALU_ex_12_port, 
                           Q => DATA_MEM_ADDR(12));
   DATA_MEM_ADDR_reg_11_inst : DLH_X1 port map( G => N14, D => ALU_ex_11_port, 
                           Q => DATA_MEM_ADDR(11));
   DATA_MEM_ADDR_reg_10_inst : DLH_X1 port map( G => N14, D => ALU_ex_10_port, 
                           Q => DATA_MEM_ADDR(10));
   DATA_MEM_ADDR_reg_9_inst : DLH_X1 port map( G => N14, D => ALU_ex_9_port, Q 
                           => DATA_MEM_ADDR(9));
   DATA_MEM_ADDR_reg_8_inst : DLH_X1 port map( G => N14, D => ALU_ex_8_port, Q 
                           => DATA_MEM_ADDR(8));
   DATA_MEM_ADDR_reg_7_inst : DLH_X1 port map( G => N14, D => ALU_ex_7_port, Q 
                           => DATA_MEM_ADDR(7));
   DATA_MEM_ADDR_reg_6_inst : DLH_X1 port map( G => N14, D => ALU_ex_6_port, Q 
                           => DATA_MEM_ADDR(6));
   DATA_MEM_ADDR_reg_5_inst : DLH_X1 port map( G => N14, D => ALU_ex_5_port, Q 
                           => DATA_MEM_ADDR(5));
   DATA_MEM_ADDR_reg_4_inst : DLH_X1 port map( G => N14, D => ALU_ex_4_port, Q 
                           => DATA_MEM_ADDR(4));
   DATA_MEM_ADDR_reg_3_inst : DLH_X1 port map( G => N14, D => ALU_ex_3_port, Q 
                           => DATA_MEM_ADDR(3));
   DATA_MEM_ADDR_reg_2_inst : DLH_X1 port map( G => N14, D => ALU_ex_2_port, Q 
                           => DATA_MEM_ADDR(2));
   DATA_MEM_ADDR_reg_1_inst : DLH_X1 port map( G => N14, D => ALU_ex_1_port, Q 
                           => DATA_MEM_ADDR(1));
   DATA_MEM_ADDR_reg_0_inst : DLH_X1 port map( G => N14, D => ALU_ex_0_port, Q 
                           => DATA_MEM_ADDR(0));
   U3 : NOR2_X1 port map( A1 => n1, A2 => jump_en, ZN => wr_signal_mem1);
   U4 : INV_X1 port map( A => wr_signal_mem, ZN => n1);
   U5 : INV_X1 port map( A => n2, ZN => wr_signal);
   U6 : OAI33_X1 port map( A1 => n3, A2 => n42, A3 => n45, B1 => n4, B2 => n5, 
                           B3 => n6, ZN => n2);
   U7 : XOR2_X1 port map( A => IR_Dec_27_port, B => n40, Z => n6);
   U8 : INV_X1 port map( A => n42, ZN => n5);
   U9 : NAND3_X1 port map( A1 => n7, A2 => n8, A3 => n45, ZN => n4);
   U10 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n3);
   U11 : INV_X1 port map( A => IR_Dec_27_port, ZN => n10);
   U12 : OAI33_X1 port map( A1 => n8, A2 => n11, A3 => n7, B1 => n12, B2 => n13
                           , B3 => n14_port, ZN => n9);
   U13 : OR4_X1 port map( A1 => IR_Dec_11_port, A2 => IR_Dec_10_port, A3 => 
                           IR_Dec_0_port, A4 => n15, ZN => n14_port);
   U14 : OR4_X1 port map( A1 => IR_Dec_13_port, A2 => IR_Dec_12_port, A3 => 
                           IR_Dec_15_port, A4 => IR_Dec_14_port, ZN => n15);
   U15 : OR4_X1 port map( A1 => IR_Dec_18_port, A2 => IR_Dec_17_port, A3 => 
                           IR_Dec_16_port, A4 => n16, ZN => n13);
   U16 : OR4_X1 port map( A1 => IR_Dec_1_port, A2 => IR_Dec_19_port, A3 => 
                           IR_Dec_21_port, A4 => IR_Dec_20_port, ZN => n16);
   U17 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           n12);
   U18 : NOR4_X1 port map( A1 => IR_Dec_9_port, A2 => IR_Dec_8_port, A3 => 
                           IR_Dec_7_port, A4 => IR_Dec_6_port, ZN => n20);
   U19 : NOR4_X1 port map( A1 => IR_Dec_5_port, A2 => IR_Dec_4_port, A3 => 
                           IR_Dec_3_port, A4 => n43, ZN => n19);
   U20 : NOR4_X1 port map( A1 => IR_Dec_2_port, A2 => IR_Dec_28_port, A3 => 
                           IR_Dec_26_port, A4 => IR_Dec_25_port, ZN => n18);
   U21 : NOR3_X1 port map( A1 => IR_Dec_22_port, A2 => IR_Dec_24_port, A3 => 
                           IR_Dec_23_port, ZN => n17);
   U22 : INV_X1 port map( A => IR_Dec_28_port, ZN => n7);
   U23 : INV_X1 port map( A => n40, ZN => n11);
   U24 : INV_X1 port map( A => n41, ZN => n8);
   U25 : AND2_X1 port map( A1 => IR_26_mem_0_port, A2 => jump_en, ZN => 
                           sel_saved_reg);
   U26 : OR2_X1 port map( A1 => cond_mem, A2 => jump_en, ZN => sel_npc);
   U27 : NAND4_X1 port map( A1 => IR_26_mem_2_port, A2 => IR_26_mem_0_port, A3 
                           => IR_26_mem_4_port, A4 => n21, ZN => N14);
   U28 : NOR3_X1 port map( A1 => IR_26_mem_1_port, A2 => IR_26_mem_5_port, A3 
                           => IR_26_mem_3_port, ZN => n21);
   U29 : AND2_X1 port map( A1 => regB_mem_9_port, A2 => n22, ZN => 
                           DATA_MEM_IN(9));
   U30 : AND2_X1 port map( A1 => regB_mem_8_port, A2 => n22, ZN => 
                           DATA_MEM_IN(8));
   U31 : INV_X1 port map( A => n23, ZN => DATA_MEM_IN(7));
   U32 : AOI22_X1 port map( A1 => n22, A2 => regB_mem_7_port, B1 => 
                           regB_mem_31_port, B2 => sb_op, ZN => n23);
   U33 : INV_X1 port map( A => n24, ZN => DATA_MEM_IN(6));
   U34 : AOI22_X1 port map( A1 => n22, A2 => regB_mem_6_port, B1 => sb_op, B2 
                           => regB_mem_30_port, ZN => n24);
   U35 : INV_X1 port map( A => n25, ZN => DATA_MEM_IN(5));
   U36 : AOI22_X1 port map( A1 => n22, A2 => regB_mem_5_port, B1 => sb_op, B2 
                           => regB_mem_29_port, ZN => n25);
   U37 : INV_X1 port map( A => n26, ZN => DATA_MEM_IN(4));
   U38 : AOI22_X1 port map( A1 => n22, A2 => regB_mem_4_port, B1 => sb_op, B2 
                           => regB_mem_28_port, ZN => n26);
   U39 : INV_X1 port map( A => n27, ZN => DATA_MEM_IN(3));
   U40 : AOI22_X1 port map( A1 => n22, A2 => regB_mem_3_port, B1 => sb_op, B2 
                           => regB_mem_27_port, ZN => n27);
   U41 : AND2_X1 port map( A1 => n22, A2 => regB_mem_31_port, ZN => 
                           DATA_MEM_IN(31));
   U42 : AND2_X1 port map( A1 => n22, A2 => regB_mem_30_port, ZN => 
                           DATA_MEM_IN(30));
   U43 : INV_X1 port map( A => n28, ZN => DATA_MEM_IN(2));
   U44 : AOI22_X1 port map( A1 => n22, A2 => regB_mem_2_port, B1 => sb_op, B2 
                           => regB_mem_26_port, ZN => n28);
   U45 : AND2_X1 port map( A1 => n22, A2 => regB_mem_29_port, ZN => 
                           DATA_MEM_IN(29));
   U46 : AND2_X1 port map( A1 => n22, A2 => regB_mem_28_port, ZN => 
                           DATA_MEM_IN(28));
   U47 : AND2_X1 port map( A1 => n22, A2 => regB_mem_27_port, ZN => 
                           DATA_MEM_IN(27));
   U48 : AND2_X1 port map( A1 => n22, A2 => regB_mem_26_port, ZN => 
                           DATA_MEM_IN(26));
   U49 : AND2_X1 port map( A1 => n22, A2 => regB_mem_25_port, ZN => 
                           DATA_MEM_IN(25));
   U50 : AND2_X1 port map( A1 => n22, A2 => regB_mem_24_port, ZN => 
                           DATA_MEM_IN(24));
   U51 : AND2_X1 port map( A1 => regB_mem_23_port, A2 => n22, ZN => 
                           DATA_MEM_IN(23));
   U52 : AND2_X1 port map( A1 => regB_mem_22_port, A2 => n22, ZN => 
                           DATA_MEM_IN(22));
   U53 : AND2_X1 port map( A1 => regB_mem_21_port, A2 => n22, ZN => 
                           DATA_MEM_IN(21));
   U54 : AND2_X1 port map( A1 => regB_mem_20_port, A2 => n22, ZN => 
                           DATA_MEM_IN(20));
   U55 : INV_X1 port map( A => n29, ZN => DATA_MEM_IN(1));
   U56 : AOI22_X1 port map( A1 => sb_op, A2 => regB_mem_25_port, B1 => n22, B2 
                           => regB_mem_1_port, ZN => n29);
   U57 : AND2_X1 port map( A1 => regB_mem_19_port, A2 => n22, ZN => 
                           DATA_MEM_IN(19));
   U58 : AND2_X1 port map( A1 => regB_mem_18_port, A2 => n22, ZN => 
                           DATA_MEM_IN(18));
   U59 : AND2_X1 port map( A1 => regB_mem_17_port, A2 => n22, ZN => 
                           DATA_MEM_IN(17));
   U60 : AND2_X1 port map( A1 => regB_mem_16_port, A2 => n22, ZN => 
                           DATA_MEM_IN(16));
   U61 : AND2_X1 port map( A1 => regB_mem_15_port, A2 => n22, ZN => 
                           DATA_MEM_IN(15));
   U62 : AND2_X1 port map( A1 => regB_mem_14_port, A2 => n22, ZN => 
                           DATA_MEM_IN(14));
   U63 : AND2_X1 port map( A1 => regB_mem_13_port, A2 => n22, ZN => 
                           DATA_MEM_IN(13));
   U64 : AND2_X1 port map( A1 => regB_mem_12_port, A2 => n22, ZN => 
                           DATA_MEM_IN(12));
   U65 : AND2_X1 port map( A1 => regB_mem_11_port, A2 => n22, ZN => 
                           DATA_MEM_IN(11));
   U66 : AND2_X1 port map( A1 => regB_mem_10_port, A2 => n22, ZN => 
                           DATA_MEM_IN(10));
   U67 : INV_X1 port map( A => n30, ZN => DATA_MEM_IN(0));
   U68 : AOI22_X1 port map( A1 => sb_op, A2 => regB_mem_24_port, B1 => n22, B2 
                           => regB_mem_0_port, ZN => n30);
   U69 : INV_X1 port map( A => sb_op, ZN => n22);
   U70 : OR4_X1 port map( A1 => n31, A2 => n32, A3 => WM, A4 => RM, ZN => 
                           DATA_MEM_ENABLE);
   U71 : NOR4_X1 port map( A1 => instruction_alu(1), A2 => n33, A3 => n34, A4 
                           => n35, ZN => n32);
   U72 : INV_X1 port map( A => instruction_alu(0), ZN => n35);
   U73 : INV_X1 port map( A => instruction_alu(2), ZN => n34);
   U74 : AOI22_X1 port map( A1 => n36, A2 => instruction_alu(4), B1 => 
                           instruction_alu(3), B2 => n37, ZN => n33);
   U75 : INV_X1 port map( A => instruction_alu(4), ZN => n37);
   U76 : NOR2_X1 port map( A1 => instruction_alu(3), A2 => n38, ZN => n36);
   U77 : NOR4_X1 port map( A1 => n39, A2 => n38, A3 => instruction_alu(0), A4 
                           => instruction_alu(2), ZN => n31);
   U78 : INV_X1 port map( A => instruction_alu(5), ZN => n38);
   U79 : NAND3_X1 port map( A1 => instruction_alu(3), A2 => instruction_alu(4),
                           A3 => instruction_alu(1), ZN => n39);
   pipeline_PCING : regFFD_NBIT32_0 port map( CK => CLK, RESET => RST, ENABLE 
                           => X_Logic1_port, D(31) => PC(31), D(30) => PC(30), 
                           D(29) => PC(29), D(28) => PC(28), D(27) => PC(27), 
                           D(26) => PC(26), D(25) => PC(25), D(24) => PC(24), 
                           D(23) => PC(23), D(22) => PC(22), D(21) => PC(21), 
                           D(20) => PC(20), D(19) => PC(19), D(18) => PC(18), 
                           D(17) => PC(17), D(16) => PC(16), D(15) => PC(15), 
                           D(14) => PC(14), D(13) => PC(13), D(12) => PC(12), 
                           D(11) => PC(11), D(10) => PC(10), D(9) => PC(9), 
                           D(8) => PC(8), D(7) => PC(7), D(6) => PC(6), D(5) =>
                           PC(5), D(4) => PC(4), D(3) => PC(3), D(2) => PC(2), 
                           D(1) => PC(1), D(0) => PC(0), Q(31) => 
                           PC_fetch0_31_port, Q(30) => PC_fetch0_30_port, Q(29)
                           => PC_fetch0_29_port, Q(28) => PC_fetch0_28_port, 
                           Q(27) => PC_fetch0_27_port, Q(26) => 
                           PC_fetch0_26_port, Q(25) => PC_fetch0_25_port, Q(24)
                           => PC_fetch0_24_port, Q(23) => PC_fetch0_23_port, 
                           Q(22) => PC_fetch0_22_port, Q(21) => 
                           PC_fetch0_21_port, Q(20) => PC_fetch0_20_port, Q(19)
                           => PC_fetch0_19_port, Q(18) => PC_fetch0_18_port, 
                           Q(17) => PC_fetch0_17_port, Q(16) => 
                           PC_fetch0_16_port, Q(15) => PC_fetch0_15_port, Q(14)
                           => PC_fetch0_14_port, Q(13) => PC_fetch0_13_port, 
                           Q(12) => PC_fetch0_12_port, Q(11) => 
                           PC_fetch0_11_port, Q(10) => PC_fetch0_10_port, Q(9) 
                           => PC_fetch0_9_port, Q(8) => PC_fetch0_8_port, Q(7) 
                           => PC_fetch0_7_port, Q(6) => PC_fetch0_6_port, Q(5) 
                           => PC_fetch0_5_port, Q(4) => PC_fetch0_4_port, Q(3) 
                           => PC_fetch0_3_port, Q(2) => PC_fetch0_2_port, Q(1) 
                           => PC_fetch0_1_port, Q(0) => PC_fetch0_0_port);
   pipeline_fetch1_NPC : regFFD_NBIT32_18 port map( CK => CLK, RESET => RST, 
                           ENABLE => NPC_LATCH_EN, D(31) => NPC_31_port, D(30) 
                           => NPC_30_port, D(29) => NPC_29_port, D(28) => 
                           NPC_28_port, D(27) => NPC_27_port, D(26) => 
                           NPC_26_port, D(25) => NPC_25_port, D(24) => 
                           NPC_24_port, D(23) => NPC_23_port, D(22) => 
                           NPC_22_port, D(21) => NPC_21_port, D(20) => 
                           NPC_20_port, D(19) => NPC_19_port, D(18) => 
                           NPC_18_port, D(17) => NPC_17_port, D(16) => 
                           NPC_16_port, D(15) => NPC_15_port, D(14) => 
                           NPC_14_port, D(13) => NPC_13_port, D(12) => 
                           NPC_12_port, D(11) => NPC_11_port, D(10) => 
                           NPC_10_port, D(9) => NPC_9_port, D(8) => NPC_8_port,
                           D(7) => NPC_7_port, D(6) => NPC_6_port, D(5) => 
                           NPC_5_port, D(4) => NPC_4_port, D(3) => NPC_3_port, 
                           D(2) => NPC_2_port, D(1) => NPC_1_port, D(0) => 
                           NPC_0_port, Q(31) => NPC_fetch1_31_port, Q(30) => 
                           NPC_fetch1_30_port, Q(29) => NPC_fetch1_29_port, 
                           Q(28) => NPC_fetch1_28_port, Q(27) => 
                           NPC_fetch1_27_port, Q(26) => NPC_fetch1_26_port, 
                           Q(25) => NPC_fetch1_25_port, Q(24) => 
                           NPC_fetch1_24_port, Q(23) => NPC_fetch1_23_port, 
                           Q(22) => NPC_fetch1_22_port, Q(21) => 
                           NPC_fetch1_21_port, Q(20) => NPC_fetch1_20_port, 
                           Q(19) => NPC_fetch1_19_port, Q(18) => 
                           NPC_fetch1_18_port, Q(17) => NPC_fetch1_17_port, 
                           Q(16) => NPC_fetch1_16_port, Q(15) => 
                           NPC_fetch1_15_port, Q(14) => NPC_fetch1_14_port, 
                           Q(13) => NPC_fetch1_13_port, Q(12) => 
                           NPC_fetch1_12_port, Q(11) => NPC_fetch1_11_port, 
                           Q(10) => NPC_fetch1_10_port, Q(9) => 
                           NPC_fetch1_9_port, Q(8) => NPC_fetch1_8_port, Q(7) 
                           => NPC_fetch1_7_port, Q(6) => NPC_fetch1_6_port, 
                           Q(5) => NPC_fetch1_5_port, Q(4) => NPC_fetch1_4_port
                           , Q(3) => NPC_fetch1_3_port, Q(2) => 
                           NPC_fetch1_2_port, Q(1) => NPC_fetch1_1_port, Q(0) 
                           => NPC_fetch1_0_port);
   pipeline_fetch1_PC : regFFD_NBIT32_17 port map( CK => CLK, RESET => RST, 
                           ENABLE => ir_LATCH_EN, D(31) => PC_fetch0_31_port, 
                           D(30) => PC_fetch0_30_port, D(29) => 
                           PC_fetch0_29_port, D(28) => PC_fetch0_28_port, D(27)
                           => PC_fetch0_27_port, D(26) => PC_fetch0_26_port, 
                           D(25) => PC_fetch0_25_port, D(24) => 
                           PC_fetch0_24_port, D(23) => PC_fetch0_23_port, D(22)
                           => PC_fetch0_22_port, D(21) => PC_fetch0_21_port, 
                           D(20) => PC_fetch0_20_port, D(19) => 
                           PC_fetch0_19_port, D(18) => PC_fetch0_18_port, D(17)
                           => PC_fetch0_17_port, D(16) => PC_fetch0_16_port, 
                           D(15) => PC_fetch0_15_port, D(14) => 
                           PC_fetch0_14_port, D(13) => PC_fetch0_13_port, D(12)
                           => PC_fetch0_12_port, D(11) => PC_fetch0_11_port, 
                           D(10) => PC_fetch0_10_port, D(9) => PC_fetch0_9_port
                           , D(8) => PC_fetch0_8_port, D(7) => PC_fetch0_7_port
                           , D(6) => PC_fetch0_6_port, D(5) => PC_fetch0_5_port
                           , D(4) => PC_fetch0_4_port, D(3) => PC_fetch0_3_port
                           , D(2) => PC_fetch0_2_port, D(1) => PC_fetch0_1_port
                           , D(0) => PC_fetch0_0_port, Q(31) => 
                           PC_fetch1_31_port, Q(30) => PC_fetch1_30_port, Q(29)
                           => PC_fetch1_29_port, Q(28) => PC_fetch1_28_port, 
                           Q(27) => PC_fetch1_27_port, Q(26) => 
                           PC_fetch1_26_port, Q(25) => PC_fetch1_25_port, Q(24)
                           => PC_fetch1_24_port, Q(23) => PC_fetch1_23_port, 
                           Q(22) => PC_fetch1_22_port, Q(21) => 
                           PC_fetch1_21_port, Q(20) => PC_fetch1_20_port, Q(19)
                           => PC_fetch1_19_port, Q(18) => PC_fetch1_18_port, 
                           Q(17) => PC_fetch1_17_port, Q(16) => 
                           PC_fetch1_16_port, Q(15) => PC_fetch1_15_port, Q(14)
                           => PC_fetch1_14_port, Q(13) => PC_fetch1_13_port, 
                           Q(12) => PC_fetch1_12_port, Q(11) => 
                           PC_fetch1_11_port, Q(10) => PC_fetch1_10_port, Q(9) 
                           => PC_fetch1_9_port, Q(8) => PC_fetch1_8_port, Q(7) 
                           => PC_fetch1_7_port, Q(6) => PC_fetch1_6_port, Q(5) 
                           => PC_fetch1_5_port, Q(4) => PC_fetch1_4_port, Q(3) 
                           => PC_fetch1_3_port, Q(2) => PC_fetch1_2_port, Q(1) 
                           => PC_fetch1_1_port, Q(0) => PC_fetch1_0_port);
   MUX_PC1 : MUX21_GENERIC_NBIT32_0 port map( A(31) => PC_OUT_i_31_port, A(30) 
                           => PC_OUT_i_30_port, A(29) => PC_OUT_i_29_port, 
                           A(28) => PC_OUT_i_28_port, A(27) => PC_OUT_i_27_port
                           , A(26) => PC_OUT_i_26_port, A(25) => 
                           PC_OUT_i_25_port, A(24) => PC_OUT_i_24_port, A(23) 
                           => PC_OUT_i_23_port, A(22) => PC_OUT_i_22_port, 
                           A(21) => PC_OUT_i_21_port, A(20) => PC_OUT_i_20_port
                           , A(19) => PC_OUT_i_19_port, A(18) => 
                           PC_OUT_i_18_port, A(17) => PC_OUT_i_17_port, A(16) 
                           => PC_OUT_i_16_port, A(15) => PC_OUT_i_15_port, 
                           A(14) => PC_OUT_i_14_port, A(13) => PC_OUT_i_13_port
                           , A(12) => PC_OUT_i_12_port, A(11) => 
                           PC_OUT_i_11_port, A(10) => PC_OUT_i_10_port, A(9) =>
                           PC_OUT_i_9_port, A(8) => PC_OUT_i_8_port, A(7) => 
                           PC_OUT_i_7_port, A(6) => PC_OUT_i_6_port, A(5) => 
                           PC_OUT_i_5_port, A(4) => PC_OUT_i_4_port, A(3) => 
                           PC_OUT_i_3_port, A(2) => PC_OUT_i_2_port, A(1) => 
                           PC_OUT_i_1_port, A(0) => PC_OUT_i_0_port, B(31) => 
                           NPC_fetch1_31_port, B(30) => NPC_fetch1_30_port, 
                           B(29) => NPC_fetch1_29_port, B(28) => 
                           NPC_fetch1_28_port, B(27) => NPC_fetch1_27_port, 
                           B(26) => NPC_fetch1_26_port, B(25) => 
                           NPC_fetch1_25_port, B(24) => NPC_fetch1_24_port, 
                           B(23) => NPC_fetch1_23_port, B(22) => 
                           NPC_fetch1_22_port, B(21) => NPC_fetch1_21_port, 
                           B(20) => NPC_fetch1_20_port, B(19) => 
                           NPC_fetch1_19_port, B(18) => NPC_fetch1_18_port, 
                           B(17) => NPC_fetch1_17_port, B(16) => 
                           NPC_fetch1_16_port, B(15) => NPC_fetch1_15_port, 
                           B(14) => NPC_fetch1_14_port, B(13) => 
                           NPC_fetch1_13_port, B(12) => NPC_fetch1_12_port, 
                           B(11) => NPC_fetch1_11_port, B(10) => 
                           NPC_fetch1_10_port, B(9) => NPC_fetch1_9_port, B(8) 
                           => NPC_fetch1_8_port, B(7) => NPC_fetch1_7_port, 
                           B(6) => NPC_fetch1_6_port, B(5) => NPC_fetch1_5_port
                           , B(4) => NPC_fetch1_4_port, B(3) => 
                           NPC_fetch1_3_port, B(2) => NPC_fetch1_2_port, B(1) 
                           => NPC_fetch1_1_port, B(0) => NPC_fetch1_0_port, SEL
                           => sel_npc, Y(31) => PC_OUT(31), Y(30) => PC_OUT(30)
                           , Y(29) => PC_OUT(29), Y(28) => PC_OUT(28), Y(27) =>
                           PC_OUT(27), Y(26) => PC_OUT(26), Y(25) => PC_OUT(25)
                           , Y(24) => PC_OUT(24), Y(23) => PC_OUT(23), Y(22) =>
                           PC_OUT(22), Y(21) => PC_OUT(21), Y(20) => PC_OUT(20)
                           , Y(19) => PC_OUT(19), Y(18) => PC_OUT(18), Y(17) =>
                           PC_OUT(17), Y(16) => PC_OUT(16), Y(15) => PC_OUT(15)
                           , Y(14) => PC_OUT(14), Y(13) => PC_OUT(13), Y(12) =>
                           PC_OUT(12), Y(11) => PC_OUT(11), Y(10) => PC_OUT(10)
                           , Y(9) => PC_OUT(9), Y(8) => PC_OUT(8), Y(7) => 
                           PC_OUT(7), Y(6) => PC_OUT(6), Y(5) => PC_OUT(5), 
                           Y(4) => PC_OUT(4), Y(3) => PC_OUT(3), Y(2) => 
                           PC_OUT(2), Y(1) => PC_OUT(1), Y(0) => PC_OUT(0));
   pipeline_fetch_NPC : regFFD_NBIT32_16 port map( CK => CLK, RESET => RST, 
                           ENABLE => NPC_LATCH_EN, D(31) => NPC_fetch1_31_port,
                           D(30) => NPC_fetch1_30_port, D(29) => 
                           NPC_fetch1_29_port, D(28) => NPC_fetch1_28_port, 
                           D(27) => NPC_fetch1_27_port, D(26) => 
                           NPC_fetch1_26_port, D(25) => NPC_fetch1_25_port, 
                           D(24) => NPC_fetch1_24_port, D(23) => 
                           NPC_fetch1_23_port, D(22) => NPC_fetch1_22_port, 
                           D(21) => NPC_fetch1_21_port, D(20) => 
                           NPC_fetch1_20_port, D(19) => NPC_fetch1_19_port, 
                           D(18) => NPC_fetch1_18_port, D(17) => 
                           NPC_fetch1_17_port, D(16) => NPC_fetch1_16_port, 
                           D(15) => NPC_fetch1_15_port, D(14) => 
                           NPC_fetch1_14_port, D(13) => NPC_fetch1_13_port, 
                           D(12) => NPC_fetch1_12_port, D(11) => 
                           NPC_fetch1_11_port, D(10) => NPC_fetch1_10_port, 
                           D(9) => NPC_fetch1_9_port, D(8) => NPC_fetch1_8_port
                           , D(7) => NPC_fetch1_7_port, D(6) => 
                           NPC_fetch1_6_port, D(5) => NPC_fetch1_5_port, D(4) 
                           => NPC_fetch1_4_port, D(3) => NPC_fetch1_3_port, 
                           D(2) => NPC_fetch1_2_port, D(1) => NPC_fetch1_1_port
                           , D(0) => NPC_fetch1_0_port, Q(31) => 
                           NPC_fetch_31_port, Q(30) => NPC_fetch_30_port, Q(29)
                           => NPC_fetch_29_port, Q(28) => NPC_fetch_28_port, 
                           Q(27) => NPC_fetch_27_port, Q(26) => 
                           NPC_fetch_26_port, Q(25) => NPC_fetch_25_port, Q(24)
                           => NPC_fetch_24_port, Q(23) => NPC_fetch_23_port, 
                           Q(22) => NPC_fetch_22_port, Q(21) => 
                           NPC_fetch_21_port, Q(20) => NPC_fetch_20_port, Q(19)
                           => NPC_fetch_19_port, Q(18) => NPC_fetch_18_port, 
                           Q(17) => NPC_fetch_17_port, Q(16) => 
                           NPC_fetch_16_port, Q(15) => NPC_fetch_15_port, Q(14)
                           => NPC_fetch_14_port, Q(13) => NPC_fetch_13_port, 
                           Q(12) => NPC_fetch_12_port, Q(11) => 
                           NPC_fetch_11_port, Q(10) => NPC_fetch_10_port, Q(9) 
                           => NPC_fetch_9_port, Q(8) => NPC_fetch_8_port, Q(7) 
                           => NPC_fetch_7_port, Q(6) => NPC_fetch_6_port, Q(5) 
                           => NPC_fetch_5_port, Q(4) => NPC_fetch_4_port, Q(3) 
                           => NPC_fetch_3_port, Q(2) => NPC_fetch_2_port, Q(1) 
                           => NPC_fetch_1_port, Q(0) => NPC_fetch_0_port);
   pipeline_fetch_PC : regFFD_NBIT32_15 port map( CK => CLK, RESET => RST, 
                           ENABLE => ir_LATCH_EN, D(31) => PC_fetch1_31_port, 
                           D(30) => PC_fetch1_30_port, D(29) => 
                           PC_fetch1_29_port, D(28) => PC_fetch1_28_port, D(27)
                           => PC_fetch1_27_port, D(26) => PC_fetch1_26_port, 
                           D(25) => PC_fetch1_25_port, D(24) => 
                           PC_fetch1_24_port, D(23) => PC_fetch1_23_port, D(22)
                           => PC_fetch1_22_port, D(21) => PC_fetch1_21_port, 
                           D(20) => PC_fetch1_20_port, D(19) => 
                           PC_fetch1_19_port, D(18) => PC_fetch1_18_port, D(17)
                           => PC_fetch1_17_port, D(16) => PC_fetch1_16_port, 
                           D(15) => PC_fetch1_15_port, D(14) => 
                           PC_fetch1_14_port, D(13) => PC_fetch1_13_port, D(12)
                           => PC_fetch1_12_port, D(11) => PC_fetch1_11_port, 
                           D(10) => PC_fetch1_10_port, D(9) => PC_fetch1_9_port
                           , D(8) => PC_fetch1_8_port, D(7) => PC_fetch1_7_port
                           , D(6) => PC_fetch1_6_port, D(5) => PC_fetch1_5_port
                           , D(4) => PC_fetch1_4_port, D(3) => PC_fetch1_3_port
                           , D(2) => PC_fetch1_2_port, D(1) => PC_fetch1_1_port
                           , D(0) => PC_fetch1_0_port, Q(31) => 
                           PC_fetch_31_port, Q(30) => PC_fetch_30_port, Q(29) 
                           => PC_fetch_29_port, Q(28) => PC_fetch_28_port, 
                           Q(27) => PC_fetch_27_port, Q(26) => PC_fetch_26_port
                           , Q(25) => PC_fetch_25_port, Q(24) => 
                           PC_fetch_24_port, Q(23) => PC_fetch_23_port, Q(22) 
                           => PC_fetch_22_port, Q(21) => PC_fetch_21_port, 
                           Q(20) => PC_fetch_20_port, Q(19) => PC_fetch_19_port
                           , Q(18) => PC_fetch_18_port, Q(17) => 
                           PC_fetch_17_port, Q(16) => PC_fetch_16_port, Q(15) 
                           => PC_fetch_15_port, Q(14) => PC_fetch_14_port, 
                           Q(13) => PC_fetch_13_port, Q(12) => PC_fetch_12_port
                           , Q(11) => PC_fetch_11_port, Q(10) => 
                           PC_fetch_10_port, Q(9) => PC_fetch_9_port, Q(8) => 
                           PC_fetch_8_port, Q(7) => PC_fetch_7_port, Q(6) => 
                           PC_fetch_6_port, Q(5) => PC_fetch_5_port, Q(4) => 
                           PC_fetch_4_port, Q(3) => PC_fetch_3_port, Q(2) => 
                           PC_fetch_2_port, Q(1) => PC_fetch_1_port, Q(0) => 
                           PC_fetch_0_port);
   pipeline_fetch_ir : regFFD_NBIT32_14 port map( CK => CLK, RESET => RST, 
                           ENABLE => ir_LATCH_EN, D(31) => IR(31), D(30) => 
                           IR(30), D(29) => IR(29), D(28) => IR(28), D(27) => 
                           IR(27), D(26) => IR(26), D(25) => IR(25), D(24) => 
                           IR(24), D(23) => IR(23), D(22) => IR(22), D(21) => 
                           IR(21), D(20) => IR(20), D(19) => IR(19), D(18) => 
                           IR(18), D(17) => IR(17), D(16) => IR(16), D(15) => 
                           IR(15), D(14) => IR(14), D(13) => IR(13), D(12) => 
                           IR(12), D(11) => IR(11), D(10) => IR(10), D(9) => 
                           IR(9), D(8) => IR(8), D(7) => IR(7), D(6) => IR(6), 
                           D(5) => IR(5), D(4) => IR(4), D(3) => IR(3), D(2) =>
                           IR(2), D(1) => IR(1), D(0) => IR(0), Q(31) => 
                           ir_fetch_31_port, Q(30) => ir_fetch_30_port, Q(29) 
                           => ir_fetch_29_port, Q(28) => ir_fetch_28_port, 
                           Q(27) => ir_fetch_27_port, Q(26) => ir_fetch_26_port
                           , Q(25) => ir_fetch_25_port, Q(24) => 
                           ir_fetch_24_port, Q(23) => ir_fetch_23_port, Q(22) 
                           => ir_fetch_22_port, Q(21) => ir_fetch_21_port, 
                           Q(20) => ir_fetch_20_port, Q(19) => ir_fetch_19_port
                           , Q(18) => ir_fetch_18_port, Q(17) => 
                           ir_fetch_17_port, Q(16) => ir_fetch_16_port, Q(15) 
                           => ir_fetch_15_port, Q(14) => ir_fetch_14_port, 
                           Q(13) => ir_fetch_13_port, Q(12) => ir_fetch_12_port
                           , Q(11) => ir_fetch_11_port, Q(10) => 
                           ir_fetch_10_port, Q(9) => ir_fetch_9_port, Q(8) => 
                           ir_fetch_8_port, Q(7) => ir_fetch_7_port, Q(6) => 
                           ir_fetch_6_port, Q(5) => ir_fetch_5_port, Q(4) => 
                           ir_fetch_4_port, Q(3) => ir_fetch_3_port, Q(2) => 
                           ir_fetch_2_port, Q(1) => ir_fetch_1_port, Q(0) => 
                           ir_fetch_0_port);
   pipeline_newpc1 : regFFD_NBIT32_13 port map( CK => CLK, RESET => RST, ENABLE
                           => NPC_LATCH_EN, D(31) => NPC_fetch_31_port, D(30) 
                           => NPC_fetch_30_port, D(29) => NPC_fetch_29_port, 
                           D(28) => NPC_fetch_28_port, D(27) => 
                           NPC_fetch_27_port, D(26) => NPC_fetch_26_port, D(25)
                           => NPC_fetch_25_port, D(24) => NPC_fetch_24_port, 
                           D(23) => NPC_fetch_23_port, D(22) => 
                           NPC_fetch_22_port, D(21) => NPC_fetch_21_port, D(20)
                           => NPC_fetch_20_port, D(19) => NPC_fetch_19_port, 
                           D(18) => NPC_fetch_18_port, D(17) => 
                           NPC_fetch_17_port, D(16) => NPC_fetch_16_port, D(15)
                           => NPC_fetch_15_port, D(14) => NPC_fetch_14_port, 
                           D(13) => NPC_fetch_13_port, D(12) => 
                           NPC_fetch_12_port, D(11) => NPC_fetch_11_port, D(10)
                           => NPC_fetch_10_port, D(9) => NPC_fetch_9_port, D(8)
                           => NPC_fetch_8_port, D(7) => NPC_fetch_7_port, D(6) 
                           => NPC_fetch_6_port, D(5) => NPC_fetch_5_port, D(4) 
                           => NPC_fetch_4_port, D(3) => NPC_fetch_3_port, D(2) 
                           => NPC_fetch_2_port, D(1) => NPC_fetch_1_port, D(0) 
                           => NPC_fetch_0_port, Q(31) => NPC_Dec_31_port, Q(30)
                           => NPC_Dec_30_port, Q(29) => NPC_Dec_29_port, Q(28) 
                           => NPC_Dec_28_port, Q(27) => NPC_Dec_27_port, Q(26) 
                           => NPC_Dec_26_port, Q(25) => NPC_Dec_25_port, Q(24) 
                           => NPC_Dec_24_port, Q(23) => NPC_Dec_23_port, Q(22) 
                           => NPC_Dec_22_port, Q(21) => NPC_Dec_21_port, Q(20) 
                           => NPC_Dec_20_port, Q(19) => NPC_Dec_19_port, Q(18) 
                           => NPC_Dec_18_port, Q(17) => NPC_Dec_17_port, Q(16) 
                           => NPC_Dec_16_port, Q(15) => NPC_Dec_15_port, Q(14) 
                           => NPC_Dec_14_port, Q(13) => NPC_Dec_13_port, Q(12) 
                           => NPC_Dec_12_port, Q(11) => NPC_Dec_11_port, Q(10) 
                           => NPC_Dec_10_port, Q(9) => NPC_Dec_9_port, Q(8) => 
                           NPC_Dec_8_port, Q(7) => NPC_Dec_7_port, Q(6) => 
                           NPC_Dec_6_port, Q(5) => NPC_Dec_5_port, Q(4) => 
                           NPC_Dec_4_port, Q(3) => NPC_Dec_3_port, Q(2) => 
                           NPC_Dec_2_port, Q(1) => NPC_Dec_1_port, Q(0) => 
                           NPC_Dec_0_port);
   pipeline_pc1 : regFFD_NBIT32_12 port map( CK => CLK, RESET => RST, ENABLE =>
                           ir_LATCH_EN, D(31) => PC_fetch_31_port, D(30) => 
                           PC_fetch_30_port, D(29) => PC_fetch_29_port, D(28) 
                           => PC_fetch_28_port, D(27) => PC_fetch_27_port, 
                           D(26) => PC_fetch_26_port, D(25) => PC_fetch_25_port
                           , D(24) => PC_fetch_24_port, D(23) => 
                           PC_fetch_23_port, D(22) => PC_fetch_22_port, D(21) 
                           => PC_fetch_21_port, D(20) => PC_fetch_20_port, 
                           D(19) => PC_fetch_19_port, D(18) => PC_fetch_18_port
                           , D(17) => PC_fetch_17_port, D(16) => 
                           PC_fetch_16_port, D(15) => PC_fetch_15_port, D(14) 
                           => PC_fetch_14_port, D(13) => PC_fetch_13_port, 
                           D(12) => PC_fetch_12_port, D(11) => PC_fetch_11_port
                           , D(10) => PC_fetch_10_port, D(9) => PC_fetch_9_port
                           , D(8) => PC_fetch_8_port, D(7) => PC_fetch_7_port, 
                           D(6) => PC_fetch_6_port, D(5) => PC_fetch_5_port, 
                           D(4) => PC_fetch_4_port, D(3) => PC_fetch_3_port, 
                           D(2) => PC_fetch_2_port, D(1) => PC_fetch_1_port, 
                           D(0) => PC_fetch_0_port, Q(31) => n_2244, Q(30) => 
                           n_2245, Q(29) => n_2246, Q(28) => n_2247, Q(27) => 
                           n_2248, Q(26) => n_2249, Q(25) => n_2250, Q(24) => 
                           n_2251, Q(23) => n_2252, Q(22) => n_2253, Q(21) => 
                           n_2254, Q(20) => n_2255, Q(19) => n_2256, Q(18) => 
                           n_2257, Q(17) => n_2258, Q(16) => n_2259, Q(15) => 
                           n_2260, Q(14) => n_2261, Q(13) => n_2262, Q(12) => 
                           n_2263, Q(11) => n_2264, Q(10) => n_2265, Q(9) => 
                           n_2266, Q(8) => n_2267, Q(7) => n_2268, Q(6) => 
                           n_2269, Q(5) => n_2270, Q(4) => n_2271, Q(3) => 
                           n_2272, Q(2) => n_2273, Q(1) => n_2274, Q(0) => 
                           n_2275);
   pipeline_IR1 : regFFD_NBIT32_11 port map( CK => CLK, RESET => RST, ENABLE =>
                           ir_LATCH_EN, D(31) => ir_fetch_31_port, D(30) => 
                           ir_fetch_30_port, D(29) => ir_fetch_29_port, D(28) 
                           => ir_fetch_28_port, D(27) => ir_fetch_27_port, 
                           D(26) => ir_fetch_26_port, D(25) => ir_fetch_25_port
                           , D(24) => ir_fetch_24_port, D(23) => 
                           ir_fetch_23_port, D(22) => ir_fetch_22_port, D(21) 
                           => ir_fetch_21_port, D(20) => ir_fetch_20_port, 
                           D(19) => ir_fetch_19_port, D(18) => ir_fetch_18_port
                           , D(17) => ir_fetch_17_port, D(16) => 
                           ir_fetch_16_port, D(15) => ir_fetch_15_port, D(14) 
                           => ir_fetch_14_port, D(13) => ir_fetch_13_port, 
                           D(12) => ir_fetch_12_port, D(11) => ir_fetch_11_port
                           , D(10) => ir_fetch_10_port, D(9) => ir_fetch_9_port
                           , D(8) => ir_fetch_8_port, D(7) => ir_fetch_7_port, 
                           D(6) => ir_fetch_6_port, D(5) => ir_fetch_5_port, 
                           D(4) => ir_fetch_4_port, D(3) => ir_fetch_3_port, 
                           D(2) => ir_fetch_2_port, D(1) => ir_fetch_1_port, 
                           D(0) => ir_fetch_0_port, Q(31) => IR_Dec_31_port, 
                           Q(30) => IR_Dec_30_port, Q(29) => IR_Dec_29_port, 
                           Q(28) => IR_Dec_28_port, Q(27) => IR_Dec_27_port, 
                           Q(26) => IR_Dec_26_port, Q(25) => IR_Dec_25_port, 
                           Q(24) => IR_Dec_24_port, Q(23) => IR_Dec_23_port, 
                           Q(22) => IR_Dec_22_port, Q(21) => IR_Dec_21_port, 
                           Q(20) => IR_Dec_20_port, Q(19) => IR_Dec_19_port, 
                           Q(18) => IR_Dec_18_port, Q(17) => IR_Dec_17_port, 
                           Q(16) => IR_Dec_16_port, Q(15) => IR_Dec_15_port, 
                           Q(14) => IR_Dec_14_port, Q(13) => IR_Dec_13_port, 
                           Q(12) => IR_Dec_12_port, Q(11) => IR_Dec_11_port, 
                           Q(10) => IR_Dec_10_port, Q(9) => IR_Dec_9_port, Q(8)
                           => IR_Dec_8_port, Q(7) => IR_Dec_7_port, Q(6) => 
                           IR_Dec_6_port, Q(5) => IR_Dec_5_port, Q(4) => 
                           IR_Dec_4_port, Q(3) => IR_Dec_3_port, Q(2) => 
                           IR_Dec_2_port, Q(1) => IR_Dec_1_port, Q(0) => 
                           IR_Dec_0_port);
   IR_OP : IR_DECODE_NBIT32_opBIT6_regBIT5 port map( CLK => CLK, IR_26(25) => 
                           IR_Dec_25_port, IR_26(24) => IR_Dec_24_port, 
                           IR_26(23) => IR_Dec_23_port, IR_26(22) => 
                           IR_Dec_22_port, IR_26(21) => IR_Dec_21_port, 
                           IR_26(20) => IR_Dec_20_port, IR_26(19) => 
                           IR_Dec_19_port, IR_26(18) => IR_Dec_18_port, 
                           IR_26(17) => IR_Dec_17_port, IR_26(16) => 
                           IR_Dec_16_port, IR_26(15) => IR_Dec_15_port, 
                           IR_26(14) => IR_Dec_14_port, IR_26(13) => 
                           IR_Dec_13_port, IR_26(12) => IR_Dec_12_port, 
                           IR_26(11) => IR_Dec_11_port, IR_26(10) => 
                           IR_Dec_10_port, IR_26(9) => IR_Dec_9_port, IR_26(8) 
                           => IR_Dec_8_port, IR_26(7) => IR_Dec_7_port, 
                           IR_26(6) => IR_Dec_6_port, IR_26(5) => IR_Dec_5_port
                           , IR_26(4) => IR_Dec_4_port, IR_26(3) => 
                           IR_Dec_3_port, IR_26(2) => IR_Dec_2_port, IR_26(1) 
                           => IR_Dec_1_port, IR_26(0) => IR_Dec_0_port, 
                           OPCODE(5) => IR_Dec_31_port, OPCODE(4) => 
                           IR_Dec_30_port, OPCODE(3) => IR_Dec_29_port, 
                           OPCODE(2) => IR_Dec_28_port, OPCODE(1) => 
                           IR_Dec_27_port, OPCODE(0) => IR_Dec_26_port, 
                           is_signed => signed_op, RS1(4) => RS1_4_port, RS1(3)
                           => RS1_3_port, RS1(2) => RS1_2_port, RS1(1) => 
                           RS1_1_port, RS1(0) => RS1_0_port, RS2(4) => 
                           RS2_4_port, RS2(3) => RS2_3_port, RS2(2) => 
                           RS2_2_port, RS2(1) => RS2_1_port, RS2(0) => 
                           RS2_0_port, RD(4) => RD_4_port, RD(3) => RD_3_port, 
                           RD(2) => RD_2_port, RD(1) => RD_1_port, RD(0) => 
                           RD_0_port, IMMEDIATE(31) => Imm_31_port, 
                           IMMEDIATE(30) => Imm_30_port, IMMEDIATE(29) => 
                           Imm_29_port, IMMEDIATE(28) => Imm_28_port, 
                           IMMEDIATE(27) => Imm_27_port, IMMEDIATE(26) => 
                           Imm_26_port, IMMEDIATE(25) => Imm_25_port, 
                           IMMEDIATE(24) => Imm_24_port, IMMEDIATE(23) => 
                           Imm_23_port, IMMEDIATE(22) => Imm_22_port, 
                           IMMEDIATE(21) => Imm_21_port, IMMEDIATE(20) => 
                           Imm_20_port, IMMEDIATE(19) => Imm_19_port, 
                           IMMEDIATE(18) => Imm_18_port, IMMEDIATE(17) => 
                           Imm_17_port, IMMEDIATE(16) => Imm_16_port, 
                           IMMEDIATE(15) => Imm_15_port, IMMEDIATE(14) => 
                           Imm_14_port, IMMEDIATE(13) => Imm_13_port, 
                           IMMEDIATE(12) => Imm_12_port, IMMEDIATE(11) => 
                           Imm_11_port, IMMEDIATE(10) => Imm_10_port, 
                           IMMEDIATE(9) => Imm_9_port, IMMEDIATE(8) => 
                           Imm_8_port, IMMEDIATE(7) => Imm_7_port, IMMEDIATE(6)
                           => Imm_6_port, IMMEDIATE(5) => Imm_5_port, 
                           IMMEDIATE(4) => Imm_4_port, IMMEDIATE(3) => 
                           Imm_3_port, IMMEDIATE(2) => Imm_2_port, IMMEDIATE(1)
                           => Imm_1_port, IMMEDIATE(0) => Imm_0_port);
   RF : register_file port map( CLK => CLK, RESET => RST, ENABLE => 
                           X_Logic1_port, RD1 => RF1, RD2 => RF2, WR => WF1, 
                           ADD_WR(4) => RD_wb_4_port, ADD_WR(3) => RD_wb_3_port
                           , ADD_WR(2) => RD_wb_2_port, ADD_WR(1) => 
                           RD_wb_1_port, ADD_WR(0) => RD_wb_0_port, ADD_RD1(4) 
                           => RS1_4_port, ADD_RD1(3) => RS1_3_port, ADD_RD1(2) 
                           => RS1_2_port, ADD_RD1(1) => RS1_1_port, ADD_RD1(0) 
                           => RS1_0_port, ADD_RD2(4) => RS2_4_port, ADD_RD2(3) 
                           => RS2_3_port, ADD_RD2(2) => RS2_2_port, ADD_RD2(1) 
                           => RS2_1_port, ADD_RD2(0) => RS2_0_port, DATAIN(31) 
                           => OUT_data_31_port, DATAIN(30) => OUT_data_30_port,
                           DATAIN(29) => OUT_data_29_port, DATAIN(28) => 
                           OUT_data_28_port, DATAIN(27) => OUT_data_27_port, 
                           DATAIN(26) => OUT_data_26_port, DATAIN(25) => 
                           OUT_data_25_port, DATAIN(24) => OUT_data_24_port, 
                           DATAIN(23) => OUT_data_23_port, DATAIN(22) => 
                           OUT_data_22_port, DATAIN(21) => OUT_data_21_port, 
                           DATAIN(20) => OUT_data_20_port, DATAIN(19) => 
                           OUT_data_19_port, DATAIN(18) => OUT_data_18_port, 
                           DATAIN(17) => OUT_data_17_port, DATAIN(16) => 
                           OUT_data_16_port, DATAIN(15) => OUT_data_15_port, 
                           DATAIN(14) => OUT_data_14_port, DATAIN(13) => 
                           OUT_data_13_port, DATAIN(12) => OUT_data_12_port, 
                           DATAIN(11) => OUT_data_11_port, DATAIN(10) => 
                           OUT_data_10_port, DATAIN(9) => OUT_data_9_port, 
                           DATAIN(8) => OUT_data_8_port, DATAIN(7) => 
                           OUT_data_7_port, DATAIN(6) => OUT_data_6_port, 
                           DATAIN(5) => OUT_data_5_port, DATAIN(4) => 
                           OUT_data_4_port, DATAIN(3) => OUT_data_3_port, 
                           DATAIN(2) => OUT_data_2_port, DATAIN(1) => 
                           OUT_data_1_port, DATAIN(0) => OUT_data_0_port, 
                           OUT1(31) => regA_31_port, OUT1(30) => regA_30_port, 
                           OUT1(29) => regA_29_port, OUT1(28) => regA_28_port, 
                           OUT1(27) => regA_27_port, OUT1(26) => regA_26_port, 
                           OUT1(25) => regA_25_port, OUT1(24) => regA_24_port, 
                           OUT1(23) => regA_23_port, OUT1(22) => regA_22_port, 
                           OUT1(21) => regA_21_port, OUT1(20) => regA_20_port, 
                           OUT1(19) => regA_19_port, OUT1(18) => regA_18_port, 
                           OUT1(17) => regA_17_port, OUT1(16) => regA_16_port, 
                           OUT1(15) => regA_15_port, OUT1(14) => regA_14_port, 
                           OUT1(13) => regA_13_port, OUT1(12) => regA_12_port, 
                           OUT1(11) => regA_11_port, OUT1(10) => regA_10_port, 
                           OUT1(9) => regA_9_port, OUT1(8) => regA_8_port, 
                           OUT1(7) => regA_7_port, OUT1(6) => regA_6_port, 
                           OUT1(5) => regA_5_port, OUT1(4) => regA_4_port, 
                           OUT1(3) => regA_3_port, OUT1(2) => regA_2_port, 
                           OUT1(1) => regA_1_port, OUT1(0) => regA_0_port, 
                           OUT2(31) => regB_31_port, OUT2(30) => regB_30_port, 
                           OUT2(29) => regB_29_port, OUT2(28) => regB_28_port, 
                           OUT2(27) => regB_27_port, OUT2(26) => regB_26_port, 
                           OUT2(25) => regB_25_port, OUT2(24) => regB_24_port, 
                           OUT2(23) => regB_23_port, OUT2(22) => regB_22_port, 
                           OUT2(21) => regB_21_port, OUT2(20) => regB_20_port, 
                           OUT2(19) => regB_19_port, OUT2(18) => regB_18_port, 
                           OUT2(17) => regB_17_port, OUT2(16) => regB_16_port, 
                           OUT2(15) => regB_15_port, OUT2(14) => regB_14_port, 
                           OUT2(13) => regB_13_port, OUT2(12) => regB_12_port, 
                           OUT2(11) => regB_11_port, OUT2(10) => regB_10_port, 
                           OUT2(9) => regB_9_port, OUT2(8) => regB_8_port, 
                           OUT2(7) => regB_7_port, OUT2(6) => regB_6_port, 
                           OUT2(5) => regB_5_port, OUT2(4) => regB_4_port, 
                           OUT2(3) => regB_3_port, OUT2(2) => regB_2_port, 
                           OUT2(1) => regB_1_port, OUT2(0) => regB_0_port, 
                           wr_signal => wr_signal_wb);
   pipeline_sign2 : FF_0 port map( CLK => CLK, RESET => RST, EN => 
                           X_Logic1_port, D => signed_op, Q => signed_op_ex);
   pipeline_newpc2 : regFFD_NBIT32_10 port map( CK => CLK, RESET => RST, ENABLE
                           => X_Logic1_port, D(31) => NPC_Dec_31_port, D(30) =>
                           NPC_Dec_30_port, D(29) => NPC_Dec_29_port, D(28) => 
                           NPC_Dec_28_port, D(27) => NPC_Dec_27_port, D(26) => 
                           NPC_Dec_26_port, D(25) => NPC_Dec_25_port, D(24) => 
                           NPC_Dec_24_port, D(23) => NPC_Dec_23_port, D(22) => 
                           NPC_Dec_22_port, D(21) => NPC_Dec_21_port, D(20) => 
                           NPC_Dec_20_port, D(19) => NPC_Dec_19_port, D(18) => 
                           NPC_Dec_18_port, D(17) => NPC_Dec_17_port, D(16) => 
                           NPC_Dec_16_port, D(15) => NPC_Dec_15_port, D(14) => 
                           NPC_Dec_14_port, D(13) => NPC_Dec_13_port, D(12) => 
                           NPC_Dec_12_port, D(11) => NPC_Dec_11_port, D(10) => 
                           NPC_Dec_10_port, D(9) => NPC_Dec_9_port, D(8) => 
                           NPC_Dec_8_port, D(7) => NPC_Dec_7_port, D(6) => 
                           NPC_Dec_6_port, D(5) => NPC_Dec_5_port, D(4) => 
                           NPC_Dec_4_port, D(3) => NPC_Dec_3_port, D(2) => 
                           NPC_Dec_2_port, D(1) => NPC_Dec_1_port, D(0) => 
                           NPC_Dec_0_port, Q(31) => NPC_ex_31_port, Q(30) => 
                           NPC_ex_30_port, Q(29) => NPC_ex_29_port, Q(28) => 
                           NPC_ex_28_port, Q(27) => NPC_ex_27_port, Q(26) => 
                           NPC_ex_26_port, Q(25) => NPC_ex_25_port, Q(24) => 
                           NPC_ex_24_port, Q(23) => NPC_ex_23_port, Q(22) => 
                           NPC_ex_22_port, Q(21) => NPC_ex_21_port, Q(20) => 
                           NPC_ex_20_port, Q(19) => NPC_ex_19_port, Q(18) => 
                           NPC_ex_18_port, Q(17) => NPC_ex_17_port, Q(16) => 
                           NPC_ex_16_port, Q(15) => NPC_ex_15_port, Q(14) => 
                           NPC_ex_14_port, Q(13) => NPC_ex_13_port, Q(12) => 
                           NPC_ex_12_port, Q(11) => NPC_ex_11_port, Q(10) => 
                           NPC_ex_10_port, Q(9) => NPC_ex_9_port, Q(8) => 
                           NPC_ex_8_port, Q(7) => NPC_ex_7_port, Q(6) => 
                           NPC_ex_6_port, Q(5) => NPC_ex_5_port, Q(4) => 
                           NPC_ex_4_port, Q(3) => NPC_ex_3_port, Q(2) => 
                           NPC_ex_2_port, Q(1) => NPC_ex_1_port, Q(0) => 
                           NPC_ex_0_port);
   pipeline_A2 : regFFD_NBIT32_9 port map( CK => CLK, RESET => RST, ENABLE => 
                           RF1, D(31) => regA_31_port, D(30) => regA_30_port, 
                           D(29) => regA_29_port, D(28) => regA_28_port, D(27) 
                           => regA_27_port, D(26) => regA_26_port, D(25) => 
                           regA_25_port, D(24) => regA_24_port, D(23) => 
                           regA_23_port, D(22) => regA_22_port, D(21) => 
                           regA_21_port, D(20) => regA_20_port, D(19) => 
                           regA_19_port, D(18) => regA_18_port, D(17) => 
                           regA_17_port, D(16) => regA_16_port, D(15) => 
                           regA_15_port, D(14) => regA_14_port, D(13) => 
                           regA_13_port, D(12) => regA_12_port, D(11) => 
                           regA_11_port, D(10) => regA_10_port, D(9) => 
                           regA_9_port, D(8) => regA_8_port, D(7) => 
                           regA_7_port, D(6) => regA_6_port, D(5) => 
                           regA_5_port, D(4) => regA_4_port, D(3) => 
                           regA_3_port, D(2) => regA_2_port, D(1) => 
                           regA_1_port, D(0) => regA_0_port, Q(31) => 
                           regA_ex_31_port, Q(30) => regA_ex_30_port, Q(29) => 
                           regA_ex_29_port, Q(28) => regA_ex_28_port, Q(27) => 
                           regA_ex_27_port, Q(26) => regA_ex_26_port, Q(25) => 
                           regA_ex_25_port, Q(24) => regA_ex_24_port, Q(23) => 
                           regA_ex_23_port, Q(22) => regA_ex_22_port, Q(21) => 
                           regA_ex_21_port, Q(20) => regA_ex_20_port, Q(19) => 
                           regA_ex_19_port, Q(18) => regA_ex_18_port, Q(17) => 
                           regA_ex_17_port, Q(16) => regA_ex_16_port, Q(15) => 
                           regA_ex_15_port, Q(14) => regA_ex_14_port, Q(13) => 
                           regA_ex_13_port, Q(12) => regA_ex_12_port, Q(11) => 
                           regA_ex_11_port, Q(10) => regA_ex_10_port, Q(9) => 
                           regA_ex_9_port, Q(8) => regA_ex_8_port, Q(7) => 
                           regA_ex_7_port, Q(6) => regA_ex_6_port, Q(5) => 
                           regA_ex_5_port, Q(4) => regA_ex_4_port, Q(3) => 
                           regA_ex_3_port, Q(2) => regA_ex_2_port, Q(1) => 
                           regA_ex_1_port, Q(0) => regA_ex_0_port);
   pipeline_B2 : regFFD_NBIT32_8 port map( CK => CLK, RESET => RST, ENABLE => 
                           RF2, D(31) => regB_31_port, D(30) => regB_30_port, 
                           D(29) => regB_29_port, D(28) => regB_28_port, D(27) 
                           => regB_27_port, D(26) => regB_26_port, D(25) => 
                           regB_25_port, D(24) => regB_24_port, D(23) => 
                           regB_23_port, D(22) => regB_22_port, D(21) => 
                           regB_21_port, D(20) => regB_20_port, D(19) => 
                           regB_19_port, D(18) => regB_18_port, D(17) => 
                           regB_17_port, D(16) => regB_16_port, D(15) => 
                           regB_15_port, D(14) => regB_14_port, D(13) => 
                           regB_13_port, D(12) => regB_12_port, D(11) => 
                           regB_11_port, D(10) => regB_10_port, D(9) => 
                           regB_9_port, D(8) => regB_8_port, D(7) => 
                           regB_7_port, D(6) => regB_6_port, D(5) => 
                           regB_5_port, D(4) => regB_4_port, D(3) => 
                           regB_3_port, D(2) => regB_2_port, D(1) => 
                           regB_1_port, D(0) => regB_0_port, Q(31) => 
                           regB_ex_31_port, Q(30) => regB_ex_30_port, Q(29) => 
                           regB_ex_29_port, Q(28) => regB_ex_28_port, Q(27) => 
                           regB_ex_27_port, Q(26) => regB_ex_26_port, Q(25) => 
                           regB_ex_25_port, Q(24) => regB_ex_24_port, Q(23) => 
                           regB_ex_23_port, Q(22) => regB_ex_22_port, Q(21) => 
                           regB_ex_21_port, Q(20) => regB_ex_20_port, Q(19) => 
                           regB_ex_19_port, Q(18) => regB_ex_18_port, Q(17) => 
                           regB_ex_17_port, Q(16) => regB_ex_16_port, Q(15) => 
                           regB_ex_15_port, Q(14) => regB_ex_14_port, Q(13) => 
                           regB_ex_13_port, Q(12) => regB_ex_12_port, Q(11) => 
                           regB_ex_11_port, Q(10) => regB_ex_10_port, Q(9) => 
                           regB_ex_9_port, Q(8) => regB_ex_8_port, Q(7) => 
                           regB_ex_7_port, Q(6) => regB_ex_6_port, Q(5) => 
                           regB_ex_5_port, Q(4) => regB_ex_4_port, Q(3) => 
                           regB_ex_3_port, Q(2) => regB_ex_2_port, Q(1) => 
                           regB_ex_1_port, Q(0) => regB_ex_0_port);
   pipeline_IMM2 : regFFD_NBIT32_7 port map( CK => CLK, RESET => RST, ENABLE =>
                           regImm_LATCH_EN, D(31) => Imm_31_port, D(30) => 
                           Imm_30_port, D(29) => Imm_29_port, D(28) => 
                           Imm_28_port, D(27) => Imm_27_port, D(26) => 
                           Imm_26_port, D(25) => Imm_25_port, D(24) => 
                           Imm_24_port, D(23) => Imm_23_port, D(22) => 
                           Imm_22_port, D(21) => Imm_21_port, D(20) => 
                           Imm_20_port, D(19) => Imm_19_port, D(18) => 
                           Imm_18_port, D(17) => Imm_17_port, D(16) => 
                           Imm_16_port, D(15) => Imm_15_port, D(14) => 
                           Imm_14_port, D(13) => Imm_13_port, D(12) => 
                           Imm_12_port, D(11) => Imm_11_port, D(10) => 
                           Imm_10_port, D(9) => Imm_9_port, D(8) => Imm_8_port,
                           D(7) => Imm_7_port, D(6) => Imm_6_port, D(5) => 
                           Imm_5_port, D(4) => Imm_4_port, D(3) => Imm_3_port, 
                           D(2) => Imm_2_port, D(1) => Imm_1_port, D(0) => 
                           Imm_0_port, Q(31) => Imm_ex_31_port, Q(30) => 
                           Imm_ex_30_port, Q(29) => Imm_ex_29_port, Q(28) => 
                           Imm_ex_28_port, Q(27) => Imm_ex_27_port, Q(26) => 
                           Imm_ex_26_port, Q(25) => Imm_ex_25_port, Q(24) => 
                           Imm_ex_24_port, Q(23) => Imm_ex_23_port, Q(22) => 
                           Imm_ex_22_port, Q(21) => Imm_ex_21_port, Q(20) => 
                           Imm_ex_20_port, Q(19) => Imm_ex_19_port, Q(18) => 
                           Imm_ex_18_port, Q(17) => Imm_ex_17_port, Q(16) => 
                           Imm_ex_16_port, Q(15) => Imm_ex_15_port, Q(14) => 
                           Imm_ex_14_port, Q(13) => Imm_ex_13_port, Q(12) => 
                           Imm_ex_12_port, Q(11) => Imm_ex_11_port, Q(10) => 
                           Imm_ex_10_port, Q(9) => Imm_ex_9_port, Q(8) => 
                           Imm_ex_8_port, Q(7) => Imm_ex_7_port, Q(6) => 
                           Imm_ex_6_port, Q(5) => Imm_ex_5_port, Q(4) => 
                           Imm_ex_4_port, Q(3) => Imm_ex_3_port, Q(2) => 
                           Imm_ex_2_port, Q(1) => Imm_ex_1_port, Q(0) => 
                           Imm_ex_0_port);
   pipeline_RD2 : regFFD_NBIT5_0 port map( CK => CLK, RESET => RST, ENABLE => 
                           X_Logic1_port, D(4) => RD_4_port, D(3) => RD_3_port,
                           D(2) => RD_2_port, D(1) => RD_1_port, D(0) => 
                           RD_0_port, Q(4) => RD_ex_4_port, Q(3) => 
                           RD_ex_3_port, Q(2) => RD_ex_2_port, Q(1) => 
                           RD_ex_1_port, Q(0) => RD_ex_0_port);
   pipeline_wr_signal : FF_7 port map( CLK => CLK, RESET => RST, EN => 
                           X_Logic1_port, D => wr_signal, Q => wr_signal_exe);
   pipeline_IR2 : regFFD_NBIT6_0 port map( CK => CLK, RESET => RST, ENABLE => 
                           X_Logic1_port, D(5) => n42, D(4) => n44, D(3) => n45
                           , D(2) => IR_Dec_28_port, D(1) => IR_Dec_27_port, 
                           D(0) => n40, Q(5) => IR_26_ex_5_port, Q(4) => 
                           IR_26_ex_4_port, Q(3) => IR_26_ex_3_port, Q(2) => 
                           IR_26_ex_2_port, Q(1) => IR_26_ex_1_port, Q(0) => 
                           IR_26_ex_0_port);
   pipeline_LHI2 : regFFD_NBIT32_6 port map( CK => CLK, RESET => RST, ENABLE =>
                           X_Logic1_port, D(31) => Imm_15_port, D(30) => 
                           Imm_14_port, D(29) => Imm_13_port, D(28) => 
                           Imm_12_port, D(27) => Imm_11_port, D(26) => 
                           Imm_10_port, D(25) => Imm_9_port, D(24) => 
                           Imm_8_port, D(23) => Imm_7_port, D(22) => Imm_6_port
                           , D(21) => Imm_5_port, D(20) => Imm_4_port, D(19) =>
                           Imm_3_port, D(18) => Imm_2_port, D(17) => Imm_1_port
                           , D(16) => Imm_0_port, D(15) => X_Logic0_port, D(14)
                           => X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, Q(31) => LHI_ex_31_port, Q(30) => 
                           LHI_ex_30_port, Q(29) => LHI_ex_29_port, Q(28) => 
                           LHI_ex_28_port, Q(27) => LHI_ex_27_port, Q(26) => 
                           LHI_ex_26_port, Q(25) => LHI_ex_25_port, Q(24) => 
                           LHI_ex_24_port, Q(23) => LHI_ex_23_port, Q(22) => 
                           LHI_ex_22_port, Q(21) => LHI_ex_21_port, Q(20) => 
                           LHI_ex_20_port, Q(19) => LHI_ex_19_port, Q(18) => 
                           LHI_ex_18_port, Q(17) => LHI_ex_17_port, Q(16) => 
                           LHI_ex_16_port, Q(15) => LHI_ex_15_port, Q(14) => 
                           LHI_ex_14_port, Q(13) => LHI_ex_13_port, Q(12) => 
                           LHI_ex_12_port, Q(11) => LHI_ex_11_port, Q(10) => 
                           LHI_ex_10_port, Q(9) => LHI_ex_9_port, Q(8) => 
                           LHI_ex_8_port, Q(7) => LHI_ex_7_port, Q(6) => 
                           LHI_ex_6_port, Q(5) => LHI_ex_5_port, Q(4) => 
                           LHI_ex_4_port, Q(3) => LHI_ex_3_port, Q(2) => 
                           LHI_ex_2_port, Q(1) => LHI_ex_1_port, Q(0) => 
                           LHI_ex_0_port);
   MUX_ALU_A : MUX21_GENERIC_NBIT32_6 port map( A(31) => NPC_ex_31_port, A(30) 
                           => NPC_ex_30_port, A(29) => NPC_ex_29_port, A(28) =>
                           NPC_ex_28_port, A(27) => NPC_ex_27_port, A(26) => 
                           NPC_ex_26_port, A(25) => NPC_ex_25_port, A(24) => 
                           NPC_ex_24_port, A(23) => NPC_ex_23_port, A(22) => 
                           NPC_ex_22_port, A(21) => NPC_ex_21_port, A(20) => 
                           NPC_ex_20_port, A(19) => NPC_ex_19_port, A(18) => 
                           NPC_ex_18_port, A(17) => NPC_ex_17_port, A(16) => 
                           NPC_ex_16_port, A(15) => NPC_ex_15_port, A(14) => 
                           NPC_ex_14_port, A(13) => NPC_ex_13_port, A(12) => 
                           NPC_ex_12_port, A(11) => NPC_ex_11_port, A(10) => 
                           NPC_ex_10_port, A(9) => NPC_ex_9_port, A(8) => 
                           NPC_ex_8_port, A(7) => NPC_ex_7_port, A(6) => 
                           NPC_ex_6_port, A(5) => NPC_ex_5_port, A(4) => 
                           NPC_ex_4_port, A(3) => NPC_ex_3_port, A(2) => 
                           NPC_ex_2_port, A(1) => NPC_ex_1_port, A(0) => 
                           NPC_ex_0_port, B(31) => regA_ex_31_port, B(30) => 
                           regA_ex_30_port, B(29) => regA_ex_29_port, B(28) => 
                           regA_ex_28_port, B(27) => regA_ex_27_port, B(26) => 
                           regA_ex_26_port, B(25) => regA_ex_25_port, B(24) => 
                           regA_ex_24_port, B(23) => regA_ex_23_port, B(22) => 
                           regA_ex_22_port, B(21) => regA_ex_21_port, B(20) => 
                           regA_ex_20_port, B(19) => regA_ex_19_port, B(18) => 
                           regA_ex_18_port, B(17) => regA_ex_17_port, B(16) => 
                           regA_ex_16_port, B(15) => regA_ex_15_port, B(14) => 
                           regA_ex_14_port, B(13) => regA_ex_13_port, B(12) => 
                           regA_ex_12_port, B(11) => regA_ex_11_port, B(10) => 
                           regA_ex_10_port, B(9) => regA_ex_9_port, B(8) => 
                           regA_ex_8_port, B(7) => regA_ex_7_port, B(6) => 
                           regA_ex_6_port, B(5) => regA_ex_5_port, B(4) => 
                           regA_ex_4_port, B(3) => regA_ex_3_port, B(2) => 
                           regA_ex_2_port, B(1) => regA_ex_1_port, B(0) => 
                           regA_ex_0_port, SEL => S1, Y(31) => 
                           input1_ALU_31_port, Y(30) => input1_ALU_30_port, 
                           Y(29) => input1_ALU_29_port, Y(28) => 
                           input1_ALU_28_port, Y(27) => input1_ALU_27_port, 
                           Y(26) => input1_ALU_26_port, Y(25) => 
                           input1_ALU_25_port, Y(24) => input1_ALU_24_port, 
                           Y(23) => input1_ALU_23_port, Y(22) => 
                           input1_ALU_22_port, Y(21) => input1_ALU_21_port, 
                           Y(20) => input1_ALU_20_port, Y(19) => 
                           input1_ALU_19_port, Y(18) => input1_ALU_18_port, 
                           Y(17) => input1_ALU_17_port, Y(16) => 
                           input1_ALU_16_port, Y(15) => input1_ALU_15_port, 
                           Y(14) => input1_ALU_14_port, Y(13) => 
                           input1_ALU_13_port, Y(12) => input1_ALU_12_port, 
                           Y(11) => input1_ALU_11_port, Y(10) => 
                           input1_ALU_10_port, Y(9) => input1_ALU_9_port, Y(8) 
                           => input1_ALU_8_port, Y(7) => input1_ALU_7_port, 
                           Y(6) => input1_ALU_6_port, Y(5) => input1_ALU_5_port
                           , Y(4) => input1_ALU_4_port, Y(3) => 
                           input1_ALU_3_port, Y(2) => input1_ALU_2_port, Y(1) 
                           => input1_ALU_1_port, Y(0) => input1_ALU_0_port);
   MUX_ALU_B : MUX21_GENERIC_NBIT32_5 port map( A(31) => Imm_ex_31_port, A(30) 
                           => Imm_ex_30_port, A(29) => Imm_ex_29_port, A(28) =>
                           Imm_ex_28_port, A(27) => Imm_ex_27_port, A(26) => 
                           Imm_ex_26_port, A(25) => Imm_ex_25_port, A(24) => 
                           Imm_ex_24_port, A(23) => Imm_ex_23_port, A(22) => 
                           Imm_ex_22_port, A(21) => Imm_ex_21_port, A(20) => 
                           Imm_ex_20_port, A(19) => Imm_ex_19_port, A(18) => 
                           Imm_ex_18_port, A(17) => Imm_ex_17_port, A(16) => 
                           Imm_ex_16_port, A(15) => Imm_ex_15_port, A(14) => 
                           Imm_ex_14_port, A(13) => Imm_ex_13_port, A(12) => 
                           Imm_ex_12_port, A(11) => Imm_ex_11_port, A(10) => 
                           Imm_ex_10_port, A(9) => Imm_ex_9_port, A(8) => 
                           Imm_ex_8_port, A(7) => Imm_ex_7_port, A(6) => 
                           Imm_ex_6_port, A(5) => Imm_ex_5_port, A(4) => 
                           Imm_ex_4_port, A(3) => Imm_ex_3_port, A(2) => 
                           Imm_ex_2_port, A(1) => Imm_ex_1_port, A(0) => 
                           Imm_ex_0_port, B(31) => regB_ex_31_port, B(30) => 
                           regB_ex_30_port, B(29) => regB_ex_29_port, B(28) => 
                           regB_ex_28_port, B(27) => regB_ex_27_port, B(26) => 
                           regB_ex_26_port, B(25) => regB_ex_25_port, B(24) => 
                           regB_ex_24_port, B(23) => regB_ex_23_port, B(22) => 
                           regB_ex_22_port, B(21) => regB_ex_21_port, B(20) => 
                           regB_ex_20_port, B(19) => regB_ex_19_port, B(18) => 
                           regB_ex_18_port, B(17) => regB_ex_17_port, B(16) => 
                           regB_ex_16_port, B(15) => regB_ex_15_port, B(14) => 
                           regB_ex_14_port, B(13) => regB_ex_13_port, B(12) => 
                           regB_ex_12_port, B(11) => regB_ex_11_port, B(10) => 
                           regB_ex_10_port, B(9) => regB_ex_9_port, B(8) => 
                           regB_ex_8_port, B(7) => regB_ex_7_port, B(6) => 
                           regB_ex_6_port, B(5) => regB_ex_5_port, B(4) => 
                           regB_ex_4_port, B(3) => regB_ex_3_port, B(2) => 
                           regB_ex_2_port, B(1) => regB_ex_1_port, B(0) => 
                           regB_ex_0_port, SEL => S2, Y(31) => 
                           input2_ALU_31_port, Y(30) => input2_ALU_30_port, 
                           Y(29) => input2_ALU_29_port, Y(28) => 
                           input2_ALU_28_port, Y(27) => input2_ALU_27_port, 
                           Y(26) => input2_ALU_26_port, Y(25) => 
                           input2_ALU_25_port, Y(24) => input2_ALU_24_port, 
                           Y(23) => input2_ALU_23_port, Y(22) => 
                           input2_ALU_22_port, Y(21) => input2_ALU_21_port, 
                           Y(20) => input2_ALU_20_port, Y(19) => 
                           input2_ALU_19_port, Y(18) => input2_ALU_18_port, 
                           Y(17) => input2_ALU_17_port, Y(16) => 
                           input2_ALU_16_port, Y(15) => input2_ALU_15_port, 
                           Y(14) => input2_ALU_14_port, Y(13) => 
                           input2_ALU_13_port, Y(12) => input2_ALU_12_port, 
                           Y(11) => input2_ALU_11_port, Y(10) => 
                           input2_ALU_10_port, Y(9) => input2_ALU_9_port, Y(8) 
                           => input2_ALU_8_port, Y(7) => input2_ALU_7_port, 
                           Y(6) => input2_ALU_6_port, Y(5) => input2_ALU_5_port
                           , Y(4) => input2_ALU_4_port, Y(3) => 
                           input2_ALU_3_port, Y(2) => input2_ALU_2_port, Y(1) 
                           => input2_ALU_1_port, Y(0) => input2_ALU_0_port);
   ALU_OP : ALU_N32 port map( CLK => CLK, FUNC(0) => instruction_alu(0), 
                           FUNC(1) => instruction_alu(1), FUNC(2) => 
                           instruction_alu(2), FUNC(3) => instruction_alu(3), 
                           FUNC(4) => instruction_alu(4), FUNC(5) => 
                           instruction_alu(5), DATA1(31) => input1_ALU_31_port,
                           DATA1(30) => input1_ALU_30_port, DATA1(29) => 
                           input1_ALU_29_port, DATA1(28) => input1_ALU_28_port,
                           DATA1(27) => input1_ALU_27_port, DATA1(26) => 
                           input1_ALU_26_port, DATA1(25) => input1_ALU_25_port,
                           DATA1(24) => input1_ALU_24_port, DATA1(23) => 
                           input1_ALU_23_port, DATA1(22) => input1_ALU_22_port,
                           DATA1(21) => input1_ALU_21_port, DATA1(20) => 
                           input1_ALU_20_port, DATA1(19) => input1_ALU_19_port,
                           DATA1(18) => input1_ALU_18_port, DATA1(17) => 
                           input1_ALU_17_port, DATA1(16) => input1_ALU_16_port,
                           DATA1(15) => input1_ALU_15_port, DATA1(14) => 
                           input1_ALU_14_port, DATA1(13) => input1_ALU_13_port,
                           DATA1(12) => input1_ALU_12_port, DATA1(11) => 
                           input1_ALU_11_port, DATA1(10) => input1_ALU_10_port,
                           DATA1(9) => input1_ALU_9_port, DATA1(8) => 
                           input1_ALU_8_port, DATA1(7) => input1_ALU_7_port, 
                           DATA1(6) => input1_ALU_6_port, DATA1(5) => 
                           input1_ALU_5_port, DATA1(4) => input1_ALU_4_port, 
                           DATA1(3) => input1_ALU_3_port, DATA1(2) => 
                           input1_ALU_2_port, DATA1(1) => input1_ALU_1_port, 
                           DATA1(0) => input1_ALU_0_port, DATA2(31) => 
                           input2_ALU_31_port, DATA2(30) => input2_ALU_30_port,
                           DATA2(29) => input2_ALU_29_port, DATA2(28) => 
                           input2_ALU_28_port, DATA2(27) => input2_ALU_27_port,
                           DATA2(26) => input2_ALU_26_port, DATA2(25) => 
                           input2_ALU_25_port, DATA2(24) => input2_ALU_24_port,
                           DATA2(23) => input2_ALU_23_port, DATA2(22) => 
                           input2_ALU_22_port, DATA2(21) => input2_ALU_21_port,
                           DATA2(20) => input2_ALU_20_port, DATA2(19) => 
                           input2_ALU_19_port, DATA2(18) => input2_ALU_18_port,
                           DATA2(17) => input2_ALU_17_port, DATA2(16) => 
                           input2_ALU_16_port, DATA2(15) => input2_ALU_15_port,
                           DATA2(14) => input2_ALU_14_port, DATA2(13) => 
                           input2_ALU_13_port, DATA2(12) => input2_ALU_12_port,
                           DATA2(11) => input2_ALU_11_port, DATA2(10) => 
                           input2_ALU_10_port, DATA2(9) => input2_ALU_9_port, 
                           DATA2(8) => input2_ALU_8_port, DATA2(7) => 
                           input2_ALU_7_port, DATA2(6) => input2_ALU_6_port, 
                           DATA2(5) => input2_ALU_5_port, DATA2(4) => 
                           input2_ALU_4_port, DATA2(3) => input2_ALU_3_port, 
                           DATA2(2) => input2_ALU_2_port, DATA2(1) => 
                           input2_ALU_1_port, DATA2(0) => input2_ALU_0_port, 
                           OUT_ALU(31) => ALU_out_31_port, OUT_ALU(30) => 
                           ALU_out_30_port, OUT_ALU(29) => ALU_out_29_port, 
                           OUT_ALU(28) => ALU_out_28_port, OUT_ALU(27) => 
                           ALU_out_27_port, OUT_ALU(26) => ALU_out_26_port, 
                           OUT_ALU(25) => ALU_out_25_port, OUT_ALU(24) => 
                           ALU_out_24_port, OUT_ALU(23) => ALU_out_23_port, 
                           OUT_ALU(22) => ALU_out_22_port, OUT_ALU(21) => 
                           ALU_out_21_port, OUT_ALU(20) => ALU_out_20_port, 
                           OUT_ALU(19) => ALU_out_19_port, OUT_ALU(18) => 
                           ALU_out_18_port, OUT_ALU(17) => ALU_out_17_port, 
                           OUT_ALU(16) => ALU_out_16_port, OUT_ALU(15) => 
                           ALU_out_15_port, OUT_ALU(14) => ALU_out_14_port, 
                           OUT_ALU(13) => ALU_out_13_port, OUT_ALU(12) => 
                           ALU_out_12_port, OUT_ALU(11) => ALU_out_11_port, 
                           OUT_ALU(10) => ALU_out_10_port, OUT_ALU(9) => 
                           ALU_out_9_port, OUT_ALU(8) => ALU_out_8_port, 
                           OUT_ALU(7) => ALU_out_7_port, OUT_ALU(6) => 
                           ALU_out_6_port, OUT_ALU(5) => ALU_out_5_port, 
                           OUT_ALU(4) => ALU_out_4_port, OUT_ALU(3) => 
                           ALU_out_3_port, OUT_ALU(2) => ALU_out_2_port, 
                           OUT_ALU(1) => ALU_out_1_port, OUT_ALU(0) => 
                           ALU_out_0_port);
   ZERO_OP : zero_eval_NBIT32 port map( input(31) => regA_ex_31_port, input(30)
                           => regA_ex_30_port, input(29) => regA_ex_29_port, 
                           input(28) => regA_ex_28_port, input(27) => 
                           regA_ex_27_port, input(26) => regA_ex_26_port, 
                           input(25) => regA_ex_25_port, input(24) => 
                           regA_ex_24_port, input(23) => regA_ex_23_port, 
                           input(22) => regA_ex_22_port, input(21) => 
                           regA_ex_21_port, input(20) => regA_ex_20_port, 
                           input(19) => regA_ex_19_port, input(18) => 
                           regA_ex_18_port, input(17) => regA_ex_17_port, 
                           input(16) => regA_ex_16_port, input(15) => 
                           regA_ex_15_port, input(14) => regA_ex_14_port, 
                           input(13) => regA_ex_13_port, input(12) => 
                           regA_ex_12_port, input(11) => regA_ex_11_port, 
                           input(10) => regA_ex_10_port, input(9) => 
                           regA_ex_9_port, input(8) => regA_ex_8_port, input(7)
                           => regA_ex_7_port, input(6) => regA_ex_6_port, 
                           input(5) => regA_ex_5_port, input(4) => 
                           regA_ex_4_port, input(3) => regA_ex_3_port, input(2)
                           => regA_ex_2_port, input(1) => regA_ex_1_port, 
                           input(0) => regA_ex_0_port, res => is_zero);
   COND_OP : COND_BT_NBIT32 port map( ZERO_BIT => is_zero, OPCODE_0 => 
                           IR_26_ex_0_port, branch_op => branch_cond, con_sign 
                           => cond);
   MUX_alu_out : MUX21_GENERIC_NBIT32_4 port map( A(31) => LHI_ex_31_port, 
                           A(30) => LHI_ex_30_port, A(29) => LHI_ex_29_port, 
                           A(28) => LHI_ex_28_port, A(27) => LHI_ex_27_port, 
                           A(26) => LHI_ex_26_port, A(25) => LHI_ex_25_port, 
                           A(24) => LHI_ex_24_port, A(23) => LHI_ex_23_port, 
                           A(22) => LHI_ex_22_port, A(21) => LHI_ex_21_port, 
                           A(20) => LHI_ex_20_port, A(19) => LHI_ex_19_port, 
                           A(18) => LHI_ex_18_port, A(17) => LHI_ex_17_port, 
                           A(16) => LHI_ex_16_port, A(15) => LHI_ex_15_port, 
                           A(14) => LHI_ex_14_port, A(13) => LHI_ex_13_port, 
                           A(12) => LHI_ex_12_port, A(11) => LHI_ex_11_port, 
                           A(10) => LHI_ex_10_port, A(9) => LHI_ex_9_port, A(8)
                           => LHI_ex_8_port, A(7) => LHI_ex_7_port, A(6) => 
                           LHI_ex_6_port, A(5) => LHI_ex_5_port, A(4) => 
                           LHI_ex_4_port, A(3) => LHI_ex_3_port, A(2) => 
                           LHI_ex_2_port, A(1) => LHI_ex_1_port, A(0) => 
                           LHI_ex_0_port, B(31) => ALU_out_31_port, B(30) => 
                           ALU_out_30_port, B(29) => ALU_out_29_port, B(28) => 
                           ALU_out_28_port, B(27) => ALU_out_27_port, B(26) => 
                           ALU_out_26_port, B(25) => ALU_out_25_port, B(24) => 
                           ALU_out_24_port, B(23) => ALU_out_23_port, B(22) => 
                           ALU_out_22_port, B(21) => ALU_out_21_port, B(20) => 
                           ALU_out_20_port, B(19) => ALU_out_19_port, B(18) => 
                           ALU_out_18_port, B(17) => ALU_out_17_port, B(16) => 
                           ALU_out_16_port, B(15) => ALU_out_15_port, B(14) => 
                           ALU_out_14_port, B(13) => ALU_out_13_port, B(12) => 
                           ALU_out_12_port, B(11) => ALU_out_11_port, B(10) => 
                           ALU_out_10_port, B(9) => ALU_out_9_port, B(8) => 
                           ALU_out_8_port, B(7) => ALU_out_7_port, B(6) => 
                           ALU_out_6_port, B(5) => ALU_out_5_port, B(4) => 
                           ALU_out_4_port, B(3) => ALU_out_3_port, B(2) => 
                           ALU_out_2_port, B(1) => ALU_out_1_port, B(0) => 
                           ALU_out_0_port, SEL => lhi_sel, Y(31) => 
                           ALU_ex_31_port, Y(30) => ALU_ex_30_port, Y(29) => 
                           ALU_ex_29_port, Y(28) => ALU_ex_28_port, Y(27) => 
                           ALU_ex_27_port, Y(26) => ALU_ex_26_port, Y(25) => 
                           ALU_ex_25_port, Y(24) => ALU_ex_24_port, Y(23) => 
                           ALU_ex_23_port, Y(22) => ALU_ex_22_port, Y(21) => 
                           ALU_ex_21_port, Y(20) => ALU_ex_20_port, Y(19) => 
                           ALU_ex_19_port, Y(18) => ALU_ex_18_port, Y(17) => 
                           ALU_ex_17_port, Y(16) => ALU_ex_16_port, Y(15) => 
                           ALU_ex_15_port, Y(14) => ALU_ex_14_port, Y(13) => 
                           ALU_ex_13_port, Y(12) => ALU_ex_12_port, Y(11) => 
                           ALU_ex_11_port, Y(10) => ALU_ex_10_port, Y(9) => 
                           ALU_ex_9_port, Y(8) => ALU_ex_8_port, Y(7) => 
                           ALU_ex_7_port, Y(6) => ALU_ex_6_port, Y(5) => 
                           ALU_ex_5_port, Y(4) => ALU_ex_4_port, Y(3) => 
                           ALU_ex_3_port, Y(2) => ALU_ex_2_port, Y(1) => 
                           ALU_ex_1_port, Y(0) => ALU_ex_0_port);
   pipeline_sign3 : FF_6 port map( CLK => CLK, RESET => RST, EN => 
                           X_Logic1_port, D => signed_op_ex, Q => signed_op_mem
                           );
   pipeline_newpc3 : regFFD_NBIT32_5 port map( CK => CLK, RESET => RST, ENABLE 
                           => X_Logic1_port, D(31) => NPC_ex_31_port, D(30) => 
                           NPC_ex_30_port, D(29) => NPC_ex_29_port, D(28) => 
                           NPC_ex_28_port, D(27) => NPC_ex_27_port, D(26) => 
                           NPC_ex_26_port, D(25) => NPC_ex_25_port, D(24) => 
                           NPC_ex_24_port, D(23) => NPC_ex_23_port, D(22) => 
                           NPC_ex_22_port, D(21) => NPC_ex_21_port, D(20) => 
                           NPC_ex_20_port, D(19) => NPC_ex_19_port, D(18) => 
                           NPC_ex_18_port, D(17) => NPC_ex_17_port, D(16) => 
                           NPC_ex_16_port, D(15) => NPC_ex_15_port, D(14) => 
                           NPC_ex_14_port, D(13) => NPC_ex_13_port, D(12) => 
                           NPC_ex_12_port, D(11) => NPC_ex_11_port, D(10) => 
                           NPC_ex_10_port, D(9) => NPC_ex_9_port, D(8) => 
                           NPC_ex_8_port, D(7) => NPC_ex_7_port, D(6) => 
                           NPC_ex_6_port, D(5) => NPC_ex_5_port, D(4) => 
                           NPC_ex_4_port, D(3) => NPC_ex_3_port, D(2) => 
                           NPC_ex_2_port, D(1) => NPC_ex_1_port, D(0) => 
                           NPC_ex_0_port, Q(31) => NPC_mem_31_port, Q(30) => 
                           NPC_mem_30_port, Q(29) => NPC_mem_29_port, Q(28) => 
                           NPC_mem_28_port, Q(27) => NPC_mem_27_port, Q(26) => 
                           NPC_mem_26_port, Q(25) => NPC_mem_25_port, Q(24) => 
                           NPC_mem_24_port, Q(23) => NPC_mem_23_port, Q(22) => 
                           NPC_mem_22_port, Q(21) => NPC_mem_21_port, Q(20) => 
                           NPC_mem_20_port, Q(19) => NPC_mem_19_port, Q(18) => 
                           NPC_mem_18_port, Q(17) => NPC_mem_17_port, Q(16) => 
                           NPC_mem_16_port, Q(15) => NPC_mem_15_port, Q(14) => 
                           NPC_mem_14_port, Q(13) => NPC_mem_13_port, Q(12) => 
                           NPC_mem_12_port, Q(11) => NPC_mem_11_port, Q(10) => 
                           NPC_mem_10_port, Q(9) => NPC_mem_9_port, Q(8) => 
                           NPC_mem_8_port, Q(7) => NPC_mem_7_port, Q(6) => 
                           NPC_mem_6_port, Q(5) => NPC_mem_5_port, Q(4) => 
                           NPC_mem_4_port, Q(3) => NPC_mem_3_port, Q(2) => 
                           NPC_mem_2_port, Q(1) => NPC_mem_1_port, Q(0) => 
                           NPC_mem_0_port);
   pipeline_cond3 : FF_5 port map( CLK => CLK, RESET => RST, EN => 
                           X_Logic1_port, D => cond, Q => cond_mem);
   pipeline_B3 : regFFD_NBIT32_4 port map( CK => CLK, RESET => RST, ENABLE => 
                           X_Logic1_port, D(31) => regB_ex_31_port, D(30) => 
                           regB_ex_30_port, D(29) => regB_ex_29_port, D(28) => 
                           regB_ex_28_port, D(27) => regB_ex_27_port, D(26) => 
                           regB_ex_26_port, D(25) => regB_ex_25_port, D(24) => 
                           regB_ex_24_port, D(23) => regB_ex_23_port, D(22) => 
                           regB_ex_22_port, D(21) => regB_ex_21_port, D(20) => 
                           regB_ex_20_port, D(19) => regB_ex_19_port, D(18) => 
                           regB_ex_18_port, D(17) => regB_ex_17_port, D(16) => 
                           regB_ex_16_port, D(15) => regB_ex_15_port, D(14) => 
                           regB_ex_14_port, D(13) => regB_ex_13_port, D(12) => 
                           regB_ex_12_port, D(11) => regB_ex_11_port, D(10) => 
                           regB_ex_10_port, D(9) => regB_ex_9_port, D(8) => 
                           regB_ex_8_port, D(7) => regB_ex_7_port, D(6) => 
                           regB_ex_6_port, D(5) => regB_ex_5_port, D(4) => 
                           regB_ex_4_port, D(3) => regB_ex_3_port, D(2) => 
                           regB_ex_2_port, D(1) => regB_ex_1_port, D(0) => 
                           regB_ex_0_port, Q(31) => regB_mem_31_port, Q(30) => 
                           regB_mem_30_port, Q(29) => regB_mem_29_port, Q(28) 
                           => regB_mem_28_port, Q(27) => regB_mem_27_port, 
                           Q(26) => regB_mem_26_port, Q(25) => regB_mem_25_port
                           , Q(24) => regB_mem_24_port, Q(23) => 
                           regB_mem_23_port, Q(22) => regB_mem_22_port, Q(21) 
                           => regB_mem_21_port, Q(20) => regB_mem_20_port, 
                           Q(19) => regB_mem_19_port, Q(18) => regB_mem_18_port
                           , Q(17) => regB_mem_17_port, Q(16) => 
                           regB_mem_16_port, Q(15) => regB_mem_15_port, Q(14) 
                           => regB_mem_14_port, Q(13) => regB_mem_13_port, 
                           Q(12) => regB_mem_12_port, Q(11) => regB_mem_11_port
                           , Q(10) => regB_mem_10_port, Q(9) => regB_mem_9_port
                           , Q(8) => regB_mem_8_port, Q(7) => regB_mem_7_port, 
                           Q(6) => regB_mem_6_port, Q(5) => regB_mem_5_port, 
                           Q(4) => regB_mem_4_port, Q(3) => regB_mem_3_port, 
                           Q(2) => regB_mem_2_port, Q(1) => regB_mem_1_port, 
                           Q(0) => regB_mem_0_port);
   pipeline_RD3 : regFFD_NBIT5_2 port map( CK => CLK, RESET => RST, ENABLE => 
                           X_Logic1_port, D(4) => RD_ex_4_port, D(3) => 
                           RD_ex_3_port, D(2) => RD_ex_2_port, D(1) => 
                           RD_ex_1_port, D(0) => RD_ex_0_port, Q(4) => 
                           RD_mem_4_port, Q(3) => RD_mem_3_port, Q(2) => 
                           RD_mem_2_port, Q(1) => RD_mem_1_port, Q(0) => 
                           RD_mem_0_port);
   pipeline_wr_signal2 : FF_4 port map( CLK => CLK, RESET => RST, EN => 
                           X_Logic1_port, D => wr_signal_exe, Q => 
                           wr_signal_mem);
   pipeline_IR3 : regFFD_NBIT6_1 port map( CK => CLK, RESET => RST, ENABLE => 
                           X_Logic1_port, D(5) => IR_26_ex_5_port, D(4) => 
                           IR_26_ex_4_port, D(3) => IR_26_ex_3_port, D(2) => 
                           IR_26_ex_2_port, D(1) => IR_26_ex_1_port, D(0) => 
                           IR_26_ex_0_port, Q(5) => IR_26_mem_5_port, Q(4) => 
                           IR_26_mem_4_port, Q(3) => IR_26_mem_3_port, Q(2) => 
                           IR_26_mem_2_port, Q(1) => IR_26_mem_1_port, Q(0) => 
                           IR_26_mem_0_port);
   MUX_PC : MUX21_GENERIC_NBIT32_3 port map( A(31) => ALU_ex_31_port, A(30) => 
                           ALU_ex_30_port, A(29) => ALU_ex_29_port, A(28) => 
                           ALU_ex_28_port, A(27) => ALU_ex_27_port, A(26) => 
                           ALU_ex_26_port, A(25) => ALU_ex_25_port, A(24) => 
                           ALU_ex_24_port, A(23) => ALU_ex_23_port, A(22) => 
                           ALU_ex_22_port, A(21) => ALU_ex_21_port, A(20) => 
                           ALU_ex_20_port, A(19) => ALU_ex_19_port, A(18) => 
                           ALU_ex_18_port, A(17) => ALU_ex_17_port, A(16) => 
                           ALU_ex_16_port, A(15) => ALU_ex_15_port, A(14) => 
                           ALU_ex_14_port, A(13) => ALU_ex_13_port, A(12) => 
                           ALU_ex_12_port, A(11) => ALU_ex_11_port, A(10) => 
                           ALU_ex_10_port, A(9) => ALU_ex_9_port, A(8) => 
                           ALU_ex_8_port, A(7) => ALU_ex_7_port, A(6) => 
                           ALU_ex_6_port, A(5) => ALU_ex_5_port, A(4) => 
                           ALU_ex_4_port, A(3) => ALU_ex_3_port, A(2) => 
                           ALU_ex_2_port, A(1) => ALU_ex_1_port, A(0) => 
                           ALU_ex_0_port, B(31) => NPC_mem_31_port, B(30) => 
                           NPC_mem_30_port, B(29) => NPC_mem_29_port, B(28) => 
                           NPC_mem_28_port, B(27) => NPC_mem_27_port, B(26) => 
                           NPC_mem_26_port, B(25) => NPC_mem_25_port, B(24) => 
                           NPC_mem_24_port, B(23) => NPC_mem_23_port, B(22) => 
                           NPC_mem_22_port, B(21) => NPC_mem_21_port, B(20) => 
                           NPC_mem_20_port, B(19) => NPC_mem_19_port, B(18) => 
                           NPC_mem_18_port, B(17) => NPC_mem_17_port, B(16) => 
                           NPC_mem_16_port, B(15) => NPC_mem_15_port, B(14) => 
                           NPC_mem_14_port, B(13) => NPC_mem_13_port, B(12) => 
                           NPC_mem_12_port, B(11) => NPC_mem_11_port, B(10) => 
                           NPC_mem_10_port, B(9) => NPC_mem_9_port, B(8) => 
                           NPC_mem_8_port, B(7) => NPC_mem_7_port, B(6) => 
                           NPC_mem_6_port, B(5) => NPC_mem_5_port, B(4) => 
                           NPC_mem_4_port, B(3) => NPC_mem_3_port, B(2) => 
                           NPC_mem_2_port, B(1) => NPC_mem_1_port, B(0) => 
                           NPC_mem_0_port, SEL => sel_npc, Y(31) => 
                           PC_OUT_i_31_port, Y(30) => PC_OUT_i_30_port, Y(29) 
                           => PC_OUT_i_29_port, Y(28) => PC_OUT_i_28_port, 
                           Y(27) => PC_OUT_i_27_port, Y(26) => PC_OUT_i_26_port
                           , Y(25) => PC_OUT_i_25_port, Y(24) => 
                           PC_OUT_i_24_port, Y(23) => PC_OUT_i_23_port, Y(22) 
                           => PC_OUT_i_22_port, Y(21) => PC_OUT_i_21_port, 
                           Y(20) => PC_OUT_i_20_port, Y(19) => PC_OUT_i_19_port
                           , Y(18) => PC_OUT_i_18_port, Y(17) => 
                           PC_OUT_i_17_port, Y(16) => PC_OUT_i_16_port, Y(15) 
                           => PC_OUT_i_15_port, Y(14) => PC_OUT_i_14_port, 
                           Y(13) => PC_OUT_i_13_port, Y(12) => PC_OUT_i_12_port
                           , Y(11) => PC_OUT_i_11_port, Y(10) => 
                           PC_OUT_i_10_port, Y(9) => PC_OUT_i_9_port, Y(8) => 
                           PC_OUT_i_8_port, Y(7) => PC_OUT_i_7_port, Y(6) => 
                           PC_OUT_i_6_port, Y(5) => PC_OUT_i_5_port, Y(4) => 
                           PC_OUT_i_4_port, Y(3) => PC_OUT_i_3_port, Y(2) => 
                           PC_OUT_i_2_port, Y(1) => PC_OUT_i_1_port, Y(0) => 
                           PC_OUT_i_0_port);
   LOAD_DATA_OUT : load_data port map( data_in(31) => DATA_MEM_OUT(31), 
                           data_in(30) => DATA_MEM_OUT(30), data_in(29) => 
                           DATA_MEM_OUT(29), data_in(28) => DATA_MEM_OUT(28), 
                           data_in(27) => DATA_MEM_OUT(27), data_in(26) => 
                           DATA_MEM_OUT(26), data_in(25) => DATA_MEM_OUT(25), 
                           data_in(24) => DATA_MEM_OUT(24), data_in(23) => 
                           DATA_MEM_OUT(23), data_in(22) => DATA_MEM_OUT(22), 
                           data_in(21) => DATA_MEM_OUT(21), data_in(20) => 
                           DATA_MEM_OUT(20), data_in(19) => DATA_MEM_OUT(19), 
                           data_in(18) => DATA_MEM_OUT(18), data_in(17) => 
                           DATA_MEM_OUT(17), data_in(16) => DATA_MEM_OUT(16), 
                           data_in(15) => DATA_MEM_OUT(15), data_in(14) => 
                           DATA_MEM_OUT(14), data_in(13) => DATA_MEM_OUT(13), 
                           data_in(12) => DATA_MEM_OUT(12), data_in(11) => 
                           DATA_MEM_OUT(11), data_in(10) => DATA_MEM_OUT(10), 
                           data_in(9) => DATA_MEM_OUT(9), data_in(8) => 
                           DATA_MEM_OUT(8), data_in(7) => DATA_MEM_OUT(7), 
                           data_in(6) => DATA_MEM_OUT(6), data_in(5) => 
                           DATA_MEM_OUT(5), data_in(4) => DATA_MEM_OUT(4), 
                           data_in(3) => DATA_MEM_OUT(3), data_in(2) => 
                           DATA_MEM_OUT(2), data_in(1) => DATA_MEM_OUT(1), 
                           data_in(0) => DATA_MEM_OUT(0), signed_val => 
                           signed_op_mem, load_op => RM, load_type(1) => 
                           IR_26_mem_1_port, load_type(0) => IR_26_mem_0_port, 
                           data_out(31) => LMD_out_31_port, data_out(30) => 
                           LMD_out_30_port, data_out(29) => LMD_out_29_port, 
                           data_out(28) => LMD_out_28_port, data_out(27) => 
                           LMD_out_27_port, data_out(26) => LMD_out_26_port, 
                           data_out(25) => LMD_out_25_port, data_out(24) => 
                           LMD_out_24_port, data_out(23) => LMD_out_23_port, 
                           data_out(22) => LMD_out_22_port, data_out(21) => 
                           LMD_out_21_port, data_out(20) => LMD_out_20_port, 
                           data_out(19) => LMD_out_19_port, data_out(18) => 
                           LMD_out_18_port, data_out(17) => LMD_out_17_port, 
                           data_out(16) => LMD_out_16_port, data_out(15) => 
                           LMD_out_15_port, data_out(14) => LMD_out_14_port, 
                           data_out(13) => LMD_out_13_port, data_out(12) => 
                           LMD_out_12_port, data_out(11) => LMD_out_11_port, 
                           data_out(10) => LMD_out_10_port, data_out(9) => 
                           LMD_out_9_port, data_out(8) => LMD_out_8_port, 
                           data_out(7) => LMD_out_7_port, data_out(6) => 
                           LMD_out_6_port, data_out(5) => LMD_out_5_port, 
                           data_out(4) => LMD_out_4_port, data_out(3) => 
                           LMD_out_3_port, data_out(2) => LMD_out_2_port, 
                           data_out(1) => LMD_out_1_port, data_out(0) => 
                           LMD_out_0_port);
   pipeline_alu4 : regFFD_NBIT32_3 port map( CK => CLK, RESET => RST, ENABLE =>
                           X_Logic1_port, D(31) => ALU_ex_31_port, D(30) => 
                           ALU_ex_30_port, D(29) => ALU_ex_29_port, D(28) => 
                           ALU_ex_28_port, D(27) => ALU_ex_27_port, D(26) => 
                           ALU_ex_26_port, D(25) => ALU_ex_25_port, D(24) => 
                           ALU_ex_24_port, D(23) => ALU_ex_23_port, D(22) => 
                           ALU_ex_22_port, D(21) => ALU_ex_21_port, D(20) => 
                           ALU_ex_20_port, D(19) => ALU_ex_19_port, D(18) => 
                           ALU_ex_18_port, D(17) => ALU_ex_17_port, D(16) => 
                           ALU_ex_16_port, D(15) => ALU_ex_15_port, D(14) => 
                           ALU_ex_14_port, D(13) => ALU_ex_13_port, D(12) => 
                           ALU_ex_12_port, D(11) => ALU_ex_11_port, D(10) => 
                           ALU_ex_10_port, D(9) => ALU_ex_9_port, D(8) => 
                           ALU_ex_8_port, D(7) => ALU_ex_7_port, D(6) => 
                           ALU_ex_6_port, D(5) => ALU_ex_5_port, D(4) => 
                           ALU_ex_4_port, D(3) => ALU_ex_3_port, D(2) => 
                           ALU_ex_2_port, D(1) => ALU_ex_1_port, D(0) => 
                           ALU_ex_0_port, Q(31) => ALU_wb_31_port, Q(30) => 
                           ALU_wb_30_port, Q(29) => ALU_wb_29_port, Q(28) => 
                           ALU_wb_28_port, Q(27) => ALU_wb_27_port, Q(26) => 
                           ALU_wb_26_port, Q(25) => ALU_wb_25_port, Q(24) => 
                           ALU_wb_24_port, Q(23) => ALU_wb_23_port, Q(22) => 
                           ALU_wb_22_port, Q(21) => ALU_wb_21_port, Q(20) => 
                           ALU_wb_20_port, Q(19) => ALU_wb_19_port, Q(18) => 
                           ALU_wb_18_port, Q(17) => ALU_wb_17_port, Q(16) => 
                           ALU_wb_16_port, Q(15) => ALU_wb_15_port, Q(14) => 
                           ALU_wb_14_port, Q(13) => ALU_wb_13_port, Q(12) => 
                           ALU_wb_12_port, Q(11) => ALU_wb_11_port, Q(10) => 
                           ALU_wb_10_port, Q(9) => ALU_wb_9_port, Q(8) => 
                           ALU_wb_8_port, Q(7) => ALU_wb_7_port, Q(6) => 
                           ALU_wb_6_port, Q(5) => ALU_wb_5_port, Q(4) => 
                           ALU_wb_4_port, Q(3) => ALU_wb_3_port, Q(2) => 
                           ALU_wb_2_port, Q(1) => ALU_wb_1_port, Q(0) => 
                           ALU_wb_0_port);
   pipeline_LMD4 : regFFD_NBIT32_2 port map( CK => CLK, RESET => RST, ENABLE =>
                           RM, D(31) => LMD_out_31_port, D(30) => 
                           LMD_out_30_port, D(29) => LMD_out_29_port, D(28) => 
                           LMD_out_28_port, D(27) => LMD_out_27_port, D(26) => 
                           LMD_out_26_port, D(25) => LMD_out_25_port, D(24) => 
                           LMD_out_24_port, D(23) => LMD_out_23_port, D(22) => 
                           LMD_out_22_port, D(21) => LMD_out_21_port, D(20) => 
                           LMD_out_20_port, D(19) => LMD_out_19_port, D(18) => 
                           LMD_out_18_port, D(17) => LMD_out_17_port, D(16) => 
                           LMD_out_16_port, D(15) => LMD_out_15_port, D(14) => 
                           LMD_out_14_port, D(13) => LMD_out_13_port, D(12) => 
                           LMD_out_12_port, D(11) => LMD_out_11_port, D(10) => 
                           LMD_out_10_port, D(9) => LMD_out_9_port, D(8) => 
                           LMD_out_8_port, D(7) => LMD_out_7_port, D(6) => 
                           LMD_out_6_port, D(5) => LMD_out_5_port, D(4) => 
                           LMD_out_4_port, D(3) => LMD_out_3_port, D(2) => 
                           LMD_out_2_port, D(1) => LMD_out_1_port, D(0) => 
                           LMD_out_0_port, Q(31) => LMD_wb_31_port, Q(30) => 
                           LMD_wb_30_port, Q(29) => LMD_wb_29_port, Q(28) => 
                           LMD_wb_28_port, Q(27) => LMD_wb_27_port, Q(26) => 
                           LMD_wb_26_port, Q(25) => LMD_wb_25_port, Q(24) => 
                           LMD_wb_24_port, Q(23) => LMD_wb_23_port, Q(22) => 
                           LMD_wb_22_port, Q(21) => LMD_wb_21_port, Q(20) => 
                           LMD_wb_20_port, Q(19) => LMD_wb_19_port, Q(18) => 
                           LMD_wb_18_port, Q(17) => LMD_wb_17_port, Q(16) => 
                           LMD_wb_16_port, Q(15) => LMD_wb_15_port, Q(14) => 
                           LMD_wb_14_port, Q(13) => LMD_wb_13_port, Q(12) => 
                           LMD_wb_12_port, Q(11) => LMD_wb_11_port, Q(10) => 
                           LMD_wb_10_port, Q(9) => LMD_wb_9_port, Q(8) => 
                           LMD_wb_8_port, Q(7) => LMD_wb_7_port, Q(6) => 
                           LMD_wb_6_port, Q(5) => LMD_wb_5_port, Q(4) => 
                           LMD_wb_4_port, Q(3) => LMD_wb_3_port, Q(2) => 
                           LMD_wb_2_port, Q(1) => LMD_wb_1_port, Q(0) => 
                           LMD_wb_0_port);
   pipeline_RD4 : regFFD_NBIT5_1 port map( CK => CLK, RESET => RST, ENABLE => 
                           X_Logic1_port, D(4) => RD_mem_4_port, D(3) => 
                           RD_mem_3_port, D(2) => RD_mem_2_port, D(1) => 
                           RD_mem_1_port, D(0) => RD_mem_0_port, Q(4) => 
                           RD_wb_4_port, Q(3) => RD_wb_3_port, Q(2) => 
                           RD_wb_2_port, Q(1) => RD_wb_1_port, Q(0) => 
                           RD_wb_0_port);
   pipeline_wr_signal3 : FF_3 port map( CLK => CLK, RESET => RST, EN => 
                           X_Logic1_port, D => wr_signal_mem1, Q => 
                           wr_signal_wb);
   pipeline_WM : FF_2 port map( CLK => CLK, RESET => RST, EN => X_Logic1_port, 
                           D => WM, Q => n_2276);
   pipeline_JAL : FF_1 port map( CLK => CLK, RESET => RST, EN => X_Logic1_port,
                           D => sel_saved_reg, Q => sel_saved_reg_wb);
   pipeline_NPC_wb : regFFD_NBIT32_1 port map( CK => CLK, RESET => RST, ENABLE 
                           => X_Logic1_port, D(31) => NPC_mem_31_port, D(30) =>
                           NPC_mem_30_port, D(29) => NPC_mem_29_port, D(28) => 
                           NPC_mem_28_port, D(27) => NPC_mem_27_port, D(26) => 
                           NPC_mem_26_port, D(25) => NPC_mem_25_port, D(24) => 
                           NPC_mem_24_port, D(23) => NPC_mem_23_port, D(22) => 
                           NPC_mem_22_port, D(21) => NPC_mem_21_port, D(20) => 
                           NPC_mem_20_port, D(19) => NPC_mem_19_port, D(18) => 
                           NPC_mem_18_port, D(17) => NPC_mem_17_port, D(16) => 
                           NPC_mem_16_port, D(15) => NPC_mem_15_port, D(14) => 
                           NPC_mem_14_port, D(13) => NPC_mem_13_port, D(12) => 
                           NPC_mem_12_port, D(11) => NPC_mem_11_port, D(10) => 
                           NPC_mem_10_port, D(9) => NPC_mem_9_port, D(8) => 
                           NPC_mem_8_port, D(7) => NPC_mem_7_port, D(6) => 
                           NPC_mem_6_port, D(5) => NPC_mem_5_port, D(4) => 
                           NPC_mem_4_port, D(3) => NPC_mem_3_port, D(2) => 
                           NPC_mem_2_port, D(1) => NPC_mem_1_port, D(0) => 
                           NPC_mem_0_port, Q(31) => NPC_wb_31_port, Q(30) => 
                           NPC_wb_30_port, Q(29) => NPC_wb_29_port, Q(28) => 
                           NPC_wb_28_port, Q(27) => NPC_wb_27_port, Q(26) => 
                           NPC_wb_26_port, Q(25) => NPC_wb_25_port, Q(24) => 
                           NPC_wb_24_port, Q(23) => NPC_wb_23_port, Q(22) => 
                           NPC_wb_22_port, Q(21) => NPC_wb_21_port, Q(20) => 
                           NPC_wb_20_port, Q(19) => NPC_wb_19_port, Q(18) => 
                           NPC_wb_18_port, Q(17) => NPC_wb_17_port, Q(16) => 
                           NPC_wb_16_port, Q(15) => NPC_wb_15_port, Q(14) => 
                           NPC_wb_14_port, Q(13) => NPC_wb_13_port, Q(12) => 
                           NPC_wb_12_port, Q(11) => NPC_wb_11_port, Q(10) => 
                           NPC_wb_10_port, Q(9) => NPC_wb_9_port, Q(8) => 
                           NPC_wb_8_port, Q(7) => NPC_wb_7_port, Q(6) => 
                           NPC_wb_6_port, Q(5) => NPC_wb_5_port, Q(4) => 
                           NPC_wb_4_port, Q(3) => NPC_wb_3_port, Q(2) => 
                           NPC_wb_2_port, Q(1) => NPC_wb_1_port, Q(0) => 
                           NPC_wb_0_port);
   MUX_WB : MUX21_GENERIC_NBIT32_2 port map( A(31) => ALU_wb_31_port, A(30) => 
                           ALU_wb_30_port, A(29) => ALU_wb_29_port, A(28) => 
                           ALU_wb_28_port, A(27) => ALU_wb_27_port, A(26) => 
                           ALU_wb_26_port, A(25) => ALU_wb_25_port, A(24) => 
                           ALU_wb_24_port, A(23) => ALU_wb_23_port, A(22) => 
                           ALU_wb_22_port, A(21) => ALU_wb_21_port, A(20) => 
                           ALU_wb_20_port, A(19) => ALU_wb_19_port, A(18) => 
                           ALU_wb_18_port, A(17) => ALU_wb_17_port, A(16) => 
                           ALU_wb_16_port, A(15) => ALU_wb_15_port, A(14) => 
                           ALU_wb_14_port, A(13) => ALU_wb_13_port, A(12) => 
                           ALU_wb_12_port, A(11) => ALU_wb_11_port, A(10) => 
                           ALU_wb_10_port, A(9) => ALU_wb_9_port, A(8) => 
                           ALU_wb_8_port, A(7) => ALU_wb_7_port, A(6) => 
                           ALU_wb_6_port, A(5) => ALU_wb_5_port, A(4) => 
                           ALU_wb_4_port, A(3) => ALU_wb_3_port, A(2) => 
                           ALU_wb_2_port, A(1) => ALU_wb_1_port, A(0) => 
                           ALU_wb_0_port, B(31) => LMD_wb_31_port, B(30) => 
                           LMD_wb_30_port, B(29) => LMD_wb_29_port, B(28) => 
                           LMD_wb_28_port, B(27) => LMD_wb_27_port, B(26) => 
                           LMD_wb_26_port, B(25) => LMD_wb_25_port, B(24) => 
                           LMD_wb_24_port, B(23) => LMD_wb_23_port, B(22) => 
                           LMD_wb_22_port, B(21) => LMD_wb_21_port, B(20) => 
                           LMD_wb_20_port, B(19) => LMD_wb_19_port, B(18) => 
                           LMD_wb_18_port, B(17) => LMD_wb_17_port, B(16) => 
                           LMD_wb_16_port, B(15) => LMD_wb_15_port, B(14) => 
                           LMD_wb_14_port, B(13) => LMD_wb_13_port, B(12) => 
                           LMD_wb_12_port, B(11) => LMD_wb_11_port, B(10) => 
                           LMD_wb_10_port, B(9) => LMD_wb_9_port, B(8) => 
                           LMD_wb_8_port, B(7) => LMD_wb_7_port, B(6) => 
                           LMD_wb_6_port, B(5) => LMD_wb_5_port, B(4) => 
                           LMD_wb_4_port, B(3) => LMD_wb_3_port, B(2) => 
                           LMD_wb_2_port, B(1) => LMD_wb_1_port, B(0) => 
                           LMD_wb_0_port, SEL => S3, Y(31) => OUT_data_31_port,
                           Y(30) => OUT_data_30_port, Y(29) => OUT_data_29_port
                           , Y(28) => OUT_data_28_port, Y(27) => 
                           OUT_data_27_port, Y(26) => OUT_data_26_port, Y(25) 
                           => OUT_data_25_port, Y(24) => OUT_data_24_port, 
                           Y(23) => OUT_data_23_port, Y(22) => OUT_data_22_port
                           , Y(21) => OUT_data_21_port, Y(20) => 
                           OUT_data_20_port, Y(19) => OUT_data_19_port, Y(18) 
                           => OUT_data_18_port, Y(17) => OUT_data_17_port, 
                           Y(16) => OUT_data_16_port, Y(15) => OUT_data_15_port
                           , Y(14) => OUT_data_14_port, Y(13) => 
                           OUT_data_13_port, Y(12) => OUT_data_12_port, Y(11) 
                           => OUT_data_11_port, Y(10) => OUT_data_10_port, Y(9)
                           => OUT_data_9_port, Y(8) => OUT_data_8_port, Y(7) =>
                           OUT_data_7_port, Y(6) => OUT_data_6_port, Y(5) => 
                           OUT_data_5_port, Y(4) => OUT_data_4_port, Y(3) => 
                           OUT_data_3_port, Y(2) => OUT_data_2_port, Y(1) => 
                           OUT_data_1_port, Y(0) => OUT_data_0_port);
   MUX_jal : MUX21_GENERIC_NBIT32_1 port map( A(31) => NPC_wb_31_port, A(30) =>
                           NPC_wb_30_port, A(29) => NPC_wb_29_port, A(28) => 
                           NPC_wb_28_port, A(27) => NPC_wb_27_port, A(26) => 
                           NPC_wb_26_port, A(25) => NPC_wb_25_port, A(24) => 
                           NPC_wb_24_port, A(23) => NPC_wb_23_port, A(22) => 
                           NPC_wb_22_port, A(21) => NPC_wb_21_port, A(20) => 
                           NPC_wb_20_port, A(19) => NPC_wb_19_port, A(18) => 
                           NPC_wb_18_port, A(17) => NPC_wb_17_port, A(16) => 
                           NPC_wb_16_port, A(15) => NPC_wb_15_port, A(14) => 
                           NPC_wb_14_port, A(13) => NPC_wb_13_port, A(12) => 
                           NPC_wb_12_port, A(11) => NPC_wb_11_port, A(10) => 
                           NPC_wb_10_port, A(9) => NPC_wb_9_port, A(8) => 
                           NPC_wb_8_port, A(7) => NPC_wb_7_port, A(6) => 
                           NPC_wb_6_port, A(5) => NPC_wb_5_port, A(4) => 
                           NPC_wb_4_port, A(3) => NPC_wb_3_port, A(2) => 
                           NPC_wb_2_port, A(1) => NPC_wb_1_port, A(0) => 
                           NPC_wb_0_port, B(31) => OUT_data_31_port, B(30) => 
                           OUT_data_30_port, B(29) => OUT_data_29_port, B(28) 
                           => OUT_data_28_port, B(27) => OUT_data_27_port, 
                           B(26) => OUT_data_26_port, B(25) => OUT_data_25_port
                           , B(24) => OUT_data_24_port, B(23) => 
                           OUT_data_23_port, B(22) => OUT_data_22_port, B(21) 
                           => OUT_data_21_port, B(20) => OUT_data_20_port, 
                           B(19) => OUT_data_19_port, B(18) => OUT_data_18_port
                           , B(17) => OUT_data_17_port, B(16) => 
                           OUT_data_16_port, B(15) => OUT_data_15_port, B(14) 
                           => OUT_data_14_port, B(13) => OUT_data_13_port, 
                           B(12) => OUT_data_12_port, B(11) => OUT_data_11_port
                           , B(10) => OUT_data_10_port, B(9) => OUT_data_9_port
                           , B(8) => OUT_data_8_port, B(7) => OUT_data_7_port, 
                           B(6) => OUT_data_6_port, B(5) => OUT_data_5_port, 
                           B(4) => OUT_data_4_port, B(3) => OUT_data_3_port, 
                           B(2) => OUT_data_2_port, B(1) => OUT_data_1_port, 
                           B(0) => OUT_data_0_port, SEL => sel_saved_reg_wb, 
                           Y(31) => n_2277, Y(30) => n_2278, Y(29) => n_2279, 
                           Y(28) => n_2280, Y(27) => n_2281, Y(26) => n_2282, 
                           Y(25) => n_2283, Y(24) => n_2284, Y(23) => n_2285, 
                           Y(22) => n_2286, Y(21) => n_2287, Y(20) => n_2288, 
                           Y(19) => n_2289, Y(18) => n_2290, Y(17) => n_2291, 
                           Y(16) => n_2292, Y(15) => n_2293, Y(14) => n_2294, 
                           Y(13) => n_2295, Y(12) => n_2296, Y(11) => n_2297, 
                           Y(10) => n_2298, Y(9) => n_2299, Y(8) => n_2300, 
                           Y(7) => n_2301, Y(6) => n_2302, Y(5) => n_2303, Y(4)
                           => n_2304, Y(3) => n_2305, Y(2) => n_2306, Y(1) => 
                           n_2307, Y(0) => n_2308);
   add_254 : DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 port map( A(31) => 
                           PC_fetch0_31_port, A(30) => PC_fetch0_30_port, A(29)
                           => PC_fetch0_29_port, A(28) => PC_fetch0_28_port, 
                           A(27) => PC_fetch0_27_port, A(26) => 
                           PC_fetch0_26_port, A(25) => PC_fetch0_25_port, A(24)
                           => PC_fetch0_24_port, A(23) => PC_fetch0_23_port, 
                           A(22) => PC_fetch0_22_port, A(21) => 
                           PC_fetch0_21_port, A(20) => PC_fetch0_20_port, A(19)
                           => PC_fetch0_19_port, A(18) => PC_fetch0_18_port, 
                           A(17) => PC_fetch0_17_port, A(16) => 
                           PC_fetch0_16_port, A(15) => PC_fetch0_15_port, A(14)
                           => PC_fetch0_14_port, A(13) => PC_fetch0_13_port, 
                           A(12) => PC_fetch0_12_port, A(11) => 
                           PC_fetch0_11_port, A(10) => PC_fetch0_10_port, A(9) 
                           => PC_fetch0_9_port, A(8) => PC_fetch0_8_port, A(7) 
                           => PC_fetch0_7_port, A(6) => PC_fetch0_6_port, A(5) 
                           => PC_fetch0_5_port, A(4) => PC_fetch0_4_port, A(3) 
                           => PC_fetch0_3_port, A(2) => PC_fetch0_2_port, A(1) 
                           => PC_fetch0_1_port, A(0) => PC_fetch0_0_port, 
                           SUM(31) => NPC_31_port, SUM(30) => NPC_30_port, 
                           SUM(29) => NPC_29_port, SUM(28) => NPC_28_port, 
                           SUM(27) => NPC_27_port, SUM(26) => NPC_26_port, 
                           SUM(25) => NPC_25_port, SUM(24) => NPC_24_port, 
                           SUM(23) => NPC_23_port, SUM(22) => NPC_22_port, 
                           SUM(21) => NPC_21_port, SUM(20) => NPC_20_port, 
                           SUM(19) => NPC_19_port, SUM(18) => NPC_18_port, 
                           SUM(17) => NPC_17_port, SUM(16) => NPC_16_port, 
                           SUM(15) => NPC_15_port, SUM(14) => NPC_14_port, 
                           SUM(13) => NPC_13_port, SUM(12) => NPC_12_port, 
                           SUM(11) => NPC_11_port, SUM(10) => NPC_10_port, 
                           SUM(9) => NPC_9_port, SUM(8) => NPC_8_port, SUM(7) 
                           => NPC_7_port, SUM(6) => NPC_6_port, SUM(5) => 
                           NPC_5_port, SUM(4) => NPC_4_port, SUM(3) => 
                           NPC_3_port, SUM(2) => NPC_2_port, SUM(1) => 
                           NPC_1_port, SUM(0) => NPC_0_port);
   U80 : CLKBUF_X1 port map( A => IR_Dec_26_port, Z => n40);
   U81 : CLKBUF_X1 port map( A => IR_Dec_30_port, Z => n41);
   U82 : CLKBUF_X1 port map( A => IR_Dec_31_port, Z => n42);
   U83 : INV_X1 port map( A => n8, ZN => n43);
   U84 : INV_X1 port map( A => n8, ZN => n44);
   U85 : CLKBUF_X1 port map( A => IR_Dec_29_port, Z => n45);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
         std_logic;  ALU_OPCODE : out std_logic_vector (0 to 5);  
         signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
         WB_MUX_SEL, RF_WE, lhi_sel, sb_op : out std_logic);

end dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3, aluOpcode1_5_port, aluOpcode1_4_port, aluOpcode1_3_port, 
      aluOpcode1_2_port, aluOpcode1_1_port, aluOpcode1_0_port, 
      aluOpcode2_5_port, aluOpcode2_4_port, aluOpcode2_3_port, 
      aluOpcode2_2_port, aluOpcode2_1_port, aluOpcode2_0_port, 
      aluOpcode_i_5_port, aluOpcode_i_4_port, aluOpcode_i_3_port, 
      aluOpcode_i_2_port, aluOpcode_i_1_port, aluOpcode_i_0_port, 
      signed_unsigned_i, N393, N394, n9, n10, n11, n12, n13, n14, n15, n16, n17
      , n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n145, n146, n147, n148, n149, n150, n1, n_2309, 
      n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, 
      n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327 : 
      std_logic;

begin
   
   aluOpcode1_reg_5_inst : DFFR_X1 port map( D => aluOpcode_i_5_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_5_port, QN => n_2309);
   aluOpcode1_reg_4_inst : DFFR_X1 port map( D => aluOpcode_i_4_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_4_port, QN => n_2310);
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_3_port, QN => n_2311);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_2_port, QN => n_2312);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_1_port, QN => n_2313);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_0_port, QN => n_2314);
   aluOpcode2_reg_5_inst : DFFR_X1 port map( D => aluOpcode1_5_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_5_port, QN => n_2315);
   aluOpcode2_reg_4_inst : DFFR_X1 port map( D => aluOpcode1_4_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_4_port, QN => n_2316);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => aluOpcode1_3_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_3_port, QN => n_2317);
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => aluOpcode1_2_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_2_port, QN => n_2318);
   aluOpcode2_reg_1_inst : DFFR_X1 port map( D => aluOpcode1_1_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_1_port, QN => n_2319);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => aluOpcode1_0_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_0_port, QN => n_2320);
   aluOpcode3_reg_5_inst : DFFR_X1 port map( D => aluOpcode2_5_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(0), QN => n_2321);
   aluOpcode3_reg_4_inst : DFFR_X1 port map( D => aluOpcode2_4_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(1), QN => n_2322);
   aluOpcode3_reg_3_inst : DFFR_X1 port map( D => aluOpcode2_3_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(2), QN => n_2323);
   aluOpcode3_reg_2_inst : DFFR_X1 port map( D => aluOpcode2_2_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(3), QN => n_2324);
   aluOpcode3_reg_1_inst : DFFR_X1 port map( D => aluOpcode2_1_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(4), QN => n_2325);
   aluOpcode3_reg_0_inst : DFFR_X1 port map( D => aluOpcode2_0_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(5), QN => n_2326);
   signed_unsigned_i_reg : DLH_X1 port map( G => N393, D => N394, Q => 
                           signed_unsigned_i);
   signed_unsigned_2_reg : DFF_X1 port map( D => n149, CK => Clk, Q => 
                           signed_unsigned, QN => n145);
   lhi_sel_reg : DFF_X1 port map( D => n148, CK => Clk, Q => n3, QN => n143);
   sb_op_reg : DFF_X1 port map( D => n147, CK => Clk, Q => sb_op, QN => n146);
   U3 : NOR2_X1 port map( A1 => Rst, A2 => n146, ZN => n147);
   U4 : NOR2_X1 port map( A1 => n143, A2 => Rst, ZN => n148);
   U5 : OAI22_X1 port map( A1 => n9, A2 => n10, B1 => Rst, B2 => n145, ZN => 
                           n149);
   U6 : INV_X1 port map( A => Rst, ZN => n9);
   U7 : OAI21_X1 port map( B1 => Rst, B2 => n10, A => n11, ZN => n150);
   U8 : NAND2_X1 port map( A1 => signed_unsigned_i, A2 => Rst, ZN => n11);
   U10 : OAI211_X1 port map( C1 => n12, C2 => n13, A => n14, B => n15, ZN => 
                           aluOpcode_i_5_port);
   U11 : INV_X1 port map( A => n16, ZN => n15);
   U12 : OAI211_X1 port map( C1 => n17, C2 => n18, A => n19, B => n20, ZN => 
                           n16);
   U13 : AND3_X1 port map( A1 => n21, A2 => n22, A3 => n23, ZN => n18);
   U14 : NAND3_X1 port map( A1 => IR_IN(0), A2 => n24, A3 => IR_IN(1), ZN => 
                           n22);
   U15 : OAI211_X1 port map( C1 => n25, C2 => n17, A => n26, B => n27, ZN => 
                           aluOpcode_i_4_port);
   U16 : OAI211_X1 port map( C1 => n28, C2 => n17, A => n14, B => n29, ZN => 
                           aluOpcode_i_3_port);
   U17 : NOR2_X1 port map( A1 => n30, A2 => n31, ZN => n29);
   U18 : NOR3_X1 port map( A1 => n32, A2 => n33, A3 => n34, ZN => n28);
   U19 : INV_X1 port map( A => n25, ZN => n33);
   U20 : NOR2_X1 port map( A1 => n35, A2 => n36, ZN => n25);
   U21 : INV_X1 port map( A => n37, ZN => n36);
   U22 : OAI21_X1 port map( B1 => n38, B2 => n39, A => n40, ZN => n32);
   U23 : NAND3_X1 port map( A1 => n41, A2 => n42, A3 => n43, ZN => 
                           aluOpcode_i_2_port);
   U24 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U25 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => n47);
   U26 : AOI21_X1 port map( B1 => n51, B2 => n52, A => n53, ZN => n41);
   U27 : OAI211_X1 port map( C1 => n54, C2 => n17, A => n55, B => n56, ZN => 
                           aluOpcode_i_1_port);
   U28 : AOI221_X1 port map( B1 => n51, B2 => n57, C1 => n58, C2 => n59, A => 
                           n60, ZN => n56);
   U29 : NOR2_X1 port map( A1 => n61, A2 => n62, ZN => n55);
   U30 : AOI21_X1 port map( B1 => n13, B2 => n63, A => n64, ZN => n62);
   U31 : AND3_X1 port map( A1 => n65, A2 => n66, A3 => n67, ZN => n54);
   U32 : NAND3_X1 port map( A1 => n68, A2 => n69, A3 => n70, ZN => 
                           aluOpcode_i_0_port);
   U33 : AOI211_X1 port map( C1 => n51, C2 => n45, A => n60, B => n71, ZN => 
                           n70);
   U34 : OAI211_X1 port map( C1 => n72, C2 => n13, A => n73, B => n74, ZN => 
                           n60);
   U35 : NOR2_X1 port map( A1 => n48, A2 => n75, ZN => n74);
   U36 : NOR3_X1 port map( A1 => n76, A2 => IR_IN(29), A3 => n64, ZN => n75);
   U37 : INV_X1 port map( A => n57, ZN => n72);
   U38 : INV_X1 port map( A => n77, ZN => n51);
   U39 : AOI21_X1 port map( B1 => n46, B2 => n78, A => n79, ZN => n69);
   U40 : NAND4_X1 port map( A1 => n80, A2 => n81, A3 => n82, A4 => n83, ZN => 
                           n78);
   U41 : AND4_X1 port map( A1 => n21, A2 => n84, A3 => n37, A4 => n85, ZN => 
                           n83);
   U42 : OAI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n82);
   U43 : OAI21_X1 port map( B1 => n89, B2 => n87, A => n90, ZN => n80);
   U44 : INV_X1 port map( A => n38, ZN => n87);
   U45 : NOR2_X1 port map( A1 => n91, A2 => n24, ZN => n38);
   U46 : AOI22_X1 port map( A1 => n92, A2 => n52, B1 => n58, B2 => n93, ZN => 
                           n68);
   U47 : INV_X1 port map( A => n94, ZN => n92);
   U48 : OAI211_X1 port map( C1 => n95, C2 => n96, A => n27, B => n73, ZN => 
                           N394);
   U49 : INV_X1 port map( A => n97, ZN => n73);
   U50 : OAI21_X1 port map( B1 => n64, B2 => n98, A => n99, ZN => n97);
   U51 : AOI22_X1 port map( A1 => n100, A2 => n45, B1 => n93, B2 => IR_IN(30), 
                           ZN => n95);
   U52 : NOR2_X1 port map( A1 => IR_IN(30), A2 => n101, ZN => n100);
   U53 : NAND4_X1 port map( A1 => n42, A2 => n27, A3 => n102, A4 => n103, ZN =>
                           N393);
   U54 : AOI211_X1 port map( C1 => n104, C2 => n57, A => n105, B => n106, ZN =>
                           n103);
   U55 : NAND2_X1 port map( A1 => n77, A2 => n13, ZN => n105);
   U56 : AOI21_X1 port map( B1 => n46, B2 => n107, A => n108, ZN => n102);
   U57 : INV_X1 port map( A => n14, ZN => n108);
   U58 : AOI211_X1 port map( C1 => n57, C2 => n58, A => n109, B => n53, ZN => 
                           n14);
   U59 : NAND2_X1 port map( A1 => n99, A2 => n110, ZN => n53);
   U60 : OR3_X1 port map( A1 => n111, A2 => n112, A3 => n94, ZN => n110);
   U61 : NAND3_X1 port map( A1 => n113, A2 => n114, A3 => n93, ZN => n99);
   U62 : AOI21_X1 port map( B1 => n76, B2 => n115, A => n64, ZN => n109);
   U63 : NAND2_X1 port map( A1 => n12, A2 => n116, ZN => n57);
   U64 : NAND4_X1 port map( A1 => n101, A2 => n49, A3 => n67, A4 => n117, ZN =>
                           n107);
   U65 : INV_X1 port map( A => n24, ZN => n117);
   U66 : INV_X1 port map( A => n34, ZN => n67);
   U67 : NAND2_X1 port map( A1 => n81, A2 => n118, ZN => n34);
   U68 : NAND3_X1 port map( A1 => n119, A2 => IR_IN(3), A3 => n120, ZN => n118)
                           ;
   U69 : NAND3_X1 port map( A1 => n90, A2 => IR_IN(3), A3 => n119, ZN => n81);
   U70 : AOI21_X1 port map( B1 => n121, B2 => n91, A => n35, ZN => n49);
   U71 : NAND2_X1 port map( A1 => n85, A2 => n66, ZN => n35);
   U72 : OAI21_X1 port map( B1 => n120, B2 => n88, A => n24, ZN => n66);
   U73 : NOR4_X1 port map( A1 => n122, A2 => n123, A3 => IR_IN(2), A4 => 
                           IR_IN(4), ZN => n24);
   U74 : NAND3_X1 port map( A1 => IR_IN(1), A2 => IR_IN(0), A3 => n86, ZN => 
                           n85);
   U75 : AND4_X1 port map( A1 => n65, A2 => n40, A3 => n37, A4 => n21, ZN => 
                           n101);
   U76 : NAND3_X1 port map( A1 => n124, A2 => n125, A3 => n88, ZN => n21);
   U77 : NAND2_X1 port map( A1 => n91, A2 => IR_IN(0), ZN => n37);
   U78 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => n40);
   U79 : AOI211_X1 port map( C1 => n121, C2 => n86, A => n126, B => n127, ZN =>
                           n65);
   U80 : OAI21_X1 port map( B1 => n128, B2 => n39, A => n23, ZN => n127);
   U81 : AND2_X1 port map( A1 => n84, A2 => n129, ZN => n23);
   U82 : NAND4_X1 port map( A1 => n124, A2 => IR_IN(1), A3 => IR_IN(0), A4 => 
                           n125, ZN => n129);
   U83 : NAND3_X1 port map( A1 => n90, A2 => n124, A3 => IR_IN(2), ZN => n84);
   U84 : AND3_X1 port map( A1 => IR_IN(5), A2 => IR_IN(3), A3 => IR_IN(4), ZN 
                           => n124);
   U85 : INV_X1 port map( A => n91, ZN => n128);
   U86 : NOR4_X1 port map( A1 => n122, A2 => IR_IN(2), A3 => IR_IN(3), A4 => 
                           IR_IN(4), ZN => n91);
   U87 : INV_X1 port map( A => n50, ZN => n126);
   U88 : OAI21_X1 port map( B1 => n120, B2 => n90, A => n89, ZN => n50);
   U89 : AND2_X1 port map( A1 => n119, A2 => n123, ZN => n89);
   U90 : INV_X1 port map( A => IR_IN(3), ZN => n123);
   U91 : NOR3_X1 port map( A1 => n122, A2 => IR_IN(4), A3 => n125, ZN => n119);
   U92 : INV_X1 port map( A => IR_IN(5), ZN => n122);
   U93 : INV_X1 port map( A => n39, ZN => n90);
   U94 : NAND2_X1 port map( A1 => IR_IN(0), A2 => n130, ZN => n39);
   U95 : NOR4_X1 port map( A1 => n125, A2 => IR_IN(3), A3 => IR_IN(4), A4 => 
                           IR_IN(5), ZN => n86);
   U96 : INV_X1 port map( A => IR_IN(2), ZN => n125);
   U97 : OR2_X1 port map( A1 => n88, A2 => n120, ZN => n121);
   U98 : NOR2_X1 port map( A1 => IR_IN(0), A2 => IR_IN(1), ZN => n120);
   U99 : NOR2_X1 port map( A1 => n130, A2 => IR_IN(0), ZN => n88);
   U100 : INV_X1 port map( A => IR_IN(1), ZN => n130);
   U101 : INV_X1 port map( A => n17, ZN => n46);
   U102 : NAND4_X1 port map( A1 => n104, A2 => n45, A3 => n131, A4 => n132, ZN 
                           => n17);
   U103 : NOR4_X1 port map( A1 => IR_IN(30), A2 => IR_IN(9), A3 => IR_IN(8), A4
                           => IR_IN(7), ZN => n132);
   U104 : NOR2_X1 port map( A1 => IR_IN(6), A2 => IR_IN(10), ZN => n131);
   U105 : INV_X1 port map( A => n96, ZN => n104);
   U106 : NAND3_X1 port map( A1 => n133, A2 => n111, A3 => n114, ZN => n96);
   U107 : AND4_X1 port map( A1 => n134, A2 => n19, A3 => n135, A4 => n136, ZN 
                           => n27);
   U108 : AOI211_X1 port map( C1 => n106, C2 => n52, A => n71, B => n30, ZN => 
                           n136);
   U109 : OAI22_X1 port map( A1 => n12, A2 => n63, B1 => n137, B2 => n77, ZN =>
                           n30);
   U110 : NOR2_X1 port map( A1 => n52, A2 => n59, ZN => n137);
   U111 : INV_X1 port map( A => n44, ZN => n63);
   U112 : NOR2_X1 port map( A1 => n76, A2 => n133, ZN => n44);
   U113 : OAI21_X1 port map( B1 => n116, B2 => n98, A => n20, ZN => n71);
   U114 : NAND3_X1 port map( A1 => n52, A2 => n113, A3 => IR_IN(28), ZN => n20)
                           ;
   U115 : INV_X1 port map( A => n98, ZN => n106);
   U116 : OAI21_X1 port map( B1 => n93, B2 => n45, A => n138, ZN => n135);
   U117 : INV_X1 port map( A => n116, ZN => n93);
   U118 : NAND3_X1 port map( A1 => n59, A2 => n114, A3 => n113, ZN => n19);
   U119 : NOR3_X1 port map( A1 => n139, A2 => n133, A3 => n111, ZN => n113);
   U120 : INV_X1 port map( A => n48, ZN => n134);
   U121 : NOR3_X1 port map( A1 => n12, A2 => IR_IN(29), A3 => n76, ZN => n48);
   U122 : NAND3_X1 port map( A1 => n114, A2 => n139, A3 => IR_IN(31), ZN => n76
                           );
   U123 : AOI211_X1 port map( C1 => n59, C2 => n138, A => n140, B => n31, ZN =>
                           n42);
   U124 : OAI222_X1 port map( A1 => n116, A2 => n77, B1 => n112, B2 => n94, C1 
                           => n64, C2 => n98, ZN => n31);
   U125 : NAND3_X1 port map( A1 => IR_IN(28), A2 => n139, A3 => n141, ZN => n98
                           );
   U126 : INV_X1 port map( A => n45, ZN => n64);
   U127 : NAND3_X1 port map( A1 => n133, A2 => n139, A3 => IR_IN(28), ZN => n94
                           );
   U128 : NOR2_X1 port map( A1 => n45, A2 => n52, ZN => n112);
   U129 : NAND3_X1 port map( A1 => n114, A2 => n139, A3 => n141, ZN => n77);
   U130 : INV_X1 port map( A => IR_IN(30), ZN => n139);
   U131 : NAND2_X1 port map( A1 => IR_IN(27), A2 => n142, ZN => n116);
   U132 : INV_X1 port map( A => n26, ZN => n140);
   U133 : AOI211_X1 port map( C1 => n52, C2 => n58, A => n79, B => n61, ZN => 
                           n26);
   U134 : AND4_X1 port map( A1 => n141, A2 => IR_IN(28), A3 => n52, A4 => 
                           IR_IN(30), ZN => n61);
   U135 : AND4_X1 port map( A1 => n45, A2 => n141, A3 => IR_IN(28), A4 => 
                           IR_IN(30), ZN => n79);
   U136 : NOR2_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), ZN => n45);
   U137 : INV_X1 port map( A => n115, ZN => n58);
   U138 : NAND3_X1 port map( A1 => IR_IN(30), A2 => n114, A3 => n141, ZN => 
                           n115);
   U139 : NOR2_X1 port map( A1 => n133, A2 => IR_IN(31), ZN => n141);
   U140 : INV_X1 port map( A => IR_IN(28), ZN => n114);
   U141 : NOR2_X1 port map( A1 => n142, A2 => IR_IN(27), ZN => n52);
   U142 : INV_X1 port map( A => IR_IN(26), ZN => n142);
   U143 : INV_X1 port map( A => n13, ZN => n138);
   U144 : NAND4_X1 port map( A1 => IR_IN(28), A2 => IR_IN(30), A3 => n133, A4 
                           => n111, ZN => n13);
   U145 : INV_X1 port map( A => IR_IN(31), ZN => n111);
   U146 : INV_X1 port map( A => IR_IN(29), ZN => n133);
   U147 : INV_X1 port map( A => n12, ZN => n59);
   U148 : NAND2_X1 port map( A1 => IR_IN(27), A2 => IR_IN(26), ZN => n12);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   PC_LATCH_EN <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   NPC_LATCH_EN <= '0';
   IR_LATCH_EN <= '0';
   signed_unsigned_1_reg : DFF_X1 port map( D => n150, CK => Clk, Q => n_2327, 
                           QN => n10);
   U9 : INV_X1 port map( A => n3, ZN => n1);
   U164 : INV_X4 port map( A => n1, ZN => lhi_sel);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ISSUE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (63 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ISSUE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (63 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DATAPTH_NBIT32_REG_BIT5
      port( CLK, RST : in std_logic;  PC, IR : in std_logic_vector (31 downto 
            0);  PC_OUT : out std_logic_vector (31 downto 0);  NPC_LATCH_EN, 
            ir_LATCH_EN, signed_op, RF1, RF2, WF1, regImm_LATCH_EN, S1, S2, EN2
            , lhi_sel, jump_en, branch_cond, sb_op, RM, WM, EN3, S3 : in 
            std_logic;  instruction_alu : in std_logic_vector (0 to 5);  
            DATA_MEM_ADDR, DATA_MEM_IN : out std_logic_vector (31 downto 0);  
            DATA_MEM_OUT : in std_logic_vector (31 downto 0);  DATA_MEM_ENABLE,
            DATA_MEM_RM, DATA_MEM_WM : out std_logic);
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
            std_logic;  ALU_OPCODE : out std_logic_vector (0 to 5);  
            signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
            WB_MUX_SEL, RF_WE, lhi_sel, sb_op : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X2
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N9, IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_25_port, IR_24_port, IR_23_port, IR_22_port, IR_21_port, 
      IR_20_port, IR_19_port, IR_18_port, IR_17_port, IR_16_port, IR_15_port, 
      IR_14_port, IR_13_port, IR_12_port, IR_11_port, IR_10_port, IR_9_port, 
      IR_8_port, IR_7_port, IR_6_port, IR_5_port, IR_4_port, IR_3_port, 
      IR_2_port, IR_1_port, IR_0_port, IR_LATCH_EN_i, PC_31_port, PC_30_port, 
      PC_29_port, PC_28_port, PC_27_port, PC_26_port, PC_25_port, PC_24_port, 
      PC_23_port, PC_22_port, PC_21_port, PC_20_port, PC_19_port, PC_18_port, 
      PC_17_port, PC_16_port, PC_15_port, PC_14_port, PC_13_port, PC_12_port, 
      PC_11_port, PC_10_port, PC_9_port, PC_8_port, PC_7_port, PC_6_port, 
      PC_5_port, PC_4_port, PC_3_port, PC_2_port, PC_1_port, PC_0_port, 
      PC_LATCH_EN_i, NPC_LATCH_EN_i, RegA_LATCH_EN_i, RegB_LATCH_EN_i, 
      RegIMM_LATCH_EN_i, MUXA_SEL_i, MUXB_SEL_i, ALU_OUTREG_EN_i, EQ_COND_i, 
      ALU_OPCODE_i_5_port, ALU_OPCODE_i_4_port, ALU_OPCODE_i_3_port, 
      ALU_OPCODE_i_2_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_0_port, 
      signed_unsigned_i, DRAM_WE_i, LMD_LATCH_EN_i, JUMP_EN_i, WB_MUX_SEL_i, 
      RF_WE_i, lhi_sel_i, sb_op_i, DATA_MEM_IN_i_31_port, DATA_MEM_IN_i_30_port
      , DATA_MEM_IN_i_29_port, DATA_MEM_IN_i_28_port, DATA_MEM_IN_i_27_port, 
      DATA_MEM_IN_i_26_port, DATA_MEM_IN_i_25_port, DATA_MEM_IN_i_24_port, 
      DATA_MEM_IN_i_23_port, DATA_MEM_IN_i_22_port, DATA_MEM_IN_i_21_port, 
      DATA_MEM_IN_i_20_port, DATA_MEM_IN_i_19_port, DATA_MEM_IN_i_18_port, 
      DATA_MEM_IN_i_17_port, DATA_MEM_IN_i_16_port, DATA_MEM_IN_i_15_port, 
      DATA_MEM_IN_i_14_port, DATA_MEM_IN_i_13_port, DATA_MEM_IN_i_12_port, 
      DATA_MEM_IN_i_11_port, DATA_MEM_IN_i_10_port, DATA_MEM_IN_i_9_port, 
      DATA_MEM_IN_i_8_port, DATA_MEM_IN_i_7_port, DATA_MEM_IN_i_6_port, 
      DATA_MEM_IN_i_5_port, DATA_MEM_IN_i_4_port, DATA_MEM_IN_i_3_port, 
      DATA_MEM_IN_i_2_port, DATA_MEM_IN_i_1_port, DATA_MEM_IN_i_0_port, 
      dram_data_i_31_port, dram_data_i_30_port, dram_data_i_29_port, 
      dram_data_i_28_port, dram_data_i_27_port, dram_data_i_26_port, 
      dram_data_i_25_port, dram_data_i_24_port, dram_data_i_23_port, 
      dram_data_i_22_port, dram_data_i_21_port, dram_data_i_20_port, 
      dram_data_i_19_port, dram_data_i_18_port, dram_data_i_17_port, 
      dram_data_i_16_port, dram_data_i_15_port, dram_data_i_14_port, 
      dram_data_i_13_port, dram_data_i_12_port, dram_data_i_11_port, 
      dram_data_i_10_port, dram_data_i_9_port, dram_data_i_8_port, 
      dram_data_i_7_port, dram_data_i_6_port, dram_data_i_5_port, 
      dram_data_i_4_port, dram_data_i_3_port, dram_data_i_2_port, 
      dram_data_i_1_port, dram_data_i_0_port, DATA_MEM_WM_i, n1, n_2361, n_2362
      , n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371,
      n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, 
      n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, 
      n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, 
      n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, 
      n_2408, n_2409 : std_logic;

begin
   
   DRAM_READNOTWRITE_reg : DFF_X1 port map( D => N9, CK => CLK, Q => 
                           DRAM_READNOTWRITE, QN => n_2361);
   DRAM_DATA_tri_0_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_0_port, EN => N9
                           , Z => DRAM_DATA(0));
   DRAM_DATA_tri_1_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_1_port, EN => N9
                           , Z => DRAM_DATA(1));
   DRAM_DATA_tri_2_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_2_port, EN => N9
                           , Z => DRAM_DATA(2));
   DRAM_DATA_tri_3_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_3_port, EN => N9
                           , Z => DRAM_DATA(3));
   DRAM_DATA_tri_4_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_4_port, EN => N9
                           , Z => DRAM_DATA(4));
   DRAM_DATA_tri_5_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_5_port, EN => N9
                           , Z => DRAM_DATA(5));
   DRAM_DATA_tri_6_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_6_port, EN => N9
                           , Z => DRAM_DATA(6));
   DRAM_DATA_tri_7_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_7_port, EN => N9
                           , Z => DRAM_DATA(7));
   DRAM_DATA_tri_8_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_8_port, EN => N9
                           , Z => DRAM_DATA(8));
   DRAM_DATA_tri_9_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_9_port, EN => N9
                           , Z => DRAM_DATA(9));
   DRAM_DATA_tri_10_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_10_port, EN => 
                           N9, Z => DRAM_DATA(10));
   DRAM_DATA_tri_11_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_11_port, EN => 
                           N9, Z => DRAM_DATA(11));
   DRAM_DATA_tri_12_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_12_port, EN => 
                           N9, Z => DRAM_DATA(12));
   DRAM_DATA_tri_13_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_13_port, EN => 
                           N9, Z => DRAM_DATA(13));
   DRAM_DATA_tri_14_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_14_port, EN => 
                           N9, Z => DRAM_DATA(14));
   DRAM_DATA_tri_15_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_15_port, EN => 
                           N9, Z => DRAM_DATA(15));
   DRAM_DATA_tri_16_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_16_port, EN => 
                           N9, Z => DRAM_DATA(16));
   DRAM_DATA_tri_17_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_17_port, EN => 
                           N9, Z => DRAM_DATA(17));
   DRAM_DATA_tri_18_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_18_port, EN => 
                           N9, Z => DRAM_DATA(18));
   DRAM_DATA_tri_19_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_19_port, EN => 
                           N9, Z => DRAM_DATA(19));
   DRAM_DATA_tri_20_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_20_port, EN => 
                           N9, Z => DRAM_DATA(20));
   DRAM_DATA_tri_21_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_21_port, EN => 
                           N9, Z => DRAM_DATA(21));
   DRAM_DATA_tri_22_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_22_port, EN => 
                           N9, Z => DRAM_DATA(22));
   DRAM_DATA_tri_23_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_23_port, EN => 
                           N9, Z => DRAM_DATA(23));
   DRAM_DATA_tri_24_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_24_port, EN => 
                           N9, Z => DRAM_DATA(24));
   DRAM_DATA_tri_25_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_25_port, EN => 
                           N9, Z => DRAM_DATA(25));
   DRAM_DATA_tri_26_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_26_port, EN => 
                           N9, Z => DRAM_DATA(26));
   DRAM_DATA_tri_27_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_27_port, EN => 
                           N9, Z => DRAM_DATA(27));
   DRAM_DATA_tri_28_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_28_port, EN => 
                           N9, Z => DRAM_DATA(28));
   DRAM_DATA_tri_29_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_29_port, EN => 
                           N9, Z => DRAM_DATA(29));
   DRAM_DATA_tri_30_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_30_port, EN => 
                           N9, Z => DRAM_DATA(30));
   DRAM_DATA_tri_31_inst : TBUF_X2 port map( A => DATA_MEM_IN_i_31_port, EN => 
                           N9, Z => DRAM_DATA(31));
   DRAM_DATA_tri_32_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(32));
   DRAM_DATA_tri_33_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(33));
   DRAM_DATA_tri_34_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(34));
   DRAM_DATA_tri_35_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(35));
   DRAM_DATA_tri_36_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(36));
   DRAM_DATA_tri_37_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(37));
   DRAM_DATA_tri_38_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(38));
   DRAM_DATA_tri_39_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(39));
   DRAM_DATA_tri_40_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(40));
   DRAM_DATA_tri_41_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(41));
   DRAM_DATA_tri_42_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(42));
   DRAM_DATA_tri_43_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(43));
   DRAM_DATA_tri_44_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(44));
   DRAM_DATA_tri_45_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(45));
   DRAM_DATA_tri_46_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(46));
   DRAM_DATA_tri_47_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(47));
   DRAM_DATA_tri_48_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(48));
   DRAM_DATA_tri_49_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(49));
   DRAM_DATA_tri_50_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(50));
   DRAM_DATA_tri_51_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(51));
   DRAM_DATA_tri_52_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(52));
   DRAM_DATA_tri_53_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(53));
   DRAM_DATA_tri_54_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(54));
   DRAM_DATA_tri_55_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(55));
   DRAM_DATA_tri_56_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(56));
   DRAM_DATA_tri_57_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(57));
   DRAM_DATA_tri_58_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(58));
   DRAM_DATA_tri_59_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(59));
   DRAM_DATA_tri_60_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(60));
   DRAM_DATA_tri_61_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(61));
   DRAM_DATA_tri_62_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(62));
   DRAM_DATA_tri_63_inst : TBUF_X2 port map( A => n1, EN => N9, Z => 
                           DRAM_DATA(63));
   n1 <= '0';
   U166 : AND2_X1 port map( A1 => N9, A2 => DRAM_DATA(41), ZN => 
                           dram_data_i_9_port);
   U167 : AND2_X1 port map( A1 => DRAM_DATA(40), A2 => N9, ZN => 
                           dram_data_i_8_port);
   U168 : AND2_X1 port map( A1 => DRAM_DATA(39), A2 => N9, ZN => 
                           dram_data_i_7_port);
   U169 : AND2_X1 port map( A1 => DRAM_DATA(38), A2 => N9, ZN => 
                           dram_data_i_6_port);
   U170 : AND2_X1 port map( A1 => DRAM_DATA(37), A2 => N9, ZN => 
                           dram_data_i_5_port);
   U171 : AND2_X1 port map( A1 => DRAM_DATA(36), A2 => N9, ZN => 
                           dram_data_i_4_port);
   U172 : AND2_X1 port map( A1 => DRAM_DATA(35), A2 => N9, ZN => 
                           dram_data_i_3_port);
   U173 : AND2_X1 port map( A1 => DRAM_DATA(63), A2 => N9, ZN => 
                           dram_data_i_31_port);
   U174 : AND2_X1 port map( A1 => DRAM_DATA(62), A2 => N9, ZN => 
                           dram_data_i_30_port);
   U175 : AND2_X1 port map( A1 => DRAM_DATA(34), A2 => N9, ZN => 
                           dram_data_i_2_port);
   U176 : AND2_X1 port map( A1 => DRAM_DATA(61), A2 => N9, ZN => 
                           dram_data_i_29_port);
   U177 : AND2_X1 port map( A1 => DRAM_DATA(60), A2 => N9, ZN => 
                           dram_data_i_28_port);
   U178 : AND2_X1 port map( A1 => DRAM_DATA(59), A2 => N9, ZN => 
                           dram_data_i_27_port);
   U179 : AND2_X1 port map( A1 => DRAM_DATA(58), A2 => N9, ZN => 
                           dram_data_i_26_port);
   U180 : AND2_X1 port map( A1 => DRAM_DATA(57), A2 => N9, ZN => 
                           dram_data_i_25_port);
   U181 : AND2_X1 port map( A1 => DRAM_DATA(56), A2 => N9, ZN => 
                           dram_data_i_24_port);
   U182 : AND2_X1 port map( A1 => DRAM_DATA(55), A2 => N9, ZN => 
                           dram_data_i_23_port);
   U183 : AND2_X1 port map( A1 => DRAM_DATA(54), A2 => N9, ZN => 
                           dram_data_i_22_port);
   U184 : AND2_X1 port map( A1 => DRAM_DATA(53), A2 => N9, ZN => 
                           dram_data_i_21_port);
   U185 : AND2_X1 port map( A1 => DRAM_DATA(52), A2 => N9, ZN => 
                           dram_data_i_20_port);
   U186 : AND2_X1 port map( A1 => DRAM_DATA(33), A2 => N9, ZN => 
                           dram_data_i_1_port);
   U187 : AND2_X1 port map( A1 => DRAM_DATA(51), A2 => N9, ZN => 
                           dram_data_i_19_port);
   U188 : AND2_X1 port map( A1 => DRAM_DATA(50), A2 => N9, ZN => 
                           dram_data_i_18_port);
   U189 : AND2_X1 port map( A1 => DRAM_DATA(49), A2 => N9, ZN => 
                           dram_data_i_17_port);
   U190 : AND2_X1 port map( A1 => DRAM_DATA(48), A2 => N9, ZN => 
                           dram_data_i_16_port);
   U191 : AND2_X1 port map( A1 => DRAM_DATA(47), A2 => N9, ZN => 
                           dram_data_i_15_port);
   U192 : AND2_X1 port map( A1 => DRAM_DATA(46), A2 => N9, ZN => 
                           dram_data_i_14_port);
   U193 : AND2_X1 port map( A1 => DRAM_DATA(45), A2 => N9, ZN => 
                           dram_data_i_13_port);
   U194 : AND2_X1 port map( A1 => DRAM_DATA(44), A2 => N9, ZN => 
                           dram_data_i_12_port);
   U195 : AND2_X1 port map( A1 => DRAM_DATA(43), A2 => N9, ZN => 
                           dram_data_i_11_port);
   U196 : AND2_X1 port map( A1 => DRAM_DATA(42), A2 => N9, ZN => 
                           dram_data_i_10_port);
   U197 : AND2_X1 port map( A1 => DRAM_DATA(32), A2 => N9, ZN => 
                           dram_data_i_0_port);
   CU_I : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 
                           port map( Clk => CLK, Rst => RST, IR_IN(31) => 
                           IR_31_port, IR_IN(30) => IR_30_port, IR_IN(29) => 
                           IR_29_port, IR_IN(28) => IR_28_port, IR_IN(27) => 
                           IR_27_port, IR_IN(26) => IR_26_port, IR_IN(25) => 
                           IR_25_port, IR_IN(24) => IR_24_port, IR_IN(23) => 
                           IR_23_port, IR_IN(22) => IR_22_port, IR_IN(21) => 
                           IR_21_port, IR_IN(20) => IR_20_port, IR_IN(19) => 
                           IR_19_port, IR_IN(18) => IR_18_port, IR_IN(17) => 
                           IR_17_port, IR_IN(16) => IR_16_port, IR_IN(15) => 
                           IR_15_port, IR_IN(14) => IR_14_port, IR_IN(13) => 
                           IR_13_port, IR_IN(12) => IR_12_port, IR_IN(11) => 
                           IR_11_port, IR_IN(10) => IR_10_port, IR_IN(9) => 
                           IR_9_port, IR_IN(8) => IR_8_port, IR_IN(7) => 
                           IR_7_port, IR_IN(6) => IR_6_port, IR_IN(5) => 
                           IR_5_port, IR_IN(4) => IR_4_port, IR_IN(3) => 
                           IR_3_port, IR_IN(2) => IR_2_port, IR_IN(1) => 
                           IR_1_port, IR_IN(0) => IR_0_port, IR_LATCH_EN => 
                           n_2362, NPC_LATCH_EN => n_2363, RegA_LATCH_EN => 
                           n_2364, RegB_LATCH_EN => n_2365, RegIMM_LATCH_EN => 
                           n_2366, MUXA_SEL => n_2367, MUXB_SEL => n_2368, 
                           ALU_OUTREG_EN => n_2369, EQ_COND => n_2370, 
                           ALU_OPCODE(0) => ALU_OPCODE_i_5_port, ALU_OPCODE(1) 
                           => ALU_OPCODE_i_4_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_i_0_port, signed_unsigned => 
                           signed_unsigned_i, DRAM_WE => n_2371, LMD_LATCH_EN 
                           => n_2372, JUMP_EN => n_2373, PC_LATCH_EN => n_2374,
                           WB_MUX_SEL => n_2375, RF_WE => n_2376, lhi_sel => 
                           lhi_sel_i, sb_op => sb_op_i);
   DTPTH_I : DATAPTH_NBIT32_REG_BIT5 port map( CLK => CLK, RST => RST, PC(31) 
                           => PC_31_port, PC(30) => PC_30_port, PC(29) => 
                           PC_29_port, PC(28) => PC_28_port, PC(27) => 
                           PC_27_port, PC(26) => PC_26_port, PC(25) => 
                           PC_25_port, PC(24) => PC_24_port, PC(23) => 
                           PC_23_port, PC(22) => PC_22_port, PC(21) => 
                           PC_21_port, PC(20) => PC_20_port, PC(19) => 
                           PC_19_port, PC(18) => PC_18_port, PC(17) => 
                           PC_17_port, PC(16) => PC_16_port, PC(15) => 
                           PC_15_port, PC(14) => PC_14_port, PC(13) => 
                           PC_13_port, PC(12) => PC_12_port, PC(11) => 
                           PC_11_port, PC(10) => PC_10_port, PC(9) => PC_9_port
                           , PC(8) => PC_8_port, PC(7) => PC_7_port, PC(6) => 
                           PC_6_port, PC(5) => PC_5_port, PC(4) => PC_4_port, 
                           PC(3) => PC_3_port, PC(2) => PC_2_port, PC(1) => 
                           PC_1_port, PC(0) => PC_0_port, IR(31) => IR_31_port,
                           IR(30) => IR_30_port, IR(29) => IR_29_port, IR(28) 
                           => IR_28_port, IR(27) => IR_27_port, IR(26) => 
                           IR_26_port, IR(25) => IR_25_port, IR(24) => 
                           IR_24_port, IR(23) => IR_23_port, IR(22) => 
                           IR_22_port, IR(21) => IR_21_port, IR(20) => 
                           IR_20_port, IR(19) => IR_19_port, IR(18) => 
                           IR_18_port, IR(17) => IR_17_port, IR(16) => 
                           IR_16_port, IR(15) => IR_15_port, IR(14) => 
                           IR_14_port, IR(13) => IR_13_port, IR(12) => 
                           IR_12_port, IR(11) => IR_11_port, IR(10) => 
                           IR_10_port, IR(9) => IR_9_port, IR(8) => IR_8_port, 
                           IR(7) => IR_7_port, IR(6) => IR_6_port, IR(5) => 
                           IR_5_port, IR(4) => IR_4_port, IR(3) => IR_3_port, 
                           IR(2) => IR_2_port, IR(1) => IR_1_port, IR(0) => 
                           IR_0_port, PC_OUT(31) => n_2377, PC_OUT(30) => 
                           n_2378, PC_OUT(29) => n_2379, PC_OUT(28) => n_2380, 
                           PC_OUT(27) => n_2381, PC_OUT(26) => n_2382, 
                           PC_OUT(25) => n_2383, PC_OUT(24) => n_2384, 
                           PC_OUT(23) => n_2385, PC_OUT(22) => n_2386, 
                           PC_OUT(21) => n_2387, PC_OUT(20) => n_2388, 
                           PC_OUT(19) => n_2389, PC_OUT(18) => n_2390, 
                           PC_OUT(17) => n_2391, PC_OUT(16) => n_2392, 
                           PC_OUT(15) => n_2393, PC_OUT(14) => n_2394, 
                           PC_OUT(13) => n_2395, PC_OUT(12) => n_2396, 
                           PC_OUT(11) => n_2397, PC_OUT(10) => n_2398, 
                           PC_OUT(9) => n_2399, PC_OUT(8) => n_2400, PC_OUT(7) 
                           => n_2401, PC_OUT(6) => n_2402, PC_OUT(5) => n_2403,
                           PC_OUT(4) => n_2404, PC_OUT(3) => n_2405, PC_OUT(2) 
                           => n_2406, PC_OUT(1) => n_2407, PC_OUT(0) => n_2408,
                           NPC_LATCH_EN => NPC_LATCH_EN_i, ir_LATCH_EN => 
                           IR_LATCH_EN_i, signed_op => signed_unsigned_i, RF1 
                           => RegA_LATCH_EN_i, RF2 => RegB_LATCH_EN_i, WF1 => 
                           RF_WE_i, regImm_LATCH_EN => RegIMM_LATCH_EN_i, S1 =>
                           MUXA_SEL_i, S2 => MUXB_SEL_i, EN2 => ALU_OUTREG_EN_i
                           , lhi_sel => lhi_sel_i, jump_en => JUMP_EN_i, 
                           branch_cond => EQ_COND_i, sb_op => sb_op_i, RM => 
                           LMD_LATCH_EN_i, WM => DRAM_WE_i, EN3 => 
                           PC_LATCH_EN_i, S3 => WB_MUX_SEL_i, 
                           instruction_alu(0) => ALU_OPCODE_i_5_port, 
                           instruction_alu(1) => ALU_OPCODE_i_4_port, 
                           instruction_alu(2) => ALU_OPCODE_i_3_port, 
                           instruction_alu(3) => ALU_OPCODE_i_2_port, 
                           instruction_alu(4) => ALU_OPCODE_i_1_port, 
                           instruction_alu(5) => ALU_OPCODE_i_0_port, 
                           DATA_MEM_ADDR(31) => DRAM_ADDRESS(31), 
                           DATA_MEM_ADDR(30) => DRAM_ADDRESS(30), 
                           DATA_MEM_ADDR(29) => DRAM_ADDRESS(29), 
                           DATA_MEM_ADDR(28) => DRAM_ADDRESS(28), 
                           DATA_MEM_ADDR(27) => DRAM_ADDRESS(27), 
                           DATA_MEM_ADDR(26) => DRAM_ADDRESS(26), 
                           DATA_MEM_ADDR(25) => DRAM_ADDRESS(25), 
                           DATA_MEM_ADDR(24) => DRAM_ADDRESS(24), 
                           DATA_MEM_ADDR(23) => DRAM_ADDRESS(23), 
                           DATA_MEM_ADDR(22) => DRAM_ADDRESS(22), 
                           DATA_MEM_ADDR(21) => DRAM_ADDRESS(21), 
                           DATA_MEM_ADDR(20) => DRAM_ADDRESS(20), 
                           DATA_MEM_ADDR(19) => DRAM_ADDRESS(19), 
                           DATA_MEM_ADDR(18) => DRAM_ADDRESS(18), 
                           DATA_MEM_ADDR(17) => DRAM_ADDRESS(17), 
                           DATA_MEM_ADDR(16) => DRAM_ADDRESS(16), 
                           DATA_MEM_ADDR(15) => DRAM_ADDRESS(15), 
                           DATA_MEM_ADDR(14) => DRAM_ADDRESS(14), 
                           DATA_MEM_ADDR(13) => DRAM_ADDRESS(13), 
                           DATA_MEM_ADDR(12) => DRAM_ADDRESS(12), 
                           DATA_MEM_ADDR(11) => DRAM_ADDRESS(11), 
                           DATA_MEM_ADDR(10) => DRAM_ADDRESS(10), 
                           DATA_MEM_ADDR(9) => DRAM_ADDRESS(9), 
                           DATA_MEM_ADDR(8) => DRAM_ADDRESS(8), 
                           DATA_MEM_ADDR(7) => DRAM_ADDRESS(7), 
                           DATA_MEM_ADDR(6) => DRAM_ADDRESS(6), 
                           DATA_MEM_ADDR(5) => DRAM_ADDRESS(5), 
                           DATA_MEM_ADDR(4) => DRAM_ADDRESS(4), 
                           DATA_MEM_ADDR(3) => DRAM_ADDRESS(3), 
                           DATA_MEM_ADDR(2) => DRAM_ADDRESS(2), 
                           DATA_MEM_ADDR(1) => DRAM_ADDRESS(1), 
                           DATA_MEM_ADDR(0) => DRAM_ADDRESS(0), DATA_MEM_IN(31)
                           => DATA_MEM_IN_i_31_port, DATA_MEM_IN(30) => 
                           DATA_MEM_IN_i_30_port, DATA_MEM_IN(29) => 
                           DATA_MEM_IN_i_29_port, DATA_MEM_IN(28) => 
                           DATA_MEM_IN_i_28_port, DATA_MEM_IN(27) => 
                           DATA_MEM_IN_i_27_port, DATA_MEM_IN(26) => 
                           DATA_MEM_IN_i_26_port, DATA_MEM_IN(25) => 
                           DATA_MEM_IN_i_25_port, DATA_MEM_IN(24) => 
                           DATA_MEM_IN_i_24_port, DATA_MEM_IN(23) => 
                           DATA_MEM_IN_i_23_port, DATA_MEM_IN(22) => 
                           DATA_MEM_IN_i_22_port, DATA_MEM_IN(21) => 
                           DATA_MEM_IN_i_21_port, DATA_MEM_IN(20) => 
                           DATA_MEM_IN_i_20_port, DATA_MEM_IN(19) => 
                           DATA_MEM_IN_i_19_port, DATA_MEM_IN(18) => 
                           DATA_MEM_IN_i_18_port, DATA_MEM_IN(17) => 
                           DATA_MEM_IN_i_17_port, DATA_MEM_IN(16) => 
                           DATA_MEM_IN_i_16_port, DATA_MEM_IN(15) => 
                           DATA_MEM_IN_i_15_port, DATA_MEM_IN(14) => 
                           DATA_MEM_IN_i_14_port, DATA_MEM_IN(13) => 
                           DATA_MEM_IN_i_13_port, DATA_MEM_IN(12) => 
                           DATA_MEM_IN_i_12_port, DATA_MEM_IN(11) => 
                           DATA_MEM_IN_i_11_port, DATA_MEM_IN(10) => 
                           DATA_MEM_IN_i_10_port, DATA_MEM_IN(9) => 
                           DATA_MEM_IN_i_9_port, DATA_MEM_IN(8) => 
                           DATA_MEM_IN_i_8_port, DATA_MEM_IN(7) => 
                           DATA_MEM_IN_i_7_port, DATA_MEM_IN(6) => 
                           DATA_MEM_IN_i_6_port, DATA_MEM_IN(5) => 
                           DATA_MEM_IN_i_5_port, DATA_MEM_IN(4) => 
                           DATA_MEM_IN_i_4_port, DATA_MEM_IN(3) => 
                           DATA_MEM_IN_i_3_port, DATA_MEM_IN(2) => 
                           DATA_MEM_IN_i_2_port, DATA_MEM_IN(1) => 
                           DATA_MEM_IN_i_1_port, DATA_MEM_IN(0) => 
                           DATA_MEM_IN_i_0_port, DATA_MEM_OUT(31) => 
                           dram_data_i_31_port, DATA_MEM_OUT(30) => 
                           dram_data_i_30_port, DATA_MEM_OUT(29) => 
                           dram_data_i_29_port, DATA_MEM_OUT(28) => 
                           dram_data_i_28_port, DATA_MEM_OUT(27) => 
                           dram_data_i_27_port, DATA_MEM_OUT(26) => 
                           dram_data_i_26_port, DATA_MEM_OUT(25) => 
                           dram_data_i_25_port, DATA_MEM_OUT(24) => 
                           dram_data_i_24_port, DATA_MEM_OUT(23) => 
                           dram_data_i_23_port, DATA_MEM_OUT(22) => 
                           dram_data_i_22_port, DATA_MEM_OUT(21) => 
                           dram_data_i_21_port, DATA_MEM_OUT(20) => 
                           dram_data_i_20_port, DATA_MEM_OUT(19) => 
                           dram_data_i_19_port, DATA_MEM_OUT(18) => 
                           dram_data_i_18_port, DATA_MEM_OUT(17) => 
                           dram_data_i_17_port, DATA_MEM_OUT(16) => 
                           dram_data_i_16_port, DATA_MEM_OUT(15) => 
                           dram_data_i_15_port, DATA_MEM_OUT(14) => 
                           dram_data_i_14_port, DATA_MEM_OUT(13) => 
                           dram_data_i_13_port, DATA_MEM_OUT(12) => 
                           dram_data_i_12_port, DATA_MEM_OUT(11) => 
                           dram_data_i_11_port, DATA_MEM_OUT(10) => 
                           dram_data_i_10_port, DATA_MEM_OUT(9) => 
                           dram_data_i_9_port, DATA_MEM_OUT(8) => 
                           dram_data_i_8_port, DATA_MEM_OUT(7) => 
                           dram_data_i_7_port, DATA_MEM_OUT(6) => 
                           dram_data_i_6_port, DATA_MEM_OUT(5) => 
                           dram_data_i_5_port, DATA_MEM_OUT(4) => 
                           dram_data_i_4_port, DATA_MEM_OUT(3) => 
                           dram_data_i_3_port, DATA_MEM_OUT(2) => 
                           dram_data_i_2_port, DATA_MEM_OUT(1) => 
                           dram_data_i_1_port, DATA_MEM_OUT(0) => 
                           dram_data_i_0_port, DATA_MEM_ENABLE => DRAM_ISSUE, 
                           DATA_MEM_RM => n_2409, DATA_MEM_WM => DATA_MEM_WM_i)
                           ;
   U198 : INV_X8 port map( A => DATA_MEM_WM_i, ZN => N9);
   IR_0_port <= '0';
   IR_1_port <= '0';
   IR_2_port <= '0';
   IR_3_port <= '0';
   IR_4_port <= '0';
   IR_5_port <= '0';
   IR_6_port <= '0';
   IR_7_port <= '0';
   IR_8_port <= '0';
   IR_9_port <= '0';
   IR_10_port <= '0';
   IR_11_port <= '0';
   IR_12_port <= '0';
   IR_13_port <= '0';
   IR_14_port <= '0';
   IR_15_port <= '0';
   IR_16_port <= '0';
   IR_17_port <= '0';
   IR_18_port <= '0';
   IR_19_port <= '0';
   IR_20_port <= '0';
   IR_21_port <= '0';
   IR_22_port <= '0';
   IR_23_port <= '0';
   IR_24_port <= '0';
   IR_25_port <= '0';
   IR_26_port <= '0';
   IR_27_port <= '0';
   IR_28_port <= '0';
   IR_29_port <= '0';
   IR_30_port <= '0';
   IR_31_port <= '0';
   PC_0_port <= '0';
   IRAM_ADDRESS(0) <= '0';
   PC_1_port <= '0';
   IRAM_ADDRESS(1) <= '0';
   PC_2_port <= '0';
   IRAM_ADDRESS(2) <= '0';
   PC_3_port <= '0';
   IRAM_ADDRESS(3) <= '0';
   PC_4_port <= '0';
   IRAM_ADDRESS(4) <= '0';
   PC_5_port <= '0';
   IRAM_ADDRESS(5) <= '0';
   PC_6_port <= '0';
   IRAM_ADDRESS(6) <= '0';
   PC_7_port <= '0';
   IRAM_ADDRESS(7) <= '0';
   PC_8_port <= '0';
   IRAM_ADDRESS(8) <= '0';
   PC_9_port <= '0';
   IRAM_ADDRESS(9) <= '0';
   PC_10_port <= '0';
   IRAM_ADDRESS(10) <= '0';
   PC_11_port <= '0';
   IRAM_ADDRESS(11) <= '0';
   PC_12_port <= '0';
   IRAM_ADDRESS(12) <= '0';
   PC_13_port <= '0';
   IRAM_ADDRESS(13) <= '0';
   PC_14_port <= '0';
   IRAM_ADDRESS(14) <= '0';
   PC_15_port <= '0';
   IRAM_ADDRESS(15) <= '0';
   PC_16_port <= '0';
   IRAM_ADDRESS(16) <= '0';
   PC_17_port <= '0';
   IRAM_ADDRESS(17) <= '0';
   PC_18_port <= '0';
   IRAM_ADDRESS(18) <= '0';
   PC_19_port <= '0';
   IRAM_ADDRESS(19) <= '0';
   PC_20_port <= '0';
   IRAM_ADDRESS(20) <= '0';
   PC_21_port <= '0';
   IRAM_ADDRESS(21) <= '0';
   PC_22_port <= '0';
   IRAM_ADDRESS(22) <= '0';
   PC_23_port <= '0';
   IRAM_ADDRESS(23) <= '0';
   PC_24_port <= '0';
   IRAM_ADDRESS(24) <= '0';
   PC_25_port <= '0';
   IRAM_ADDRESS(25) <= '0';
   PC_26_port <= '0';
   IRAM_ADDRESS(26) <= '0';
   PC_27_port <= '0';
   IRAM_ADDRESS(27) <= '0';
   PC_28_port <= '0';
   IRAM_ADDRESS(28) <= '0';
   PC_29_port <= '0';
   IRAM_ADDRESS(29) <= '0';
   PC_30_port <= '0';
   IRAM_ADDRESS(30) <= '0';
   PC_31_port <= '0';
   IRAM_ADDRESS(31) <= '0';
   RF_WE_i <= '0';
   WB_MUX_SEL_i <= '0';
   PC_LATCH_EN_i <= '0';
   JUMP_EN_i <= '0';
   LMD_LATCH_EN_i <= '0';
   DRAM_WE_i <= '0';
   EQ_COND_i <= '0';
   ALU_OUTREG_EN_i <= '0';
   MUXB_SEL_i <= '0';
   MUXA_SEL_i <= '0';
   RegIMM_LATCH_EN_i <= '0';
   RegB_LATCH_EN_i <= '0';
   RegA_LATCH_EN_i <= '0';
   NPC_LATCH_EN_i <= '0';
   IR_LATCH_EN_i <= '0';

end SYN_dlx_rtl;


library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (NOP, ADDS, LLS, LRS, ADD, SUB, ANDR, ORR, XORR, SNE, SLE, SGE, 
   BEQZ, BNEZ, SUBI, ANDI, ORI, XORI, SLLI, SRLI, SNEI, SLEI, SGEI, LW, SW, 
   SUBU, SUBUI, ADDU, ADDUI, SRA1, SEQ, SLT, SGT, SLTU, SGTU, SGEU, LHI, JR, 
   JALR, SRAI, SEQI, SLTI, SGTI, LB, LBU, LHU, SB, SLTUI, SGTUI, SGEUI, trap, 
   rfe);
attribute ENUM_ENCODING of aluOp : type is 
   "000000 000001 000010 000011 000100 000101 000110 000111 001000 001001 001010 001011 001100 001101 001110 001111 010000 010001 010010 010011 010100 010101 010110 010111 011000 011001 011010 011011 011100 011101 011110 011111 100000 100001 100010 100011 100100 100101 100110 100111 101000 101001 101010 101011 101100 101101 101110 101111 110000 110001 110010 110011";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 6 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 6 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "000000" => return NOP;
         when "000001" => return ADDS;
         when "000010" => return LLS;
         when "000011" => return LRS;
         when "000100" => return ADD;
         when "000101" => return SUB;
         when "000110" => return ANDR;
         when "000111" => return ORR;
         when "001000" => return XORR;
         when "001001" => return SNE;
         when "001010" => return SLE;
         when "001011" => return SGE;
         when "001100" => return BEQZ;
         when "001101" => return BNEZ;
         when "001110" => return SUBI;
         when "001111" => return ANDI;
         when "010000" => return ORI;
         when "010001" => return XORI;
         when "010010" => return SLLI;
         when "010011" => return SRLI;
         when "010100" => return SNEI;
         when "010101" => return SLEI;
         when "010110" => return SGEI;
         when "010111" => return LW;
         when "011000" => return SW;
         when "011001" => return SUBU;
         when "011010" => return SUBUI;
         when "011011" => return ADDU;
         when "011100" => return ADDUI;
         when "011101" => return SRA1;
         when "011110" => return SEQ;
         when "011111" => return SLT;
         when "100000" => return SGT;
         when "100001" => return SLTU;
         when "100010" => return SGTU;
         when "100011" => return SGEU;
         when "100100" => return LHI;
         when "100101" => return JR;
         when "100110" => return JALR;
         when "100111" => return SRAI;
         when "101000" => return SEQI;
         when "101001" => return SLTI;
         when "101010" => return SGTI;
         when "101011" => return LB;
         when "101100" => return LBU;
         when "101101" => return LHU;
         when "101110" => return SB;
         when "101111" => return SLTUI;
         when "110000" => return SGTUI;
         when "110001" => return SGEUI;
         when "110010" => return trap;
         when "110011" => return rfe;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "000000";
         when ADDS => return "000001";
         when LLS => return "000010";
         when LRS => return "000011";
         when ADD => return "000100";
         when SUB => return "000101";
         when ANDR => return "000110";
         when ORR => return "000111";
         when XORR => return "001000";
         when SNE => return "001001";
         when SLE => return "001010";
         when SGE => return "001011";
         when BEQZ => return "001100";
         when BNEZ => return "001101";
         when SUBI => return "001110";
         when ANDI => return "001111";
         when ORI => return "010000";
         when XORI => return "010001";
         when SLLI => return "010010";
         when SRLI => return "010011";
         when SNEI => return "010100";
         when SLEI => return "010101";
         when SGEI => return "010110";
         when LW => return "010111";
         when SW => return "011000";
         when SUBU => return "011001";
         when SUBUI => return "011010";
         when ADDU => return "011011";
         when ADDUI => return "011100";
         when SRA1 => return "011101";
         when SEQ => return "011110";
         when SLT => return "011111";
         when SGT => return "100000";
         when SLTU => return "100001";
         when SGTU => return "100010";
         when SGEU => return "100011";
         when LHI => return "100100";
         when JR => return "100101";
         when JALR => return "100110";
         when SRAI => return "100111";
         when SEQI => return "101000";
         when SLTI => return "101001";
         when SGTI => return "101010";
         when LB => return "101011";
         when LBU => return "101100";
         when LHU => return "101101";
         when SB => return "101110";
         when SLTUI => return "101111";
         when SGTUI => return "110000";
         when SGEUI => return "110001";
         when trap => return "110010";
         when rfe => return "110011";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "000000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_7 
   is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_7;

architecture SYN_cla of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_7 
   is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port );
   
   U2 : OR2_X2 port map( A1 => n100, A2 => n53, ZN => n72);
   U3 : OR2_X2 port map( A1 => n72, A2 => n73, ZN => n88);
   U4 : INV_X1 port map( A => n46, ZN => n1);
   U5 : AND2_X1 port map( A1 => n10, A2 => n21, ZN => n2);
   U6 : CLKBUF_X1 port map( A => n35, Z => n3);
   U7 : OR2_X1 port map( A1 => n76, A2 => n60, ZN => n4);
   U8 : OR2_X1 port map( A1 => n4, A2 => n57, ZN => n96);
   U9 : CLKBUF_X1 port map( A => A(7), Z => n5);
   U10 : BUF_X1 port map( A => A(2), Z => n20);
   U11 : CLKBUF_X1 port map( A => A(15), Z => n6);
   U12 : CLKBUF_X1 port map( A => A(5), Z => n7);
   U13 : CLKBUF_X1 port map( A => A(3), Z => n8);
   U14 : CLKBUF_X1 port map( A => A(12), Z => n9);
   U15 : CLKBUF_X1 port map( A => A(13), Z => n10);
   U16 : CLKBUF_X1 port map( A => A(0), Z => n11);
   U17 : CLKBUF_X1 port map( A => A(1), Z => n12);
   U18 : CLKBUF_X1 port map( A => A(8), Z => n13);
   U19 : CLKBUF_X1 port map( A => n6, Z => n14);
   U20 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => n60);
   U21 : AND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n15);
   U22 : AND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n16);
   U23 : CLKBUF_X1 port map( A => A(10), Z => n17);
   U24 : AND4_X1 port map( A1 => A(5), A2 => A(6), A3 => A(7), A4 => A(4), ZN 
                           => n18);
   U25 : AND4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(7), A4 => A(6), ZN 
                           => n109);
   U26 : CLKBUF_X1 port map( A => A(4), Z => n19);
   U27 : CLKBUF_X1 port map( A => n9, Z => n21);
   U28 : CLKBUF_X1 port map( A => A(14), Z => n22);
   U29 : CLKBUF_X1 port map( A => A(16), Z => n23);
   U30 : INV_X1 port map( A => n27, ZN => n24);
   U31 : CLKBUF_X1 port map( A => A(6), Z => n25);
   U32 : AND4_X1 port map( A1 => A(1), A2 => A(0), A3 => A(3), A4 => A(2), ZN 
                           => n26);
   U33 : AND4_X1 port map( A1 => A(1), A2 => A(0), A3 => A(3), A4 => A(2), ZN 
                           => n110);
   U34 : AND4_X1 port map( A1 => A(11), A2 => A(10), A3 => A(8), A4 => A(9), ZN
                           => n27);
   U35 : CLKBUF_X1 port map( A => n19, Z => n28);
   U36 : OR2_X1 port map( A1 => n66, A2 => n59, ZN => n57);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n18, ZN => n29);
   U38 : AND2_X1 port map( A1 => n26, A2 => n18, ZN => n30);
   U39 : INV_X1 port map( A => n43, ZN => n31);
   U40 : NAND4_X1 port map( A1 => A(11), A2 => A(10), A3 => A(8), A4 => A(9), 
                           ZN => n66);
   U41 : NAND4_X1 port map( A1 => A(13), A2 => A(14), A3 => A(15), A4 => A(12),
                           ZN => n59);
   U42 : AND4_X1 port map( A1 => n49, A2 => n48, A3 => n32, A4 => n27, ZN => 
                           n42);
   U43 : INV_X1 port map( A => n52, ZN => n32);
   U44 : XOR2_X1 port map( A => A(26), B => n3, Z => SUM_26_port);
   U45 : NAND2_X1 port map( A1 => n106, A2 => n2, ZN => n103);
   U46 : OR2_X1 port map( A1 => n72, A2 => n33, ZN => n87);
   U47 : OR2_X1 port map( A1 => n73, A2 => n70, ZN => n33);
   U48 : INV_X1 port map( A => A(31), ZN => n39);
   U49 : INV_X1 port map( A => SUM_0_port, ZN => n34);
   U50 : NOR2_X1 port map( A1 => n47, A2 => n96, ZN => n35);
   U51 : NOR2_X1 port map( A1 => n36, A2 => n46, ZN => n67);
   U52 : OR2_X1 port map( A1 => n74, A2 => n37, ZN => n36);
   U53 : INV_X1 port map( A => A(24), ZN => n37);
   U54 : OR2_X1 port map( A1 => n96, A2 => n55, ZN => n38);
   U55 : OR2_X1 port map( A1 => n96, A2 => n55, ZN => n95);
   U56 : XNOR2_X1 port map( A => n39, B => n40, ZN => SUM_31_port);
   U57 : AND2_X1 port map( A1 => A(30), A2 => n86, ZN => n40);
   U58 : XOR2_X1 port map( A => A(20), B => n1, Z => SUM_20_port);
   U59 : XOR2_X1 port map( A => A(11), B => n41, Z => SUM_11_port);
   U60 : AND2_X1 port map( A1 => n107, A2 => n17, ZN => n41);
   U61 : NAND2_X1 port map( A1 => n30, A2 => n42, ZN => n99);
   U62 : INV_X1 port map( A => n30, ZN => n43);
   U63 : INV_X1 port map( A => n101, ZN => n44);
   U64 : OR2_X1 port map( A1 => n57, A2 => n29, ZN => n100);
   U65 : BUF_X1 port map( A => n99, Z => n45);
   U66 : OR2_X1 port map( A1 => n50, A2 => n57, ZN => n46);
   U67 : OR2_X1 port map( A1 => n91, A2 => n74, ZN => n47);
   U68 : AND2_X1 port map( A1 => n6, A2 => A(14), ZN => n48);
   U69 : AND2_X1 port map( A1 => n9, A2 => A(13), ZN => n49);
   U70 : OR2_X1 port map( A1 => n76, A2 => n60, ZN => n50);
   U71 : CLKBUF_X1 port map( A => A(9), Z => n51);
   U72 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n52);
   U73 : OR2_X1 port map( A1 => n60, A2 => n74, ZN => n53);
   U74 : CLKBUF_X1 port map( A => n21, Z => n54);
   U75 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n55);
   U76 : CLKBUF_X1 port map( A => n13, Z => n56);
   U77 : OR2_X1 port map( A1 => n29, A2 => n24, ZN => n104);
   U78 : INV_X1 port map( A => A(29), ZN => n58);
   U79 : XNOR2_X1 port map( A => n61, B => n58, ZN => SUM_29_port);
   U80 : NOR2_X1 port map( A1 => n88, A2 => n89, ZN => n61);
   U81 : XOR2_X1 port map( A => A(17), B => n62, Z => SUM_17_port);
   U82 : AND2_X1 port map( A1 => n23, A2 => n101, ZN => n62);
   U83 : XOR2_X1 port map( A => n63, B => A(21), Z => SUM_21_port);
   U84 : AND2_X1 port map( A1 => n97, A2 => A(20), ZN => n63);
   U85 : XOR2_X1 port map( A => n64, B => A(23), Z => SUM_23_port);
   U86 : AND2_X1 port map( A1 => n94, A2 => A(22), ZN => n64);
   U87 : XOR2_X1 port map( A => n14, B => n65, Z => SUM_15_port);
   U88 : AND2_X1 port map( A1 => n102, A2 => n22, ZN => n65);
   U89 : XNOR2_X1 port map( A => n38, B => A(22), ZN => SUM_22_port);
   U90 : XNOR2_X1 port map( A => n22, B => n103, ZN => SUM_14_port);
   U91 : XNOR2_X1 port map( A => n51, B => n75, ZN => SUM_9_port);
   U92 : NAND2_X1 port map( A1 => n56, A2 => n31, ZN => n75);
   U93 : XOR2_X1 port map( A => n67, B => A(25), Z => SUM_25_port);
   U94 : OR2_X1 port map( A1 => n68, A2 => n80, ZN => n79);
   U95 : NAND2_X1 port map( A1 => A(5), A2 => n19, ZN => n68);
   U96 : XNOR2_X1 port map( A => n8, B => n83, ZN => SUM_3_port);
   U97 : INV_X1 port map( A => n85, ZN => n84);
   U98 : NAND2_X1 port map( A1 => A(27), A2 => A(26), ZN => n90);
   U99 : XOR2_X1 port map( A => A(19), B => n69, Z => SUM_19_port);
   U100 : AND2_X1 port map( A1 => n98, A2 => A(18), ZN => n69);
   U101 : XNOR2_X1 port map( A => n10, B => n105, ZN => SUM_13_port);
   U102 : NAND2_X1 port map( A1 => n54, A2 => n106, ZN => n105);
   U103 : XNOR2_X1 port map( A => n25, B => n79, ZN => SUM_6_port);
   U104 : XNOR2_X1 port map( A => A(18), B => n45, ZN => SUM_18_port);
   U105 : XNOR2_X1 port map( A => n7, B => n81, ZN => SUM_5_port);
   U106 : INV_X1 port map( A => n80, ZN => n82);
   U107 : XNOR2_X1 port map( A => n108, B => n17, ZN => SUM_10_port);
   U108 : NAND2_X1 port map( A1 => A(28), A2 => A(29), ZN => n70);
   U109 : NAND2_X1 port map( A1 => A(23), A2 => A(22), ZN => n92);
   U110 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n93);
   U111 : XOR2_X1 port map( A => A(27), B => n71, Z => SUM_27_port);
   U112 : AND2_X1 port map( A1 => n35, A2 => A(26), ZN => n71);
   U113 : INV_X1 port map( A => A(28), ZN => n89);
   U114 : NAND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n91);
   U115 : XNOR2_X1 port map( A => n87, B => A(30), ZN => SUM_30_port);
   U116 : XNOR2_X1 port map( A => A(28), B => n88, ZN => SUM_28_port);
   U117 : OR2_X1 port map( A1 => n90, A2 => n91, ZN => n73);
   U118 : XNOR2_X1 port map( A => n20, B => n85, ZN => SUM_2_port);
   U119 : OR2_X1 port map( A1 => n92, A2 => n93, ZN => n74);
   U120 : NAND2_X1 port map( A1 => n28, A2 => n82, ZN => n81);
   U121 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => n76);
   U122 : XNOR2_X1 port map( A => n23, B => n44, ZN => SUM_16_port);
   U123 : INV_X1 port map( A => n100, ZN => n101);
   U124 : XNOR2_X1 port map( A => n54, B => n104, ZN => SUM_12_port);
   U125 : INV_X1 port map( A => n104, ZN => n106);
   U126 : INV_X1 port map( A => n46, ZN => n97);
   U127 : XOR2_X1 port map( A => n12, B => n34, Z => SUM_1_port);
   U128 : XNOR2_X1 port map( A => n56, B => n43, ZN => SUM_8_port);
   U129 : XNOR2_X1 port map( A => A(24), B => n72, ZN => SUM_24_port);
   U130 : NAND2_X1 port map( A1 => n20, A2 => n84, ZN => n83);
   U131 : INV_X1 port map( A => n11, ZN => SUM_0_port);
   U132 : NAND2_X1 port map( A1 => n12, A2 => n34, ZN => n85);
   U133 : NAND4_X1 port map( A1 => n20, A2 => n8, A3 => A(1), A4 => n11, ZN => 
                           n80);
   U134 : XNOR2_X1 port map( A => n5, B => n77, ZN => SUM_7_port);
   U135 : NAND2_X1 port map( A1 => n78, A2 => n25, ZN => n77);
   U136 : INV_X1 port map( A => n79, ZN => n78);
   U137 : XNOR2_X1 port map( A => n28, B => n80, ZN => SUM_4_port);
   U138 : INV_X1 port map( A => n87, ZN => n86);
   U139 : INV_X1 port map( A => n95, ZN => n94);
   U140 : INV_X1 port map( A => n99, ZN => n98);
   U141 : INV_X1 port map( A => n103, ZN => n102);
   U142 : INV_X1 port map( A => n108, ZN => n107);
   U143 : NAND3_X1 port map( A1 => n13, A2 => n51, A3 => n30, ZN => n108);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_6 
   is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_6;

architecture SYN_cla of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_6 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port );
   
   U2 : CLKBUF_X1 port map( A => A(2), Z => n1);
   U3 : AND2_X1 port map( A1 => n40, A2 => n2, ZN => n34);
   U4 : AND2_X1 port map( A1 => n27, A2 => n3, ZN => n2);
   U5 : INV_X1 port map( A => n41, ZN => n3);
   U6 : AND2_X2 port map( A1 => n16, A2 => n15, ZN => n40);
   U7 : AND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n4);
   U8 : AND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n5);
   U9 : CLKBUF_X1 port map( A => A(8), Z => n6);
   U10 : NOR2_X1 port map( A1 => n55, A2 => n7, ZN => n37);
   U11 : OR2_X1 port map( A1 => n58, A2 => n76, ZN => n7);
   U12 : NAND2_X1 port map( A1 => n17, A2 => n4, ZN => n95);
   U13 : BUF_X1 port map( A => n49, Z => n8);
   U14 : AND3_X1 port map( A1 => n11, A2 => n13, A3 => n91, ZN => n9);
   U15 : AND2_X1 port map( A1 => n56, A2 => n85, ZN => n10);
   U16 : AND2_X1 port map( A1 => n56, A2 => n85, ZN => n23);
   U17 : AND4_X1 port map( A1 => A(1), A2 => A(0), A3 => A(2), A4 => A(3), ZN 
                           => n11);
   U18 : AND4_X1 port map( A1 => A(1), A2 => A(0), A3 => A(2), A4 => A(3), ZN 
                           => n97);
   U19 : NAND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n12);
   U20 : AND4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(7), A4 => A(6), ZN 
                           => n13);
   U21 : CLKBUF_X1 port map( A => A(4), Z => n14);
   U22 : AND4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(7), A4 => A(6), ZN 
                           => n96);
   U23 : NOR2_X1 port map( A1 => n92, A2 => n12, ZN => n15);
   U24 : AND2_X1 port map( A1 => n11, A2 => n13, ZN => n16);
   U25 : AND2_X1 port map( A1 => n97, A2 => n96, ZN => n17);
   U26 : AND2_X1 port map( A1 => n97, A2 => n96, ZN => n57);
   U27 : AND4_X1 port map( A1 => n85, A2 => n17, A3 => n4, A4 => n18, ZN => n49
                           );
   U28 : INV_X1 port map( A => n92, ZN => n18);
   U29 : AND3_X1 port map( A1 => n11, A2 => n13, A3 => n91, ZN => n25);
   U30 : CLKBUF_X1 port map( A => n16, Z => n19);
   U31 : XOR2_X1 port map( A => A(26), B => n20, Z => SUM_26_port);
   U32 : AND3_X1 port map( A1 => A(24), A2 => A(25), A3 => n39, ZN => n20);
   U33 : NAND2_X1 port map( A1 => n8, A2 => n21, ZN => n72);
   U34 : AND2_X1 port map( A1 => n50, A2 => n22, ZN => n21);
   U35 : INV_X1 port map( A => n47, ZN => n22);
   U36 : CLKBUF_X1 port map( A => A(1), Z => n24);
   U37 : INV_X1 port map( A => SUM_0_port, ZN => n26);
   U38 : NAND2_X1 port map( A1 => n40, A2 => n27, ZN => n82);
   U39 : AND2_X1 port map( A1 => n85, A2 => n28, ZN => n27);
   U40 : INV_X1 port map( A => n58, ZN => n28);
   U41 : XOR2_X1 port map( A => A(11), B => n29, Z => SUM_11_port);
   U42 : AND2_X1 port map( A1 => n94, A2 => A(10), ZN => n29);
   U43 : XOR2_X1 port map( A => A(15), B => n30, Z => SUM_15_port);
   U44 : AND2_X1 port map( A1 => n88, A2 => A(14), ZN => n30);
   U45 : AND2_X1 port map( A1 => n49, A2 => n50, ZN => n31);
   U46 : NOR2_X2 port map( A1 => n55, A2 => n58, ZN => n50);
   U47 : INV_X1 port map( A => n34, ZN => n81);
   U48 : AND2_X1 port map( A1 => n23, A2 => n5, ZN => n32);
   U49 : CLKBUF_X1 port map( A => n82, Z => n33);
   U50 : XOR2_X1 port map( A => A(17), B => n35, Z => SUM_17_port);
   U51 : AND2_X1 port map( A1 => A(16), A2 => n10, ZN => n35);
   U52 : AND2_X1 port map( A1 => n25, A2 => n85, ZN => n36);
   U53 : AND2_X1 port map( A1 => n36, A2 => n37, ZN => n77);
   U54 : XOR2_X1 port map( A => A(25), B => n38, Z => SUM_25_port);
   U55 : AND2_X1 port map( A1 => A(24), A2 => n31, ZN => n38);
   U56 : AND2_X1 port map( A1 => n36, A2 => n50, ZN => n39);
   U57 : NAND2_X1 port map( A1 => n10, A2 => n5, ZN => n84);
   U58 : AND2_X1 port map( A1 => n57, A2 => n15, ZN => n56);
   U59 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n41);
   U60 : CLKBUF_X1 port map( A => n1, Z => n42);
   U61 : XOR2_X1 port map( A => A(19), B => n43, Z => SUM_19_port);
   U62 : AND2_X1 port map( A1 => n32, A2 => A(18), ZN => n43);
   U63 : INV_X1 port map( A => n10, ZN => n44);
   U64 : NAND2_X1 port map( A1 => n31, A2 => n45, ZN => n71);
   U65 : NOR2_X1 port map( A1 => n52, A2 => n47, ZN => n45);
   U66 : XOR2_X1 port map( A => A(27), B => n46, Z => SUM_27_port);
   U67 : AND2_X1 port map( A1 => n77, A2 => A(26), ZN => n46);
   U68 : OR2_X1 port map( A1 => n75, A2 => n76, ZN => n47);
   U69 : XOR2_X1 port map( A => n73, B => A(29), Z => SUM_29_port);
   U70 : XOR2_X1 port map( A => n48, B => A(21), Z => SUM_21_port);
   U71 : AND2_X1 port map( A1 => A(20), A2 => n83, ZN => n48);
   U72 : NAND2_X1 port map( A1 => n8, A2 => n50, ZN => n78);
   U73 : XNOR2_X1 port map( A => n24, B => SUM_0_port, ZN => SUM_1_port);
   U74 : NAND2_X1 port map( A1 => A(27), A2 => A(26), ZN => n75);
   U75 : NAND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n76);
   U76 : XOR2_X1 port map( A => n51, B => A(23), Z => SUM_23_port);
   U77 : AND2_X1 port map( A1 => n34, A2 => A(22), ZN => n51);
   U78 : XOR2_X1 port map( A => n6, B => n19, Z => SUM_8_port);
   U79 : XNOR2_X1 port map( A => n81, B => A(22), ZN => SUM_22_port);
   U80 : XNOR2_X1 port map( A => n89, B => A(14), ZN => SUM_14_port);
   U81 : XNOR2_X1 port map( A => A(28), B => n72, ZN => SUM_28_port);
   U82 : XNOR2_X1 port map( A => A(9), B => n59, ZN => SUM_9_port);
   U83 : XNOR2_X1 port map( A => A(30), B => n71, ZN => SUM_30_port);
   U84 : NOR2_X1 port map( A1 => n72, A2 => n74, ZN => n73);
   U85 : INV_X1 port map( A => A(28), ZN => n74);
   U86 : OR2_X1 port map( A1 => n98, A2 => n63, ZN => n62);
   U87 : XNOR2_X1 port map( A => A(13), B => n90, ZN => SUM_13_port);
   U88 : NOR2_X1 port map( A1 => n86, A2 => n87, ZN => n85);
   U89 : NAND2_X1 port map( A1 => A(15), A2 => A(14), ZN => n86);
   U90 : NAND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n87);
   U91 : XNOR2_X1 port map( A => A(18), B => n84, ZN => SUM_18_port);
   U92 : NOR2_X1 port map( A1 => n92, A2 => n93, ZN => n91);
   U93 : NAND2_X1 port map( A1 => A(11), A2 => A(10), ZN => n92);
   U94 : NAND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n93);
   U95 : NAND2_X1 port map( A1 => A(28), A2 => A(29), ZN => n52);
   U96 : XOR2_X1 port map( A => A(12), B => n40, Z => SUM_12_port);
   U97 : XNOR2_X1 port map( A => A(10), B => n95, ZN => SUM_10_port);
   U98 : XNOR2_X1 port map( A => A(3), B => n66, ZN => SUM_3_port);
   U99 : INV_X1 port map( A => n68, ZN => n67);
   U100 : XNOR2_X1 port map( A => A(5), B => n64, ZN => SUM_5_port);
   U101 : INV_X1 port map( A => n63, ZN => n65);
   U102 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => n58);
   U103 : AND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n53);
   U104 : AND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n54);
   U105 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n80);
   U106 : NAND2_X1 port map( A1 => A(23), A2 => A(22), ZN => n79);
   U107 : OR2_X1 port map( A1 => n79, A2 => n80, ZN => n55);
   U108 : NAND2_X1 port map( A1 => A(12), A2 => n9, ZN => n90);
   U109 : NAND2_X1 port map( A1 => n6, A2 => n19, ZN => n59);
   U110 : XNOR2_X1 port map( A => A(6), B => n62, ZN => SUM_6_port);
   U111 : INV_X1 port map( A => n33, ZN => n83);
   U112 : XNOR2_X1 port map( A => n82, B => A(20), ZN => SUM_20_port);
   U113 : XNOR2_X1 port map( A => A(16), B => n44, ZN => SUM_16_port);
   U114 : NAND2_X1 port map( A1 => n14, A2 => n65, ZN => n64);
   U115 : NAND2_X1 port map( A1 => A(5), A2 => A(4), ZN => n98);
   U116 : XNOR2_X1 port map( A => n42, B => n68, ZN => SUM_2_port);
   U117 : NAND2_X1 port map( A1 => n1, A2 => n67, ZN => n66);
   U118 : XNOR2_X1 port map( A => A(24), B => n78, ZN => SUM_24_port);
   U119 : INV_X1 port map( A => A(0), ZN => SUM_0_port);
   U120 : NAND2_X1 port map( A1 => n24, A2 => n26, ZN => n68);
   U121 : NAND4_X1 port map( A1 => A(3), A2 => A(2), A3 => A(1), A4 => A(0), ZN
                           => n63);
   U122 : XNOR2_X1 port map( A => A(7), B => n60, ZN => SUM_7_port);
   U123 : NAND2_X1 port map( A1 => n61, A2 => A(6), ZN => n60);
   U124 : INV_X1 port map( A => n62, ZN => n61);
   U125 : XNOR2_X1 port map( A => n14, B => n63, ZN => SUM_4_port);
   U126 : XNOR2_X1 port map( A => A(31), B => n69, ZN => SUM_31_port);
   U127 : NAND2_X1 port map( A1 => A(30), A2 => n70, ZN => n69);
   U128 : INV_X1 port map( A => n71, ZN => n70);
   U129 : INV_X1 port map( A => n89, ZN => n88);
   U130 : NAND3_X1 port map( A1 => A(12), A2 => A(13), A3 => n9, ZN => n89);
   U131 : INV_X1 port map( A => n95, ZN => n94);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 
   is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5;

architecture SYN_cla of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 
   is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => n46, A2 => n36, ZN => n17);
   U3 : OR2_X1 port map( A1 => n19, A2 => n61, ZN => n43);
   U4 : INV_X1 port map( A => n68, ZN => n67);
   U5 : INV_X1 port map( A => n17, ZN => n89);
   U6 : INV_X1 port map( A => n14, ZN => n83);
   U7 : AND2_X1 port map( A1 => n13, A2 => A(17), ZN => n1);
   U8 : AND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n2);
   U9 : AND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n3);
   U10 : NOR2_X1 port map( A1 => n80, A2 => n61, ZN => n4);
   U11 : AND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n5);
   U12 : AND2_X1 port map( A1 => n27, A2 => n24, ZN => n6);
   U13 : AND2_X1 port map( A1 => n94, A2 => n95, ZN => n7);
   U14 : AND2_X1 port map( A1 => n94, A2 => n95, ZN => n8);
   U15 : AND2_X1 port map( A1 => n94, A2 => n95, ZN => n59);
   U16 : BUF_X1 port map( A => n12, Z => n39);
   U17 : AND4_X1 port map( A1 => A(15), A2 => A(14), A3 => A(12), A4 => A(13), 
                           ZN => n9);
   U18 : AND4_X1 port map( A1 => A(15), A2 => A(14), A3 => A(12), A4 => A(13), 
                           ZN => n30);
   U19 : AND4_X2 port map( A1 => A(8), A2 => A(9), A3 => A(10), A4 => A(11), ZN
                           => n90);
   U20 : CLKBUF_X1 port map( A => A(2), Z => n10);
   U21 : CLKBUF_X1 port map( A => A(1), Z => n11);
   U22 : NAND2_X1 port map( A1 => n15, A2 => n7, ZN => n12);
   U23 : CLKBUF_X1 port map( A => A(16), Z => n13);
   U24 : AND4_X2 port map( A1 => n9, A2 => n90, A3 => n3, A4 => n2, ZN => n15);
   U25 : AND2_X2 port map( A1 => n50, A2 => n8, ZN => n14);
   U26 : AND4_X1 port map( A1 => n90, A2 => n30, A3 => n3, A4 => n2, ZN => n40)
                           ;
   U27 : CLKBUF_X1 port map( A => A(4), Z => n16);
   U28 : XOR2_X1 port map( A => n29, B => n18, Z => SUM(13));
   U29 : AND2_X1 port map( A1 => n35, A2 => n17, ZN => n18);
   U30 : AND2_X1 port map( A1 => n46, A2 => n6, ZN => n92);
   U31 : NAND2_X1 port map( A1 => n15, A2 => n7, ZN => n19);
   U32 : AND3_X1 port map( A1 => A(18), A2 => n14, A3 => n1, ZN => n57);
   U33 : NOR2_X1 port map( A1 => n71, A2 => n70, ZN => n69);
   U34 : AND4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(7), A4 => A(6), ZN 
                           => n37);
   U35 : NOR3_X1 port map( A1 => n20, A2 => n21, A3 => n43, ZN => n41);
   U36 : INV_X1 port map( A => A(24), ZN => n20);
   U37 : INV_X1 port map( A => A(25), ZN => n21);
   U38 : NOR2_X1 port map( A1 => n79, A2 => n22, ZN => n56);
   U39 : INV_X1 port map( A => A(22), ZN => n22);
   U40 : AND4_X1 port map( A1 => A(11), A2 => A(9), A3 => A(8), A4 => A(10), ZN
                           => n36);
   U41 : AND4_X1 port map( A1 => A(5), A2 => A(4), A3 => A(7), A4 => A(6), ZN 
                           => n94);
   U42 : AND4_X1 port map( A1 => A(1), A2 => A(0), A3 => A(3), A4 => A(2), ZN 
                           => n38);
   U43 : AND4_X1 port map( A1 => A(1), A2 => A(0), A3 => A(3), A4 => A(2), ZN 
                           => n95);
   U44 : NAND3_X1 port map( A1 => n23, A2 => n66, A3 => A(6), ZN => n62);
   U45 : INV_X1 port map( A => n55, ZN => n23);
   U46 : CLKBUF_X1 port map( A => A(8), Z => n24);
   U47 : CLKBUF_X1 port map( A => A(11), Z => n25);
   U48 : CLKBUF_X1 port map( A => A(14), Z => n26);
   U49 : CLKBUF_X1 port map( A => A(9), Z => n27);
   U50 : CLKBUF_X1 port map( A => A(10), Z => n28);
   U51 : CLKBUF_X1 port map( A => A(13), Z => n29);
   U52 : CLKBUF_X1 port map( A => n24, Z => n31);
   U53 : AND2_X1 port map( A1 => n4, A2 => n32, ZN => n60);
   U54 : AND2_X1 port map( A1 => n5, A2 => A(26), ZN => n32);
   U55 : AND2_X2 port map( A1 => n37, A2 => n38, ZN => n46);
   U56 : INV_X1 port map( A => n39, ZN => n33);
   U57 : AND2_X1 port map( A1 => n33, A2 => n34, ZN => n74);
   U58 : AND2_X1 port map( A1 => n42, A2 => A(28), ZN => n34);
   U59 : CLKBUF_X1 port map( A => A(12), Z => n35);
   U60 : NAND2_X1 port map( A1 => n14, A2 => n1, ZN => n82);
   U61 : OR2_X1 port map( A1 => n44, A2 => n12, ZN => n79);
   U62 : NAND2_X1 port map( A1 => n40, A2 => n59, ZN => n80);
   U63 : XOR2_X1 port map( A => n41, B => A(26), Z => SUM(26));
   U64 : NAND2_X1 port map( A1 => n81, A2 => n42, ZN => n71);
   U65 : NOR2_X1 port map( A1 => n61, A2 => n45, ZN => n42);
   U66 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n44);
   U67 : OR2_X1 port map( A1 => n75, A2 => n76, ZN => n45);
   U68 : INV_X1 port map( A => A(31), ZN => n49);
   U69 : CLKBUF_X1 port map( A => A(0), Z => n47);
   U70 : NOR2_X1 port map( A1 => n85, A2 => n86, ZN => n48);
   U71 : XNOR2_X1 port map( A => n69, B => n49, ZN => SUM(31));
   U72 : AND2_X1 port map( A1 => n36, A2 => n48, ZN => n50);
   U73 : XOR2_X1 port map( A => A(25), B => n51, Z => SUM(25));
   U74 : AND2_X1 port map( A1 => A(24), A2 => n4, ZN => n51);
   U75 : XOR2_X1 port map( A => A(21), B => n52, Z => SUM(21));
   U76 : AND2_X1 port map( A1 => n81, A2 => A(20), ZN => n52);
   U77 : XOR2_X1 port map( A => A(15), B => n53, Z => SUM(15));
   U78 : AND2_X1 port map( A1 => n87, A2 => n26, ZN => n53);
   U79 : NAND2_X1 port map( A1 => A(27), A2 => A(26), ZN => n75);
   U80 : NAND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n76);
   U81 : XNOR2_X1 port map( A => n28, B => n93, ZN => SUM(10));
   U82 : XNOR2_X1 port map( A => n26, B => n88, ZN => SUM(14));
   U83 : XOR2_X1 port map( A => n27, B => n54, Z => SUM(9));
   U84 : AND2_X1 port map( A1 => n31, A2 => n46, ZN => n54);
   U85 : OR2_X1 port map( A1 => n55, A2 => n64, ZN => n63);
   U86 : NAND2_X1 port map( A1 => A(5), A2 => A(4), ZN => n55);
   U87 : XNOR2_X1 port map( A => A(17), B => n84, ZN => SUM(17));
   U88 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => n84);
   U89 : XOR2_X1 port map( A => n74, B => A(29), Z => SUM(29));
   U90 : NAND2_X1 port map( A1 => A(15), A2 => A(14), ZN => n85);
   U91 : NAND2_X1 port map( A1 => A(13), A2 => A(12), ZN => n86);
   U92 : XOR2_X1 port map( A => n56, B => A(23), Z => SUM(23));
   U93 : XOR2_X1 port map( A => A(19), B => n57, Z => SUM(19));
   U94 : XNOR2_X1 port map( A => n79, B => A(22), ZN => SUM(22));
   U95 : XNOR2_X1 port map( A => A(18), B => n82, ZN => SUM(18));
   U96 : XOR2_X1 port map( A => n72, B => A(30), Z => SUM(30));
   U97 : XNOR2_X1 port map( A => A(5), B => n65, ZN => SUM(5));
   U98 : INV_X1 port map( A => n64, ZN => n66);
   U99 : XOR2_X1 port map( A => n31, B => n46, Z => SUM(8));
   U100 : NAND2_X1 port map( A1 => A(23), A2 => A(22), ZN => n77);
   U101 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n78);
   U102 : NAND2_X1 port map( A1 => A(28), A2 => A(29), ZN => n73);
   U103 : XOR2_X1 port map( A => A(3), B => n58, Z => SUM(3));
   U104 : AND2_X1 port map( A1 => n10, A2 => n67, ZN => n58);
   U105 : NOR2_X1 port map( A1 => n71, A2 => n73, ZN => n72);
   U106 : XNOR2_X1 port map( A => n71, B => A(28), ZN => SUM(28));
   U107 : XOR2_X1 port map( A => n60, B => A(27), Z => SUM(27));
   U108 : XNOR2_X1 port map( A => A(6), B => n63, ZN => SUM(6));
   U109 : NAND2_X1 port map( A1 => n16, A2 => n66, ZN => n65);
   U110 : OR2_X1 port map( A1 => n77, A2 => n78, ZN => n61);
   U111 : XNOR2_X1 port map( A => n43, B => A(24), ZN => SUM(24));
   U112 : XNOR2_X1 port map( A => A(20), B => n39, ZN => SUM(20));
   U113 : INV_X1 port map( A => n80, ZN => n81);
   U114 : XNOR2_X1 port map( A => n13, B => n83, ZN => SUM(16));
   U115 : XNOR2_X1 port map( A => n35, B => n89, ZN => SUM(12));
   U116 : XNOR2_X1 port map( A => n10, B => n68, ZN => SUM(2));
   U117 : INV_X1 port map( A => n47, ZN => SUM(0));
   U118 : NAND2_X1 port map( A1 => n11, A2 => n47, ZN => n68);
   U119 : NAND4_X1 port map( A1 => A(3), A2 => A(2), A3 => A(1), A4 => A(0), ZN
                           => n64);
   U120 : XNOR2_X1 port map( A => A(7), B => n62, ZN => SUM(7));
   U121 : XNOR2_X1 port map( A => n16, B => n64, ZN => SUM(4));
   U122 : NAND3_X1 port map( A1 => A(30), A2 => A(29), A3 => A(28), ZN => n70);
   U123 : XOR2_X1 port map( A => n11, B => n47, Z => SUM(1));
   U124 : INV_X1 port map( A => n88, ZN => n87);
   U125 : NAND3_X1 port map( A1 => n35, A2 => n29, A3 => n17, ZN => n88);
   U126 : XNOR2_X1 port map( A => n25, B => n91, ZN => SUM(11));
   U127 : NAND2_X1 port map( A1 => n92, A2 => n28, ZN => n91);
   U128 : NAND3_X1 port map( A1 => n24, A2 => n27, A3 => n46, ZN => n93);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 
   is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4;

architecture SYN_cla of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 
   is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port );
   
   U2 : INV_X1 port map( A => A(2), ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => n2);
   U4 : AND2_X2 port map( A1 => n29, A2 => n78, ZN => n26);
   U5 : AND2_X2 port map( A1 => n85, A2 => n84, ZN => n12);
   U6 : AND2_X2 port map( A1 => n12, A2 => n78, ZN => n15);
   U7 : AND2_X1 port map( A1 => n15, A2 => n72, ZN => n22);
   U8 : AND2_X1 port map( A1 => n25, A2 => n24, ZN => n30);
   U9 : AND3_X1 port map( A1 => n8, A2 => A(17), A3 => n22, ZN => n3);
   U10 : AND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n4);
   U11 : AND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n5);
   U12 : NOR2_X1 port map( A1 => n69, A2 => n70, ZN => n6);
   U13 : AND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n7);
   U14 : CLKBUF_X1 port map( A => A(16), Z => n8);
   U15 : AND4_X1 port map( A1 => A(1), A2 => A(0), A3 => A(3), A4 => A(2), ZN 
                           => n9);
   U16 : AND4_X1 port map( A1 => A(1), A2 => A(0), A3 => A(3), A4 => A(2), ZN 
                           => n85);
   U17 : XOR2_X1 port map( A => A(18), B => n3, Z => SUM_18_port);
   U18 : AND2_X1 port map( A1 => n5, A2 => n24, ZN => n10);
   U19 : XOR2_X1 port map( A => A(7), B => n11, Z => SUM_7_port);
   U20 : AND2_X1 port map( A1 => n40, A2 => A(6), ZN => n11);
   U21 : AND2_X2 port map( A1 => n23, A2 => n26, ZN => n28);
   U22 : AND2_X1 port map( A1 => n15, A2 => n4, ZN => n13);
   U23 : CLKBUF_X1 port map( A => n26, Z => n14);
   U24 : INV_X1 port map( A => n14, ZN => n27);
   U25 : CLKBUF_X1 port map( A => A(4), Z => n16);
   U26 : AND4_X2 port map( A1 => A(5), A2 => A(4), A3 => A(7), A4 => A(6), ZN 
                           => n84);
   U27 : AND3_X1 port map( A1 => n64, A2 => n72, A3 => n6, ZN => n23);
   U28 : AND2_X1 port map( A1 => n58, A2 => n26, ZN => n17);
   U29 : XOR2_X1 port map( A => A(25), B => n18, Z => SUM_25_port);
   U30 : AND2_X1 port map( A1 => A(24), A2 => n28, ZN => n18);
   U31 : AND2_X1 port map( A1 => n9, A2 => n84, ZN => n19);
   U32 : CLKBUF_X1 port map( A => n2, Z => n20);
   U33 : AND2_X1 port map( A1 => n9, A2 => n84, ZN => n29);
   U34 : AND2_X1 port map( A1 => n28, A2 => n7, ZN => n61);
   U35 : INV_X1 port map( A => n22, ZN => n71);
   U36 : AND2_X1 port map( A1 => n10, A2 => n25, ZN => n21);
   U37 : NAND2_X1 port map( A1 => n26, A2 => n4, ZN => n76);
   U38 : NAND2_X1 port map( A1 => n30, A2 => n5, ZN => n67);
   U39 : INV_X1 port map( A => n28, ZN => n63);
   U40 : INV_X1 port map( A => n19, ZN => n39);
   U41 : AND2_X1 port map( A1 => n29, A2 => n78, ZN => n24);
   U42 : AND2_X1 port map( A1 => n72, A2 => n6, ZN => n25);
   U43 : INV_X1 port map( A => n30, ZN => n68);
   U44 : INV_X1 port map( A => SUM_0_port, ZN => n31);
   U45 : XOR2_X1 port map( A => A(9), B => n32, Z => SUM_9_port);
   U46 : AND2_X1 port map( A1 => A(8), A2 => n19, ZN => n32);
   U47 : XOR2_X1 port map( A => A(21), B => n33, Z => SUM_21_port);
   U48 : AND2_X1 port map( A1 => A(20), A2 => n30, ZN => n33);
   U49 : XOR2_X1 port map( A => A(17), B => n34, Z => SUM_17_port);
   U50 : AND2_X1 port map( A1 => A(16), A2 => n22, ZN => n34);
   U51 : NOR2_X1 port map( A1 => n73, A2 => n74, ZN => n72);
   U52 : NAND2_X1 port map( A1 => A(15), A2 => A(14), ZN => n73);
   U53 : NAND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n74);
   U54 : NAND2_X1 port map( A1 => n17, A2 => n23, ZN => n51);
   U55 : NOR2_X1 port map( A1 => n59, A2 => n60, ZN => n58);
   U56 : NAND2_X1 port map( A1 => A(27), A2 => A(26), ZN => n59);
   U57 : NAND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n60);
   U58 : INV_X1 port map( A => A(30), ZN => n53);
   U59 : NOR2_X1 port map( A1 => n51, A2 => n54, ZN => n52);
   U60 : NOR2_X1 port map( A1 => n79, A2 => n80, ZN => n78);
   U61 : NAND2_X1 port map( A1 => A(11), A2 => A(10), ZN => n79);
   U62 : NAND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n80);
   U63 : NOR2_X1 port map( A1 => n65, A2 => n66, ZN => n64);
   U64 : NAND2_X1 port map( A1 => A(23), A2 => A(22), ZN => n65);
   U65 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n66);
   U66 : XOR2_X1 port map( A => A(19), B => n35, Z => SUM_19_port);
   U67 : AND2_X1 port map( A1 => n3, A2 => A(18), ZN => n35);
   U68 : XOR2_X1 port map( A => A(23), B => n36, Z => SUM_23_port);
   U69 : AND2_X1 port map( A1 => n21, A2 => A(22), ZN => n36);
   U70 : XNOR2_X1 port map( A => A(14), B => n76, ZN => SUM_14_port);
   U71 : XNOR2_X1 port map( A => A(10), B => n83, ZN => SUM_10_port);
   U72 : XNOR2_X1 port map( A => A(22), B => n67, ZN => SUM_22_port);
   U73 : XNOR2_X1 port map( A => A(3), B => n45, ZN => SUM_3_port);
   U74 : INV_X1 port map( A => n47, ZN => n46);
   U75 : NAND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n69);
   U76 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n70);
   U77 : XNOR2_X1 port map( A => A(5), B => n43, ZN => SUM_5_port);
   U78 : INV_X1 port map( A => n42, ZN => n44);
   U79 : XNOR2_X1 port map( A => A(13), B => n77, ZN => SUM_13_port);
   U80 : NAND2_X1 port map( A1 => A(12), A2 => n15, ZN => n77);
   U81 : OR2_X1 port map( A1 => n37, A2 => n42, ZN => n41);
   U82 : NAND2_X1 port map( A1 => A(5), A2 => A(4), ZN => n37);
   U83 : NAND2_X1 port map( A1 => A(28), A2 => A(29), ZN => n54);
   U84 : INV_X1 port map( A => A(31), ZN => n49);
   U85 : NOR2_X1 port map( A1 => n51, A2 => n50, ZN => n48);
   U86 : INV_X1 port map( A => A(29), ZN => n56);
   U87 : NOR2_X1 port map( A1 => n51, A2 => n57, ZN => n55);
   U88 : INV_X1 port map( A => A(28), ZN => n57);
   U89 : XNOR2_X1 port map( A => n55, B => n56, ZN => SUM_29_port);
   U90 : XNOR2_X1 port map( A => n52, B => n53, ZN => SUM_30_port);
   U91 : XNOR2_X1 port map( A => n48, B => n49, ZN => SUM_31_port);
   U92 : XNOR2_X1 port map( A => A(26), B => n62, ZN => SUM_26_port);
   U93 : XNOR2_X1 port map( A => n51, B => A(28), ZN => SUM_28_port);
   U94 : XNOR2_X1 port map( A => A(6), B => n41, ZN => SUM_6_port);
   U95 : XOR2_X1 port map( A => A(27), B => n38, Z => SUM_27_port);
   U96 : AND2_X1 port map( A1 => n61, A2 => A(26), ZN => n38);
   U97 : NAND2_X1 port map( A1 => n16, A2 => n44, ZN => n43);
   U98 : XNOR2_X1 port map( A => A(20), B => n68, ZN => SUM_20_port);
   U99 : XNOR2_X1 port map( A => n20, B => n47, ZN => SUM_2_port);
   U100 : XNOR2_X1 port map( A => n8, B => n71, ZN => SUM_16_port);
   U101 : NAND2_X1 port map( A1 => n2, A2 => n46, ZN => n45);
   U102 : INV_X1 port map( A => A(0), ZN => SUM_0_port);
   U103 : XNOR2_X1 port map( A => A(12), B => n27, ZN => SUM_12_port);
   U104 : NAND2_X1 port map( A1 => A(1), A2 => n31, ZN => n47);
   U105 : NAND4_X1 port map( A1 => A(3), A2 => A(2), A3 => A(1), A4 => A(0), ZN
                           => n42);
   U106 : XNOR2_X1 port map( A => A(24), B => n63, ZN => SUM_24_port);
   U107 : XNOR2_X1 port map( A => A(8), B => n39, ZN => SUM_8_port);
   U108 : INV_X1 port map( A => n41, ZN => n40);
   U109 : XNOR2_X1 port map( A => n16, B => n42, ZN => SUM_4_port);
   U110 : NAND3_X1 port map( A1 => A(30), A2 => A(29), A3 => A(28), ZN => n50);
   U111 : NAND3_X1 port map( A1 => A(24), A2 => A(25), A3 => n28, ZN => n62);
   U112 : XOR2_X1 port map( A => A(1), B => n31, Z => SUM_1_port);
   U113 : XNOR2_X1 port map( A => A(15), B => n75, ZN => SUM_15_port);
   U114 : NAND2_X1 port map( A1 => n13, A2 => A(14), ZN => n75);
   U115 : XNOR2_X1 port map( A => A(11), B => n81, ZN => SUM_11_port);
   U116 : NAND2_X1 port map( A1 => n82, A2 => A(10), ZN => n81);
   U117 : INV_X1 port map( A => n83, ZN => n82);
   U118 : NAND3_X1 port map( A1 => A(8), A2 => A(9), A3 => n12, ZN => n83);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_15;

architecture SYN_BEHAVIORAL of RCA_NBIT4_15 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_14;

architecture SYN_BEHAVIORAL of RCA_NBIT4_14 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_13;

architecture SYN_BEHAVIORAL of RCA_NBIT4_13 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_12;

architecture SYN_BEHAVIORAL of RCA_NBIT4_12 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_11;

architecture SYN_BEHAVIORAL of RCA_NBIT4_11 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_10;

architecture SYN_BEHAVIORAL of RCA_NBIT4_10 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_9;

architecture SYN_BEHAVIORAL of RCA_NBIT4_9 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_8;

architecture SYN_BEHAVIORAL of RCA_NBIT4_8 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_7;

architecture SYN_BEHAVIORAL of RCA_NBIT4_7 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_6;

architecture SYN_BEHAVIORAL of RCA_NBIT4_6 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_5;

architecture SYN_BEHAVIORAL of RCA_NBIT4_5 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_4;

architecture SYN_BEHAVIORAL of RCA_NBIT4_4 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_3;

architecture SYN_BEHAVIORAL of RCA_NBIT4_3 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_2;

architecture SYN_BEHAVIORAL of RCA_NBIT4_2 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_1;

architecture SYN_BEHAVIORAL of RCA_NBIT4_1 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_42 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_42;

architecture SYN_behave of P_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_41 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_41;

architecture SYN_behave of P_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_40 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_40;

architecture SYN_behave of P_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_39 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_39;

architecture SYN_behave of P_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_38 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_38;

architecture SYN_behave of P_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_37 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_37;

architecture SYN_behave of P_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_36 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_36;

architecture SYN_behave of P_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_35 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_35;

architecture SYN_behave of P_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_34 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_34;

architecture SYN_behave of P_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_33 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_33;

architecture SYN_behave of P_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_32 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_32;

architecture SYN_behave of P_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_31 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_31;

architecture SYN_behave of P_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_30 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_30;

architecture SYN_behave of P_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_29 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_29;

architecture SYN_behave of P_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_28 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_28;

architecture SYN_behave of P_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_27 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_27;

architecture SYN_behave of P_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_26 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_26;

architecture SYN_behave of P_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_25 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_25;

architecture SYN_behave of P_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_24 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_24;

architecture SYN_behave of P_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_23 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_23;

architecture SYN_behave of P_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_22 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_22;

architecture SYN_behave of P_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_21 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_21;

architecture SYN_behave of P_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_20 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_20;

architecture SYN_behave of P_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_19 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_19;

architecture SYN_behave of P_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_18 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_18;

architecture SYN_behave of P_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_17 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_17;

architecture SYN_behave of P_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_16 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_16;

architecture SYN_behave of P_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_15 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_15;

architecture SYN_behave of P_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_14 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_14;

architecture SYN_behave of P_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_13 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_13;

architecture SYN_behave of P_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_12 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_12;

architecture SYN_behave of P_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_11 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_11;

architecture SYN_behave of P_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_10 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_10;

architecture SYN_behave of P_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_9 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_9;

architecture SYN_behave of P_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_8 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_8;

architecture SYN_behave of P_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_7 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_7;

architecture SYN_behave of P_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_6 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_6;

architecture SYN_behave of P_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_5 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_5;

architecture SYN_behave of P_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_4 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_4;

architecture SYN_behave of P_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_3 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_3;

architecture SYN_behave of P_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_2 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_2;

architecture SYN_behave of P_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_1 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_1;

architecture SYN_behave of P_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_41 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_41;

architecture SYN_arch of PG_41 is

   component P_41
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_41
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_41 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_41 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_40 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_40;

architecture SYN_arch of PG_40 is

   component P_40
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_40
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_40 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_40 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_39 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_39;

architecture SYN_arch of PG_39 is

   component P_39
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_39
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_39 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_39 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_38 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_38;

architecture SYN_arch of PG_38 is

   component P_38
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_38
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_38 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_38 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_37 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_37;

architecture SYN_arch of PG_37 is

   component P_37
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_37
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_37 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_37 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_36 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_36;

architecture SYN_arch of PG_36 is

   component P_36
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_36
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_36 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_36 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_35 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_35;

architecture SYN_arch of PG_35 is

   component P_35
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_35
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_35 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_35 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_34 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_34;

architecture SYN_arch of PG_34 is

   component P_34
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_34
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_34 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_34 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_33 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_33;

architecture SYN_arch of PG_33 is

   component P_33
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_33
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_33 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_33 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_32 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_32;

architecture SYN_arch of PG_32 is

   component P_32
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_32
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_32 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_32 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_31 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_31;

architecture SYN_arch of PG_31 is

   component P_31
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_31
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_31 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_31 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_30 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_30;

architecture SYN_arch of PG_30 is

   component P_30
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_30
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_30 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_30 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_29 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_29;

architecture SYN_arch of PG_29 is

   component P_29
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_29
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_29 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_29 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_28 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_28;

architecture SYN_arch of PG_28 is

   component P_28
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_28
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_28 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_28 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_27 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_27;

architecture SYN_arch of PG_27 is

   component P_27
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_27
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_27 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_27 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_26 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_26;

architecture SYN_arch of PG_26 is

   component P_26
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_26
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_26 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_26 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_25 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_25;

architecture SYN_arch of PG_25 is

   component P_25
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_25
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_25 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_25 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_24 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_24;

architecture SYN_arch of PG_24 is

   component P_24
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_24
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_24 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_24 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_23 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_23;

architecture SYN_arch of PG_23 is

   component P_23
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_23
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_23 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_23 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_22 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_22;

architecture SYN_arch of PG_22 is

   component P_22
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_22
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_22 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_22 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_21 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_21;

architecture SYN_arch of PG_21 is

   component P_21
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_21
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_21 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_21 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_20 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_20;

architecture SYN_arch of PG_20 is

   component P_20
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_20
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_20 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_20 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_19 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_19;

architecture SYN_arch of PG_19 is

   component P_19
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_19
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_19 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_19 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_18 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_18;

architecture SYN_arch of PG_18 is

   component P_18
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_18
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_18 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_18 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_17 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_17;

architecture SYN_arch of PG_17 is

   component P_17
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_17
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_17 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_17 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_16 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_16;

architecture SYN_arch of PG_16 is

   component P_16
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_16
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_16 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_16 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_15 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_15;

architecture SYN_arch of PG_15 is

   component P_15
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_15
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_15 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_15 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_14 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_14;

architecture SYN_arch of PG_14 is

   component P_14
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_14
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_14 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_14 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_13 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_13;

architecture SYN_arch of PG_13 is

   component P_13
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_13
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_13 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_13 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_12 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_12;

architecture SYN_arch of PG_12 is

   component P_12
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_12
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_12 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_12 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_11 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_11;

architecture SYN_arch of PG_11 is

   component P_11
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_11
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_11 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_11 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_10 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_10;

architecture SYN_arch of PG_10 is

   component P_10
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_10
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_10 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_10 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_9 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_9;

architecture SYN_arch of PG_9 is

   component P_9
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_9
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_9 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_9 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_8 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_8;

architecture SYN_arch of PG_8 is

   component P_8
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_8
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_8 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_8 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_7 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_7;

architecture SYN_arch of PG_7 is

   component P_7
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_7
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_7 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_7 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_6 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_6;

architecture SYN_arch of PG_6 is

   component P_6
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_6
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_6 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_6 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_5 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_5;

architecture SYN_arch of PG_5 is

   component P_5
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_5
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_5 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_5 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_4 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_4;

architecture SYN_arch of PG_4 is

   component P_4
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_4
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_4 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_4 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_3 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_3;

architecture SYN_arch of PG_3 is

   component P_3
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_3
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_3 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_3 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_2 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_2;

architecture SYN_arch of PG_2 is

   component P_2
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_2
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_2 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_2 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_1 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_1;

architecture SYN_arch of PG_1 is

   component P_1
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_1
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_1 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_1 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_52 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_52;

architecture SYN_behave of G_52 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_51 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_51;

architecture SYN_behave of G_51 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_50 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_50;

architecture SYN_behave of G_50 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_49 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_49;

architecture SYN_behave of G_49 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_48 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_48;

architecture SYN_behave of G_48 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_47 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_47;

architecture SYN_behave of G_47 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_46 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_46;

architecture SYN_behave of G_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_45 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_45;

architecture SYN_behave of G_45 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_44 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_44;

architecture SYN_behave of G_44 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_43 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_43;

architecture SYN_behave of G_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_42 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_42;

architecture SYN_behave of G_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_41 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_41;

architecture SYN_behave of G_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_40 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_40;

architecture SYN_behave of G_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_39 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_39;

architecture SYN_behave of G_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_38 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_38;

architecture SYN_behave of G_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_37 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_37;

architecture SYN_behave of G_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_36 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_36;

architecture SYN_behave of G_36 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_35 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_35;

architecture SYN_behave of G_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_34 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_34;

architecture SYN_behave of G_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_33 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_33;

architecture SYN_behave of G_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_32 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_32;

architecture SYN_behave of G_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_31 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_31;

architecture SYN_behave of G_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_30 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_30;

architecture SYN_behave of G_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_29 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_29;

architecture SYN_behave of G_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_28 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_28;

architecture SYN_behave of G_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_27 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_27;

architecture SYN_behave of G_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_26 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_26;

architecture SYN_behave of G_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_25 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_25;

architecture SYN_behave of G_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_24 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_24;

architecture SYN_behave of G_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_23 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_23;

architecture SYN_behave of G_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_22 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_22;

architecture SYN_behave of G_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_21 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_21;

architecture SYN_behave of G_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_20 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_20;

architecture SYN_behave of G_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_19 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_19;

architecture SYN_behave of G_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_18 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_18;

architecture SYN_behave of G_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_17 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_17;

architecture SYN_behave of G_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_16 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_16;

architecture SYN_behave of G_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_15 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_15;

architecture SYN_behave of G_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_14 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_14;

architecture SYN_behave of G_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_13 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_13;

architecture SYN_behave of G_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_12 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_12;

architecture SYN_behave of G_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_11 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_11;

architecture SYN_behave of G_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_10 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_10;

architecture SYN_behave of G_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_9 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_9;

architecture SYN_behave of G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_8 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_8;

architecture SYN_behave of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_7 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_7;

architecture SYN_behave of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_6 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_6;

architecture SYN_behave of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_5 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_5;

architecture SYN_behave of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_4 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_4;

architecture SYN_behave of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_3 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_3;

architecture SYN_behave of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_2 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_2;

architecture SYN_behave of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_1 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_1;

architecture SYN_behave of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n4);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_571 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_571;

architecture SYN_ARCH2 of ND2_571 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_568 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_568;

architecture SYN_ARCH2 of ND2_568 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_565 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_565;

architecture SYN_ARCH2 of ND2_565 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_767 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_767;

architecture SYN_ARCH2 of ND2_767 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_766 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_766;

architecture SYN_ARCH2 of ND2_766 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_765 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_765;

architecture SYN_ARCH2 of ND2_765 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_764 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_764;

architecture SYN_ARCH2 of ND2_764 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_763 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_763;

architecture SYN_ARCH2 of ND2_763 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_762 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_762;

architecture SYN_ARCH2 of ND2_762 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_761 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_761;

architecture SYN_ARCH2 of ND2_761 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_760 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_760;

architecture SYN_ARCH2 of ND2_760 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_759 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_759;

architecture SYN_ARCH2 of ND2_759 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_758 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_758;

architecture SYN_ARCH2 of ND2_758 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_757 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_757;

architecture SYN_ARCH2 of ND2_757 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_756 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_756;

architecture SYN_ARCH2 of ND2_756 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_755 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_755;

architecture SYN_ARCH2 of ND2_755 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_754 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_754;

architecture SYN_ARCH2 of ND2_754 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_753 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_753;

architecture SYN_ARCH2 of ND2_753 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_752 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_752;

architecture SYN_ARCH2 of ND2_752 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_751 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_751;

architecture SYN_ARCH2 of ND2_751 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_750 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_750;

architecture SYN_ARCH2 of ND2_750 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_749 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_749;

architecture SYN_ARCH2 of ND2_749 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_748 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_748;

architecture SYN_ARCH2 of ND2_748 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_747 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_747;

architecture SYN_ARCH2 of ND2_747 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_746 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_746;

architecture SYN_ARCH2 of ND2_746 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_745 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_745;

architecture SYN_ARCH2 of ND2_745 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_744 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_744;

architecture SYN_ARCH2 of ND2_744 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_743 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_743;

architecture SYN_ARCH2 of ND2_743 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_742 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_742;

architecture SYN_ARCH2 of ND2_742 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_741 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_741;

architecture SYN_ARCH2 of ND2_741 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_740 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_740;

architecture SYN_ARCH2 of ND2_740 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_739 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_739;

architecture SYN_ARCH2 of ND2_739 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_738 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_738;

architecture SYN_ARCH2 of ND2_738 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_737 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_737;

architecture SYN_ARCH2 of ND2_737 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_736 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_736;

architecture SYN_ARCH2 of ND2_736 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_735 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_735;

architecture SYN_ARCH2 of ND2_735 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_734 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_734;

architecture SYN_ARCH2 of ND2_734 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_733 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_733;

architecture SYN_ARCH2 of ND2_733 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_732 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_732;

architecture SYN_ARCH2 of ND2_732 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_731 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_731;

architecture SYN_ARCH2 of ND2_731 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_730 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_730;

architecture SYN_ARCH2 of ND2_730 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_729 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_729;

architecture SYN_ARCH2 of ND2_729 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_728 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_728;

architecture SYN_ARCH2 of ND2_728 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_727 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_727;

architecture SYN_ARCH2 of ND2_727 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_726 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_726;

architecture SYN_ARCH2 of ND2_726 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_725 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_725;

architecture SYN_ARCH2 of ND2_725 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_724 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_724;

architecture SYN_ARCH2 of ND2_724 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_723 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_723;

architecture SYN_ARCH2 of ND2_723 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_722 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_722;

architecture SYN_ARCH2 of ND2_722 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_721 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_721;

architecture SYN_ARCH2 of ND2_721 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_720 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_720;

architecture SYN_ARCH2 of ND2_720 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_719 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_719;

architecture SYN_ARCH2 of ND2_719 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_718 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_718;

architecture SYN_ARCH2 of ND2_718 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_717 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_717;

architecture SYN_ARCH2 of ND2_717 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_716 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_716;

architecture SYN_ARCH2 of ND2_716 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_715 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_715;

architecture SYN_ARCH2 of ND2_715 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_714 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_714;

architecture SYN_ARCH2 of ND2_714 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_713 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_713;

architecture SYN_ARCH2 of ND2_713 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_712 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_712;

architecture SYN_ARCH2 of ND2_712 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_711 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_711;

architecture SYN_ARCH2 of ND2_711 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_710 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_710;

architecture SYN_ARCH2 of ND2_710 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_709 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_709;

architecture SYN_ARCH2 of ND2_709 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_708 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_708;

architecture SYN_ARCH2 of ND2_708 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_707 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_707;

architecture SYN_ARCH2 of ND2_707 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_706 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_706;

architecture SYN_ARCH2 of ND2_706 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_705 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_705;

architecture SYN_ARCH2 of ND2_705 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_704 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_704;

architecture SYN_ARCH2 of ND2_704 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_703 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_703;

architecture SYN_ARCH2 of ND2_703 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_702 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_702;

architecture SYN_ARCH2 of ND2_702 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_701 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_701;

architecture SYN_ARCH2 of ND2_701 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_700 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_700;

architecture SYN_ARCH2 of ND2_700 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_699 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_699;

architecture SYN_ARCH2 of ND2_699 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_698 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_698;

architecture SYN_ARCH2 of ND2_698 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_697 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_697;

architecture SYN_ARCH2 of ND2_697 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_696 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_696;

architecture SYN_ARCH2 of ND2_696 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_695 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_695;

architecture SYN_ARCH2 of ND2_695 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_694 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_694;

architecture SYN_ARCH2 of ND2_694 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_693 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_693;

architecture SYN_ARCH2 of ND2_693 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_692 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_692;

architecture SYN_ARCH2 of ND2_692 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_691 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_691;

architecture SYN_ARCH2 of ND2_691 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_690 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_690;

architecture SYN_ARCH2 of ND2_690 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_689 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_689;

architecture SYN_ARCH2 of ND2_689 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_688 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_688;

architecture SYN_ARCH2 of ND2_688 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_687 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_687;

architecture SYN_ARCH2 of ND2_687 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_686 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_686;

architecture SYN_ARCH2 of ND2_686 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_685 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_685;

architecture SYN_ARCH2 of ND2_685 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_684 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_684;

architecture SYN_ARCH2 of ND2_684 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_683 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_683;

architecture SYN_ARCH2 of ND2_683 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_682 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_682;

architecture SYN_ARCH2 of ND2_682 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_681 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_681;

architecture SYN_ARCH2 of ND2_681 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_680 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_680;

architecture SYN_ARCH2 of ND2_680 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_679 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_679;

architecture SYN_ARCH2 of ND2_679 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_678 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_678;

architecture SYN_ARCH2 of ND2_678 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_677 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_677;

architecture SYN_ARCH2 of ND2_677 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_676 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_676;

architecture SYN_ARCH2 of ND2_676 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_675 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_675;

architecture SYN_ARCH2 of ND2_675 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_674 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_674;

architecture SYN_ARCH2 of ND2_674 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_673 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_673;

architecture SYN_ARCH2 of ND2_673 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_672 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_672;

architecture SYN_ARCH2 of ND2_672 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_671 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_671;

architecture SYN_ARCH2 of ND2_671 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_670 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_670;

architecture SYN_ARCH2 of ND2_670 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_669 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_669;

architecture SYN_ARCH2 of ND2_669 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_668 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_668;

architecture SYN_ARCH2 of ND2_668 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_667 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_667;

architecture SYN_ARCH2 of ND2_667 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_666 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_666;

architecture SYN_ARCH2 of ND2_666 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_665 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_665;

architecture SYN_ARCH2 of ND2_665 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_664 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_664;

architecture SYN_ARCH2 of ND2_664 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_663 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_663;

architecture SYN_ARCH2 of ND2_663 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_662 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_662;

architecture SYN_ARCH2 of ND2_662 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_661 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_661;

architecture SYN_ARCH2 of ND2_661 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_660 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_660;

architecture SYN_ARCH2 of ND2_660 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_659 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_659;

architecture SYN_ARCH2 of ND2_659 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_658 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_658;

architecture SYN_ARCH2 of ND2_658 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_657 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_657;

architecture SYN_ARCH2 of ND2_657 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_656 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_656;

architecture SYN_ARCH2 of ND2_656 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_655 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_655;

architecture SYN_ARCH2 of ND2_655 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_654 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_654;

architecture SYN_ARCH2 of ND2_654 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_653 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_653;

architecture SYN_ARCH2 of ND2_653 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_652 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_652;

architecture SYN_ARCH2 of ND2_652 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_651 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_651;

architecture SYN_ARCH2 of ND2_651 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_650 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_650;

architecture SYN_ARCH2 of ND2_650 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_649 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_649;

architecture SYN_ARCH2 of ND2_649 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_648 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_648;

architecture SYN_ARCH2 of ND2_648 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_647 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_647;

architecture SYN_ARCH2 of ND2_647 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_646 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_646;

architecture SYN_ARCH2 of ND2_646 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_645 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_645;

architecture SYN_ARCH2 of ND2_645 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_644 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_644;

architecture SYN_ARCH2 of ND2_644 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_643 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_643;

architecture SYN_ARCH2 of ND2_643 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_642 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_642;

architecture SYN_ARCH2 of ND2_642 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_641 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_641;

architecture SYN_ARCH2 of ND2_641 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_640 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_640;

architecture SYN_ARCH2 of ND2_640 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_639 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_639;

architecture SYN_ARCH2 of ND2_639 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_638 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_638;

architecture SYN_ARCH2 of ND2_638 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_637 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_637;

architecture SYN_ARCH2 of ND2_637 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_636 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_636;

architecture SYN_ARCH2 of ND2_636 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_635 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_635;

architecture SYN_ARCH2 of ND2_635 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_634 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_634;

architecture SYN_ARCH2 of ND2_634 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_633 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_633;

architecture SYN_ARCH2 of ND2_633 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_632 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_632;

architecture SYN_ARCH2 of ND2_632 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_631 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_631;

architecture SYN_ARCH2 of ND2_631 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_630 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_630;

architecture SYN_ARCH2 of ND2_630 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_629 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_629;

architecture SYN_ARCH2 of ND2_629 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_628 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_628;

architecture SYN_ARCH2 of ND2_628 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_627 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_627;

architecture SYN_ARCH2 of ND2_627 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_626 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_626;

architecture SYN_ARCH2 of ND2_626 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_625 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_625;

architecture SYN_ARCH2 of ND2_625 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_624 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_624;

architecture SYN_ARCH2 of ND2_624 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_623 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_623;

architecture SYN_ARCH2 of ND2_623 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_622 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_622;

architecture SYN_ARCH2 of ND2_622 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_621 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_621;

architecture SYN_ARCH2 of ND2_621 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_620 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_620;

architecture SYN_ARCH2 of ND2_620 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_619 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_619;

architecture SYN_ARCH2 of ND2_619 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_618 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_618;

architecture SYN_ARCH2 of ND2_618 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_617 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_617;

architecture SYN_ARCH2 of ND2_617 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_616 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_616;

architecture SYN_ARCH2 of ND2_616 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_615 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_615;

architecture SYN_ARCH2 of ND2_615 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_614 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_614;

architecture SYN_ARCH2 of ND2_614 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_613 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_613;

architecture SYN_ARCH2 of ND2_613 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_612 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_612;

architecture SYN_ARCH2 of ND2_612 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_611 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_611;

architecture SYN_ARCH2 of ND2_611 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_610 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_610;

architecture SYN_ARCH2 of ND2_610 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_609 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_609;

architecture SYN_ARCH2 of ND2_609 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_608 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_608;

architecture SYN_ARCH2 of ND2_608 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_607 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_607;

architecture SYN_ARCH2 of ND2_607 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_606 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_606;

architecture SYN_ARCH2 of ND2_606 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_605 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_605;

architecture SYN_ARCH2 of ND2_605 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_604 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_604;

architecture SYN_ARCH2 of ND2_604 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_603 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_603;

architecture SYN_ARCH2 of ND2_603 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_602 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_602;

architecture SYN_ARCH2 of ND2_602 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_601 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_601;

architecture SYN_ARCH2 of ND2_601 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_600 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_600;

architecture SYN_ARCH2 of ND2_600 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_599 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_599;

architecture SYN_ARCH2 of ND2_599 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_598 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_598;

architecture SYN_ARCH2 of ND2_598 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_597 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_597;

architecture SYN_ARCH2 of ND2_597 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_596 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_596;

architecture SYN_ARCH2 of ND2_596 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_595 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_595;

architecture SYN_ARCH2 of ND2_595 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_594 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_594;

architecture SYN_ARCH2 of ND2_594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_593 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_593;

architecture SYN_ARCH2 of ND2_593 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_592 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_592;

architecture SYN_ARCH2 of ND2_592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_591 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_591;

architecture SYN_ARCH2 of ND2_591 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_590 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_590;

architecture SYN_ARCH2 of ND2_590 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_589 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_589;

architecture SYN_ARCH2 of ND2_589 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_588 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_588;

architecture SYN_ARCH2 of ND2_588 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_587 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_587;

architecture SYN_ARCH2 of ND2_587 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_586 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_586;

architecture SYN_ARCH2 of ND2_586 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_585 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_585;

architecture SYN_ARCH2 of ND2_585 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_584 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_584;

architecture SYN_ARCH2 of ND2_584 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_583 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_583;

architecture SYN_ARCH2 of ND2_583 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_582 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_582;

architecture SYN_ARCH2 of ND2_582 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_581 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_581;

architecture SYN_ARCH2 of ND2_581 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_580 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_580;

architecture SYN_ARCH2 of ND2_580 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_579 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_579;

architecture SYN_ARCH2 of ND2_579 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_578 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_578;

architecture SYN_ARCH2 of ND2_578 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_577 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_577;

architecture SYN_ARCH2 of ND2_577 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_576 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_576;

architecture SYN_ARCH2 of ND2_576 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_575 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_575;

architecture SYN_ARCH2 of ND2_575 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_573 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_573;

architecture SYN_ARCH2 of ND2_573 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_572 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_572;

architecture SYN_ARCH2 of ND2_572 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_570 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_570;

architecture SYN_ARCH2 of ND2_570 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_569 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_569;

architecture SYN_ARCH2 of ND2_569 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_567 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_567;

architecture SYN_ARCH2 of ND2_567 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_566 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_566;

architecture SYN_ARCH2 of ND2_566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_564 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_564;

architecture SYN_ARCH2 of ND2_564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_563 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_563;

architecture SYN_ARCH2 of ND2_563 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_562 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_562;

architecture SYN_ARCH2 of ND2_562 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_561 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_561;

architecture SYN_ARCH2 of ND2_561 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_560 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_560;

architecture SYN_ARCH2 of ND2_560 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_559 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_559;

architecture SYN_ARCH2 of ND2_559 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_558 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_558;

architecture SYN_ARCH2 of ND2_558 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_557 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_557;

architecture SYN_ARCH2 of ND2_557 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_556 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_556;

architecture SYN_ARCH2 of ND2_556 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_555 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_555;

architecture SYN_ARCH2 of ND2_555 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_554 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_554;

architecture SYN_ARCH2 of ND2_554 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_553 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_553;

architecture SYN_ARCH2 of ND2_553 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_552 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_552;

architecture SYN_ARCH2 of ND2_552 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_551 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_551;

architecture SYN_ARCH2 of ND2_551 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_550 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_550;

architecture SYN_ARCH2 of ND2_550 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_549 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_549;

architecture SYN_ARCH2 of ND2_549 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_548 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_548;

architecture SYN_ARCH2 of ND2_548 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_547 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_547;

architecture SYN_ARCH2 of ND2_547 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_546 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_546;

architecture SYN_ARCH2 of ND2_546 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_545 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_545;

architecture SYN_ARCH2 of ND2_545 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_544 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_544;

architecture SYN_ARCH2 of ND2_544 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_543 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_543;

architecture SYN_ARCH2 of ND2_543 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_542 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_542;

architecture SYN_ARCH2 of ND2_542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_541 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_541;

architecture SYN_ARCH2 of ND2_541 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_540 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_540;

architecture SYN_ARCH2 of ND2_540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_539 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_539;

architecture SYN_ARCH2 of ND2_539 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_538 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_538;

architecture SYN_ARCH2 of ND2_538 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_537 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_537;

architecture SYN_ARCH2 of ND2_537 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_536 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_536;

architecture SYN_ARCH2 of ND2_536 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_535 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_535;

architecture SYN_ARCH2 of ND2_535 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_534 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_534;

architecture SYN_ARCH2 of ND2_534 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_533 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_533;

architecture SYN_ARCH2 of ND2_533 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_532 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_532;

architecture SYN_ARCH2 of ND2_532 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_531 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_531;

architecture SYN_ARCH2 of ND2_531 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_530 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_530;

architecture SYN_ARCH2 of ND2_530 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_529 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_529;

architecture SYN_ARCH2 of ND2_529 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_528 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_528;

architecture SYN_ARCH2 of ND2_528 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_527 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_527;

architecture SYN_ARCH2 of ND2_527 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_526 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_526;

architecture SYN_ARCH2 of ND2_526 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_525 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_525;

architecture SYN_ARCH2 of ND2_525 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_524 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_524;

architecture SYN_ARCH2 of ND2_524 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_523 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_523;

architecture SYN_ARCH2 of ND2_523 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_522 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_522;

architecture SYN_ARCH2 of ND2_522 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_521 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_521;

architecture SYN_ARCH2 of ND2_521 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_520 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_520;

architecture SYN_ARCH2 of ND2_520 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_519 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_519;

architecture SYN_ARCH2 of ND2_519 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_518 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_518;

architecture SYN_ARCH2 of ND2_518 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_517 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_517;

architecture SYN_ARCH2 of ND2_517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_516 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_516;

architecture SYN_ARCH2 of ND2_516 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_515 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_515;

architecture SYN_ARCH2 of ND2_515 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_514 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_514;

architecture SYN_ARCH2 of ND2_514 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_513 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_513;

architecture SYN_ARCH2 of ND2_513 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_512 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_512;

architecture SYN_ARCH2 of ND2_512 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_511 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_511;

architecture SYN_ARCH2 of ND2_511 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_510 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_510;

architecture SYN_ARCH2 of ND2_510 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_509 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_509;

architecture SYN_ARCH2 of ND2_509 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_508 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_508;

architecture SYN_ARCH2 of ND2_508 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_507 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_507;

architecture SYN_ARCH2 of ND2_507 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_506 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_506;

architecture SYN_ARCH2 of ND2_506 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_505 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_505;

architecture SYN_ARCH2 of ND2_505 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_504 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_504;

architecture SYN_ARCH2 of ND2_504 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_503 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_503;

architecture SYN_ARCH2 of ND2_503 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_502 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_502;

architecture SYN_ARCH2 of ND2_502 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_501 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_501;

architecture SYN_ARCH2 of ND2_501 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_500 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_500;

architecture SYN_ARCH2 of ND2_500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_499 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_499;

architecture SYN_ARCH2 of ND2_499 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_498 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_498;

architecture SYN_ARCH2 of ND2_498 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_497 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_497;

architecture SYN_ARCH2 of ND2_497 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_496 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_496;

architecture SYN_ARCH2 of ND2_496 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_495 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_495;

architecture SYN_ARCH2 of ND2_495 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_494 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_494;

architecture SYN_ARCH2 of ND2_494 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_493 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_493;

architecture SYN_ARCH2 of ND2_493 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_492 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_492;

architecture SYN_ARCH2 of ND2_492 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_491 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_491;

architecture SYN_ARCH2 of ND2_491 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_490 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_490;

architecture SYN_ARCH2 of ND2_490 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_489 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_489;

architecture SYN_ARCH2 of ND2_489 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_488 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_488;

architecture SYN_ARCH2 of ND2_488 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_487 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_487;

architecture SYN_ARCH2 of ND2_487 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_486 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_486;

architecture SYN_ARCH2 of ND2_486 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_485 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_485;

architecture SYN_ARCH2 of ND2_485 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_484 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_484;

architecture SYN_ARCH2 of ND2_484 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_483 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_483;

architecture SYN_ARCH2 of ND2_483 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_482 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_482;

architecture SYN_ARCH2 of ND2_482 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_481 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_481;

architecture SYN_ARCH2 of ND2_481 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_480 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_480;

architecture SYN_ARCH2 of ND2_480 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_479 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_479;

architecture SYN_ARCH2 of ND2_479 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_478 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_478;

architecture SYN_ARCH2 of ND2_478 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_477 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_477;

architecture SYN_ARCH2 of ND2_477 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_476 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_476;

architecture SYN_ARCH2 of ND2_476 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_475 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_475;

architecture SYN_ARCH2 of ND2_475 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_474 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_474;

architecture SYN_ARCH2 of ND2_474 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_473 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_473;

architecture SYN_ARCH2 of ND2_473 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_472 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_472;

architecture SYN_ARCH2 of ND2_472 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_471 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_471;

architecture SYN_ARCH2 of ND2_471 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_470 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_470;

architecture SYN_ARCH2 of ND2_470 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_469 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_469;

architecture SYN_ARCH2 of ND2_469 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_468 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_468;

architecture SYN_ARCH2 of ND2_468 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_467 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_467;

architecture SYN_ARCH2 of ND2_467 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_466 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_466;

architecture SYN_ARCH2 of ND2_466 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_465 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_465;

architecture SYN_ARCH2 of ND2_465 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_464 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_464;

architecture SYN_ARCH2 of ND2_464 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_463 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_463;

architecture SYN_ARCH2 of ND2_463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_462 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_462;

architecture SYN_ARCH2 of ND2_462 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_461 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_461;

architecture SYN_ARCH2 of ND2_461 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_460 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_460;

architecture SYN_ARCH2 of ND2_460 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_459 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_459;

architecture SYN_ARCH2 of ND2_459 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_458 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_458;

architecture SYN_ARCH2 of ND2_458 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_457 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_457;

architecture SYN_ARCH2 of ND2_457 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_456 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_456;

architecture SYN_ARCH2 of ND2_456 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_455 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_455;

architecture SYN_ARCH2 of ND2_455 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_454 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_454;

architecture SYN_ARCH2 of ND2_454 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_453 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_453;

architecture SYN_ARCH2 of ND2_453 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_452 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_452;

architecture SYN_ARCH2 of ND2_452 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_451 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_451;

architecture SYN_ARCH2 of ND2_451 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_450 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_450;

architecture SYN_ARCH2 of ND2_450 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_449 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_449;

architecture SYN_ARCH2 of ND2_449 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_448 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_448;

architecture SYN_ARCH2 of ND2_448 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_447 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_447;

architecture SYN_ARCH2 of ND2_447 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_446 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_446;

architecture SYN_ARCH2 of ND2_446 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_445 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_445;

architecture SYN_ARCH2 of ND2_445 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_444 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_444;

architecture SYN_ARCH2 of ND2_444 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_443 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_443;

architecture SYN_ARCH2 of ND2_443 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_442 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_442;

architecture SYN_ARCH2 of ND2_442 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_441 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_441;

architecture SYN_ARCH2 of ND2_441 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_440 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_440;

architecture SYN_ARCH2 of ND2_440 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_439 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_439;

architecture SYN_ARCH2 of ND2_439 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_438 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_438;

architecture SYN_ARCH2 of ND2_438 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_437 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_437;

architecture SYN_ARCH2 of ND2_437 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_436 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_436;

architecture SYN_ARCH2 of ND2_436 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_435 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_435;

architecture SYN_ARCH2 of ND2_435 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_434 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_434;

architecture SYN_ARCH2 of ND2_434 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_433 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_433;

architecture SYN_ARCH2 of ND2_433 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_432 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_432;

architecture SYN_ARCH2 of ND2_432 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_431 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_431;

architecture SYN_ARCH2 of ND2_431 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_430 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_430;

architecture SYN_ARCH2 of ND2_430 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_429 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_429;

architecture SYN_ARCH2 of ND2_429 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_428 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_428;

architecture SYN_ARCH2 of ND2_428 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_427 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_427;

architecture SYN_ARCH2 of ND2_427 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_426 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_426;

architecture SYN_ARCH2 of ND2_426 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_425 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_425;

architecture SYN_ARCH2 of ND2_425 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_424 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_424;

architecture SYN_ARCH2 of ND2_424 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_423 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_423;

architecture SYN_ARCH2 of ND2_423 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_422 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_422;

architecture SYN_ARCH2 of ND2_422 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_421 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_421;

architecture SYN_ARCH2 of ND2_421 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_420 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_420;

architecture SYN_ARCH2 of ND2_420 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_419 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_419;

architecture SYN_ARCH2 of ND2_419 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_418 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_418;

architecture SYN_ARCH2 of ND2_418 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_417 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_417;

architecture SYN_ARCH2 of ND2_417 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_416 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_416;

architecture SYN_ARCH2 of ND2_416 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_415 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_415;

architecture SYN_ARCH2 of ND2_415 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_414 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_414;

architecture SYN_ARCH2 of ND2_414 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_413 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_413;

architecture SYN_ARCH2 of ND2_413 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_412 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_412;

architecture SYN_ARCH2 of ND2_412 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_411 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_411;

architecture SYN_ARCH2 of ND2_411 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_410 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_410;

architecture SYN_ARCH2 of ND2_410 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_409 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_409;

architecture SYN_ARCH2 of ND2_409 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_408 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_408;

architecture SYN_ARCH2 of ND2_408 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_407 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_407;

architecture SYN_ARCH2 of ND2_407 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_406 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_406;

architecture SYN_ARCH2 of ND2_406 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_405 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_405;

architecture SYN_ARCH2 of ND2_405 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_404 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_404;

architecture SYN_ARCH2 of ND2_404 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_403 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_403;

architecture SYN_ARCH2 of ND2_403 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_402 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_402;

architecture SYN_ARCH2 of ND2_402 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_401 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_401;

architecture SYN_ARCH2 of ND2_401 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_400 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_400;

architecture SYN_ARCH2 of ND2_400 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_399 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_399;

architecture SYN_ARCH2 of ND2_399 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_398 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_398;

architecture SYN_ARCH2 of ND2_398 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_397 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_397;

architecture SYN_ARCH2 of ND2_397 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_396 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_396;

architecture SYN_ARCH2 of ND2_396 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_395 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_395;

architecture SYN_ARCH2 of ND2_395 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_394 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_394;

architecture SYN_ARCH2 of ND2_394 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_393 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_393;

architecture SYN_ARCH2 of ND2_393 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_392 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_392;

architecture SYN_ARCH2 of ND2_392 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_391 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_391;

architecture SYN_ARCH2 of ND2_391 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_390 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_390;

architecture SYN_ARCH2 of ND2_390 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_389 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_389;

architecture SYN_ARCH2 of ND2_389 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_388 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_388;

architecture SYN_ARCH2 of ND2_388 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_387 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_387;

architecture SYN_ARCH2 of ND2_387 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_386 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_386;

architecture SYN_ARCH2 of ND2_386 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_385 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_385;

architecture SYN_ARCH2 of ND2_385 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_384 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_384;

architecture SYN_ARCH2 of ND2_384 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_383 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_383;

architecture SYN_ARCH2 of ND2_383 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_382 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_382;

architecture SYN_ARCH2 of ND2_382 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_381 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_381;

architecture SYN_ARCH2 of ND2_381 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_380 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_380;

architecture SYN_ARCH2 of ND2_380 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_379 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_379;

architecture SYN_ARCH2 of ND2_379 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_378 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_378;

architecture SYN_ARCH2 of ND2_378 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_377 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_377;

architecture SYN_ARCH2 of ND2_377 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_376 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_376;

architecture SYN_ARCH2 of ND2_376 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_375 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_375;

architecture SYN_ARCH2 of ND2_375 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_374 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_374;

architecture SYN_ARCH2 of ND2_374 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_373 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_373;

architecture SYN_ARCH2 of ND2_373 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_372 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_372;

architecture SYN_ARCH2 of ND2_372 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_371 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_371;

architecture SYN_ARCH2 of ND2_371 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_370 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_370;

architecture SYN_ARCH2 of ND2_370 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_369 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_369;

architecture SYN_ARCH2 of ND2_369 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_368 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_368;

architecture SYN_ARCH2 of ND2_368 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_367 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_367;

architecture SYN_ARCH2 of ND2_367 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_366 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_366;

architecture SYN_ARCH2 of ND2_366 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_365 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_365;

architecture SYN_ARCH2 of ND2_365 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_364 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_364;

architecture SYN_ARCH2 of ND2_364 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_363 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_363;

architecture SYN_ARCH2 of ND2_363 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_362 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_362;

architecture SYN_ARCH2 of ND2_362 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_361 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_361;

architecture SYN_ARCH2 of ND2_361 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_360 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_360;

architecture SYN_ARCH2 of ND2_360 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_359 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_359;

architecture SYN_ARCH2 of ND2_359 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_358 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_358;

architecture SYN_ARCH2 of ND2_358 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_357 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_357;

architecture SYN_ARCH2 of ND2_357 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_356 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_356;

architecture SYN_ARCH2 of ND2_356 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_355 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_355;

architecture SYN_ARCH2 of ND2_355 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_354 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_354;

architecture SYN_ARCH2 of ND2_354 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_353 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_353;

architecture SYN_ARCH2 of ND2_353 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_352 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_352;

architecture SYN_ARCH2 of ND2_352 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_351 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_351;

architecture SYN_ARCH2 of ND2_351 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_350 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_350;

architecture SYN_ARCH2 of ND2_350 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_349 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_349;

architecture SYN_ARCH2 of ND2_349 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_348 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_348;

architecture SYN_ARCH2 of ND2_348 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_347 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_347;

architecture SYN_ARCH2 of ND2_347 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_346 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_346;

architecture SYN_ARCH2 of ND2_346 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_345 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_345;

architecture SYN_ARCH2 of ND2_345 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_344 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_344;

architecture SYN_ARCH2 of ND2_344 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_343 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_343;

architecture SYN_ARCH2 of ND2_343 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_342 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_342;

architecture SYN_ARCH2 of ND2_342 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_341 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_341;

architecture SYN_ARCH2 of ND2_341 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_340 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_340;

architecture SYN_ARCH2 of ND2_340 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_339 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_339;

architecture SYN_ARCH2 of ND2_339 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_338 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_338;

architecture SYN_ARCH2 of ND2_338 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_337 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_337;

architecture SYN_ARCH2 of ND2_337 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_336 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_336;

architecture SYN_ARCH2 of ND2_336 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_335 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_335;

architecture SYN_ARCH2 of ND2_335 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_334 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_334;

architecture SYN_ARCH2 of ND2_334 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_333 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_333;

architecture SYN_ARCH2 of ND2_333 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_332 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_332;

architecture SYN_ARCH2 of ND2_332 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_331 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_331;

architecture SYN_ARCH2 of ND2_331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_330 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_330;

architecture SYN_ARCH2 of ND2_330 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_329 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_329;

architecture SYN_ARCH2 of ND2_329 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_328 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_328;

architecture SYN_ARCH2 of ND2_328 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_327 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_327;

architecture SYN_ARCH2 of ND2_327 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_326 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_326;

architecture SYN_ARCH2 of ND2_326 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_325 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_325;

architecture SYN_ARCH2 of ND2_325 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_324 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_324;

architecture SYN_ARCH2 of ND2_324 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_323 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_323;

architecture SYN_ARCH2 of ND2_323 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_322 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_322;

architecture SYN_ARCH2 of ND2_322 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_321 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_321;

architecture SYN_ARCH2 of ND2_321 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_320 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_320;

architecture SYN_ARCH2 of ND2_320 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_319 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_319;

architecture SYN_ARCH2 of ND2_319 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_318 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_318;

architecture SYN_ARCH2 of ND2_318 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_317 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_317;

architecture SYN_ARCH2 of ND2_317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_316 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_316;

architecture SYN_ARCH2 of ND2_316 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_315 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_315;

architecture SYN_ARCH2 of ND2_315 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_314 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_314;

architecture SYN_ARCH2 of ND2_314 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_313 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_313;

architecture SYN_ARCH2 of ND2_313 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_312 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_312;

architecture SYN_ARCH2 of ND2_312 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_311 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_311;

architecture SYN_ARCH2 of ND2_311 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_310 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_310;

architecture SYN_ARCH2 of ND2_310 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_309 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_309;

architecture SYN_ARCH2 of ND2_309 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_308 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_308;

architecture SYN_ARCH2 of ND2_308 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_307 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_307;

architecture SYN_ARCH2 of ND2_307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_306 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_306;

architecture SYN_ARCH2 of ND2_306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_305 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_305;

architecture SYN_ARCH2 of ND2_305 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_304 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_304;

architecture SYN_ARCH2 of ND2_304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_303 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_303;

architecture SYN_ARCH2 of ND2_303 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_302 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_302;

architecture SYN_ARCH2 of ND2_302 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_301 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_301;

architecture SYN_ARCH2 of ND2_301 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_300 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_300;

architecture SYN_ARCH2 of ND2_300 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_299 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_299;

architecture SYN_ARCH2 of ND2_299 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_298 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_298;

architecture SYN_ARCH2 of ND2_298 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_297 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_297;

architecture SYN_ARCH2 of ND2_297 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_296 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_296;

architecture SYN_ARCH2 of ND2_296 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_295 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_295;

architecture SYN_ARCH2 of ND2_295 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_294 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_294;

architecture SYN_ARCH2 of ND2_294 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_293 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_293;

architecture SYN_ARCH2 of ND2_293 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_292 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_292;

architecture SYN_ARCH2 of ND2_292 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_291 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_291;

architecture SYN_ARCH2 of ND2_291 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_290 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_290;

architecture SYN_ARCH2 of ND2_290 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_289 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_289;

architecture SYN_ARCH2 of ND2_289 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_288 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_288;

architecture SYN_ARCH2 of ND2_288 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_287 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_287;

architecture SYN_ARCH2 of ND2_287 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_286 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_286;

architecture SYN_ARCH2 of ND2_286 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_285 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_285;

architecture SYN_ARCH2 of ND2_285 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_284 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_284;

architecture SYN_ARCH2 of ND2_284 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_283 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_283;

architecture SYN_ARCH2 of ND2_283 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_282 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_282;

architecture SYN_ARCH2 of ND2_282 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_281 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_281;

architecture SYN_ARCH2 of ND2_281 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_280 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_280;

architecture SYN_ARCH2 of ND2_280 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_279 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_279;

architecture SYN_ARCH2 of ND2_279 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_278 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_278;

architecture SYN_ARCH2 of ND2_278 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_277 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_277;

architecture SYN_ARCH2 of ND2_277 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_276 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_276;

architecture SYN_ARCH2 of ND2_276 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_275 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_275;

architecture SYN_ARCH2 of ND2_275 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_274 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_274;

architecture SYN_ARCH2 of ND2_274 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_273 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_273;

architecture SYN_ARCH2 of ND2_273 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_272 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_272;

architecture SYN_ARCH2 of ND2_272 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_271 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_271;

architecture SYN_ARCH2 of ND2_271 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_270 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_270;

architecture SYN_ARCH2 of ND2_270 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_269 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_269;

architecture SYN_ARCH2 of ND2_269 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_268 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_268;

architecture SYN_ARCH2 of ND2_268 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_267 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_267;

architecture SYN_ARCH2 of ND2_267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_266 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_266;

architecture SYN_ARCH2 of ND2_266 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_265 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_265;

architecture SYN_ARCH2 of ND2_265 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_264 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_264;

architecture SYN_ARCH2 of ND2_264 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_263 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_263;

architecture SYN_ARCH2 of ND2_263 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_262 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_262;

architecture SYN_ARCH2 of ND2_262 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_261 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_261;

architecture SYN_ARCH2 of ND2_261 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_260 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_260;

architecture SYN_ARCH2 of ND2_260 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_259 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_259;

architecture SYN_ARCH2 of ND2_259 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_258 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_258;

architecture SYN_ARCH2 of ND2_258 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_257 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_257;

architecture SYN_ARCH2 of ND2_257 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_256 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_256;

architecture SYN_ARCH2 of ND2_256 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_255 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_255;

architecture SYN_ARCH2 of ND2_255 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_254 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_254;

architecture SYN_ARCH2 of ND2_254 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_253 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_253;

architecture SYN_ARCH2 of ND2_253 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_252 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_252;

architecture SYN_ARCH2 of ND2_252 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_251 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_251;

architecture SYN_ARCH2 of ND2_251 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_250 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_250;

architecture SYN_ARCH2 of ND2_250 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_249 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_249;

architecture SYN_ARCH2 of ND2_249 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_248 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_248;

architecture SYN_ARCH2 of ND2_248 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_247 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_247;

architecture SYN_ARCH2 of ND2_247 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_246 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_246;

architecture SYN_ARCH2 of ND2_246 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_245 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_245;

architecture SYN_ARCH2 of ND2_245 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_244 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_244;

architecture SYN_ARCH2 of ND2_244 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_243 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_243;

architecture SYN_ARCH2 of ND2_243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_242 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_242;

architecture SYN_ARCH2 of ND2_242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_241 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_241;

architecture SYN_ARCH2 of ND2_241 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_240 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_240;

architecture SYN_ARCH2 of ND2_240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_239 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_239;

architecture SYN_ARCH2 of ND2_239 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_238 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_238;

architecture SYN_ARCH2 of ND2_238 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_237 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_237;

architecture SYN_ARCH2 of ND2_237 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_236 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_236;

architecture SYN_ARCH2 of ND2_236 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_235 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_235;

architecture SYN_ARCH2 of ND2_235 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_234 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_234;

architecture SYN_ARCH2 of ND2_234 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_233 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_233;

architecture SYN_ARCH2 of ND2_233 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_232 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_232;

architecture SYN_ARCH2 of ND2_232 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_231 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_231;

architecture SYN_ARCH2 of ND2_231 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_230 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_230;

architecture SYN_ARCH2 of ND2_230 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_229 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_229;

architecture SYN_ARCH2 of ND2_229 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_228 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_228;

architecture SYN_ARCH2 of ND2_228 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_227 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_227;

architecture SYN_ARCH2 of ND2_227 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_226 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_226;

architecture SYN_ARCH2 of ND2_226 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_225 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_225;

architecture SYN_ARCH2 of ND2_225 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_224 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_224;

architecture SYN_ARCH2 of ND2_224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_223 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_223;

architecture SYN_ARCH2 of ND2_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_222 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_222;

architecture SYN_ARCH2 of ND2_222 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_221 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_221;

architecture SYN_ARCH2 of ND2_221 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_220 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_220;

architecture SYN_ARCH2 of ND2_220 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_219 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_219;

architecture SYN_ARCH2 of ND2_219 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_218 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_218;

architecture SYN_ARCH2 of ND2_218 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_217 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_217;

architecture SYN_ARCH2 of ND2_217 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_216 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_216;

architecture SYN_ARCH2 of ND2_216 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_215 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_215;

architecture SYN_ARCH2 of ND2_215 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_214 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_214;

architecture SYN_ARCH2 of ND2_214 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_213 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_213;

architecture SYN_ARCH2 of ND2_213 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_212 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_212;

architecture SYN_ARCH2 of ND2_212 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_211 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_211;

architecture SYN_ARCH2 of ND2_211 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_210 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_210;

architecture SYN_ARCH2 of ND2_210 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_209 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_209;

architecture SYN_ARCH2 of ND2_209 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_208 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_208;

architecture SYN_ARCH2 of ND2_208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_207 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_207;

architecture SYN_ARCH2 of ND2_207 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_206 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_206;

architecture SYN_ARCH2 of ND2_206 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_205 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_205;

architecture SYN_ARCH2 of ND2_205 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_204 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_204;

architecture SYN_ARCH2 of ND2_204 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_203 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_203;

architecture SYN_ARCH2 of ND2_203 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_202 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_202;

architecture SYN_ARCH2 of ND2_202 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_201 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_201;

architecture SYN_ARCH2 of ND2_201 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_200 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_200;

architecture SYN_ARCH2 of ND2_200 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_199 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_199;

architecture SYN_ARCH2 of ND2_199 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_198 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_198;

architecture SYN_ARCH2 of ND2_198 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_197 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_197;

architecture SYN_ARCH2 of ND2_197 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_196 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_196;

architecture SYN_ARCH2 of ND2_196 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_195 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_195;

architecture SYN_ARCH2 of ND2_195 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_194 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_194;

architecture SYN_ARCH2 of ND2_194 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_193 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_193;

architecture SYN_ARCH2 of ND2_193 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_192 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_192;

architecture SYN_ARCH2 of ND2_192 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_191;

architecture SYN_ARCH2 of ND2_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_189;

architecture SYN_ARCH2 of ND2_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_188;

architecture SYN_ARCH2 of ND2_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_186;

architecture SYN_ARCH2 of ND2_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_185;

architecture SYN_ARCH2 of ND2_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_183;

architecture SYN_ARCH2 of ND2_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_182;

architecture SYN_ARCH2 of ND2_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_180;

architecture SYN_ARCH2 of ND2_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_179;

architecture SYN_ARCH2 of ND2_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_177;

architecture SYN_ARCH2 of ND2_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_176;

architecture SYN_ARCH2 of ND2_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_174;

architecture SYN_ARCH2 of ND2_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_173;

architecture SYN_ARCH2 of ND2_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_171;

architecture SYN_ARCH2 of ND2_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_170;

architecture SYN_ARCH2 of ND2_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_168;

architecture SYN_ARCH2 of ND2_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_167;

architecture SYN_ARCH2 of ND2_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_165;

architecture SYN_ARCH2 of ND2_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_164;

architecture SYN_ARCH2 of ND2_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_162;

architecture SYN_ARCH2 of ND2_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_161;

architecture SYN_ARCH2 of ND2_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_159;

architecture SYN_ARCH2 of ND2_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_158;

architecture SYN_ARCH2 of ND2_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_156;

architecture SYN_ARCH2 of ND2_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_155;

architecture SYN_ARCH2 of ND2_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_153;

architecture SYN_ARCH2 of ND2_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_152;

architecture SYN_ARCH2 of ND2_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_150;

architecture SYN_ARCH2 of ND2_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_149;

architecture SYN_ARCH2 of ND2_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_147;

architecture SYN_ARCH2 of ND2_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_146;

architecture SYN_ARCH2 of ND2_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_144;

architecture SYN_ARCH2 of ND2_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_143;

architecture SYN_ARCH2 of ND2_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_141;

architecture SYN_ARCH2 of ND2_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_140;

architecture SYN_ARCH2 of ND2_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_138;

architecture SYN_ARCH2 of ND2_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_137;

architecture SYN_ARCH2 of ND2_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_135;

architecture SYN_ARCH2 of ND2_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_134;

architecture SYN_ARCH2 of ND2_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_132;

architecture SYN_ARCH2 of ND2_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_131;

architecture SYN_ARCH2 of ND2_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_129;

architecture SYN_ARCH2 of ND2_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_128;

architecture SYN_ARCH2 of ND2_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_126;

architecture SYN_ARCH2 of ND2_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_125;

architecture SYN_ARCH2 of ND2_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_123;

architecture SYN_ARCH2 of ND2_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_122;

architecture SYN_ARCH2 of ND2_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_120;

architecture SYN_ARCH2 of ND2_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_119;

architecture SYN_ARCH2 of ND2_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_117;

architecture SYN_ARCH2 of ND2_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_116;

architecture SYN_ARCH2 of ND2_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_114;

architecture SYN_ARCH2 of ND2_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_113;

architecture SYN_ARCH2 of ND2_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_111;

architecture SYN_ARCH2 of ND2_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_110;

architecture SYN_ARCH2 of ND2_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_108;

architecture SYN_ARCH2 of ND2_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_107;

architecture SYN_ARCH2 of ND2_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_105;

architecture SYN_ARCH2 of ND2_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_104;

architecture SYN_ARCH2 of ND2_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_102;

architecture SYN_ARCH2 of ND2_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_101;

architecture SYN_ARCH2 of ND2_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_99;

architecture SYN_ARCH2 of ND2_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_98;

architecture SYN_ARCH2 of ND2_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_96;

architecture SYN_ARCH2 of ND2_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95;

architecture SYN_ARCH2 of ND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94;

architecture SYN_ARCH2 of ND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH2 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH2 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH2 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH2 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH2 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH2 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH2 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH2 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH2 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH2 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH2 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH2 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH2 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH2 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH2 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH2 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH2 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH2 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH2 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH2 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH2 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH2 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH2 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH2 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH2 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH2 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH2 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH2 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH2 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH2 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH2 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH2 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH2 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH2 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH2 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH2 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH2 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH2 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH2 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH2 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH2 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH2 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH2 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH2 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH2 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH2 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH2 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH2 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH2 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH2 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH2 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH2 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH2 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH2 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH2 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH2 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH2 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH2 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH2 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH2 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH2 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH2 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH2 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH2 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH2 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH2 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH2 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH2 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH2 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH2 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH2 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH2 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH2 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH2 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH2 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH2 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH2 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH2 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH2 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH2 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH2 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH2 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH2 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH2 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH2 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH2 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH2 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH2 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH2 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH2 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH2 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH2 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH2 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_187;

architecture SYN_ARCH2 of ND2_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_184;

architecture SYN_ARCH2 of ND2_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_181;

architecture SYN_ARCH2 of ND2_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_178;

architecture SYN_ARCH2 of ND2_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_175;

architecture SYN_ARCH2 of ND2_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_172;

architecture SYN_ARCH2 of ND2_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_169;

architecture SYN_ARCH2 of ND2_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_166;

architecture SYN_ARCH2 of ND2_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_163;

architecture SYN_ARCH2 of ND2_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_160;

architecture SYN_ARCH2 of ND2_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_157;

architecture SYN_ARCH2 of ND2_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_154;

architecture SYN_ARCH2 of ND2_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_151;

architecture SYN_ARCH2 of ND2_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_148;

architecture SYN_ARCH2 of ND2_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_145;

architecture SYN_ARCH2 of ND2_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_142;

architecture SYN_ARCH2 of ND2_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_139;

architecture SYN_ARCH2 of ND2_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_136;

architecture SYN_ARCH2 of ND2_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_133;

architecture SYN_ARCH2 of ND2_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_130;

architecture SYN_ARCH2 of ND2_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_127;

architecture SYN_ARCH2 of ND2_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_124;

architecture SYN_ARCH2 of ND2_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_121;

architecture SYN_ARCH2 of ND2_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_118;

architecture SYN_ARCH2 of ND2_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_115;

architecture SYN_ARCH2 of ND2_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_112;

architecture SYN_ARCH2 of ND2_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_109;

architecture SYN_ARCH2 of ND2_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_106;

architecture SYN_ARCH2 of ND2_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_103;

architecture SYN_ARCH2 of ND2_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_100;

architecture SYN_ARCH2 of ND2_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_97;

architecture SYN_ARCH2 of ND2_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_255 is

   port( A : in std_logic;  Y : out std_logic);

end IV_255;

architecture SYN_BEHAVIORAL of IV_255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_254 is

   port( A : in std_logic;  Y : out std_logic);

end IV_254;

architecture SYN_BEHAVIORAL of IV_254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_253 is

   port( A : in std_logic;  Y : out std_logic);

end IV_253;

architecture SYN_BEHAVIORAL of IV_253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_252 is

   port( A : in std_logic;  Y : out std_logic);

end IV_252;

architecture SYN_BEHAVIORAL of IV_252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_251 is

   port( A : in std_logic;  Y : out std_logic);

end IV_251;

architecture SYN_BEHAVIORAL of IV_251 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_250 is

   port( A : in std_logic;  Y : out std_logic);

end IV_250;

architecture SYN_BEHAVIORAL of IV_250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_249 is

   port( A : in std_logic;  Y : out std_logic);

end IV_249;

architecture SYN_BEHAVIORAL of IV_249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_248 is

   port( A : in std_logic;  Y : out std_logic);

end IV_248;

architecture SYN_BEHAVIORAL of IV_248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_247 is

   port( A : in std_logic;  Y : out std_logic);

end IV_247;

architecture SYN_BEHAVIORAL of IV_247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_246 is

   port( A : in std_logic;  Y : out std_logic);

end IV_246;

architecture SYN_BEHAVIORAL of IV_246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_245 is

   port( A : in std_logic;  Y : out std_logic);

end IV_245;

architecture SYN_BEHAVIORAL of IV_245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_244 is

   port( A : in std_logic;  Y : out std_logic);

end IV_244;

architecture SYN_BEHAVIORAL of IV_244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_243 is

   port( A : in std_logic;  Y : out std_logic);

end IV_243;

architecture SYN_BEHAVIORAL of IV_243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_242 is

   port( A : in std_logic;  Y : out std_logic);

end IV_242;

architecture SYN_BEHAVIORAL of IV_242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_241 is

   port( A : in std_logic;  Y : out std_logic);

end IV_241;

architecture SYN_BEHAVIORAL of IV_241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_240 is

   port( A : in std_logic;  Y : out std_logic);

end IV_240;

architecture SYN_BEHAVIORAL of IV_240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_239 is

   port( A : in std_logic;  Y : out std_logic);

end IV_239;

architecture SYN_BEHAVIORAL of IV_239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_238 is

   port( A : in std_logic;  Y : out std_logic);

end IV_238;

architecture SYN_BEHAVIORAL of IV_238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_237 is

   port( A : in std_logic;  Y : out std_logic);

end IV_237;

architecture SYN_BEHAVIORAL of IV_237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_236 is

   port( A : in std_logic;  Y : out std_logic);

end IV_236;

architecture SYN_BEHAVIORAL of IV_236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_235 is

   port( A : in std_logic;  Y : out std_logic);

end IV_235;

architecture SYN_BEHAVIORAL of IV_235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_234 is

   port( A : in std_logic;  Y : out std_logic);

end IV_234;

architecture SYN_BEHAVIORAL of IV_234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_233 is

   port( A : in std_logic;  Y : out std_logic);

end IV_233;

architecture SYN_BEHAVIORAL of IV_233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_232 is

   port( A : in std_logic;  Y : out std_logic);

end IV_232;

architecture SYN_BEHAVIORAL of IV_232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_231 is

   port( A : in std_logic;  Y : out std_logic);

end IV_231;

architecture SYN_BEHAVIORAL of IV_231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_230 is

   port( A : in std_logic;  Y : out std_logic);

end IV_230;

architecture SYN_BEHAVIORAL of IV_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_229 is

   port( A : in std_logic;  Y : out std_logic);

end IV_229;

architecture SYN_BEHAVIORAL of IV_229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_228 is

   port( A : in std_logic;  Y : out std_logic);

end IV_228;

architecture SYN_BEHAVIORAL of IV_228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_227 is

   port( A : in std_logic;  Y : out std_logic);

end IV_227;

architecture SYN_BEHAVIORAL of IV_227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_226 is

   port( A : in std_logic;  Y : out std_logic);

end IV_226;

architecture SYN_BEHAVIORAL of IV_226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_225 is

   port( A : in std_logic;  Y : out std_logic);

end IV_225;

architecture SYN_BEHAVIORAL of IV_225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_224 is

   port( A : in std_logic;  Y : out std_logic);

end IV_224;

architecture SYN_BEHAVIORAL of IV_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_223 is

   port( A : in std_logic;  Y : out std_logic);

end IV_223;

architecture SYN_BEHAVIORAL of IV_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_222 is

   port( A : in std_logic;  Y : out std_logic);

end IV_222;

architecture SYN_BEHAVIORAL of IV_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_221 is

   port( A : in std_logic;  Y : out std_logic);

end IV_221;

architecture SYN_BEHAVIORAL of IV_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_220 is

   port( A : in std_logic;  Y : out std_logic);

end IV_220;

architecture SYN_BEHAVIORAL of IV_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_219 is

   port( A : in std_logic;  Y : out std_logic);

end IV_219;

architecture SYN_BEHAVIORAL of IV_219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_218 is

   port( A : in std_logic;  Y : out std_logic);

end IV_218;

architecture SYN_BEHAVIORAL of IV_218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_217 is

   port( A : in std_logic;  Y : out std_logic);

end IV_217;

architecture SYN_BEHAVIORAL of IV_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_216 is

   port( A : in std_logic;  Y : out std_logic);

end IV_216;

architecture SYN_BEHAVIORAL of IV_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_215 is

   port( A : in std_logic;  Y : out std_logic);

end IV_215;

architecture SYN_BEHAVIORAL of IV_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_214 is

   port( A : in std_logic;  Y : out std_logic);

end IV_214;

architecture SYN_BEHAVIORAL of IV_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_213 is

   port( A : in std_logic;  Y : out std_logic);

end IV_213;

architecture SYN_BEHAVIORAL of IV_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_212 is

   port( A : in std_logic;  Y : out std_logic);

end IV_212;

architecture SYN_BEHAVIORAL of IV_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_211 is

   port( A : in std_logic;  Y : out std_logic);

end IV_211;

architecture SYN_BEHAVIORAL of IV_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_210 is

   port( A : in std_logic;  Y : out std_logic);

end IV_210;

architecture SYN_BEHAVIORAL of IV_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_209 is

   port( A : in std_logic;  Y : out std_logic);

end IV_209;

architecture SYN_BEHAVIORAL of IV_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_208 is

   port( A : in std_logic;  Y : out std_logic);

end IV_208;

architecture SYN_BEHAVIORAL of IV_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_207 is

   port( A : in std_logic;  Y : out std_logic);

end IV_207;

architecture SYN_BEHAVIORAL of IV_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_206 is

   port( A : in std_logic;  Y : out std_logic);

end IV_206;

architecture SYN_BEHAVIORAL of IV_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_205 is

   port( A : in std_logic;  Y : out std_logic);

end IV_205;

architecture SYN_BEHAVIORAL of IV_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_204 is

   port( A : in std_logic;  Y : out std_logic);

end IV_204;

architecture SYN_BEHAVIORAL of IV_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_203 is

   port( A : in std_logic;  Y : out std_logic);

end IV_203;

architecture SYN_BEHAVIORAL of IV_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_202 is

   port( A : in std_logic;  Y : out std_logic);

end IV_202;

architecture SYN_BEHAVIORAL of IV_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_201 is

   port( A : in std_logic;  Y : out std_logic);

end IV_201;

architecture SYN_BEHAVIORAL of IV_201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_200 is

   port( A : in std_logic;  Y : out std_logic);

end IV_200;

architecture SYN_BEHAVIORAL of IV_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_199 is

   port( A : in std_logic;  Y : out std_logic);

end IV_199;

architecture SYN_BEHAVIORAL of IV_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_198 is

   port( A : in std_logic;  Y : out std_logic);

end IV_198;

architecture SYN_BEHAVIORAL of IV_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_197 is

   port( A : in std_logic;  Y : out std_logic);

end IV_197;

architecture SYN_BEHAVIORAL of IV_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_196 is

   port( A : in std_logic;  Y : out std_logic);

end IV_196;

architecture SYN_BEHAVIORAL of IV_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_195 is

   port( A : in std_logic;  Y : out std_logic);

end IV_195;

architecture SYN_BEHAVIORAL of IV_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_194 is

   port( A : in std_logic;  Y : out std_logic);

end IV_194;

architecture SYN_BEHAVIORAL of IV_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_193 is

   port( A : in std_logic;  Y : out std_logic);

end IV_193;

architecture SYN_BEHAVIORAL of IV_193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_192 is

   port( A : in std_logic;  Y : out std_logic);

end IV_192;

architecture SYN_BEHAVIORAL of IV_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_191 is

   port( A : in std_logic;  Y : out std_logic);

end IV_191;

architecture SYN_BEHAVIORAL of IV_191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_190 is

   port( A : in std_logic;  Y : out std_logic);

end IV_190;

architecture SYN_BEHAVIORAL of IV_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_189 is

   port( A : in std_logic;  Y : out std_logic);

end IV_189;

architecture SYN_BEHAVIORAL of IV_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_188 is

   port( A : in std_logic;  Y : out std_logic);

end IV_188;

architecture SYN_BEHAVIORAL of IV_188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_187 is

   port( A : in std_logic;  Y : out std_logic);

end IV_187;

architecture SYN_BEHAVIORAL of IV_187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_186 is

   port( A : in std_logic;  Y : out std_logic);

end IV_186;

architecture SYN_BEHAVIORAL of IV_186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_185 is

   port( A : in std_logic;  Y : out std_logic);

end IV_185;

architecture SYN_BEHAVIORAL of IV_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_184 is

   port( A : in std_logic;  Y : out std_logic);

end IV_184;

architecture SYN_BEHAVIORAL of IV_184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_183 is

   port( A : in std_logic;  Y : out std_logic);

end IV_183;

architecture SYN_BEHAVIORAL of IV_183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_182 is

   port( A : in std_logic;  Y : out std_logic);

end IV_182;

architecture SYN_BEHAVIORAL of IV_182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_181 is

   port( A : in std_logic;  Y : out std_logic);

end IV_181;

architecture SYN_BEHAVIORAL of IV_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_180 is

   port( A : in std_logic;  Y : out std_logic);

end IV_180;

architecture SYN_BEHAVIORAL of IV_180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_179 is

   port( A : in std_logic;  Y : out std_logic);

end IV_179;

architecture SYN_BEHAVIORAL of IV_179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_178 is

   port( A : in std_logic;  Y : out std_logic);

end IV_178;

architecture SYN_BEHAVIORAL of IV_178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_177 is

   port( A : in std_logic;  Y : out std_logic);

end IV_177;

architecture SYN_BEHAVIORAL of IV_177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_176 is

   port( A : in std_logic;  Y : out std_logic);

end IV_176;

architecture SYN_BEHAVIORAL of IV_176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_175 is

   port( A : in std_logic;  Y : out std_logic);

end IV_175;

architecture SYN_BEHAVIORAL of IV_175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_174 is

   port( A : in std_logic;  Y : out std_logic);

end IV_174;

architecture SYN_BEHAVIORAL of IV_174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_173 is

   port( A : in std_logic;  Y : out std_logic);

end IV_173;

architecture SYN_BEHAVIORAL of IV_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_172 is

   port( A : in std_logic;  Y : out std_logic);

end IV_172;

architecture SYN_BEHAVIORAL of IV_172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_171 is

   port( A : in std_logic;  Y : out std_logic);

end IV_171;

architecture SYN_BEHAVIORAL of IV_171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_170 is

   port( A : in std_logic;  Y : out std_logic);

end IV_170;

architecture SYN_BEHAVIORAL of IV_170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_169 is

   port( A : in std_logic;  Y : out std_logic);

end IV_169;

architecture SYN_BEHAVIORAL of IV_169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_168 is

   port( A : in std_logic;  Y : out std_logic);

end IV_168;

architecture SYN_BEHAVIORAL of IV_168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_167 is

   port( A : in std_logic;  Y : out std_logic);

end IV_167;

architecture SYN_BEHAVIORAL of IV_167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_166 is

   port( A : in std_logic;  Y : out std_logic);

end IV_166;

architecture SYN_BEHAVIORAL of IV_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_165 is

   port( A : in std_logic;  Y : out std_logic);

end IV_165;

architecture SYN_BEHAVIORAL of IV_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_164 is

   port( A : in std_logic;  Y : out std_logic);

end IV_164;

architecture SYN_BEHAVIORAL of IV_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_163 is

   port( A : in std_logic;  Y : out std_logic);

end IV_163;

architecture SYN_BEHAVIORAL of IV_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_162 is

   port( A : in std_logic;  Y : out std_logic);

end IV_162;

architecture SYN_BEHAVIORAL of IV_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_161 is

   port( A : in std_logic;  Y : out std_logic);

end IV_161;

architecture SYN_BEHAVIORAL of IV_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_160 is

   port( A : in std_logic;  Y : out std_logic);

end IV_160;

architecture SYN_BEHAVIORAL of IV_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_159 is

   port( A : in std_logic;  Y : out std_logic);

end IV_159;

architecture SYN_BEHAVIORAL of IV_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_158 is

   port( A : in std_logic;  Y : out std_logic);

end IV_158;

architecture SYN_BEHAVIORAL of IV_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_157 is

   port( A : in std_logic;  Y : out std_logic);

end IV_157;

architecture SYN_BEHAVIORAL of IV_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_156 is

   port( A : in std_logic;  Y : out std_logic);

end IV_156;

architecture SYN_BEHAVIORAL of IV_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_155 is

   port( A : in std_logic;  Y : out std_logic);

end IV_155;

architecture SYN_BEHAVIORAL of IV_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_154 is

   port( A : in std_logic;  Y : out std_logic);

end IV_154;

architecture SYN_BEHAVIORAL of IV_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_153 is

   port( A : in std_logic;  Y : out std_logic);

end IV_153;

architecture SYN_BEHAVIORAL of IV_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_152 is

   port( A : in std_logic;  Y : out std_logic);

end IV_152;

architecture SYN_BEHAVIORAL of IV_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_151 is

   port( A : in std_logic;  Y : out std_logic);

end IV_151;

architecture SYN_BEHAVIORAL of IV_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_150 is

   port( A : in std_logic;  Y : out std_logic);

end IV_150;

architecture SYN_BEHAVIORAL of IV_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_149 is

   port( A : in std_logic;  Y : out std_logic);

end IV_149;

architecture SYN_BEHAVIORAL of IV_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_148 is

   port( A : in std_logic;  Y : out std_logic);

end IV_148;

architecture SYN_BEHAVIORAL of IV_148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_147 is

   port( A : in std_logic;  Y : out std_logic);

end IV_147;

architecture SYN_BEHAVIORAL of IV_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_146 is

   port( A : in std_logic;  Y : out std_logic);

end IV_146;

architecture SYN_BEHAVIORAL of IV_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_145 is

   port( A : in std_logic;  Y : out std_logic);

end IV_145;

architecture SYN_BEHAVIORAL of IV_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_144 is

   port( A : in std_logic;  Y : out std_logic);

end IV_144;

architecture SYN_BEHAVIORAL of IV_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_143 is

   port( A : in std_logic;  Y : out std_logic);

end IV_143;

architecture SYN_BEHAVIORAL of IV_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_142 is

   port( A : in std_logic;  Y : out std_logic);

end IV_142;

architecture SYN_BEHAVIORAL of IV_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_141 is

   port( A : in std_logic;  Y : out std_logic);

end IV_141;

architecture SYN_BEHAVIORAL of IV_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_140 is

   port( A : in std_logic;  Y : out std_logic);

end IV_140;

architecture SYN_BEHAVIORAL of IV_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_139 is

   port( A : in std_logic;  Y : out std_logic);

end IV_139;

architecture SYN_BEHAVIORAL of IV_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_138 is

   port( A : in std_logic;  Y : out std_logic);

end IV_138;

architecture SYN_BEHAVIORAL of IV_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_137 is

   port( A : in std_logic;  Y : out std_logic);

end IV_137;

architecture SYN_BEHAVIORAL of IV_137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_136 is

   port( A : in std_logic;  Y : out std_logic);

end IV_136;

architecture SYN_BEHAVIORAL of IV_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_135 is

   port( A : in std_logic;  Y : out std_logic);

end IV_135;

architecture SYN_BEHAVIORAL of IV_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_134 is

   port( A : in std_logic;  Y : out std_logic);

end IV_134;

architecture SYN_BEHAVIORAL of IV_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_133 is

   port( A : in std_logic;  Y : out std_logic);

end IV_133;

architecture SYN_BEHAVIORAL of IV_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_132 is

   port( A : in std_logic;  Y : out std_logic);

end IV_132;

architecture SYN_BEHAVIORAL of IV_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_131 is

   port( A : in std_logic;  Y : out std_logic);

end IV_131;

architecture SYN_BEHAVIORAL of IV_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_130 is

   port( A : in std_logic;  Y : out std_logic);

end IV_130;

architecture SYN_BEHAVIORAL of IV_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_129 is

   port( A : in std_logic;  Y : out std_logic);

end IV_129;

architecture SYN_BEHAVIORAL of IV_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_128 is

   port( A : in std_logic;  Y : out std_logic);

end IV_128;

architecture SYN_BEHAVIORAL of IV_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_127 is

   port( A : in std_logic;  Y : out std_logic);

end IV_127;

architecture SYN_BEHAVIORAL of IV_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_126 is

   port( A : in std_logic;  Y : out std_logic);

end IV_126;

architecture SYN_BEHAVIORAL of IV_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_125 is

   port( A : in std_logic;  Y : out std_logic);

end IV_125;

architecture SYN_BEHAVIORAL of IV_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_124 is

   port( A : in std_logic;  Y : out std_logic);

end IV_124;

architecture SYN_BEHAVIORAL of IV_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_123 is

   port( A : in std_logic;  Y : out std_logic);

end IV_123;

architecture SYN_BEHAVIORAL of IV_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_122 is

   port( A : in std_logic;  Y : out std_logic);

end IV_122;

architecture SYN_BEHAVIORAL of IV_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_121 is

   port( A : in std_logic;  Y : out std_logic);

end IV_121;

architecture SYN_BEHAVIORAL of IV_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_120 is

   port( A : in std_logic;  Y : out std_logic);

end IV_120;

architecture SYN_BEHAVIORAL of IV_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_119 is

   port( A : in std_logic;  Y : out std_logic);

end IV_119;

architecture SYN_BEHAVIORAL of IV_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_118 is

   port( A : in std_logic;  Y : out std_logic);

end IV_118;

architecture SYN_BEHAVIORAL of IV_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_117 is

   port( A : in std_logic;  Y : out std_logic);

end IV_117;

architecture SYN_BEHAVIORAL of IV_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_116 is

   port( A : in std_logic;  Y : out std_logic);

end IV_116;

architecture SYN_BEHAVIORAL of IV_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_115 is

   port( A : in std_logic;  Y : out std_logic);

end IV_115;

architecture SYN_BEHAVIORAL of IV_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_114 is

   port( A : in std_logic;  Y : out std_logic);

end IV_114;

architecture SYN_BEHAVIORAL of IV_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_113 is

   port( A : in std_logic;  Y : out std_logic);

end IV_113;

architecture SYN_BEHAVIORAL of IV_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_112 is

   port( A : in std_logic;  Y : out std_logic);

end IV_112;

architecture SYN_BEHAVIORAL of IV_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_111 is

   port( A : in std_logic;  Y : out std_logic);

end IV_111;

architecture SYN_BEHAVIORAL of IV_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_110 is

   port( A : in std_logic;  Y : out std_logic);

end IV_110;

architecture SYN_BEHAVIORAL of IV_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_109 is

   port( A : in std_logic;  Y : out std_logic);

end IV_109;

architecture SYN_BEHAVIORAL of IV_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_108 is

   port( A : in std_logic;  Y : out std_logic);

end IV_108;

architecture SYN_BEHAVIORAL of IV_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_107 is

   port( A : in std_logic;  Y : out std_logic);

end IV_107;

architecture SYN_BEHAVIORAL of IV_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_106 is

   port( A : in std_logic;  Y : out std_logic);

end IV_106;

architecture SYN_BEHAVIORAL of IV_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_105 is

   port( A : in std_logic;  Y : out std_logic);

end IV_105;

architecture SYN_BEHAVIORAL of IV_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_104 is

   port( A : in std_logic;  Y : out std_logic);

end IV_104;

architecture SYN_BEHAVIORAL of IV_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_103 is

   port( A : in std_logic;  Y : out std_logic);

end IV_103;

architecture SYN_BEHAVIORAL of IV_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_102 is

   port( A : in std_logic;  Y : out std_logic);

end IV_102;

architecture SYN_BEHAVIORAL of IV_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_101 is

   port( A : in std_logic;  Y : out std_logic);

end IV_101;

architecture SYN_BEHAVIORAL of IV_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_100 is

   port( A : in std_logic;  Y : out std_logic);

end IV_100;

architecture SYN_BEHAVIORAL of IV_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_99 is

   port( A : in std_logic;  Y : out std_logic);

end IV_99;

architecture SYN_BEHAVIORAL of IV_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_98 is

   port( A : in std_logic;  Y : out std_logic);

end IV_98;

architecture SYN_BEHAVIORAL of IV_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_97 is

   port( A : in std_logic;  Y : out std_logic);

end IV_97;

architecture SYN_BEHAVIORAL of IV_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_96 is

   port( A : in std_logic;  Y : out std_logic);

end IV_96;

architecture SYN_BEHAVIORAL of IV_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_95 is

   port( A : in std_logic;  Y : out std_logic);

end IV_95;

architecture SYN_BEHAVIORAL of IV_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_94 is

   port( A : in std_logic;  Y : out std_logic);

end IV_94;

architecture SYN_BEHAVIORAL of IV_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_93 is

   port( A : in std_logic;  Y : out std_logic);

end IV_93;

architecture SYN_BEHAVIORAL of IV_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_92 is

   port( A : in std_logic;  Y : out std_logic);

end IV_92;

architecture SYN_BEHAVIORAL of IV_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_91 is

   port( A : in std_logic;  Y : out std_logic);

end IV_91;

architecture SYN_BEHAVIORAL of IV_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_90 is

   port( A : in std_logic;  Y : out std_logic);

end IV_90;

architecture SYN_BEHAVIORAL of IV_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_89 is

   port( A : in std_logic;  Y : out std_logic);

end IV_89;

architecture SYN_BEHAVIORAL of IV_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_88 is

   port( A : in std_logic;  Y : out std_logic);

end IV_88;

architecture SYN_BEHAVIORAL of IV_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_87 is

   port( A : in std_logic;  Y : out std_logic);

end IV_87;

architecture SYN_BEHAVIORAL of IV_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_86 is

   port( A : in std_logic;  Y : out std_logic);

end IV_86;

architecture SYN_BEHAVIORAL of IV_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_85 is

   port( A : in std_logic;  Y : out std_logic);

end IV_85;

architecture SYN_BEHAVIORAL of IV_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_84 is

   port( A : in std_logic;  Y : out std_logic);

end IV_84;

architecture SYN_BEHAVIORAL of IV_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_83 is

   port( A : in std_logic;  Y : out std_logic);

end IV_83;

architecture SYN_BEHAVIORAL of IV_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_82 is

   port( A : in std_logic;  Y : out std_logic);

end IV_82;

architecture SYN_BEHAVIORAL of IV_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_81 is

   port( A : in std_logic;  Y : out std_logic);

end IV_81;

architecture SYN_BEHAVIORAL of IV_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_80 is

   port( A : in std_logic;  Y : out std_logic);

end IV_80;

architecture SYN_BEHAVIORAL of IV_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_79 is

   port( A : in std_logic;  Y : out std_logic);

end IV_79;

architecture SYN_BEHAVIORAL of IV_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_78 is

   port( A : in std_logic;  Y : out std_logic);

end IV_78;

architecture SYN_BEHAVIORAL of IV_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_77 is

   port( A : in std_logic;  Y : out std_logic);

end IV_77;

architecture SYN_BEHAVIORAL of IV_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_76 is

   port( A : in std_logic;  Y : out std_logic);

end IV_76;

architecture SYN_BEHAVIORAL of IV_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_75 is

   port( A : in std_logic;  Y : out std_logic);

end IV_75;

architecture SYN_BEHAVIORAL of IV_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_74 is

   port( A : in std_logic;  Y : out std_logic);

end IV_74;

architecture SYN_BEHAVIORAL of IV_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_73 is

   port( A : in std_logic;  Y : out std_logic);

end IV_73;

architecture SYN_BEHAVIORAL of IV_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_72 is

   port( A : in std_logic;  Y : out std_logic);

end IV_72;

architecture SYN_BEHAVIORAL of IV_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_71 is

   port( A : in std_logic;  Y : out std_logic);

end IV_71;

architecture SYN_BEHAVIORAL of IV_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_70 is

   port( A : in std_logic;  Y : out std_logic);

end IV_70;

architecture SYN_BEHAVIORAL of IV_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_69 is

   port( A : in std_logic;  Y : out std_logic);

end IV_69;

architecture SYN_BEHAVIORAL of IV_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_68 is

   port( A : in std_logic;  Y : out std_logic);

end IV_68;

architecture SYN_BEHAVIORAL of IV_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_67 is

   port( A : in std_logic;  Y : out std_logic);

end IV_67;

architecture SYN_BEHAVIORAL of IV_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_66 is

   port( A : in std_logic;  Y : out std_logic);

end IV_66;

architecture SYN_BEHAVIORAL of IV_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_65 is

   port( A : in std_logic;  Y : out std_logic);

end IV_65;

architecture SYN_BEHAVIORAL of IV_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_64 is

   port( A : in std_logic;  Y : out std_logic);

end IV_64;

architecture SYN_BEHAVIORAL of IV_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_191;

architecture SYN_STRUCTURAL of MUX21_191 is

   component ND2_571
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_572
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_573
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_191
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_191 port map( A => S, Y => SB);
   UND1 : ND2_573 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_572 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_571 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_190;

architecture SYN_STRUCTURAL of MUX21_190 is

   component ND2_568
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_569
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_570
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_190
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_190 port map( A => S, Y => SB);
   UND1 : ND2_570 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_569 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_568 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_189;

architecture SYN_STRUCTURAL of MUX21_189 is

   component ND2_565
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_566
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_567
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_189
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_189 port map( A => S, Y => SB);
   UND1 : ND2_567 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_566 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_565 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_255 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_255;

architecture SYN_STRUCTURAL of MUX21_255 is

   component ND2_763
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_764
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_765
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_255
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_255 port map( A => S, Y => SB);
   UND1 : ND2_765 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_764 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_763 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_254 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_254;

architecture SYN_STRUCTURAL of MUX21_254 is

   component ND2_760
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_761
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_762
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_254
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_254 port map( A => S, Y => SB);
   UND1 : ND2_762 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_761 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_760 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_253 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_253;

architecture SYN_STRUCTURAL of MUX21_253 is

   component ND2_757
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_758
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_759
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_253
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_253 port map( A => S, Y => SB);
   UND1 : ND2_759 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_758 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_757 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_252 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_252;

architecture SYN_STRUCTURAL of MUX21_252 is

   component ND2_754
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_755
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_756
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_252
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_252 port map( A => S, Y => SB);
   UND1 : ND2_756 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_755 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_754 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_251 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_251;

architecture SYN_STRUCTURAL of MUX21_251 is

   component ND2_751
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_752
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_753
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_251
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_251 port map( A => S, Y => SB);
   UND1 : ND2_753 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_752 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_751 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_250 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_250;

architecture SYN_STRUCTURAL of MUX21_250 is

   component ND2_748
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_749
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_750
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_250
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_250 port map( A => S, Y => SB);
   UND1 : ND2_750 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_749 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_748 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_249 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_249;

architecture SYN_STRUCTURAL of MUX21_249 is

   component ND2_745
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_746
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_747
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_249
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_249 port map( A => S, Y => SB);
   UND1 : ND2_747 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_746 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_745 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_248 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_248;

architecture SYN_STRUCTURAL of MUX21_248 is

   component ND2_742
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_743
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_744
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_248
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_248 port map( A => S, Y => SB);
   UND1 : ND2_744 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_743 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_742 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_247 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_247;

architecture SYN_STRUCTURAL of MUX21_247 is

   component ND2_739
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_740
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_741
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_247
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_247 port map( A => S, Y => SB);
   UND1 : ND2_741 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_740 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_739 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_246 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_246;

architecture SYN_STRUCTURAL of MUX21_246 is

   component ND2_736
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_737
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_738
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_246
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_246 port map( A => S, Y => SB);
   UND1 : ND2_738 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_737 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_736 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_245 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_245;

architecture SYN_STRUCTURAL of MUX21_245 is

   component ND2_733
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_734
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_735
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_245
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_245 port map( A => S, Y => SB);
   UND1 : ND2_735 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_734 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_733 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_244 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_244;

architecture SYN_STRUCTURAL of MUX21_244 is

   component ND2_730
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_731
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_732
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_244
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_244 port map( A => S, Y => SB);
   UND1 : ND2_732 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_731 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_730 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_243 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_243;

architecture SYN_STRUCTURAL of MUX21_243 is

   component ND2_727
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_728
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_729
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_243
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_243 port map( A => S, Y => SB);
   UND1 : ND2_729 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_728 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_727 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_242 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_242;

architecture SYN_STRUCTURAL of MUX21_242 is

   component ND2_724
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_725
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_726
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_242
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_242 port map( A => S, Y => SB);
   UND1 : ND2_726 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_725 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_724 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_241 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_241;

architecture SYN_STRUCTURAL of MUX21_241 is

   component ND2_721
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_722
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_723
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_241
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_241 port map( A => S, Y => SB);
   UND1 : ND2_723 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_722 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_721 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_240 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_240;

architecture SYN_STRUCTURAL of MUX21_240 is

   component ND2_718
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_719
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_720
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_240
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_240 port map( A => S, Y => SB);
   UND1 : ND2_720 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_719 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_718 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_239 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_239;

architecture SYN_STRUCTURAL of MUX21_239 is

   component ND2_715
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_716
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_717
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_239
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_239 port map( A => S, Y => SB);
   UND1 : ND2_717 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_716 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_715 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_238 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_238;

architecture SYN_STRUCTURAL of MUX21_238 is

   component ND2_712
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_713
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_714
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_238
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_238 port map( A => S, Y => SB);
   UND1 : ND2_714 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_713 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_712 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_237 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_237;

architecture SYN_STRUCTURAL of MUX21_237 is

   component ND2_709
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_710
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_711
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_237
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_237 port map( A => S, Y => SB);
   UND1 : ND2_711 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_710 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_709 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_236 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_236;

architecture SYN_STRUCTURAL of MUX21_236 is

   component ND2_706
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_707
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_708
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_236
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_236 port map( A => S, Y => SB);
   UND1 : ND2_708 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_707 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_706 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_235 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_235;

architecture SYN_STRUCTURAL of MUX21_235 is

   component ND2_703
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_704
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_705
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_235
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_235 port map( A => S, Y => SB);
   UND1 : ND2_705 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_704 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_703 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_234 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_234;

architecture SYN_STRUCTURAL of MUX21_234 is

   component ND2_700
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_701
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_702
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_234
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_234 port map( A => S, Y => SB);
   UND1 : ND2_702 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_701 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_700 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_233 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_233;

architecture SYN_STRUCTURAL of MUX21_233 is

   component ND2_697
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_698
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_699
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_233
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_233 port map( A => S, Y => SB);
   UND1 : ND2_699 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_698 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_697 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_232 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_232;

architecture SYN_STRUCTURAL of MUX21_232 is

   component ND2_694
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_695
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_696
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_232
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_232 port map( A => S, Y => SB);
   UND1 : ND2_696 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_695 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_694 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_231 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_231;

architecture SYN_STRUCTURAL of MUX21_231 is

   component ND2_691
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_692
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_693
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_231
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_231 port map( A => S, Y => SB);
   UND1 : ND2_693 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_692 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_691 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_230 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_230;

architecture SYN_STRUCTURAL of MUX21_230 is

   component ND2_688
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_689
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_690
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_230
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_230 port map( A => S, Y => SB);
   UND1 : ND2_690 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_689 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_688 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_229 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_229;

architecture SYN_STRUCTURAL of MUX21_229 is

   component ND2_685
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_686
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_687
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_229
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_229 port map( A => S, Y => SB);
   UND1 : ND2_687 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_686 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_685 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_228 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_228;

architecture SYN_STRUCTURAL of MUX21_228 is

   component ND2_682
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_683
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_684
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_228
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_228 port map( A => S, Y => SB);
   UND1 : ND2_684 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_683 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_682 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_227 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_227;

architecture SYN_STRUCTURAL of MUX21_227 is

   component ND2_679
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_680
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_681
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_227
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_227 port map( A => S, Y => SB);
   UND1 : ND2_681 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_680 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_679 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_226 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_226;

architecture SYN_STRUCTURAL of MUX21_226 is

   component ND2_676
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_677
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_678
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_226
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_226 port map( A => S, Y => SB);
   UND1 : ND2_678 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_677 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_676 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_225 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_225;

architecture SYN_STRUCTURAL of MUX21_225 is

   component ND2_673
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_674
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_675
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_225
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_225 port map( A => S, Y => SB);
   UND1 : ND2_675 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_674 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_673 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_224 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_224;

architecture SYN_STRUCTURAL of MUX21_224 is

   component ND2_670
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_671
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_672
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_224
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_224 port map( A => S, Y => SB);
   UND1 : ND2_672 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_671 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_670 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_223 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_223;

architecture SYN_STRUCTURAL of MUX21_223 is

   component ND2_667
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_668
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_669
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_223
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_223 port map( A => S, Y => SB);
   UND1 : ND2_669 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_668 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_667 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_222 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_222;

architecture SYN_STRUCTURAL of MUX21_222 is

   component ND2_664
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_665
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_666
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_222
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_222 port map( A => S, Y => SB);
   UND1 : ND2_666 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_665 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_664 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_221 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_221;

architecture SYN_STRUCTURAL of MUX21_221 is

   component ND2_661
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_662
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_663
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_221
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_221 port map( A => S, Y => SB);
   UND1 : ND2_663 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_662 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_661 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_220 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_220;

architecture SYN_STRUCTURAL of MUX21_220 is

   component ND2_658
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_659
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_660
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_220
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_220 port map( A => S, Y => SB);
   UND1 : ND2_660 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_659 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_658 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_219 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_219;

architecture SYN_STRUCTURAL of MUX21_219 is

   component ND2_655
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_656
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_657
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_219
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_219 port map( A => S, Y => SB);
   UND1 : ND2_657 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_656 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_655 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_218 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_218;

architecture SYN_STRUCTURAL of MUX21_218 is

   component ND2_652
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_653
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_654
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_218
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_218 port map( A => S, Y => SB);
   UND1 : ND2_654 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_653 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_652 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_217;

architecture SYN_STRUCTURAL of MUX21_217 is

   component ND2_649
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_650
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_651
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_217
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_217 port map( A => S, Y => SB);
   UND1 : ND2_651 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_650 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_649 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_216;

architecture SYN_STRUCTURAL of MUX21_216 is

   component ND2_646
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_647
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_648
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_216
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_216 port map( A => S, Y => SB);
   UND1 : ND2_648 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_647 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_646 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_215;

architecture SYN_STRUCTURAL of MUX21_215 is

   component ND2_643
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_644
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_645
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_215
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_215 port map( A => S, Y => SB);
   UND1 : ND2_645 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_644 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_643 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_214;

architecture SYN_STRUCTURAL of MUX21_214 is

   component ND2_640
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_641
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_642
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_214
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_214 port map( A => S, Y => SB);
   UND1 : ND2_642 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_641 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_640 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_213;

architecture SYN_STRUCTURAL of MUX21_213 is

   component ND2_637
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_638
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_639
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_213
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_213 port map( A => S, Y => SB);
   UND1 : ND2_639 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_638 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_637 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_212;

architecture SYN_STRUCTURAL of MUX21_212 is

   component ND2_634
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_635
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_636
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_212
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_212 port map( A => S, Y => SB);
   UND1 : ND2_636 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_635 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_634 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_211;

architecture SYN_STRUCTURAL of MUX21_211 is

   component ND2_631
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_632
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_633
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_211
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_211 port map( A => S, Y => SB);
   UND1 : ND2_633 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_632 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_631 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_210;

architecture SYN_STRUCTURAL of MUX21_210 is

   component ND2_628
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_629
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_630
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_210
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_210 port map( A => S, Y => SB);
   UND1 : ND2_630 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_629 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_628 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_209;

architecture SYN_STRUCTURAL of MUX21_209 is

   component ND2_625
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_626
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_627
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_209
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_209 port map( A => S, Y => SB);
   UND1 : ND2_627 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_626 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_625 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_208;

architecture SYN_STRUCTURAL of MUX21_208 is

   component ND2_622
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_623
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_624
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_208
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_208 port map( A => S, Y => SB);
   UND1 : ND2_624 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_623 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_622 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_207;

architecture SYN_STRUCTURAL of MUX21_207 is

   component ND2_619
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_620
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_621
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_207
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_207 port map( A => S, Y => SB);
   UND1 : ND2_621 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_620 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_619 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_206;

architecture SYN_STRUCTURAL of MUX21_206 is

   component ND2_616
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_617
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_618
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_206
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_206 port map( A => S, Y => SB);
   UND1 : ND2_618 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_617 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_616 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_205;

architecture SYN_STRUCTURAL of MUX21_205 is

   component ND2_613
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_614
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_615
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_205
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_205 port map( A => S, Y => SB);
   UND1 : ND2_615 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_614 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_613 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_204;

architecture SYN_STRUCTURAL of MUX21_204 is

   component ND2_610
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_611
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_612
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_204
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_204 port map( A => S, Y => SB);
   UND1 : ND2_612 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_611 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_610 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_203;

architecture SYN_STRUCTURAL of MUX21_203 is

   component ND2_607
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_608
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_609
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_203
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_203 port map( A => S, Y => SB);
   UND1 : ND2_609 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_608 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_607 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_202;

architecture SYN_STRUCTURAL of MUX21_202 is

   component ND2_604
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_605
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_606
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_202
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_202 port map( A => S, Y => SB);
   UND1 : ND2_606 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_605 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_604 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_201;

architecture SYN_STRUCTURAL of MUX21_201 is

   component ND2_601
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_602
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_603
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_201
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_201 port map( A => S, Y => SB);
   UND1 : ND2_603 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_602 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_601 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_200;

architecture SYN_STRUCTURAL of MUX21_200 is

   component ND2_598
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_599
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_600
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_200
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_200 port map( A => S, Y => SB);
   UND1 : ND2_600 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_599 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_598 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_199;

architecture SYN_STRUCTURAL of MUX21_199 is

   component ND2_595
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_596
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_597
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_199
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_199 port map( A => S, Y => SB);
   UND1 : ND2_597 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_596 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_595 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_198;

architecture SYN_STRUCTURAL of MUX21_198 is

   component ND2_592
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_593
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_594
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_198
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_198 port map( A => S, Y => SB);
   UND1 : ND2_594 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_593 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_592 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_197;

architecture SYN_STRUCTURAL of MUX21_197 is

   component ND2_589
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_590
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_591
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_197
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_197 port map( A => S, Y => SB);
   UND1 : ND2_591 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_590 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_589 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_196;

architecture SYN_STRUCTURAL of MUX21_196 is

   component ND2_586
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_587
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_588
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_196
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_196 port map( A => S, Y => SB);
   UND1 : ND2_588 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_587 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_586 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_195;

architecture SYN_STRUCTURAL of MUX21_195 is

   component ND2_583
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_584
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_585
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_195
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_195 port map( A => S, Y => SB);
   UND1 : ND2_585 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_584 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_583 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_194;

architecture SYN_STRUCTURAL of MUX21_194 is

   component ND2_580
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_581
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_582
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_194
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_194 port map( A => S, Y => SB);
   UND1 : ND2_582 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_581 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_580 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_193;

architecture SYN_STRUCTURAL of MUX21_193 is

   component ND2_577
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_578
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_579
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_193
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_193 port map( A => S, Y => SB);
   UND1 : ND2_579 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_578 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_577 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_188;

architecture SYN_STRUCTURAL of MUX21_188 is

   component ND2_562
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_563
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_564
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_188
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_188 port map( A => S, Y => SB);
   UND1 : ND2_564 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_563 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_562 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_187;

architecture SYN_STRUCTURAL of MUX21_187 is

   component ND2_559
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_560
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_561
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_187
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_187 port map( A => S, Y => SB);
   UND1 : ND2_561 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_560 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_559 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_186;

architecture SYN_STRUCTURAL of MUX21_186 is

   component ND2_556
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_557
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_558
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_186
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_186 port map( A => S, Y => SB);
   UND1 : ND2_558 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_557 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_556 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_185;

architecture SYN_STRUCTURAL of MUX21_185 is

   component ND2_553
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_554
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_555
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_185
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_185 port map( A => S, Y => SB);
   UND1 : ND2_555 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_554 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_553 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_184;

architecture SYN_STRUCTURAL of MUX21_184 is

   component ND2_550
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_551
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_552
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_184
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_184 port map( A => S, Y => SB);
   UND1 : ND2_552 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_551 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_550 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_183;

architecture SYN_STRUCTURAL of MUX21_183 is

   component ND2_547
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_548
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_549
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_183
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_183 port map( A => S, Y => SB);
   UND1 : ND2_549 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_548 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_547 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_182;

architecture SYN_STRUCTURAL of MUX21_182 is

   component ND2_544
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_545
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_546
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_182
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_182 port map( A => S, Y => SB);
   UND1 : ND2_546 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_545 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_544 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_181;

architecture SYN_STRUCTURAL of MUX21_181 is

   component ND2_541
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_542
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_543
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_181
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_181 port map( A => S, Y => SB);
   UND1 : ND2_543 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_542 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_541 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_180;

architecture SYN_STRUCTURAL of MUX21_180 is

   component ND2_538
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_539
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_540
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_180
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_180 port map( A => S, Y => SB);
   UND1 : ND2_540 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_539 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_538 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_179;

architecture SYN_STRUCTURAL of MUX21_179 is

   component ND2_535
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_536
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_537
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_179
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_179 port map( A => S, Y => SB);
   UND1 : ND2_537 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_536 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_535 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_178;

architecture SYN_STRUCTURAL of MUX21_178 is

   component ND2_532
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_533
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_534
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_178
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_178 port map( A => S, Y => SB);
   UND1 : ND2_534 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_533 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_532 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_177;

architecture SYN_STRUCTURAL of MUX21_177 is

   component ND2_529
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_530
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_531
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_177
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_177 port map( A => S, Y => SB);
   UND1 : ND2_531 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_530 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_529 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_176;

architecture SYN_STRUCTURAL of MUX21_176 is

   component ND2_526
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_527
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_528
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_176
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_176 port map( A => S, Y => SB);
   UND1 : ND2_528 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_527 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_526 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_175;

architecture SYN_STRUCTURAL of MUX21_175 is

   component ND2_523
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_524
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_525
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_175
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_175 port map( A => S, Y => SB);
   UND1 : ND2_525 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_524 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_523 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_174;

architecture SYN_STRUCTURAL of MUX21_174 is

   component ND2_520
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_521
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_522
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_174
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_174 port map( A => S, Y => SB);
   UND1 : ND2_522 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_521 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_520 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_173;

architecture SYN_STRUCTURAL of MUX21_173 is

   component ND2_517
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_518
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_519
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_173
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_173 port map( A => S, Y => SB);
   UND1 : ND2_519 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_518 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_517 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_172;

architecture SYN_STRUCTURAL of MUX21_172 is

   component ND2_514
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_515
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_516
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_172
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_172 port map( A => S, Y => SB);
   UND1 : ND2_516 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_515 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_514 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_171;

architecture SYN_STRUCTURAL of MUX21_171 is

   component ND2_511
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_512
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_513
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_171
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_171 port map( A => S, Y => SB);
   UND1 : ND2_513 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_512 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_511 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_170;

architecture SYN_STRUCTURAL of MUX21_170 is

   component ND2_508
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_509
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_510
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_170
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_170 port map( A => S, Y => SB);
   UND1 : ND2_510 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_509 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_508 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_169;

architecture SYN_STRUCTURAL of MUX21_169 is

   component ND2_505
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_506
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_507
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_169
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_169 port map( A => S, Y => SB);
   UND1 : ND2_507 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_506 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_505 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_168;

architecture SYN_STRUCTURAL of MUX21_168 is

   component ND2_502
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_503
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_504
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_168
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_168 port map( A => S, Y => SB);
   UND1 : ND2_504 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_503 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_502 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_167;

architecture SYN_STRUCTURAL of MUX21_167 is

   component ND2_499
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_500
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_501
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_167
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_167 port map( A => S, Y => SB);
   UND1 : ND2_501 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_500 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_499 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_166;

architecture SYN_STRUCTURAL of MUX21_166 is

   component ND2_496
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_497
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_498
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_166
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_166 port map( A => S, Y => SB);
   UND1 : ND2_498 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_497 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_496 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_165;

architecture SYN_STRUCTURAL of MUX21_165 is

   component ND2_493
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_494
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_495
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_165
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_165 port map( A => S, Y => SB);
   UND1 : ND2_495 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_494 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_493 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_164;

architecture SYN_STRUCTURAL of MUX21_164 is

   component ND2_490
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_491
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_492
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_164
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_164 port map( A => S, Y => SB);
   UND1 : ND2_492 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_491 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_490 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_163;

architecture SYN_STRUCTURAL of MUX21_163 is

   component ND2_487
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_488
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_489
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_163
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_163 port map( A => S, Y => SB);
   UND1 : ND2_489 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_488 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_487 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_162;

architecture SYN_STRUCTURAL of MUX21_162 is

   component ND2_484
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_485
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_486
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_162
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_162 port map( A => S, Y => SB);
   UND1 : ND2_486 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_485 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_484 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_161;

architecture SYN_STRUCTURAL of MUX21_161 is

   component ND2_481
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_482
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_483
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_161
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_161 port map( A => S, Y => SB);
   UND1 : ND2_483 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_482 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_481 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_160;

architecture SYN_STRUCTURAL of MUX21_160 is

   component ND2_478
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_479
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_480
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_160
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_160 port map( A => S, Y => SB);
   UND1 : ND2_480 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_479 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_478 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_159;

architecture SYN_STRUCTURAL of MUX21_159 is

   component ND2_475
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_476
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_477
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_159
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_159 port map( A => S, Y => SB);
   UND1 : ND2_477 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_476 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_475 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_158;

architecture SYN_STRUCTURAL of MUX21_158 is

   component ND2_472
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_473
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_474
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_158
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_158 port map( A => S, Y => SB);
   UND1 : ND2_474 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_473 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_472 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_157;

architecture SYN_STRUCTURAL of MUX21_157 is

   component ND2_469
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_470
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_471
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_157
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_157 port map( A => S, Y => SB);
   UND1 : ND2_471 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_470 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_469 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_156;

architecture SYN_STRUCTURAL of MUX21_156 is

   component ND2_466
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_467
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_468
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_156
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_156 port map( A => S, Y => SB);
   UND1 : ND2_468 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_467 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_466 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_155;

architecture SYN_STRUCTURAL of MUX21_155 is

   component ND2_463
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_464
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_465
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_155
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_155 port map( A => S, Y => SB);
   UND1 : ND2_465 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_464 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_463 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_154;

architecture SYN_STRUCTURAL of MUX21_154 is

   component ND2_460
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_461
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_462
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_154
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_154 port map( A => S, Y => SB);
   UND1 : ND2_462 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_461 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_460 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_153;

architecture SYN_STRUCTURAL of MUX21_153 is

   component ND2_457
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_458
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_459
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_153
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_153 port map( A => S, Y => SB);
   UND1 : ND2_459 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_458 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_457 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_152;

architecture SYN_STRUCTURAL of MUX21_152 is

   component ND2_454
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_455
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_456
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_152
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_152 port map( A => S, Y => SB);
   UND1 : ND2_456 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_455 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_454 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_151;

architecture SYN_STRUCTURAL of MUX21_151 is

   component ND2_451
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_452
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_453
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_151
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_151 port map( A => S, Y => SB);
   UND1 : ND2_453 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_452 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_451 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_150;

architecture SYN_STRUCTURAL of MUX21_150 is

   component ND2_448
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_449
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_450
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_150
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_150 port map( A => S, Y => SB);
   UND1 : ND2_450 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_449 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_448 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_149;

architecture SYN_STRUCTURAL of MUX21_149 is

   component ND2_445
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_446
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_447
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_149
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_149 port map( A => S, Y => SB);
   UND1 : ND2_447 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_446 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_445 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_148;

architecture SYN_STRUCTURAL of MUX21_148 is

   component ND2_442
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_443
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_444
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_148
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_148 port map( A => S, Y => SB);
   UND1 : ND2_444 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_443 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_442 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_147;

architecture SYN_STRUCTURAL of MUX21_147 is

   component ND2_439
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_440
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_441
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_147
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_147 port map( A => S, Y => SB);
   UND1 : ND2_441 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_440 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_439 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_146;

architecture SYN_STRUCTURAL of MUX21_146 is

   component ND2_436
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_437
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_438
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_146
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_146 port map( A => S, Y => SB);
   UND1 : ND2_438 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_437 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_436 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_145;

architecture SYN_STRUCTURAL of MUX21_145 is

   component ND2_433
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_434
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_435
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_145
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_145 port map( A => S, Y => SB);
   UND1 : ND2_435 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_434 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_433 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_144;

architecture SYN_STRUCTURAL of MUX21_144 is

   component ND2_430
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_431
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_432
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_144
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_144 port map( A => S, Y => SB);
   UND1 : ND2_432 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_431 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_430 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_143;

architecture SYN_STRUCTURAL of MUX21_143 is

   component ND2_427
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_428
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_429
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_143
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_143 port map( A => S, Y => SB);
   UND1 : ND2_429 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_428 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_427 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_142;

architecture SYN_STRUCTURAL of MUX21_142 is

   component ND2_424
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_425
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_426
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_142
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_142 port map( A => S, Y => SB);
   UND1 : ND2_426 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_425 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_424 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_141;

architecture SYN_STRUCTURAL of MUX21_141 is

   component ND2_421
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_422
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_423
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_141
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_141 port map( A => S, Y => SB);
   UND1 : ND2_423 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_422 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_421 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_140;

architecture SYN_STRUCTURAL of MUX21_140 is

   component ND2_418
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_419
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_420
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_140
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_140 port map( A => S, Y => SB);
   UND1 : ND2_420 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_419 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_418 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_139;

architecture SYN_STRUCTURAL of MUX21_139 is

   component ND2_415
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_416
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_417
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_139
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_139 port map( A => S, Y => SB);
   UND1 : ND2_417 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_416 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_415 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_138;

architecture SYN_STRUCTURAL of MUX21_138 is

   component ND2_412
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_413
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_414
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_138
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_138 port map( A => S, Y => SB);
   UND1 : ND2_414 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_413 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_412 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_137;

architecture SYN_STRUCTURAL of MUX21_137 is

   component ND2_409
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_410
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_411
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_137
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_137 port map( A => S, Y => SB);
   UND1 : ND2_411 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_410 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_409 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_136;

architecture SYN_STRUCTURAL of MUX21_136 is

   component ND2_406
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_407
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_408
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_136
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_136 port map( A => S, Y => SB);
   UND1 : ND2_408 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_407 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_406 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_135;

architecture SYN_STRUCTURAL of MUX21_135 is

   component ND2_403
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_404
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_405
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_135
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_135 port map( A => S, Y => SB);
   UND1 : ND2_405 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_404 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_403 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_134;

architecture SYN_STRUCTURAL of MUX21_134 is

   component ND2_400
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_401
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_402
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_134
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_134 port map( A => S, Y => SB);
   UND1 : ND2_402 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_401 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_400 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_133;

architecture SYN_STRUCTURAL of MUX21_133 is

   component ND2_397
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_398
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_399
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_133
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_133 port map( A => S, Y => SB);
   UND1 : ND2_399 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_398 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_397 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_132;

architecture SYN_STRUCTURAL of MUX21_132 is

   component ND2_394
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_395
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_396
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_132
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_132 port map( A => S, Y => SB);
   UND1 : ND2_396 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_395 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_394 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_131;

architecture SYN_STRUCTURAL of MUX21_131 is

   component ND2_391
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_392
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_393
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_131
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_131 port map( A => S, Y => SB);
   UND1 : ND2_393 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_392 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_391 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_130;

architecture SYN_STRUCTURAL of MUX21_130 is

   component ND2_388
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_389
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_390
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_130
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_130 port map( A => S, Y => SB);
   UND1 : ND2_390 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_389 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_388 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_129;

architecture SYN_STRUCTURAL of MUX21_129 is

   component ND2_385
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_386
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_387
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_129
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_129 port map( A => S, Y => SB);
   UND1 : ND2_387 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_386 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_385 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_128;

architecture SYN_STRUCTURAL of MUX21_128 is

   component ND2_382
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_383
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_384
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_128
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_128 port map( A => S, Y => SB);
   UND1 : ND2_384 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_383 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_382 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_127 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_127;

architecture SYN_STRUCTURAL of MUX21_127 is

   component ND2_379
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_380
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_381
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_127
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_127 port map( A => S, Y => SB);
   UND1 : ND2_381 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_380 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_379 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_126 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_126;

architecture SYN_STRUCTURAL of MUX21_126 is

   component ND2_376
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_377
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_378
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_126
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_126 port map( A => S, Y => SB);
   UND1 : ND2_378 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_377 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_376 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_125 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_125;

architecture SYN_STRUCTURAL of MUX21_125 is

   component ND2_373
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_374
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_375
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_125
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_125 port map( A => S, Y => SB);
   UND1 : ND2_375 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_374 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_373 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_124 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_124;

architecture SYN_STRUCTURAL of MUX21_124 is

   component ND2_370
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_371
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_372
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_124
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_124 port map( A => S, Y => SB);
   UND1 : ND2_372 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_371 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_370 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_123 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_123;

architecture SYN_STRUCTURAL of MUX21_123 is

   component ND2_367
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_368
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_369
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_123
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_123 port map( A => S, Y => SB);
   UND1 : ND2_369 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_368 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_367 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_122 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_122;

architecture SYN_STRUCTURAL of MUX21_122 is

   component ND2_364
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_365
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_366
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_122
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_122 port map( A => S, Y => SB);
   UND1 : ND2_366 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_365 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_364 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_121 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_121;

architecture SYN_STRUCTURAL of MUX21_121 is

   component ND2_361
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_362
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_363
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_121
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_121 port map( A => S, Y => SB);
   UND1 : ND2_363 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_362 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_361 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_120 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_120;

architecture SYN_STRUCTURAL of MUX21_120 is

   component ND2_358
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_359
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_360
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_120
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_120 port map( A => S, Y => SB);
   UND1 : ND2_360 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_359 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_358 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_119 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_119;

architecture SYN_STRUCTURAL of MUX21_119 is

   component ND2_355
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_356
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_357
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_119
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_119 port map( A => S, Y => SB);
   UND1 : ND2_357 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_356 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_355 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_118 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_118;

architecture SYN_STRUCTURAL of MUX21_118 is

   component ND2_352
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_353
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_354
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_118
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_118 port map( A => S, Y => SB);
   UND1 : ND2_354 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_353 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_352 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_117 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_117;

architecture SYN_STRUCTURAL of MUX21_117 is

   component ND2_349
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_350
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_351
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_117
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_117 port map( A => S, Y => SB);
   UND1 : ND2_351 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_350 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_349 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_116 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_116;

architecture SYN_STRUCTURAL of MUX21_116 is

   component ND2_346
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_347
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_348
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_116
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_116 port map( A => S, Y => SB);
   UND1 : ND2_348 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_347 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_346 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_115 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_115;

architecture SYN_STRUCTURAL of MUX21_115 is

   component ND2_343
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_344
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_345
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_115
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_115 port map( A => S, Y => SB);
   UND1 : ND2_345 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_344 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_343 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_114 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_114;

architecture SYN_STRUCTURAL of MUX21_114 is

   component ND2_340
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_341
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_342
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_114
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_114 port map( A => S, Y => SB);
   UND1 : ND2_342 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_341 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_340 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_113 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_113;

architecture SYN_STRUCTURAL of MUX21_113 is

   component ND2_337
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_338
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_339
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_113
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_113 port map( A => S, Y => SB);
   UND1 : ND2_339 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_338 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_337 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_112 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_112;

architecture SYN_STRUCTURAL of MUX21_112 is

   component ND2_334
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_335
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_336
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_112
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_112 port map( A => S, Y => SB);
   UND1 : ND2_336 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_335 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_334 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_111 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_111;

architecture SYN_STRUCTURAL of MUX21_111 is

   component ND2_331
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_332
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_333
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_111
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_111 port map( A => S, Y => SB);
   UND1 : ND2_333 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_332 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_331 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_110 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_110;

architecture SYN_STRUCTURAL of MUX21_110 is

   component ND2_328
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_329
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_330
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_110
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_110 port map( A => S, Y => SB);
   UND1 : ND2_330 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_329 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_328 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_109 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_109;

architecture SYN_STRUCTURAL of MUX21_109 is

   component ND2_325
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_326
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_327
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_109
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_109 port map( A => S, Y => SB);
   UND1 : ND2_327 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_326 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_325 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_108 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_108;

architecture SYN_STRUCTURAL of MUX21_108 is

   component ND2_322
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_323
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_324
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_108
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_108 port map( A => S, Y => SB);
   UND1 : ND2_324 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_323 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_322 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_107 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_107;

architecture SYN_STRUCTURAL of MUX21_107 is

   component ND2_319
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_320
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_321
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_107
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_107 port map( A => S, Y => SB);
   UND1 : ND2_321 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_320 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_319 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_106 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_106;

architecture SYN_STRUCTURAL of MUX21_106 is

   component ND2_316
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_317
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_318
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_106
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_106 port map( A => S, Y => SB);
   UND1 : ND2_318 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_317 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_316 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_105 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_105;

architecture SYN_STRUCTURAL of MUX21_105 is

   component ND2_313
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_314
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_315
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_105
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_105 port map( A => S, Y => SB);
   UND1 : ND2_315 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_314 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_313 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_104 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_104;

architecture SYN_STRUCTURAL of MUX21_104 is

   component ND2_310
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_311
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_312
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_104
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_104 port map( A => S, Y => SB);
   UND1 : ND2_312 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_311 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_310 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_103 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_103;

architecture SYN_STRUCTURAL of MUX21_103 is

   component ND2_307
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_308
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_309
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_103
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_103 port map( A => S, Y => SB);
   UND1 : ND2_309 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_308 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_307 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_102 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_102;

architecture SYN_STRUCTURAL of MUX21_102 is

   component ND2_304
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_305
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_306
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_102
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_102 port map( A => S, Y => SB);
   UND1 : ND2_306 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_305 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_304 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_101 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_101;

architecture SYN_STRUCTURAL of MUX21_101 is

   component ND2_301
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_302
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_303
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_101
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_101 port map( A => S, Y => SB);
   UND1 : ND2_303 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_302 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_301 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_100 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_100;

architecture SYN_STRUCTURAL of MUX21_100 is

   component ND2_298
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_299
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_300
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_100
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_100 port map( A => S, Y => SB);
   UND1 : ND2_300 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_299 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_298 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_99 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_99;

architecture SYN_STRUCTURAL of MUX21_99 is

   component ND2_295
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_296
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_297
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_99
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_99 port map( A => S, Y => SB);
   UND1 : ND2_297 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_296 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_295 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_98 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_98;

architecture SYN_STRUCTURAL of MUX21_98 is

   component ND2_292
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_293
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_294
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_98
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_98 port map( A => S, Y => SB);
   UND1 : ND2_294 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_293 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_292 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_97 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_97;

architecture SYN_STRUCTURAL of MUX21_97 is

   component ND2_289
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_290
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_291
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_97
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_97 port map( A => S, Y => SB);
   UND1 : ND2_291 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_290 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_289 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_96 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_96;

architecture SYN_STRUCTURAL of MUX21_96 is

   component ND2_286
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_287
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_288
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_96
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_96 port map( A => S, Y => SB);
   UND1 : ND2_288 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_287 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_286 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_95 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_95;

architecture SYN_STRUCTURAL of MUX21_95 is

   component ND2_283
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_284
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_285
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_95
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_95 port map( A => S, Y => SB);
   UND1 : ND2_285 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_284 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_283 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_94 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_94;

architecture SYN_STRUCTURAL of MUX21_94 is

   component ND2_280
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_281
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_282
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_94
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_94 port map( A => S, Y => SB);
   UND1 : ND2_282 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_281 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_280 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_93 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_93;

architecture SYN_STRUCTURAL of MUX21_93 is

   component ND2_277
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_278
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_279
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_93
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_93 port map( A => S, Y => SB);
   UND1 : ND2_279 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_278 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_277 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_92 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_92;

architecture SYN_STRUCTURAL of MUX21_92 is

   component ND2_274
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_275
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_276
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_92
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_92 port map( A => S, Y => SB);
   UND1 : ND2_276 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_275 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_274 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_91 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_91;

architecture SYN_STRUCTURAL of MUX21_91 is

   component ND2_271
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_272
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_273
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_91
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_91 port map( A => S, Y => SB);
   UND1 : ND2_273 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_272 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_271 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_90 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_90;

architecture SYN_STRUCTURAL of MUX21_90 is

   component ND2_268
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_269
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_270
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_90
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_90 port map( A => S, Y => SB);
   UND1 : ND2_270 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_269 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_268 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_89 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_89;

architecture SYN_STRUCTURAL of MUX21_89 is

   component ND2_265
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_266
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_267
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_89
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_89 port map( A => S, Y => SB);
   UND1 : ND2_267 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_266 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_265 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_88 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_88;

architecture SYN_STRUCTURAL of MUX21_88 is

   component ND2_262
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_263
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_264
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_88
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_88 port map( A => S, Y => SB);
   UND1 : ND2_264 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_263 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_262 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_87 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_87;

architecture SYN_STRUCTURAL of MUX21_87 is

   component ND2_259
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_260
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_261
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_87
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_87 port map( A => S, Y => SB);
   UND1 : ND2_261 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_260 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_259 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_86 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_86;

architecture SYN_STRUCTURAL of MUX21_86 is

   component ND2_256
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_257
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_258
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_86
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_86 port map( A => S, Y => SB);
   UND1 : ND2_258 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_257 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_256 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_85 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_85;

architecture SYN_STRUCTURAL of MUX21_85 is

   component ND2_253
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_254
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_255
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_85
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_85 port map( A => S, Y => SB);
   UND1 : ND2_255 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_254 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_253 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_84 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_84;

architecture SYN_STRUCTURAL of MUX21_84 is

   component ND2_250
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_251
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_252
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_84
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_84 port map( A => S, Y => SB);
   UND1 : ND2_252 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_251 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_250 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_83 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_83;

architecture SYN_STRUCTURAL of MUX21_83 is

   component ND2_247
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_248
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_249
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_83
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_83 port map( A => S, Y => SB);
   UND1 : ND2_249 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_248 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_247 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_82 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_82;

architecture SYN_STRUCTURAL of MUX21_82 is

   component ND2_244
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_245
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_246
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_82
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_82 port map( A => S, Y => SB);
   UND1 : ND2_246 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_245 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_244 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_81 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_81;

architecture SYN_STRUCTURAL of MUX21_81 is

   component ND2_241
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_242
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_243
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_81
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_81 port map( A => S, Y => SB);
   UND1 : ND2_243 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_242 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_241 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_80 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_80;

architecture SYN_STRUCTURAL of MUX21_80 is

   component ND2_238
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_239
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_240
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_80
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_80 port map( A => S, Y => SB);
   UND1 : ND2_240 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_239 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_238 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_79 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_79;

architecture SYN_STRUCTURAL of MUX21_79 is

   component ND2_235
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_236
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_237
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_79
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_79 port map( A => S, Y => SB);
   UND1 : ND2_237 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_236 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_235 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_78 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_78;

architecture SYN_STRUCTURAL of MUX21_78 is

   component ND2_232
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_233
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_234
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_78
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_78 port map( A => S, Y => SB);
   UND1 : ND2_234 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_233 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_232 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_77 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_77;

architecture SYN_STRUCTURAL of MUX21_77 is

   component ND2_229
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_230
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_231
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_77
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_77 port map( A => S, Y => SB);
   UND1 : ND2_231 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_230 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_229 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_76 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_76;

architecture SYN_STRUCTURAL of MUX21_76 is

   component ND2_226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_76
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_76 port map( A => S, Y => SB);
   UND1 : ND2_228 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_227 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_226 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_75 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_75;

architecture SYN_STRUCTURAL of MUX21_75 is

   component ND2_223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_75
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_75 port map( A => S, Y => SB);
   UND1 : ND2_225 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_224 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_223 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_74 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_74;

architecture SYN_STRUCTURAL of MUX21_74 is

   component ND2_220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_74
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_74 port map( A => S, Y => SB);
   UND1 : ND2_222 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_221 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_220 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_73 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_73;

architecture SYN_STRUCTURAL of MUX21_73 is

   component ND2_217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_73
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_73 port map( A => S, Y => SB);
   UND1 : ND2_219 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_218 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_217 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_72 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_72;

architecture SYN_STRUCTURAL of MUX21_72 is

   component ND2_214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_72
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_72 port map( A => S, Y => SB);
   UND1 : ND2_216 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_215 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_214 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_71 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_71;

architecture SYN_STRUCTURAL of MUX21_71 is

   component ND2_211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_71
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_71 port map( A => S, Y => SB);
   UND1 : ND2_213 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_212 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_211 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_70 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_70;

architecture SYN_STRUCTURAL of MUX21_70 is

   component ND2_208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_70
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_70 port map( A => S, Y => SB);
   UND1 : ND2_210 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_209 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_208 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_69 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_69;

architecture SYN_STRUCTURAL of MUX21_69 is

   component ND2_205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_69
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_69 port map( A => S, Y => SB);
   UND1 : ND2_207 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_206 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_205 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_68 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_68;

architecture SYN_STRUCTURAL of MUX21_68 is

   component ND2_202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_68
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_68 port map( A => S, Y => SB);
   UND1 : ND2_204 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_203 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_202 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_67 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_67;

architecture SYN_STRUCTURAL of MUX21_67 is

   component ND2_199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_67
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_67 port map( A => S, Y => SB);
   UND1 : ND2_201 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_200 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_199 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_66 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_66;

architecture SYN_STRUCTURAL of MUX21_66 is

   component ND2_196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_66
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_66 port map( A => S, Y => SB);
   UND1 : ND2_198 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_197 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_196 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_65 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_65;

architecture SYN_STRUCTURAL of MUX21_65 is

   component ND2_193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_65
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_65 port map( A => S, Y => SB);
   UND1 : ND2_195 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_194 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_193 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_32;

architecture SYN_STRUCTURAL of MUX21_32 is

   component ND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_32 port map( A => S, Y => SB);
   UND1 : ND2_96 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31;

architecture SYN_STRUCTURAL of MUX21_31 is

   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31 port map( A => S, Y => SB);
   UND1 : ND2_93 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_92 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_91 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30;

architecture SYN_STRUCTURAL of MUX21_30 is

   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30 port map( A => S, Y => SB);
   UND1 : ND2_90 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_89 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_88 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_29;

architecture SYN_STRUCTURAL of MUX21_29 is

   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_29 port map( A => S, Y => SB);
   UND1 : ND2_87 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_86 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_85 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_63 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_63;

architecture SYN_STRUCTURAL of MUX21_63 is

   component ND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_63 port map( A => S, Y => SB);
   UND1 : ND2_189 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_188 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_187 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_62 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_62;

architecture SYN_STRUCTURAL of MUX21_62 is

   component ND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_62 port map( A => S, Y => SB);
   UND1 : ND2_186 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_185 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_184 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_61 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_61;

architecture SYN_STRUCTURAL of MUX21_61 is

   component ND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_61 port map( A => S, Y => SB);
   UND1 : ND2_183 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_182 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_181 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_60;

architecture SYN_STRUCTURAL of MUX21_60 is

   component ND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_60 port map( A => S, Y => SB);
   UND1 : ND2_180 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_179 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_178 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_59;

architecture SYN_STRUCTURAL of MUX21_59 is

   component ND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_59 port map( A => S, Y => SB);
   UND1 : ND2_177 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_176 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_175 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_58;

architecture SYN_STRUCTURAL of MUX21_58 is

   component ND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_58 port map( A => S, Y => SB);
   UND1 : ND2_174 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_173 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_172 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_57;

architecture SYN_STRUCTURAL of MUX21_57 is

   component ND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_57 port map( A => S, Y => SB);
   UND1 : ND2_171 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_170 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_169 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_56;

architecture SYN_STRUCTURAL of MUX21_56 is

   component ND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_56 port map( A => S, Y => SB);
   UND1 : ND2_168 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_167 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_166 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_55;

architecture SYN_STRUCTURAL of MUX21_55 is

   component ND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_55 port map( A => S, Y => SB);
   UND1 : ND2_165 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_164 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_163 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_54;

architecture SYN_STRUCTURAL of MUX21_54 is

   component ND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_54 port map( A => S, Y => SB);
   UND1 : ND2_162 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_161 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_160 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_53;

architecture SYN_STRUCTURAL of MUX21_53 is

   component ND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_53 port map( A => S, Y => SB);
   UND1 : ND2_159 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_158 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_157 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_52;

architecture SYN_STRUCTURAL of MUX21_52 is

   component ND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_52 port map( A => S, Y => SB);
   UND1 : ND2_156 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_155 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_154 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_51;

architecture SYN_STRUCTURAL of MUX21_51 is

   component ND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_51 port map( A => S, Y => SB);
   UND1 : ND2_153 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_152 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_151 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_50;

architecture SYN_STRUCTURAL of MUX21_50 is

   component ND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_50 port map( A => S, Y => SB);
   UND1 : ND2_150 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_149 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_148 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_49;

architecture SYN_STRUCTURAL of MUX21_49 is

   component ND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_49 port map( A => S, Y => SB);
   UND1 : ND2_147 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_146 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_145 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_48;

architecture SYN_STRUCTURAL of MUX21_48 is

   component ND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_48 port map( A => S, Y => SB);
   UND1 : ND2_144 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_143 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_142 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_47;

architecture SYN_STRUCTURAL of MUX21_47 is

   component ND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_47 port map( A => S, Y => SB);
   UND1 : ND2_141 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_140 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_139 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_46;

architecture SYN_STRUCTURAL of MUX21_46 is

   component ND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_46 port map( A => S, Y => SB);
   UND1 : ND2_138 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_137 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_136 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_45;

architecture SYN_STRUCTURAL of MUX21_45 is

   component ND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_45 port map( A => S, Y => SB);
   UND1 : ND2_135 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_134 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_133 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_44;

architecture SYN_STRUCTURAL of MUX21_44 is

   component ND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_44 port map( A => S, Y => SB);
   UND1 : ND2_132 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_131 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_130 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_43;

architecture SYN_STRUCTURAL of MUX21_43 is

   component ND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_43 port map( A => S, Y => SB);
   UND1 : ND2_129 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_128 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_127 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_42;

architecture SYN_STRUCTURAL of MUX21_42 is

   component ND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_42 port map( A => S, Y => SB);
   UND1 : ND2_126 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_125 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_124 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_41;

architecture SYN_STRUCTURAL of MUX21_41 is

   component ND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_41 port map( A => S, Y => SB);
   UND1 : ND2_123 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_122 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_121 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_40;

architecture SYN_STRUCTURAL of MUX21_40 is

   component ND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_40 port map( A => S, Y => SB);
   UND1 : ND2_120 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_119 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_118 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_39;

architecture SYN_STRUCTURAL of MUX21_39 is

   component ND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_39 port map( A => S, Y => SB);
   UND1 : ND2_117 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_116 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_115 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_38;

architecture SYN_STRUCTURAL of MUX21_38 is

   component ND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_38 port map( A => S, Y => SB);
   UND1 : ND2_114 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_113 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_112 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_37;

architecture SYN_STRUCTURAL of MUX21_37 is

   component ND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_37 port map( A => S, Y => SB);
   UND1 : ND2_111 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_110 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_109 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_36;

architecture SYN_STRUCTURAL of MUX21_36 is

   component ND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_36 port map( A => S, Y => SB);
   UND1 : ND2_108 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_107 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_106 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_35;

architecture SYN_STRUCTURAL of MUX21_35 is

   component ND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_35 port map( A => S, Y => SB);
   UND1 : ND2_105 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_104 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_103 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_34;

architecture SYN_STRUCTURAL of MUX21_34 is

   component ND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_34 port map( A => S, Y => SB);
   UND1 : ND2_102 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_101 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_100 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_33;

architecture SYN_STRUCTURAL of MUX21_33 is

   component ND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_33 port map( A => S, Y => SB);
   UND1 : ND2_99 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_98 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_97 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_27;

architecture SYN_STRUCTURAL of MUX21_27 is

   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_27 port map( A => S, Y => SB);
   UND1 : ND2_81 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_80 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_79 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_26;

architecture SYN_STRUCTURAL of MUX21_26 is

   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_26 port map( A => S, Y => SB);
   UND1 : ND2_78 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_77 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_76 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_25;

architecture SYN_STRUCTURAL of MUX21_25 is

   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_25 port map( A => S, Y => SB);
   UND1 : ND2_75 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_74 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_73 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_24;

architecture SYN_STRUCTURAL of MUX21_24 is

   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_24 port map( A => S, Y => SB);
   UND1 : ND2_72 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_71 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_70 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_23;

architecture SYN_STRUCTURAL of MUX21_23 is

   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_23 port map( A => S, Y => SB);
   UND1 : ND2_69 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_68 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_67 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_22;

architecture SYN_STRUCTURAL of MUX21_22 is

   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_22 port map( A => S, Y => SB);
   UND1 : ND2_66 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_65 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_64 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_21;

architecture SYN_STRUCTURAL of MUX21_21 is

   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_21 port map( A => S, Y => SB);
   UND1 : ND2_63 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_62 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_61 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_20;

architecture SYN_STRUCTURAL of MUX21_20 is

   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_20 port map( A => S, Y => SB);
   UND1 : ND2_60 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_59 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_58 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_19;

architecture SYN_STRUCTURAL of MUX21_19 is

   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_19 port map( A => S, Y => SB);
   UND1 : ND2_57 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_56 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_55 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_18;

architecture SYN_STRUCTURAL of MUX21_18 is

   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_18 port map( A => S, Y => SB);
   UND1 : ND2_54 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_53 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_52 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_17;

architecture SYN_STRUCTURAL of MUX21_17 is

   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_17 port map( A => S, Y => SB);
   UND1 : ND2_51 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_50 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_49 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_16;

architecture SYN_STRUCTURAL of MUX21_16 is

   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_16 port map( A => S, Y => SB);
   UND1 : ND2_48 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_47 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_46 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_15;

architecture SYN_STRUCTURAL of MUX21_15 is

   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_15 port map( A => S, Y => SB);
   UND1 : ND2_45 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_44 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_43 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_14;

architecture SYN_STRUCTURAL of MUX21_14 is

   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_14 port map( A => S, Y => SB);
   UND1 : ND2_42 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_41 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_40 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_13;

architecture SYN_STRUCTURAL of MUX21_13 is

   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_13 port map( A => S, Y => SB);
   UND1 : ND2_39 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_38 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_37 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_12;

architecture SYN_STRUCTURAL of MUX21_12 is

   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_12 port map( A => S, Y => SB);
   UND1 : ND2_36 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_35 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_34 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_11;

architecture SYN_STRUCTURAL of MUX21_11 is

   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_11 port map( A => S, Y => SB);
   UND1 : ND2_33 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_32 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_31 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_10;

architecture SYN_STRUCTURAL of MUX21_10 is

   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_10 port map( A => S, Y => SB);
   UND1 : ND2_30 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_29 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_28 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_9;

architecture SYN_STRUCTURAL of MUX21_9 is

   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_9 port map( A => S, Y => SB);
   UND1 : ND2_27 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_26 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_25 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_8;

architecture SYN_STRUCTURAL of MUX21_8 is

   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_8 port map( A => S, Y => SB);
   UND1 : ND2_24 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_23 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_22 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_7;

architecture SYN_STRUCTURAL of MUX21_7 is

   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_7 port map( A => S, Y => SB);
   UND1 : ND2_21 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_20 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_19 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_6;

architecture SYN_STRUCTURAL of MUX21_6 is

   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_6 port map( A => S, Y => SB);
   UND1 : ND2_18 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_17 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_16 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_5;

architecture SYN_STRUCTURAL of MUX21_5 is

   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_5 port map( A => S, Y => SB);
   UND1 : ND2_15 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_14 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_13 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_4;

architecture SYN_STRUCTURAL of MUX21_4 is

   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_4 port map( A => S, Y => SB);
   UND1 : ND2_12 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_11 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_10 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_3;

architecture SYN_STRUCTURAL of MUX21_3 is

   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_3 port map( A => S, Y => SB);
   UND1 : ND2_9 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_8 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_7 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_2;

architecture SYN_STRUCTURAL of MUX21_2 is

   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_2 port map( A => S, Y => SB);
   UND1 : ND2_6 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_5 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_4 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_1;

architecture SYN_STRUCTURAL of MUX21_1 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_1 port map( A => S, Y => SB);
   UND1 : ND2_3 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_2 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_6;

architecture SYN_struct of MUX21_GENERIC_NBIT4_6 is

   component MUX21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_24 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_23 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_22 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_21 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_5;

architecture SYN_struct of MUX21_GENERIC_NBIT4_5 is

   component MUX21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_20 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_19 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_18 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_17 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_4;

architecture SYN_struct of MUX21_GENERIC_NBIT4_4 is

   component MUX21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_16 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_15 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_14 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_13 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_3;

architecture SYN_struct of MUX21_GENERIC_NBIT4_3 is

   component MUX21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_12 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_11 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_10 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_9 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_2;

architecture SYN_struct of MUX21_GENERIC_NBIT4_2 is

   component MUX21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_8 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_7 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_6 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_5 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_1;

architecture SYN_struct of MUX21_GENERIC_NBIT4_1 is

   component MUX21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_4 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_3 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_2 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_1 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_6;

architecture SYN_STRUCTURAL of CSB_NBIT4_6 is

   component MUX21_GENERIC_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1000, n_1001 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1000);
   RCA1 : RCA_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1001);
   MUXCin : MUX21_GENERIC_NBIT4_6 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_5;

architecture SYN_STRUCTURAL of CSB_NBIT4_5 is

   component MUX21_GENERIC_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1002, n_1003 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1002);
   RCA1 : RCA_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1003);
   MUXCin : MUX21_GENERIC_NBIT4_5 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_4;

architecture SYN_STRUCTURAL of CSB_NBIT4_4 is

   component MUX21_GENERIC_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1004, n_1005 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1004);
   RCA1 : RCA_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1005);
   MUXCin : MUX21_GENERIC_NBIT4_4 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_3;

architecture SYN_STRUCTURAL of CSB_NBIT4_3 is

   component MUX21_GENERIC_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1006, n_1007 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1006);
   RCA1 : RCA_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1007);
   MUXCin : MUX21_GENERIC_NBIT4_3 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_2;

architecture SYN_STRUCTURAL of CSB_NBIT4_2 is

   component MUX21_GENERIC_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1008, n_1009 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1008);
   RCA1 : RCA_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1009);
   MUXCin : MUX21_GENERIC_NBIT4_2 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_1;

architecture SYN_STRUCTURAL of CSB_NBIT4_1 is

   component MUX21_GENERIC_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1010, n_1011 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1010);
   RCA1 : RCA_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1011);
   MUXCin : MUX21_GENERIC_NBIT4_1 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT6_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 downto 
         0);  Q : out std_logic_vector (5 downto 0));

end regFFD_NBIT6_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT6_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n19, n20, n21, n22, n23, n24, n25, n26, n27, 
      n28, n29, n30 : std_logic;

begin
   
   Q_reg_5_inst : DFFR_X1 port map( D => n1, CK => CK, RN => RESET, Q => Q(5), 
                           QN => n24);
   Q_reg_4_inst : DFFR_X1 port map( D => n2, CK => CK, RN => RESET, Q => Q(4), 
                           QN => n23);
   Q_reg_3_inst : DFFR_X1 port map( D => n3, CK => CK, RN => RESET, Q => Q(3), 
                           QN => n22);
   Q_reg_2_inst : DFFR_X1 port map( D => n4, CK => CK, RN => RESET, Q => Q(2), 
                           QN => n21);
   Q_reg_1_inst : DFFR_X1 port map( D => n5, CK => CK, RN => RESET, Q => Q(1), 
                           QN => n20);
   Q_reg_0_inst : DFFR_X1 port map( D => n6, CK => CK, RN => RESET, Q => Q(0), 
                           QN => n19);
   U2 : OAI21_X1 port map( B1 => n19, B2 => ENABLE, A => n30, ZN => n6);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n20, B2 => ENABLE, A => n29, ZN => n5);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n21, B2 => ENABLE, A => n28, ZN => n4);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => ENABLE, A => n27, ZN => n3);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n23, B2 => ENABLE, A => n26, ZN => n2);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n26);
   U12 : OAI21_X1 port map( B1 => n24, B2 => ENABLE, A => n25, ZN => n1);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n25);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_2 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_2;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25 
      : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n1, CK => CK, RN => RESET, Q => Q(4), 
                           QN => n20);
   Q_reg_3_inst : DFFR_X1 port map( D => n2, CK => CK, RN => RESET, Q => Q(3), 
                           QN => n19);
   Q_reg_2_inst : DFFR_X1 port map( D => n3, CK => CK, RN => RESET, Q => Q(2), 
                           QN => n18);
   Q_reg_1_inst : DFFR_X1 port map( D => n4, CK => CK, RN => RESET, Q => Q(1), 
                           QN => n17);
   Q_reg_0_inst : DFFR_X1 port map( D => n5, CK => CK, RN => RESET, Q => Q(0), 
                           QN => n16);
   U2 : OAI21_X1 port map( B1 => n16, B2 => ENABLE, A => n25, ZN => n5);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n25);
   U4 : OAI21_X1 port map( B1 => n17, B2 => ENABLE, A => n24, ZN => n4);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n24);
   U6 : OAI21_X1 port map( B1 => n18, B2 => ENABLE, A => n23, ZN => n3);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n23);
   U8 : OAI21_X1 port map( B1 => n19, B2 => ENABLE, A => n22, ZN => n2);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n22);
   U10 : OAI21_X1 port map( B1 => n20, B2 => ENABLE, A => n21, ZN => n1);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n21);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25 
      : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n1, CK => CK, RN => RESET, Q => Q(4), 
                           QN => n20);
   Q_reg_3_inst : DFFR_X1 port map( D => n2, CK => CK, RN => RESET, Q => Q(3), 
                           QN => n19);
   Q_reg_2_inst : DFFR_X1 port map( D => n3, CK => CK, RN => RESET, Q => Q(2), 
                           QN => n18);
   Q_reg_1_inst : DFFR_X1 port map( D => n4, CK => CK, RN => RESET, Q => Q(1), 
                           QN => n17);
   Q_reg_0_inst : DFFR_X1 port map( D => n5, CK => CK, RN => RESET, Q => Q(0), 
                           QN => n16);
   U2 : OAI21_X1 port map( B1 => n16, B2 => ENABLE, A => n25, ZN => n5);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n25);
   U4 : OAI21_X1 port map( B1 => n17, B2 => ENABLE, A => n24, ZN => n4);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n24);
   U6 : OAI21_X1 port map( B1 => n18, B2 => ENABLE, A => n23, ZN => n3);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n23);
   U8 : OAI21_X1 port map( B1 => n19, B2 => ENABLE, A => n22, ZN => n2);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n22);
   U10 : OAI21_X1 port map( B1 => n20, B2 => ENABLE, A => n21, ZN => n1);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n21);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_7 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_7;

architecture SYN_SYNC_BHV of FF_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n2, n3, n5, n6, n_1012 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1012);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n3, ZN => n2);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => n5, B2 => Q_port, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n5);
   U6 : INV_X1 port map( A => RESET, ZN => n3);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_6 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_6;

architecture SYN_SYNC_BHV of FF_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n2, n3, n5, n6, n_1013 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1013);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n3, ZN => n2);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => n5, B2 => Q_port, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n5);
   U6 : INV_X1 port map( A => RESET, ZN => n3);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_5 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_5;

architecture SYN_SYNC_BHV of FF_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n2, n3, n5, n6, n_1014 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1014);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n3, ZN => n2);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => n5, B2 => Q_port, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n5);
   U6 : INV_X1 port map( A => RESET, ZN => n3);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_4 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_4;

architecture SYN_SYNC_BHV of FF_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n3, n5, n6, n_1015 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : SDFF_X1 port map( D => RESET, SI => n3, SE => n6, CK => CLK, Q => 
                           Q_port, QN => n_1015);
   n3 <= '0';
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => n5, B2 => Q_port, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n5);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_3 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_3;

architecture SYN_SYNC_BHV of FF_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n2, n3, n5, n6, n_1016 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1016);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n3, ZN => n2);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => n5, B2 => Q_port, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n5);
   U6 : INV_X1 port map( A => RESET, ZN => n3);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_2 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_2;

architecture SYN_SYNC_BHV of FF_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n2, n3, n5, n6, n_1017 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1017);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n3, ZN => n2);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => n5, B2 => Q_port, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n5);
   U6 : INV_X1 port map( A => RESET, ZN => n3);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_4;

architecture SYN_struct of MUX21_GENERIC_NBIT32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   gen1_0 : MUX21_160 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   gen1_1 : MUX21_159 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   gen1_2 : MUX21_158 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   gen1_3 : MUX21_157 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   gen1_4 : MUX21_156 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   gen1_5 : MUX21_155 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   gen1_6 : MUX21_154 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   gen1_7 : MUX21_153 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   gen1_8 : MUX21_152 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   gen1_9 : MUX21_151 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   gen1_10 : MUX21_150 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   gen1_11 : MUX21_149 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   gen1_12 : MUX21_148 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   gen1_13 : MUX21_147 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   gen1_14 : MUX21_146 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   gen1_15 : MUX21_145 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   gen1_16 : MUX21_144 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   gen1_17 : MUX21_143 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   gen1_18 : MUX21_142 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   gen1_19 : MUX21_141 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   gen1_20 : MUX21_140 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   gen1_21 : MUX21_139 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   gen1_22 : MUX21_138 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   gen1_23 : MUX21_137 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   gen1_24 : MUX21_136 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   gen1_25 : MUX21_135 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   gen1_26 : MUX21_134 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   gen1_27 : MUX21_133 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   gen1_28 : MUX21_132 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   gen1_29 : MUX21_131 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   gen1_30 : MUX21_130 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   gen1_31 : MUX21_129 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_2;

architecture SYN_struct of MUX21_GENERIC_NBIT32_2 is

   component MUX21_65
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_66
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_67
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_68
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_69
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_70
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_71
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_72
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_73
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_74
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_75
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_76
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_77
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_78
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_79
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_80
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_81
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_82
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_83
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_84
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_85
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_86
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_87
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_88
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_89
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_90
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_91
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_92
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_93
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_94
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_95
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_96
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_96 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_95 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_94 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_93 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_92 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_91 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_90 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_89 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_88 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_87 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_86 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_85 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_84 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_83 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_82 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_81 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_80 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_79 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_78 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_77 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_76 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_75 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_74 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_73 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_72 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_71 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_70 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_69 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_68 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_67 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_66 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_65 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_3 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_3;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n99, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n99, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n99, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n99, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n98, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n98, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n98, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n98, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n99, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n98, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n98, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n97, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n99, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n97, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n97, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n97, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n99, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n97, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n97, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n97, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n98, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n98, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n97, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n97, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n98, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n97, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n97, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U7 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U8 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U9 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U10 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U11 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U12 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U13 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U14 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U15 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U16 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U17 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U18 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U19 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U20 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U21 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U22 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);
   U23 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U24 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U25 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U26 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U27 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U28 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U29 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U30 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U31 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U32 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U33 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U34 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U35 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U36 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U37 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U38 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U39 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U40 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U41 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U42 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U43 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U44 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U45 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U46 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U47 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U48 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U49 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U50 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U51 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U52 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U53 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U54 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U55 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U56 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U57 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U58 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U59 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U60 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U61 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U62 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U63 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U64 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U65 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U66 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U67 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U68 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_19 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_19;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_18 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_18;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_17 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_17;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_16 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_16;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_15 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_15;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_14 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_14;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_13 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_13;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_12 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_12;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_11 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_11;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U7 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U8 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U9 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U10 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U11 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U12 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U13 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U14 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U15 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U16 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U17 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U18 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U19 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U20 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U21 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U22 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U23 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U24 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U25 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U26 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U27 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U28 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U29 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U30 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U31 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U32 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U33 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U34 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U35 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U36 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U37 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U38 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U39 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U40 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U41 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U42 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U43 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U44 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U45 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U46 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U47 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U48 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U49 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U50 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U51 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U52 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_7 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_7;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U7 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U8 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U9 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U10 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U11 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U12 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U13 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U14 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U15 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U16 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U17 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U18 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U19 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U20 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U21 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U22 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U23 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U24 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U25 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U26 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U27 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U28 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U29 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U30 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U31 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U32 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U33 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U34 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U35 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U36 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);
   U37 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U38 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U39 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U40 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U41 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U42 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U43 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U44 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U45 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U46 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U47 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U48 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U49 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U50 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U51 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U52 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U53 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U54 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U55 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U56 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U57 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U58 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U59 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U60 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U61 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U62 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U63 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U64 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U65 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U66 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U67 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U68 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_6 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_6;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U7 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U8 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U9 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U10 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U11 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U12 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U13 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U14 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U15 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U16 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U17 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U18 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U19 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U20 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U21 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U22 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U23 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U24 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U25 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U26 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U27 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U28 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U29 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U30 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U31 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U32 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U33 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U34 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U35 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U36 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U37 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U38 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U39 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U40 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U41 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U42 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U43 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U44 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U45 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U46 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U47 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U48 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U49 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U50 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U51 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U52 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_5 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_5;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U52 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U53 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U54 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U55 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U56 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U57 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U58 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U59 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U60 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U61 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U62 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U63 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U64 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U65 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U66 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);
   U67 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U68 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_2 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_2;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);
   U53 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U55 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U57 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U59 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U61 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U63 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U65 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U67 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n131);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n130);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n129);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n128);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n127);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n126);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n125);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n124);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n123);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n122);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n121);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n120);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n119);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n118);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n117);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n116);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n115);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n114);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n113);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n112);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n111);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n110);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n109);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n108);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n107);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n106);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n105);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n104);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n103);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n102);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n101);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n100);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n100, B2 => ENABLE, A => n157, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n157);
   U7 : OAI21_X1 port map( B1 => n101, B2 => ENABLE, A => n156, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n156);
   U9 : OAI21_X1 port map( B1 => n102, B2 => ENABLE, A => n155, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n155);
   U11 : OAI21_X1 port map( B1 => n103, B2 => ENABLE, A => n153, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n153);
   U13 : OAI21_X1 port map( B1 => n104, B2 => ENABLE, A => n152, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n152);
   U15 : OAI21_X1 port map( B1 => n105, B2 => ENABLE, A => n151, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n151);
   U17 : OAI21_X1 port map( B1 => n106, B2 => ENABLE, A => n150, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n150);
   U19 : OAI21_X1 port map( B1 => n107, B2 => ENABLE, A => n149, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n149);
   U21 : OAI21_X1 port map( B1 => n108, B2 => ENABLE, A => n148, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n148);
   U23 : OAI21_X1 port map( B1 => n109, B2 => ENABLE, A => n147, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n147);
   U25 : OAI21_X1 port map( B1 => n110, B2 => ENABLE, A => n146, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n146);
   U27 : OAI21_X1 port map( B1 => n111, B2 => ENABLE, A => n145, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n145);
   U29 : OAI21_X1 port map( B1 => n112, B2 => ENABLE, A => n144, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n144);
   U31 : OAI21_X1 port map( B1 => n113, B2 => ENABLE, A => n142, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n142);
   U33 : OAI21_X1 port map( B1 => n114, B2 => ENABLE, A => n141, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n141);
   U35 : OAI21_X1 port map( B1 => n115, B2 => ENABLE, A => n140, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n140);
   U37 : OAI21_X1 port map( B1 => n116, B2 => ENABLE, A => n139, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n139);
   U39 : OAI21_X1 port map( B1 => n117, B2 => ENABLE, A => n138, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n138);
   U41 : OAI21_X1 port map( B1 => n118, B2 => ENABLE, A => n137, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n137);
   U43 : OAI21_X1 port map( B1 => n119, B2 => ENABLE, A => n136, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n136);
   U45 : OAI21_X1 port map( B1 => n120, B2 => ENABLE, A => n135, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n135);
   U47 : OAI21_X1 port map( B1 => n121, B2 => ENABLE, A => n134, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n134);
   U49 : OAI21_X1 port map( B1 => n122, B2 => ENABLE, A => n133, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n133);
   U51 : OAI21_X1 port map( B1 => n124, B2 => ENABLE, A => n162, ZN => n8);
   U52 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n162);
   U53 : OAI21_X1 port map( B1 => n125, B2 => ENABLE, A => n161, ZN => n7);
   U54 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n161);
   U55 : OAI21_X1 port map( B1 => n126, B2 => ENABLE, A => n160, ZN => n6);
   U56 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n160);
   U57 : OAI21_X1 port map( B1 => n127, B2 => ENABLE, A => n159, ZN => n5);
   U58 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n159);
   U59 : OAI21_X1 port map( B1 => n128, B2 => ENABLE, A => n158, ZN => n4);
   U60 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n158);
   U61 : OAI21_X1 port map( B1 => n129, B2 => ENABLE, A => n154, ZN => n3);
   U62 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n154);
   U63 : OAI21_X1 port map( B1 => n130, B2 => ENABLE, A => n143, ZN => n2);
   U64 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n143);
   U65 : OAI21_X1 port map( B1 => n131, B2 => ENABLE, A => n132, ZN => n1);
   U66 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n132);
   U67 : OAI21_X1 port map( B1 => n123, B2 => ENABLE, A => n163, ZN => n9);
   U68 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n163);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_28;

architecture SYN_STRUCTURAL of MUX21_28 is

   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_28 port map( A => S, Y => SB);
   UND1 : ND2_84 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_83 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_82 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_7;

architecture SYN_struct of MUX21_GENERIC_NBIT4_7 is

   component MUX21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_28 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_27 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_26 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_25 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_0;

architecture SYN_struct of MUX21_GENERIC_NBIT4_0 is

   component MUX21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_32 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_31 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_30 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_29 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_0;

architecture SYN_BEHAVIORAL of RCA_NBIT4_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_0 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_0;

architecture SYN_behave of P_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_7;

architecture SYN_STRUCTURAL of CSB_NBIT4_7 is

   component MUX21_GENERIC_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1018, n_1019 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1018);
   RCA1 : RCA_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1019);
   MUXCin : MUX21_GENERIC_NBIT4_7 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_0;

architecture SYN_STRUCTURAL of CSB_NBIT4_0 is

   component MUX21_GENERIC_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1020, n_1021 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1020);
   RCA1 : RCA_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1021);
   MUXCin : MUX21_GENERIC_NBIT4_0 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_42 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_42;

architecture SYN_arch of PG_42 is

   component P_42
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_42
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_42 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_42 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_0 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_0;

architecture SYN_arch of PG_0 is

   component P_0
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_43
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_43 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_0 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_0 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_0;

architecture SYN_behave of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_190;

architecture SYN_ARCH2 of ND2_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_STRUCTURAL of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component CSB_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_0 : CSB_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), S(2) 
                           => S(2), S(1) => S(1), S(0) => S(0));
   CSBI_1 : CSB_NBIT4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5), 
                           A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1) => 
                           B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), S(2) 
                           => S(6), S(1) => S(5), S(0) => S(4));
   CSBI_2 : CSB_NBIT4_6 port map( A(3) => A(11), A(2) => A(10), A(1) => A(9), 
                           A(0) => A(8), B(3) => B(11), B(2) => B(10), B(1) => 
                           B(9), B(0) => B(8), Ci => Ci(2), S(3) => S(11), S(2)
                           => S(10), S(1) => S(9), S(0) => S(8));
   CSBI_3 : CSB_NBIT4_5 port map( A(3) => A(15), A(2) => A(14), A(1) => A(13), 
                           A(0) => A(12), B(3) => B(15), B(2) => B(14), B(1) =>
                           B(13), B(0) => B(12), Ci => Ci(3), S(3) => S(15), 
                           S(2) => S(14), S(1) => S(13), S(0) => S(12));
   CSBI_4 : CSB_NBIT4_4 port map( A(3) => A(19), A(2) => A(18), A(1) => A(17), 
                           A(0) => A(16), B(3) => B(19), B(2) => B(18), B(1) =>
                           B(17), B(0) => B(16), Ci => Ci(4), S(3) => S(19), 
                           S(2) => S(18), S(1) => S(17), S(0) => S(16));
   CSBI_5 : CSB_NBIT4_3 port map( A(3) => A(23), A(2) => A(22), A(1) => A(21), 
                           A(0) => A(20), B(3) => B(23), B(2) => B(22), B(1) =>
                           B(21), B(0) => B(20), Ci => Ci(5), S(3) => S(23), 
                           S(2) => S(22), S(1) => S(21), S(0) => S(20));
   CSBI_6 : CSB_NBIT4_2 port map( A(3) => A(27), A(2) => A(26), A(1) => A(25), 
                           A(0) => A(24), B(3) => B(27), B(2) => B(26), B(1) =>
                           B(25), B(0) => B(24), Ci => Ci(6), S(3) => S(27), 
                           S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CSBI_7 : CSB_NBIT4_1 port map( A(3) => A(31), A(2) => A(30), A(1) => A(29), 
                           A(0) => A(28), B(3) => B(31), B(2) => B(30), B(1) =>
                           B(29), B(0) => B(28), Ci => Ci(7), S(3) => S(31), 
                           S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_arch of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_44
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_45
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_46
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_47
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_1
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_2
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_48
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_49
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_3
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_4
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_5
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_50
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_6
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_7
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_8
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_9
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_10
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_11
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_12
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_51
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_13
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_14
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_15
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_16
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_17
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_18
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_19
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_20
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_21
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_22
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_23
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_24
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_25
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_26
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_27
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_28
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_29
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_30
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_31
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_32
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_33
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_34
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_35
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_36
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_37
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_38
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_39
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_40
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_41
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_42
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_52
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_0
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_0
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port,
      Co_2_port, Co_1_port, Co_0_port, gi_32_4_port, gi_32_3_port, gi_32_2_port
      , gi_32_1_port, gi_32_0_port, gi_31_0_port, gi_30_0_port, gi_29_0_port, 
      gi_28_4_port, gi_28_2_port, gi_28_1_port, gi_28_0_port, gi_27_0_port, 
      gi_26_0_port, gi_25_0_port, gi_24_3_port, gi_24_2_port, gi_24_1_port, 
      gi_24_0_port, gi_23_0_port, gi_22_0_port, gi_21_0_port, gi_20_2_port, 
      gi_20_1_port, gi_20_0_port, gi_19_0_port, gi_18_0_port, gi_17_0_port, 
      gi_16_3_port, gi_16_2_port, gi_16_1_port, gi_16_0_port, gi_15_0_port, 
      gi_14_0_port, gi_13_0_port, gi_12_2_port, gi_12_1_port, gi_12_0_port, 
      gi_11_0_port, gi_10_0_port, gi_9_0_port, gi_8_2_port, gi_8_1_port, 
      gi_8_0_port, gi_7_0_port, gi_6_0_port, gi_5_0_port, gi_4_1_port, 
      gi_4_0_port, gi_3_0_port, gi_2_1_port, gi_2_0_port, gi_1_0_port, 
      gi_0_0_port, pi_32_4_port, pi_32_3_port, pi_32_2_port, pi_32_1_port, 
      pi_32_0_port, pi_31_0_port, pi_30_0_port, pi_29_0_port, pi_28_4_port, 
      pi_28_2_port, pi_28_1_port, pi_28_0_port, pi_27_0_port, pi_26_0_port, 
      pi_25_0_port, pi_24_3_port, pi_24_2_port, pi_24_1_port, pi_24_0_port, 
      pi_23_0_port, pi_22_0_port, pi_21_0_port, pi_20_2_port, pi_20_1_port, 
      pi_20_0_port, pi_19_0_port, pi_18_0_port, pi_17_0_port, pi_16_3_port, 
      pi_16_2_port, pi_16_1_port, pi_16_0_port, pi_15_0_port, pi_14_0_port, 
      pi_13_0_port, pi_12_2_port, pi_12_1_port, pi_12_0_port, pi_11_0_port, 
      pi_10_0_port, pi_9_0_port, pi_8_2_port, pi_8_1_port, pi_8_0_port, 
      pi_7_0_port, pi_6_0_port, pi_5_0_port, pi_4_1_port, pi_4_0_port, 
      pi_3_0_port, pi_2_0_port, pi_0_0_port, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   X_Logic0_port <= '0';
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => pi_9_0_port);
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => pi_8_0_port);
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => pi_7_0_port);
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => pi_6_0_port);
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => pi_5_0_port);
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => pi_4_0_port);
   U40 : XOR2_X1 port map( A => B(2), B => A(2), Z => pi_3_0_port);
   U41 : XOR2_X1 port map( A => B(31), B => A(31), Z => pi_32_0_port);
   U42 : XOR2_X1 port map( A => B(30), B => A(30), Z => pi_31_0_port);
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => pi_30_0_port);
   U44 : XOR2_X1 port map( A => B(1), B => A(1), Z => pi_2_0_port);
   U45 : XOR2_X1 port map( A => B(28), B => A(28), Z => pi_29_0_port);
   U46 : XOR2_X1 port map( A => B(27), B => A(27), Z => pi_28_0_port);
   U47 : XOR2_X1 port map( A => B(26), B => A(26), Z => pi_27_0_port);
   U48 : XOR2_X1 port map( A => B(25), B => A(25), Z => pi_26_0_port);
   U49 : XOR2_X1 port map( A => B(24), B => A(24), Z => pi_25_0_port);
   U50 : XOR2_X1 port map( A => B(23), B => A(23), Z => pi_24_0_port);
   U51 : XOR2_X1 port map( A => B(22), B => A(22), Z => pi_23_0_port);
   U52 : XOR2_X1 port map( A => B(21), B => A(21), Z => pi_22_0_port);
   U53 : XOR2_X1 port map( A => B(20), B => A(20), Z => pi_21_0_port);
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => pi_20_0_port);
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => pi_19_0_port);
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => pi_18_0_port);
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => pi_17_0_port);
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => pi_16_0_port);
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => pi_15_0_port);
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => pi_14_0_port);
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => pi_13_0_port);
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => pi_12_0_port);
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => pi_11_0_port);
   U64 : XOR2_X1 port map( A => B(9), B => A(9), Z => pi_10_0_port);
   U65 : XOR2_X1 port map( A => B(0), B => A(0), Z => pi_0_0_port);
   g_port0_0_1 : G_0 port map( G1 => gi_0_0_port, P => pi_0_0_port, G2 => Cin, 
                           Co => gi_1_0_port);
   pg_port2_1_1 : PG_0 port map( G1 => gi_1_0_port, P1 => X_Logic0_port, G2 => 
                           gi_0_0_port, P2 => pi_0_0_port, gout => n_1022, pout
                           => n_1023);
   g_port1_1_2 : G_52 port map( G1 => gi_2_0_port, P => pi_2_0_port, G2 => 
                           gi_1_0_port, Co => gi_2_1_port);
   pg_port2_1_3 : PG_42 port map( G1 => gi_3_0_port, P1 => pi_3_0_port, G2 => 
                           gi_2_0_port, P2 => pi_2_0_port, gout => n_1024, pout
                           => n_1025);
   pg_port2_1_4 : PG_41 port map( G1 => gi_4_0_port, P1 => pi_4_0_port, G2 => 
                           gi_3_0_port, P2 => pi_3_0_port, gout => gi_4_1_port,
                           pout => pi_4_1_port);
   pg_port2_1_5 : PG_40 port map( G1 => gi_5_0_port, P1 => pi_5_0_port, G2 => 
                           gi_4_0_port, P2 => pi_4_0_port, gout => n_1026, pout
                           => n_1027);
   pg_port2_1_6 : PG_39 port map( G1 => gi_6_0_port, P1 => pi_6_0_port, G2 => 
                           gi_5_0_port, P2 => pi_5_0_port, gout => n_1028, pout
                           => n_1029);
   pg_port2_1_7 : PG_38 port map( G1 => gi_7_0_port, P1 => pi_7_0_port, G2 => 
                           gi_6_0_port, P2 => pi_6_0_port, gout => n_1030, pout
                           => n_1031);
   pg_port2_1_8 : PG_37 port map( G1 => gi_8_0_port, P1 => pi_8_0_port, G2 => 
                           gi_7_0_port, P2 => pi_7_0_port, gout => gi_8_1_port,
                           pout => pi_8_1_port);
   pg_port2_1_9 : PG_36 port map( G1 => gi_9_0_port, P1 => pi_9_0_port, G2 => 
                           gi_8_0_port, P2 => pi_8_0_port, gout => n_1032, pout
                           => n_1033);
   pg_port2_1_10 : PG_35 port map( G1 => gi_10_0_port, P1 => pi_10_0_port, G2 
                           => gi_9_0_port, P2 => pi_9_0_port, gout => n_1034, 
                           pout => n_1035);
   pg_port2_1_11 : PG_34 port map( G1 => gi_11_0_port, P1 => pi_11_0_port, G2 
                           => gi_10_0_port, P2 => pi_10_0_port, gout => n_1036,
                           pout => n_1037);
   pg_port2_1_12 : PG_33 port map( G1 => gi_12_0_port, P1 => pi_12_0_port, G2 
                           => gi_11_0_port, P2 => pi_11_0_port, gout => 
                           gi_12_1_port, pout => pi_12_1_port);
   pg_port2_1_13 : PG_32 port map( G1 => gi_13_0_port, P1 => pi_13_0_port, G2 
                           => gi_12_0_port, P2 => pi_12_0_port, gout => n_1038,
                           pout => n_1039);
   pg_port2_1_14 : PG_31 port map( G1 => gi_14_0_port, P1 => pi_14_0_port, G2 
                           => gi_13_0_port, P2 => pi_13_0_port, gout => n_1040,
                           pout => n_1041);
   pg_port2_1_15 : PG_30 port map( G1 => gi_15_0_port, P1 => pi_15_0_port, G2 
                           => gi_14_0_port, P2 => pi_14_0_port, gout => n_1042,
                           pout => n_1043);
   pg_port2_1_16 : PG_29 port map( G1 => gi_16_0_port, P1 => pi_16_0_port, G2 
                           => gi_15_0_port, P2 => pi_15_0_port, gout => 
                           gi_16_1_port, pout => pi_16_1_port);
   pg_port2_1_17 : PG_28 port map( G1 => gi_17_0_port, P1 => pi_17_0_port, G2 
                           => gi_16_0_port, P2 => pi_16_0_port, gout => n_1044,
                           pout => n_1045);
   pg_port2_1_18 : PG_27 port map( G1 => gi_18_0_port, P1 => pi_18_0_port, G2 
                           => gi_17_0_port, P2 => pi_17_0_port, gout => n_1046,
                           pout => n_1047);
   pg_port2_1_19 : PG_26 port map( G1 => gi_19_0_port, P1 => pi_19_0_port, G2 
                           => gi_18_0_port, P2 => pi_18_0_port, gout => n_1048,
                           pout => n_1049);
   pg_port2_1_20 : PG_25 port map( G1 => gi_20_0_port, P1 => pi_20_0_port, G2 
                           => gi_19_0_port, P2 => pi_19_0_port, gout => 
                           gi_20_1_port, pout => pi_20_1_port);
   pg_port2_1_21 : PG_24 port map( G1 => gi_21_0_port, P1 => pi_21_0_port, G2 
                           => gi_20_0_port, P2 => pi_20_0_port, gout => n_1050,
                           pout => n_1051);
   pg_port2_1_22 : PG_23 port map( G1 => gi_22_0_port, P1 => pi_22_0_port, G2 
                           => gi_21_0_port, P2 => pi_21_0_port, gout => n_1052,
                           pout => n_1053);
   pg_port2_1_23 : PG_22 port map( G1 => gi_23_0_port, P1 => pi_23_0_port, G2 
                           => gi_22_0_port, P2 => pi_22_0_port, gout => n_1054,
                           pout => n_1055);
   pg_port2_1_24 : PG_21 port map( G1 => gi_24_0_port, P1 => pi_24_0_port, G2 
                           => gi_23_0_port, P2 => pi_23_0_port, gout => 
                           gi_24_1_port, pout => pi_24_1_port);
   pg_port2_1_25 : PG_20 port map( G1 => gi_25_0_port, P1 => pi_25_0_port, G2 
                           => gi_24_0_port, P2 => pi_24_0_port, gout => n_1056,
                           pout => n_1057);
   pg_port2_1_26 : PG_19 port map( G1 => gi_26_0_port, P1 => pi_26_0_port, G2 
                           => gi_25_0_port, P2 => pi_25_0_port, gout => n_1058,
                           pout => n_1059);
   pg_port2_1_27 : PG_18 port map( G1 => gi_27_0_port, P1 => pi_27_0_port, G2 
                           => gi_26_0_port, P2 => pi_26_0_port, gout => n_1060,
                           pout => n_1061);
   pg_port2_1_28 : PG_17 port map( G1 => gi_28_0_port, P1 => pi_28_0_port, G2 
                           => gi_27_0_port, P2 => pi_27_0_port, gout => 
                           gi_28_1_port, pout => pi_28_1_port);
   pg_port2_1_29 : PG_16 port map( G1 => gi_29_0_port, P1 => pi_29_0_port, G2 
                           => gi_28_0_port, P2 => pi_28_0_port, gout => n_1062,
                           pout => n_1063);
   pg_port2_1_30 : PG_15 port map( G1 => gi_30_0_port, P1 => pi_30_0_port, G2 
                           => gi_29_0_port, P2 => pi_29_0_port, gout => n_1064,
                           pout => n_1065);
   pg_port2_1_31 : PG_14 port map( G1 => gi_31_0_port, P1 => pi_31_0_port, G2 
                           => gi_30_0_port, P2 => pi_30_0_port, gout => n_1066,
                           pout => n_1067);
   pg_port2_1_32 : PG_13 port map( G1 => gi_32_0_port, P1 => pi_32_0_port, G2 
                           => gi_31_0_port, P2 => pi_31_0_port, gout => 
                           gi_32_1_port, pout => pi_32_1_port);
   g_port_0 : G_51 port map( G1 => gi_4_1_port, P => pi_4_1_port, G2 => 
                           gi_2_1_port, Co => Co_0_port);
   pg_port2_0_1_2 : PG_12 port map( G1 => gi_8_1_port, P1 => pi_8_1_port, G2 =>
                           gi_4_1_port, P2 => pi_4_1_port, gout => gi_8_2_port,
                           pout => pi_8_2_port);
   pg_port2_0_2_3 : PG_11 port map( G1 => gi_12_1_port, P1 => pi_12_1_port, G2 
                           => gi_8_1_port, P2 => pi_8_1_port, gout => 
                           gi_12_2_port, pout => pi_12_2_port);
   pg_port2_0_3_4 : PG_10 port map( G1 => gi_16_1_port, P1 => pi_16_1_port, G2 
                           => gi_12_1_port, P2 => pi_12_1_port, gout => 
                           gi_16_2_port, pout => pi_16_2_port);
   pg_port2_0_4_5 : PG_9 port map( G1 => gi_20_1_port, P1 => pi_20_1_port, G2 
                           => gi_16_1_port, P2 => pi_16_1_port, gout => 
                           gi_20_2_port, pout => pi_20_2_port);
   pg_port2_0_5_6 : PG_8 port map( G1 => gi_24_1_port, P1 => pi_24_1_port, G2 
                           => gi_20_1_port, P2 => pi_20_1_port, gout => 
                           gi_24_2_port, pout => pi_24_2_port);
   pg_port2_0_6_7 : PG_7 port map( G1 => gi_28_1_port, P1 => pi_28_1_port, G2 
                           => gi_24_1_port, P2 => pi_24_1_port, gout => 
                           gi_28_2_port, pout => pi_28_2_port);
   pg_port2_0_7_8 : PG_6 port map( G1 => gi_32_1_port, P1 => pi_32_1_port, G2 
                           => gi_28_1_port, P2 => pi_28_1_port, gout => 
                           gi_32_2_port, pout => pi_32_2_port);
   g_port_1_2 : G_50 port map( G1 => gi_8_2_port, P => pi_8_2_port, G2 => 
                           Co_0_port, Co => Co_1_port);
   pg_port2_1_1_4 : PG_5 port map( G1 => gi_16_2_port, P1 => pi_16_2_port, G2 
                           => gi_12_2_port, P2 => pi_12_2_port, gout => 
                           gi_16_3_port, pout => pi_16_3_port);
   pg_port2_1_2_6 : PG_4 port map( G1 => gi_24_2_port, P1 => pi_24_2_port, G2 
                           => gi_20_2_port, P2 => pi_20_2_port, gout => 
                           gi_24_3_port, pout => pi_24_3_port);
   pg_port2_1_3_8 : PG_3 port map( G1 => gi_32_2_port, P1 => pi_32_2_port, G2 
                           => gi_28_2_port, P2 => pi_28_2_port, gout => 
                           gi_32_3_port, pout => pi_32_3_port);
   g_port_2_3 : G_49 port map( G1 => gi_12_2_port, P => pi_12_2_port, G2 => 
                           Co_1_port, Co => Co_2_port);
   g_port_2_4 : G_48 port map( G1 => gi_16_3_port, P => pi_16_3_port, G2 => 
                           Co_1_port, Co => Co_3_port);
   pg_port2_2_1_7 : PG_2 port map( G1 => gi_28_2_port, P1 => pi_28_2_port, G2 
                           => gi_24_3_port, P2 => pi_24_3_port, gout => 
                           gi_28_4_port, pout => pi_28_4_port);
   pg_port2_2_1_8 : PG_1 port map( G1 => gi_32_3_port, P1 => pi_32_3_port, G2 
                           => gi_24_3_port, P2 => pi_24_3_port, gout => 
                           gi_32_4_port, pout => pi_32_4_port);
   g_port_3_5 : G_47 port map( G1 => gi_20_2_port, P => pi_20_2_port, G2 => 
                           Co_3_port, Co => Co_4_port);
   g_port_3_6 : G_46 port map( G1 => gi_24_3_port, P => pi_24_3_port, G2 => 
                           Co_3_port, Co => Co_5_port);
   g_port_3_7 : G_45 port map( G1 => gi_28_4_port, P => pi_28_4_port, G2 => 
                           Co_3_port, Co => Co_6_port);
   g_port_3_8 : G_44 port map( G1 => gi_32_4_port, P => pi_32_4_port, G2 => 
                           Co_3_port, Co => Co_7_port);
   U2 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => gi_32_0_port);
   U3 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => gi_16_0_port);
   U4 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => gi_15_0_port);
   U5 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => gi_24_0_port);
   U6 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => gi_23_0_port);
   U7 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => gi_20_0_port);
   U8 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => gi_19_0_port);
   U9 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => gi_0_0_port);
   U10 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => gi_4_0_port);
   U11 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => gi_3_0_port);
   U12 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => gi_8_0_port);
   U13 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => gi_7_0_port);
   U14 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => gi_12_0_port);
   U15 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => gi_11_0_port);
   U16 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => gi_28_0_port);
   U17 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => gi_27_0_port);
   U18 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => gi_31_0_port);
   U19 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => gi_2_0_port);
   U20 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => gi_5_0_port);
   U21 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => gi_6_0_port);
   U22 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => gi_9_0_port);
   U23 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => gi_10_0_port);
   U24 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => gi_13_0_port);
   U25 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => gi_14_0_port);
   U26 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => gi_17_0_port);
   U27 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => gi_18_0_port);
   U28 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => gi_21_0_port);
   U29 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => gi_22_0_port);
   U30 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => gi_25_0_port);
   U31 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => gi_26_0_port);
   U32 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => gi_29_0_port);
   U33 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => gi_30_0_port);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_rbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_rbsh_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal MR_int_1_31_port, MR_int_1_30_port, MR_int_1_29_port, 
      MR_int_1_28_port, MR_int_1_27_port, MR_int_1_26_port, MR_int_1_25_port, 
      MR_int_1_24_port, MR_int_1_23_port, MR_int_1_22_port, MR_int_1_21_port, 
      MR_int_1_20_port, MR_int_1_19_port, MR_int_1_18_port, MR_int_1_17_port, 
      MR_int_1_16_port, MR_int_1_15_port, MR_int_1_14_port, MR_int_1_13_port, 
      MR_int_1_12_port, MR_int_1_11_port, MR_int_1_10_port, MR_int_1_9_port, 
      MR_int_1_8_port, MR_int_1_7_port, MR_int_1_6_port, MR_int_1_5_port, 
      MR_int_1_4_port, MR_int_1_3_port, MR_int_1_2_port, MR_int_1_1_port, 
      MR_int_1_0_port, MR_int_2_31_port, MR_int_2_30_port, MR_int_2_29_port, 
      MR_int_2_28_port, MR_int_2_27_port, MR_int_2_26_port, MR_int_2_25_port, 
      MR_int_2_24_port, MR_int_2_23_port, MR_int_2_22_port, MR_int_2_21_port, 
      MR_int_2_20_port, MR_int_2_19_port, MR_int_2_18_port, MR_int_2_17_port, 
      MR_int_2_16_port, MR_int_2_15_port, MR_int_2_14_port, MR_int_2_13_port, 
      MR_int_2_12_port, MR_int_2_11_port, MR_int_2_10_port, MR_int_2_9_port, 
      MR_int_2_8_port, MR_int_2_7_port, MR_int_2_6_port, MR_int_2_5_port, 
      MR_int_2_4_port, MR_int_2_3_port, MR_int_2_2_port, MR_int_2_1_port, 
      MR_int_2_0_port, MR_int_3_31_port, MR_int_3_30_port, MR_int_3_29_port, 
      MR_int_3_28_port, MR_int_3_27_port, MR_int_3_26_port, MR_int_3_25_port, 
      MR_int_3_24_port, MR_int_3_23_port, MR_int_3_22_port, MR_int_3_21_port, 
      MR_int_3_20_port, MR_int_3_19_port, MR_int_3_18_port, MR_int_3_17_port, 
      MR_int_3_16_port, MR_int_3_15_port, MR_int_3_14_port, MR_int_3_13_port, 
      MR_int_3_12_port, MR_int_3_11_port, MR_int_3_10_port, MR_int_3_9_port, 
      MR_int_3_8_port, MR_int_3_7_port, MR_int_3_6_port, MR_int_3_5_port, 
      MR_int_3_4_port, MR_int_3_3_port, MR_int_3_2_port, MR_int_3_1_port, 
      MR_int_3_0_port, MR_int_4_31_port, MR_int_4_30_port, MR_int_4_29_port, 
      MR_int_4_28_port, MR_int_4_27_port, MR_int_4_26_port, MR_int_4_25_port, 
      MR_int_4_24_port, MR_int_4_23_port, MR_int_4_22_port, MR_int_4_21_port, 
      MR_int_4_20_port, MR_int_4_19_port, MR_int_4_18_port, MR_int_4_17_port, 
      MR_int_4_16_port, MR_int_4_15_port, MR_int_4_14_port, MR_int_4_13_port, 
      MR_int_4_12_port, MR_int_4_11_port, MR_int_4_10_port, MR_int_4_9_port, 
      MR_int_4_8_port, MR_int_4_7_port, MR_int_4_6_port, MR_int_4_5_port, 
      MR_int_4_4_port, MR_int_4_3_port, MR_int_4_2_port, MR_int_4_1_port, 
      MR_int_4_0_port, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => MR_int_4_31_port, B => MR_int_4_15_port, S 
                           => n18, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => MR_int_4_30_port, B => MR_int_4_14_port, S 
                           => n18, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => MR_int_4_29_port, B => MR_int_4_13_port, S 
                           => n18, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => MR_int_4_28_port, B => MR_int_4_12_port, S 
                           => n18, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => MR_int_4_27_port, B => MR_int_4_11_port, S 
                           => n18, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => MR_int_4_26_port, B => MR_int_4_10_port, S 
                           => n18, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => MR_int_4_25_port, B => MR_int_4_9_port, S 
                           => n18, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => MR_int_4_24_port, B => MR_int_4_8_port, S 
                           => n18, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => MR_int_4_23_port, B => MR_int_4_7_port, S 
                           => n18, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => MR_int_4_22_port, B => MR_int_4_6_port, S 
                           => n18, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => MR_int_4_21_port, B => MR_int_4_5_port, S 
                           => n16, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => MR_int_4_20_port, B => MR_int_4_4_port, S 
                           => n16, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => MR_int_4_19_port, B => MR_int_4_3_port, S 
                           => n16, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => MR_int_4_18_port, B => MR_int_4_2_port, S 
                           => n16, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => MR_int_4_17_port, B => MR_int_4_1_port, S 
                           => n16, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => MR_int_4_16_port, B => MR_int_4_0_port, S 
                           => n16, Z => B(16));
   M1_4_15 : MUX2_X1 port map( A => MR_int_4_15_port, B => MR_int_4_31_port, S 
                           => n16, Z => B(15));
   M1_4_14 : MUX2_X1 port map( A => MR_int_4_14_port, B => MR_int_4_30_port, S 
                           => n16, Z => B(14));
   M1_4_13 : MUX2_X1 port map( A => MR_int_4_13_port, B => MR_int_4_29_port, S 
                           => n16, Z => B(13));
   M1_4_12 : MUX2_X1 port map( A => MR_int_4_12_port, B => MR_int_4_28_port, S 
                           => n16, Z => B(12));
   M1_4_11 : MUX2_X1 port map( A => MR_int_4_11_port, B => MR_int_4_27_port, S 
                           => n16, Z => B(11));
   M1_4_10 : MUX2_X1 port map( A => MR_int_4_10_port, B => MR_int_4_26_port, S 
                           => n17, Z => B(10));
   M1_4_9 : MUX2_X1 port map( A => MR_int_4_9_port, B => MR_int_4_25_port, S =>
                           n17, Z => B(9));
   M1_4_8 : MUX2_X1 port map( A => MR_int_4_8_port, B => MR_int_4_24_port, S =>
                           n17, Z => B(8));
   M1_4_7 : MUX2_X1 port map( A => MR_int_4_7_port, B => MR_int_4_23_port, S =>
                           n17, Z => B(7));
   M1_4_6 : MUX2_X1 port map( A => MR_int_4_6_port, B => MR_int_4_22_port, S =>
                           n17, Z => B(6));
   M1_4_5 : MUX2_X1 port map( A => MR_int_4_5_port, B => MR_int_4_21_port, S =>
                           n17, Z => B(5));
   M1_4_4 : MUX2_X1 port map( A => MR_int_4_4_port, B => MR_int_4_20_port, S =>
                           n17, Z => B(4));
   M1_4_3 : MUX2_X1 port map( A => MR_int_4_3_port, B => MR_int_4_19_port, S =>
                           n17, Z => B(3));
   M1_4_2 : MUX2_X1 port map( A => MR_int_4_2_port, B => MR_int_4_18_port, S =>
                           n17, Z => B(2));
   M1_4_1 : MUX2_X1 port map( A => MR_int_4_1_port, B => MR_int_4_17_port, S =>
                           n17, Z => B(1));
   M1_4_0 : MUX2_X1 port map( A => MR_int_4_0_port, B => MR_int_4_16_port, S =>
                           n17, Z => B(0));
   M1_3_31_0 : MUX2_X1 port map( A => MR_int_3_31_port, B => MR_int_3_7_port, S
                           => n15, Z => MR_int_4_31_port);
   M1_3_30_0 : MUX2_X1 port map( A => MR_int_3_30_port, B => MR_int_3_6_port, S
                           => n15, Z => MR_int_4_30_port);
   M1_3_29_0 : MUX2_X1 port map( A => MR_int_3_29_port, B => MR_int_3_5_port, S
                           => n15, Z => MR_int_4_29_port);
   M1_3_28_0 : MUX2_X1 port map( A => MR_int_3_28_port, B => MR_int_3_4_port, S
                           => n15, Z => MR_int_4_28_port);
   M1_3_27_0 : MUX2_X1 port map( A => MR_int_3_27_port, B => MR_int_3_3_port, S
                           => n15, Z => MR_int_4_27_port);
   M1_3_26_0 : MUX2_X1 port map( A => MR_int_3_26_port, B => MR_int_3_2_port, S
                           => n15, Z => MR_int_4_26_port);
   M1_3_25_0 : MUX2_X1 port map( A => MR_int_3_25_port, B => MR_int_3_1_port, S
                           => n15, Z => MR_int_4_25_port);
   M1_3_24_0 : MUX2_X1 port map( A => MR_int_3_24_port, B => MR_int_3_0_port, S
                           => n15, Z => MR_int_4_24_port);
   M1_3_23_0 : MUX2_X1 port map( A => MR_int_3_23_port, B => MR_int_3_31_port, 
                           S => n15, Z => MR_int_4_23_port);
   M1_3_22_0 : MUX2_X1 port map( A => MR_int_3_22_port, B => MR_int_3_30_port, 
                           S => n15, Z => MR_int_4_22_port);
   M1_3_21_0 : MUX2_X1 port map( A => MR_int_3_21_port, B => MR_int_3_29_port, 
                           S => n14, Z => MR_int_4_21_port);
   M1_3_20_0 : MUX2_X1 port map( A => MR_int_3_20_port, B => MR_int_3_28_port, 
                           S => n14, Z => MR_int_4_20_port);
   M1_3_19_0 : MUX2_X1 port map( A => MR_int_3_19_port, B => MR_int_3_27_port, 
                           S => n14, Z => MR_int_4_19_port);
   M1_3_18_0 : MUX2_X1 port map( A => MR_int_3_18_port, B => MR_int_3_26_port, 
                           S => n14, Z => MR_int_4_18_port);
   M1_3_17_0 : MUX2_X1 port map( A => MR_int_3_17_port, B => MR_int_3_25_port, 
                           S => n14, Z => MR_int_4_17_port);
   M1_3_16_0 : MUX2_X1 port map( A => MR_int_3_16_port, B => MR_int_3_24_port, 
                           S => n14, Z => MR_int_4_16_port);
   M1_3_15_0 : MUX2_X1 port map( A => MR_int_3_15_port, B => MR_int_3_23_port, 
                           S => n14, Z => MR_int_4_15_port);
   M1_3_14_0 : MUX2_X1 port map( A => MR_int_3_14_port, B => MR_int_3_22_port, 
                           S => n14, Z => MR_int_4_14_port);
   M1_3_13_0 : MUX2_X1 port map( A => MR_int_3_13_port, B => MR_int_3_21_port, 
                           S => n14, Z => MR_int_4_13_port);
   M1_3_12_0 : MUX2_X1 port map( A => MR_int_3_12_port, B => MR_int_3_20_port, 
                           S => n14, Z => MR_int_4_12_port);
   M1_3_11_0 : MUX2_X1 port map( A => MR_int_3_11_port, B => MR_int_3_19_port, 
                           S => n14, Z => MR_int_4_11_port);
   M1_3_10_0 : MUX2_X1 port map( A => MR_int_3_10_port, B => MR_int_3_18_port, 
                           S => n13, Z => MR_int_4_10_port);
   M1_3_9_0 : MUX2_X1 port map( A => MR_int_3_9_port, B => MR_int_3_17_port, S 
                           => n13, Z => MR_int_4_9_port);
   M1_3_8_0 : MUX2_X1 port map( A => MR_int_3_8_port, B => MR_int_3_16_port, S 
                           => n13, Z => MR_int_4_8_port);
   M1_3_7 : MUX2_X1 port map( A => MR_int_3_7_port, B => MR_int_3_15_port, S =>
                           n13, Z => MR_int_4_7_port);
   M1_3_6 : MUX2_X1 port map( A => MR_int_3_6_port, B => MR_int_3_14_port, S =>
                           n13, Z => MR_int_4_6_port);
   M1_3_5 : MUX2_X1 port map( A => MR_int_3_5_port, B => MR_int_3_13_port, S =>
                           n13, Z => MR_int_4_5_port);
   M1_3_4 : MUX2_X1 port map( A => MR_int_3_4_port, B => MR_int_3_12_port, S =>
                           n13, Z => MR_int_4_4_port);
   M1_3_3 : MUX2_X1 port map( A => MR_int_3_3_port, B => MR_int_3_11_port, S =>
                           n13, Z => MR_int_4_3_port);
   M1_3_2 : MUX2_X1 port map( A => MR_int_3_2_port, B => MR_int_3_10_port, S =>
                           n13, Z => MR_int_4_2_port);
   M1_3_1 : MUX2_X1 port map( A => MR_int_3_1_port, B => MR_int_3_9_port, S => 
                           n13, Z => MR_int_4_1_port);
   M1_3_0 : MUX2_X1 port map( A => MR_int_3_0_port, B => MR_int_3_8_port, S => 
                           n13, Z => MR_int_4_0_port);
   M1_2_31_0 : MUX2_X1 port map( A => MR_int_2_31_port, B => MR_int_2_3_port, S
                           => n12, Z => MR_int_3_31_port);
   M1_2_30_0 : MUX2_X1 port map( A => MR_int_2_30_port, B => MR_int_2_2_port, S
                           => n12, Z => MR_int_3_30_port);
   M1_2_29_0 : MUX2_X1 port map( A => MR_int_2_29_port, B => MR_int_2_1_port, S
                           => n12, Z => MR_int_3_29_port);
   M1_2_28_0 : MUX2_X1 port map( A => MR_int_2_28_port, B => MR_int_2_0_port, S
                           => n12, Z => MR_int_3_28_port);
   M1_2_27_0 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, 
                           S => n12, Z => MR_int_3_27_port);
   M1_2_26_0 : MUX2_X1 port map( A => MR_int_2_26_port, B => MR_int_2_30_port, 
                           S => n12, Z => MR_int_3_26_port);
   M1_2_25_0 : MUX2_X1 port map( A => MR_int_2_25_port, B => MR_int_2_29_port, 
                           S => n12, Z => MR_int_3_25_port);
   M1_2_24_0 : MUX2_X1 port map( A => MR_int_2_24_port, B => MR_int_2_28_port, 
                           S => n12, Z => MR_int_3_24_port);
   M1_2_23_0 : MUX2_X1 port map( A => MR_int_2_23_port, B => MR_int_2_27_port, 
                           S => n12, Z => MR_int_3_23_port);
   M1_2_22_0 : MUX2_X1 port map( A => MR_int_2_22_port, B => MR_int_2_26_port, 
                           S => n12, Z => MR_int_3_22_port);
   M1_2_21_0 : MUX2_X1 port map( A => MR_int_2_21_port, B => MR_int_2_25_port, 
                           S => n11, Z => MR_int_3_21_port);
   M1_2_20_0 : MUX2_X1 port map( A => MR_int_2_20_port, B => MR_int_2_24_port, 
                           S => n11, Z => MR_int_3_20_port);
   M1_2_19_0 : MUX2_X1 port map( A => MR_int_2_19_port, B => MR_int_2_23_port, 
                           S => n11, Z => MR_int_3_19_port);
   M1_2_18_0 : MUX2_X1 port map( A => MR_int_2_18_port, B => MR_int_2_22_port, 
                           S => n11, Z => MR_int_3_18_port);
   M1_2_17_0 : MUX2_X1 port map( A => MR_int_2_17_port, B => MR_int_2_21_port, 
                           S => n11, Z => MR_int_3_17_port);
   M1_2_16_0 : MUX2_X1 port map( A => MR_int_2_16_port, B => MR_int_2_20_port, 
                           S => n11, Z => MR_int_3_16_port);
   M1_2_15_0 : MUX2_X1 port map( A => MR_int_2_15_port, B => MR_int_2_19_port, 
                           S => n11, Z => MR_int_3_15_port);
   M1_2_14_0 : MUX2_X1 port map( A => MR_int_2_14_port, B => MR_int_2_18_port, 
                           S => n11, Z => MR_int_3_14_port);
   M1_2_13_0 : MUX2_X1 port map( A => MR_int_2_13_port, B => MR_int_2_17_port, 
                           S => n11, Z => MR_int_3_13_port);
   M1_2_12_0 : MUX2_X1 port map( A => MR_int_2_12_port, B => MR_int_2_16_port, 
                           S => n11, Z => MR_int_3_12_port);
   M1_2_11_0 : MUX2_X1 port map( A => MR_int_2_11_port, B => MR_int_2_15_port, 
                           S => n11, Z => MR_int_3_11_port);
   M1_2_10_0 : MUX2_X1 port map( A => MR_int_2_10_port, B => MR_int_2_14_port, 
                           S => n10, Z => MR_int_3_10_port);
   M1_2_9_0 : MUX2_X1 port map( A => MR_int_2_9_port, B => MR_int_2_13_port, S 
                           => n10, Z => MR_int_3_9_port);
   M1_2_8_0 : MUX2_X1 port map( A => MR_int_2_8_port, B => MR_int_2_12_port, S 
                           => n10, Z => MR_int_3_8_port);
   M1_2_7_0 : MUX2_X1 port map( A => MR_int_2_7_port, B => MR_int_2_11_port, S 
                           => n10, Z => MR_int_3_7_port);
   M1_2_6_0 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_10_port, S 
                           => n10, Z => MR_int_3_6_port);
   M1_2_5_0 : MUX2_X1 port map( A => MR_int_2_5_port, B => MR_int_2_9_port, S 
                           => n10, Z => MR_int_3_5_port);
   M1_2_4_0 : MUX2_X1 port map( A => MR_int_2_4_port, B => MR_int_2_8_port, S 
                           => n10, Z => MR_int_3_4_port);
   M1_2_3 : MUX2_X1 port map( A => MR_int_2_3_port, B => MR_int_2_7_port, S => 
                           n10, Z => MR_int_3_3_port);
   M1_2_2 : MUX2_X1 port map( A => MR_int_2_2_port, B => MR_int_2_6_port, S => 
                           n10, Z => MR_int_3_2_port);
   M1_2_1 : MUX2_X1 port map( A => MR_int_2_1_port, B => MR_int_2_5_port, S => 
                           n10, Z => MR_int_3_1_port);
   M1_2_0 : MUX2_X1 port map( A => MR_int_2_0_port, B => MR_int_2_4_port, S => 
                           n10, Z => MR_int_3_0_port);
   M1_1_31_0 : MUX2_X1 port map( A => MR_int_1_31_port, B => MR_int_1_1_port, S
                           => n9, Z => MR_int_2_31_port);
   M1_1_30_0 : MUX2_X1 port map( A => MR_int_1_30_port, B => MR_int_1_0_port, S
                           => n9, Z => MR_int_2_30_port);
   M1_1_29_0 : MUX2_X1 port map( A => MR_int_1_29_port, B => MR_int_1_31_port, 
                           S => n9, Z => MR_int_2_29_port);
   M1_1_28_0 : MUX2_X1 port map( A => MR_int_1_28_port, B => MR_int_1_30_port, 
                           S => n9, Z => MR_int_2_28_port);
   M1_1_27_0 : MUX2_X1 port map( A => MR_int_1_27_port, B => MR_int_1_29_port, 
                           S => n9, Z => MR_int_2_27_port);
   M1_1_26_0 : MUX2_X1 port map( A => MR_int_1_26_port, B => MR_int_1_28_port, 
                           S => n9, Z => MR_int_2_26_port);
   M1_1_25_0 : MUX2_X1 port map( A => MR_int_1_25_port, B => MR_int_1_27_port, 
                           S => n9, Z => MR_int_2_25_port);
   M1_1_24_0 : MUX2_X1 port map( A => MR_int_1_24_port, B => MR_int_1_26_port, 
                           S => n9, Z => MR_int_2_24_port);
   M1_1_23_0 : MUX2_X1 port map( A => MR_int_1_23_port, B => MR_int_1_25_port, 
                           S => n9, Z => MR_int_2_23_port);
   M1_1_22_0 : MUX2_X1 port map( A => MR_int_1_22_port, B => MR_int_1_24_port, 
                           S => n9, Z => MR_int_2_22_port);
   M1_1_21_0 : MUX2_X1 port map( A => MR_int_1_21_port, B => MR_int_1_23_port, 
                           S => n8, Z => MR_int_2_21_port);
   M1_1_20_0 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_22_port, 
                           S => n8, Z => MR_int_2_20_port);
   M1_1_19_0 : MUX2_X1 port map( A => MR_int_1_19_port, B => MR_int_1_21_port, 
                           S => n8, Z => MR_int_2_19_port);
   M1_1_18_0 : MUX2_X1 port map( A => MR_int_1_18_port, B => MR_int_1_20_port, 
                           S => n8, Z => MR_int_2_18_port);
   M1_1_17_0 : MUX2_X1 port map( A => MR_int_1_17_port, B => MR_int_1_19_port, 
                           S => n8, Z => MR_int_2_17_port);
   M1_1_16_0 : MUX2_X1 port map( A => MR_int_1_16_port, B => MR_int_1_18_port, 
                           S => n8, Z => MR_int_2_16_port);
   M1_1_15_0 : MUX2_X1 port map( A => MR_int_1_15_port, B => MR_int_1_17_port, 
                           S => n8, Z => MR_int_2_15_port);
   M1_1_14_0 : MUX2_X1 port map( A => MR_int_1_14_port, B => MR_int_1_16_port, 
                           S => n8, Z => MR_int_2_14_port);
   M1_1_13_0 : MUX2_X1 port map( A => MR_int_1_13_port, B => MR_int_1_15_port, 
                           S => n8, Z => MR_int_2_13_port);
   M1_1_12_0 : MUX2_X1 port map( A => MR_int_1_12_port, B => MR_int_1_14_port, 
                           S => n8, Z => MR_int_2_12_port);
   M1_1_11_0 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_13_port, 
                           S => n8, Z => MR_int_2_11_port);
   M1_1_10_0 : MUX2_X1 port map( A => MR_int_1_10_port, B => MR_int_1_12_port, 
                           S => n7, Z => MR_int_2_10_port);
   M1_1_9_0 : MUX2_X1 port map( A => MR_int_1_9_port, B => MR_int_1_11_port, S 
                           => n7, Z => MR_int_2_9_port);
   M1_1_8_0 : MUX2_X1 port map( A => MR_int_1_8_port, B => MR_int_1_10_port, S 
                           => n7, Z => MR_int_2_8_port);
   M1_1_7_0 : MUX2_X1 port map( A => MR_int_1_7_port, B => MR_int_1_9_port, S 
                           => n7, Z => MR_int_2_7_port);
   M1_1_6_0 : MUX2_X1 port map( A => MR_int_1_6_port, B => MR_int_1_8_port, S 
                           => n7, Z => MR_int_2_6_port);
   M1_1_5_0 : MUX2_X1 port map( A => MR_int_1_5_port, B => MR_int_1_7_port, S 
                           => n7, Z => MR_int_2_5_port);
   M1_1_4_0 : MUX2_X1 port map( A => MR_int_1_4_port, B => MR_int_1_6_port, S 
                           => n7, Z => MR_int_2_4_port);
   M1_1_3_0 : MUX2_X1 port map( A => MR_int_1_3_port, B => MR_int_1_5_port, S 
                           => n7, Z => MR_int_2_3_port);
   M1_1_2_0 : MUX2_X1 port map( A => MR_int_1_2_port, B => MR_int_1_4_port, S 
                           => n7, Z => MR_int_2_2_port);
   M1_1_1 : MUX2_X1 port map( A => MR_int_1_1_port, B => MR_int_1_3_port, S => 
                           n7, Z => MR_int_2_1_port);
   M1_1_0 : MUX2_X1 port map( A => MR_int_1_0_port, B => MR_int_1_2_port, S => 
                           n7, Z => MR_int_2_0_port);
   M1_0_31_0 : MUX2_X1 port map( A => A(31), B => A(0), S => n6, Z => 
                           MR_int_1_31_port);
   M1_0_30_0 : MUX2_X1 port map( A => A(30), B => A(31), S => n6, Z => 
                           MR_int_1_30_port);
   M1_0_29_0 : MUX2_X1 port map( A => A(29), B => A(30), S => n6, Z => 
                           MR_int_1_29_port);
   M1_0_28_0 : MUX2_X1 port map( A => A(28), B => A(29), S => n6, Z => 
                           MR_int_1_28_port);
   M1_0_27_0 : MUX2_X1 port map( A => A(27), B => A(28), S => n6, Z => 
                           MR_int_1_27_port);
   M1_0_26_0 : MUX2_X1 port map( A => A(26), B => A(27), S => n6, Z => 
                           MR_int_1_26_port);
   M1_0_25_0 : MUX2_X1 port map( A => A(25), B => A(26), S => n6, Z => 
                           MR_int_1_25_port);
   M1_0_24_0 : MUX2_X1 port map( A => A(24), B => A(25), S => n6, Z => 
                           MR_int_1_24_port);
   M1_0_23_0 : MUX2_X1 port map( A => A(23), B => A(24), S => n6, Z => 
                           MR_int_1_23_port);
   M1_0_22_0 : MUX2_X1 port map( A => A(22), B => A(23), S => n6, Z => 
                           MR_int_1_22_port);
   M1_0_21_0 : MUX2_X1 port map( A => A(21), B => A(22), S => n5, Z => 
                           MR_int_1_21_port);
   M1_0_20_0 : MUX2_X1 port map( A => A(20), B => A(21), S => n5, Z => 
                           MR_int_1_20_port);
   M1_0_19_0 : MUX2_X1 port map( A => A(19), B => A(20), S => n5, Z => 
                           MR_int_1_19_port);
   M1_0_18_0 : MUX2_X1 port map( A => A(18), B => A(19), S => n5, Z => 
                           MR_int_1_18_port);
   M1_0_17_0 : MUX2_X1 port map( A => A(17), B => A(18), S => n5, Z => 
                           MR_int_1_17_port);
   M1_0_16_0 : MUX2_X1 port map( A => A(16), B => A(17), S => n5, Z => 
                           MR_int_1_16_port);
   M1_0_15_0 : MUX2_X1 port map( A => A(15), B => A(16), S => n5, Z => 
                           MR_int_1_15_port);
   M1_0_14_0 : MUX2_X1 port map( A => A(14), B => A(15), S => n5, Z => 
                           MR_int_1_14_port);
   M1_0_13_0 : MUX2_X1 port map( A => A(13), B => A(14), S => n5, Z => 
                           MR_int_1_13_port);
   M1_0_12_0 : MUX2_X1 port map( A => A(12), B => A(13), S => n5, Z => 
                           MR_int_1_12_port);
   M1_0_11_0 : MUX2_X1 port map( A => A(11), B => A(12), S => n5, Z => 
                           MR_int_1_11_port);
   M1_0_10_0 : MUX2_X1 port map( A => A(10), B => A(11), S => n4, Z => 
                           MR_int_1_10_port);
   M1_0_9_0 : MUX2_X1 port map( A => A(9), B => A(10), S => n4, Z => 
                           MR_int_1_9_port);
   M1_0_8_0 : MUX2_X1 port map( A => A(8), B => A(9), S => n4, Z => 
                           MR_int_1_8_port);
   M1_0_7_0 : MUX2_X1 port map( A => A(7), B => A(8), S => n4, Z => 
                           MR_int_1_7_port);
   M1_0_6_0 : MUX2_X1 port map( A => A(6), B => A(7), S => n4, Z => 
                           MR_int_1_6_port);
   M1_0_5_0 : MUX2_X1 port map( A => A(5), B => A(6), S => n4, Z => 
                           MR_int_1_5_port);
   M1_0_4_0 : MUX2_X1 port map( A => A(4), B => A(5), S => n4, Z => 
                           MR_int_1_4_port);
   M1_0_3_0 : MUX2_X1 port map( A => A(3), B => A(4), S => n4, Z => 
                           MR_int_1_3_port);
   M1_0_2_0 : MUX2_X1 port map( A => A(2), B => A(3), S => n4, Z => 
                           MR_int_1_2_port);
   M1_0_1_0 : MUX2_X1 port map( A => A(1), B => A(2), S => n4, Z => 
                           MR_int_1_1_port);
   M1_0_0 : MUX2_X1 port map( A => A(0), B => A(1), S => n4, Z => 
                           MR_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(3), Z => n14);
   U3 : BUF_X1 port map( A => SH(3), Z => n13);
   U4 : BUF_X1 port map( A => SH(4), Z => n16);
   U5 : BUF_X1 port map( A => SH(4), Z => n17);
   U6 : BUF_X1 port map( A => SH(3), Z => n15);
   U7 : BUF_X1 port map( A => SH(4), Z => n18);
   U8 : BUF_X1 port map( A => SH(0), Z => n5);
   U9 : BUF_X1 port map( A => SH(0), Z => n4);
   U10 : BUF_X1 port map( A => SH(1), Z => n8);
   U11 : BUF_X1 port map( A => SH(1), Z => n7);
   U12 : BUF_X1 port map( A => SH(2), Z => n11);
   U13 : BUF_X1 port map( A => SH(2), Z => n10);
   U14 : BUF_X1 port map( A => SH(0), Z => n6);
   U15 : BUF_X1 port map( A => SH(1), Z => n9);
   U16 : BUF_X1 port map( A => SH(2), Z => n12);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_lbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_lbsh_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_lbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n18, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n18, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n18, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n18, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n18, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n18, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n18, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n18, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n18, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n18, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n16, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n16, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n16, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n16, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n16, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n16, Z => B(16));
   M0_4_15 : MUX2_X1 port map( A => ML_int_4_15_port, B => ML_int_4_31_port, S 
                           => n16, Z => B(15));
   M0_4_14 : MUX2_X1 port map( A => ML_int_4_14_port, B => ML_int_4_30_port, S 
                           => n16, Z => B(14));
   M0_4_13 : MUX2_X1 port map( A => ML_int_4_13_port, B => ML_int_4_29_port, S 
                           => n16, Z => B(13));
   M0_4_12 : MUX2_X1 port map( A => ML_int_4_12_port, B => ML_int_4_28_port, S 
                           => n16, Z => B(12));
   M0_4_11 : MUX2_X1 port map( A => ML_int_4_11_port, B => ML_int_4_27_port, S 
                           => n16, Z => B(11));
   M0_4_10 : MUX2_X1 port map( A => ML_int_4_10_port, B => ML_int_4_26_port, S 
                           => n17, Z => B(10));
   M0_4_9 : MUX2_X1 port map( A => ML_int_4_9_port, B => ML_int_4_25_port, S =>
                           n17, Z => B(9));
   M0_4_8 : MUX2_X1 port map( A => ML_int_4_8_port, B => ML_int_4_24_port, S =>
                           n17, Z => B(8));
   M0_4_7 : MUX2_X1 port map( A => ML_int_4_7_port, B => ML_int_4_23_port, S =>
                           n17, Z => B(7));
   M0_4_6 : MUX2_X1 port map( A => ML_int_4_6_port, B => ML_int_4_22_port, S =>
                           n17, Z => B(6));
   M0_4_5 : MUX2_X1 port map( A => ML_int_4_5_port, B => ML_int_4_21_port, S =>
                           n17, Z => B(5));
   M0_4_4 : MUX2_X1 port map( A => ML_int_4_4_port, B => ML_int_4_20_port, S =>
                           n17, Z => B(4));
   M0_4_3 : MUX2_X1 port map( A => ML_int_4_3_port, B => ML_int_4_19_port, S =>
                           n17, Z => B(3));
   M0_4_2 : MUX2_X1 port map( A => ML_int_4_2_port, B => ML_int_4_18_port, S =>
                           n17, Z => B(2));
   M0_4_1 : MUX2_X1 port map( A => ML_int_4_1_port, B => ML_int_4_17_port, S =>
                           n17, Z => B(1));
   M0_4_0 : MUX2_X1 port map( A => ML_int_4_0_port, B => ML_int_4_16_port, S =>
                           n17, Z => B(0));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n15, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n15, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n15, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n15, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n15, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n15, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n15, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => n15, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n15, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => n15, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n14, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n14, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n14, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n14, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n14, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n14, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n14, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n14, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n14, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n14, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n14, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n13, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n13, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n13, Z => ML_int_4_8_port);
   M0_3_7 : MUX2_X1 port map( A => ML_int_3_7_port, B => ML_int_3_31_port, S =>
                           n13, Z => ML_int_4_7_port);
   M0_3_6 : MUX2_X1 port map( A => ML_int_3_6_port, B => ML_int_3_30_port, S =>
                           n13, Z => ML_int_4_6_port);
   M0_3_5 : MUX2_X1 port map( A => ML_int_3_5_port, B => ML_int_3_29_port, S =>
                           n13, Z => ML_int_4_5_port);
   M0_3_4 : MUX2_X1 port map( A => ML_int_3_4_port, B => ML_int_3_28_port, S =>
                           n13, Z => ML_int_4_4_port);
   M0_3_3 : MUX2_X1 port map( A => ML_int_3_3_port, B => ML_int_3_27_port, S =>
                           n13, Z => ML_int_4_3_port);
   M0_3_2 : MUX2_X1 port map( A => ML_int_3_2_port, B => ML_int_3_26_port, S =>
                           n13, Z => ML_int_4_2_port);
   M0_3_1 : MUX2_X1 port map( A => ML_int_3_1_port, B => ML_int_3_25_port, S =>
                           n13, Z => ML_int_4_1_port);
   M0_3_0 : MUX2_X1 port map( A => ML_int_3_0_port, B => ML_int_3_24_port, S =>
                           n13, Z => ML_int_4_0_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => n12, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n12, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n12, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => n12, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n12, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n12, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n12, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n12, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n12, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n12, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n11, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n11, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => n11, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n11, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => n11, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n11, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n11, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n11, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n11, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n11, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => n11, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n10, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n10, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n10, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n10, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n10, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n10, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n10, Z => ML_int_3_4_port);
   M0_2_3 : MUX2_X1 port map( A => ML_int_2_3_port, B => ML_int_2_31_port, S =>
                           n10, Z => ML_int_3_3_port);
   M0_2_2 : MUX2_X1 port map( A => ML_int_2_2_port, B => ML_int_2_30_port, S =>
                           n10, Z => ML_int_3_2_port);
   M0_2_1 : MUX2_X1 port map( A => ML_int_2_1_port, B => ML_int_2_29_port, S =>
                           n10, Z => ML_int_3_1_port);
   M0_2_0 : MUX2_X1 port map( A => ML_int_2_0_port, B => ML_int_2_28_port, S =>
                           n10, Z => ML_int_3_0_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => n9, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => n9, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => n9, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => n9, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n9, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => n9, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => n9, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => n9, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => n9, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n9, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => n8, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => n8, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n8, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n8, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => n8, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n8, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => n8, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n8, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n8, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n8, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n8, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n7, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n7, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n7, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n7, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n7, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n7, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n7, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n7, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n7, Z => ML_int_2_2_port);
   M0_1_1 : MUX2_X1 port map( A => ML_int_1_1_port, B => ML_int_1_31_port, S =>
                           n7, Z => ML_int_2_1_port);
   M0_1_0 : MUX2_X1 port map( A => ML_int_1_0_port, B => ML_int_1_30_port, S =>
                           n7, Z => ML_int_2_0_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n6, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n6, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n6, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n6, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n6, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n6, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n6, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n6, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n6, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n6, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n5, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n5, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n5, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n5, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n5, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n5, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n5, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n5, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n5, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n5, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n5, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n4, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n4, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n4, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n4, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n4, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n4, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n4, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n4, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n4, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n4, Z => 
                           ML_int_1_1_port);
   M0_0_0 : MUX2_X1 port map( A => A(0), B => A(31), S => n4, Z => 
                           ML_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(3), Z => n14);
   U3 : BUF_X1 port map( A => SH(3), Z => n13);
   U4 : BUF_X1 port map( A => SH(4), Z => n16);
   U5 : BUF_X1 port map( A => SH(4), Z => n17);
   U6 : BUF_X1 port map( A => SH(3), Z => n15);
   U7 : BUF_X1 port map( A => SH(4), Z => n18);
   U8 : BUF_X1 port map( A => SH(0), Z => n4);
   U9 : BUF_X1 port map( A => SH(0), Z => n5);
   U10 : BUF_X1 port map( A => SH(1), Z => n7);
   U11 : BUF_X1 port map( A => SH(1), Z => n8);
   U12 : BUF_X1 port map( A => SH(2), Z => n11);
   U13 : BUF_X1 port map( A => SH(2), Z => n10);
   U14 : BUF_X1 port map( A => SH(0), Z => n6);
   U15 : BUF_X1 port map( A => SH(1), Z => n9);
   U16 : BUF_X1 port map( A => SH(2), Z => n12);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sra_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sra_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n57, n58, n59
      , n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102
      , n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233 : 
      std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U4 : NOR2_X2 port map( A1 => n174, A2 => SH(3), ZN => n109);
   U7 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n111);
   U174 : MUX2_X1 port map( A => A(30), B => A(31), S => n95, Z => n120);
   U2 : NAND2_X1 port map( A1 => n181, A2 => A(31), ZN => n97);
   U3 : INV_X1 port map( A => n181, ZN => n177);
   U5 : INV_X1 port map( A => n85, ZN => n228);
   U6 : INV_X1 port map( A => n94, ZN => n232);
   U8 : INV_X1 port map( A => n95, ZN => n233);
   U9 : INV_X1 port map( A => n91, ZN => n230);
   U10 : INV_X1 port map( A => n92, ZN => n231);
   U11 : NAND2_X1 port map( A1 => n109, A2 => n177, ZN => n85);
   U12 : INV_X1 port map( A => n58, ZN => n229);
   U13 : BUF_X1 port map( A => n176, Z => n180);
   U14 : BUF_X1 port map( A => n175, Z => n179);
   U15 : BUF_X1 port map( A => n175, Z => n178);
   U16 : BUF_X1 port map( A => n176, Z => n181);
   U17 : NOR2_X2 port map( A1 => n173, A2 => SH(0), ZN => n91);
   U18 : NOR2_X2 port map( A1 => n172, A2 => n173, ZN => n92);
   U19 : NAND2_X1 port map( A1 => n111, A2 => n177, ZN => n58);
   U20 : NAND2_X1 port map( A1 => n172, A2 => n173, ZN => n95);
   U21 : NAND2_X1 port map( A1 => SH(0), A2 => n173, ZN => n94);
   U22 : AND2_X1 port map( A1 => n163, A2 => n174, ZN => n61);
   U23 : AND2_X1 port map( A1 => SH(3), A2 => n174, ZN => n119);
   U24 : AOI21_X1 port map( B1 => n108, B2 => n111, A => n140, ZN => n104);
   U25 : AND2_X1 port map( A1 => SH(3), A2 => n177, ZN => n163);
   U26 : BUF_X1 port map( A => SH(4), Z => n176);
   U27 : BUF_X1 port map( A => SH(4), Z => n175);
   U28 : OAI222_X1 port map( A1 => n95, A2 => n192, B1 => n94, B2 => n191, C1 
                           => n173, C2 => n186, ZN => n108);
   U29 : AND2_X1 port map( A1 => SH(2), A2 => n163, ZN => n63);
   U30 : AOI221_X1 port map( B1 => n120, B2 => n109, C1 => n116, C2 => n111, A 
                           => n188, ZN => n107);
   U31 : AOI221_X1 port map( B1 => n108, B2 => n109, C1 => n110, C2 => n111, A 
                           => n188, ZN => n59);
   U32 : AOI221_X1 port map( B1 => n112, B2 => n109, C1 => n113, C2 => n111, A 
                           => n188, ZN => n66);
   U33 : AOI221_X1 port map( B1 => n114, B2 => n109, C1 => n115, C2 => n111, A 
                           => n188, ZN => n71);
   U34 : AOI221_X1 port map( B1 => n116, B2 => n109, C1 => n117, C2 => n111, A 
                           => n189, ZN => n76);
   U35 : INV_X1 port map( A => n118, ZN => n189);
   U36 : AOI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n118);
   U37 : AOI221_X1 port map( B1 => n110, B2 => n109, C1 => n64, C2 => n111, A 
                           => n184, ZN => n80);
   U38 : INV_X1 port map( A => n122, ZN => n184);
   U39 : AOI21_X1 port map( B1 => n119, B2 => n108, A => n121, ZN => n122);
   U40 : AOI221_X1 port map( B1 => n113, B2 => n109, C1 => n69, C2 => n111, A 
                           => n182, ZN => n83);
   U41 : INV_X1 port map( A => n123, ZN => n182);
   U42 : AOI21_X1 port map( B1 => n119, B2 => n112, A => n121, ZN => n123);
   U43 : AOI221_X1 port map( B1 => n115, B2 => n109, C1 => n74, C2 => n111, A 
                           => n190, ZN => n86);
   U44 : INV_X1 port map( A => n131, ZN => n190);
   U45 : AOI21_X1 port map( B1 => n119, B2 => n114, A => n121, ZN => n131);
   U46 : AOI221_X1 port map( B1 => n120, B2 => n133, C1 => n116, C2 => n119, A 
                           => n196, ZN => n98);
   U47 : INV_X1 port map( A => n134, ZN => n196);
   U48 : AOI22_X1 port map( A1 => n109, A2 => n117, B1 => n111, B2 => n78, ZN 
                           => n134);
   U49 : AOI221_X1 port map( B1 => n64, B2 => n109, C1 => n62, C2 => n111, A =>
                           n185, ZN => n124);
   U50 : INV_X1 port map( A => n135, ZN => n185);
   U51 : AOI22_X1 port map( A1 => n133, A2 => n108, B1 => n119, B2 => n110, ZN 
                           => n135);
   U52 : AOI221_X1 port map( B1 => n69, B2 => n109, C1 => n68, C2 => n111, A =>
                           n183, ZN => n136);
   U53 : INV_X1 port map( A => n166, ZN => n183);
   U54 : AOI22_X1 port map( A1 => n133, A2 => n112, B1 => n119, B2 => n113, ZN 
                           => n166);
   U55 : AOI222_X1 port map( A1 => n228, A2 => n68, B1 => n61, B2 => n69, C1 =>
                           n63, C2 => n113, ZN => n147);
   U56 : AOI222_X1 port map( A1 => n228, A2 => n73, B1 => n61, B2 => n74, C1 =>
                           n63, C2 => n115, ZN => n148);
   U57 : AOI222_X1 port map( A1 => n228, A2 => n207, B1 => n61, B2 => n78, C1 
                           => n63, C2 => n117, ZN => n154);
   U58 : AOI222_X1 port map( A1 => n228, A2 => n78, B1 => n61, B2 => n117, C1 
                           => n63, C2 => n116, ZN => n139);
   U59 : AOI222_X1 port map( A1 => n228, A2 => n209, B1 => n61, B2 => n68, C1 
                           => n63, C2 => n69, ZN => n67);
   U60 : AOI222_X1 port map( A1 => n228, A2 => n62, B1 => n61, B2 => n64, C1 =>
                           n63, C2 => n110, ZN => n141);
   U61 : AOI222_X1 port map( A1 => n228, A2 => n208, B1 => n61, B2 => n62, C1 
                           => n63, C2 => n64, ZN => n60);
   U62 : AOI222_X1 port map( A1 => n228, A2 => n212, B1 => n61, B2 => n73, C1 
                           => n63, C2 => n74, ZN => n72);
   U63 : AOI222_X1 port map( A1 => n228, A2 => n213, B1 => n61, B2 => n207, C1 
                           => n63, C2 => n78, ZN => n77);
   U64 : AOI222_X1 port map( A1 => n228, A2 => n216, B1 => n61, B2 => n208, C1 
                           => n63, C2 => n62, ZN => n81);
   U65 : AOI222_X1 port map( A1 => n228, A2 => n218, B1 => n61, B2 => n209, C1 
                           => n63, C2 => n68, ZN => n84);
   U66 : OAI21_X1 port map( B1 => n180, B2 => n96, A => n97, ZN => B_30_port);
   U67 : OAI21_X1 port map( B1 => n180, B2 => n104, A => n97, ZN => B_29_port);
   U68 : OAI21_X1 port map( B1 => n180, B2 => n105, A => n97, ZN => B_28_port);
   U69 : OAI21_X1 port map( B1 => n180, B2 => n106, A => n97, ZN => B_27_port);
   U70 : OAI21_X1 port map( B1 => n180, B2 => n107, A => n97, ZN => B_26_port);
   U71 : OAI21_X1 port map( B1 => n179, B2 => n59, A => n97, ZN => B_25_port);
   U72 : OAI21_X1 port map( B1 => n179, B2 => n66, A => n97, ZN => B_24_port);
   U73 : OAI21_X1 port map( B1 => n179, B2 => n71, A => n97, ZN => B_23_port);
   U74 : OAI21_X1 port map( B1 => n179, B2 => n76, A => n97, ZN => B_22_port);
   U75 : OAI21_X1 port map( B1 => n178, B2 => n80, A => n97, ZN => B_21_port);
   U76 : OAI21_X1 port map( B1 => n178, B2 => n83, A => n97, ZN => B_20_port);
   U77 : OAI21_X1 port map( B1 => n179, B2 => n86, A => n97, ZN => B_19_port);
   U78 : OAI21_X1 port map( B1 => n178, B2 => n98, A => n97, ZN => B_18_port);
   U79 : OAI21_X1 port map( B1 => n178, B2 => n124, A => n97, ZN => B_17_port);
   U80 : OAI21_X1 port map( B1 => n178, B2 => n136, A => n97, ZN => B_16_port);
   U81 : OAI221_X1 port map( B1 => n200, B2 => n85, C1 => n204, C2 => n58, A =>
                           n137, ZN => B_15_port);
   U82 : OAI221_X1 port map( B1 => n138, B2 => n58, C1 => n96, C2 => n177, A =>
                           n139, ZN => B_14_port);
   U83 : OAI221_X1 port map( B1 => n129, B2 => n58, C1 => n104, C2 => n177, A 
                           => n141, ZN => B_13_port);
   U84 : OAI221_X1 port map( B1 => n146, B2 => n58, C1 => n105, C2 => n177, A 
                           => n147, ZN => B_12_port);
   U85 : OAI221_X1 port map( B1 => n89, B2 => n58, C1 => n106, C2 => n177, A =>
                           n148, ZN => B_11_port);
   U86 : OAI221_X1 port map( B1 => n101, B2 => n58, C1 => n107, C2 => n177, A 
                           => n154, ZN => B_10_port);
   U87 : OAI221_X1 port map( B1 => n75, B2 => n85, C1 => n98, C2 => n177, A => 
                           n99, ZN => B_2_port);
   U88 : OAI221_X1 port map( B1 => n79, B2 => n85, C1 => n124, C2 => n177, A =>
                           n125, ZN => B_1_port);
   U89 : OAI221_X1 port map( B1 => n57, B2 => n58, C1 => n59, C2 => n177, A => 
                           n60, ZN => B_9_port);
   U90 : OAI221_X1 port map( B1 => n65, B2 => n58, C1 => n66, C2 => n177, A => 
                           n67, ZN => B_8_port);
   U91 : OAI221_X1 port map( B1 => n70, B2 => n58, C1 => n71, C2 => n177, A => 
                           n72, ZN => B_7_port);
   U92 : OAI221_X1 port map( B1 => n75, B2 => n58, C1 => n76, C2 => n177, A => 
                           n77, ZN => B_6_port);
   U93 : OAI221_X1 port map( B1 => n79, B2 => n58, C1 => n80, C2 => n177, A => 
                           n81, ZN => B_5_port);
   U94 : OAI221_X1 port map( B1 => n82, B2 => n58, C1 => n83, C2 => n177, A => 
                           n84, ZN => B_4_port);
   U95 : OAI221_X1 port map( B1 => n70, B2 => n85, C1 => n86, C2 => n177, A => 
                           n87, ZN => B_3_port);
   U96 : OAI21_X1 port map( B1 => n174, B2 => n186, A => n132, ZN => n140);
   U97 : AOI221_X1 port map( B1 => n63, B2 => n114, C1 => n61, C2 => n115, A =>
                           n187, ZN => n137);
   U98 : INV_X1 port map( A => n97, ZN => n187);
   U99 : NOR2_X1 port map( A1 => n132, A2 => n174, ZN => n121);
   U100 : AOI21_X1 port map( B1 => n120, B2 => n111, A => n140, ZN => n96);
   U101 : AOI21_X1 port map( B1 => n112, B2 => n111, A => n140, ZN => n105);
   U102 : AOI21_X1 port map( B1 => n114, B2 => n111, A => n140, ZN => n106);
   U103 : INV_X1 port map( A => SH(0), ZN => n172);
   U104 : INV_X1 port map( A => n132, ZN => n188);
   U105 : INV_X1 port map( A => n138, ZN => n207);
   U106 : INV_X1 port map( A => n129, ZN => n208);
   U107 : INV_X1 port map( A => n146, ZN => n209);
   U108 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n133);
   U109 : INV_X1 port map( A => n57, ZN => n216);
   U110 : INV_X1 port map( A => n101, ZN => n213);
   U111 : INV_X1 port map( A => n89, ZN => n212);
   U112 : INV_X1 port map( A => n65, ZN => n218);
   U113 : INV_X1 port map( A => n74, ZN => n200);
   U114 : INV_X1 port map( A => n73, ZN => n204);
   U115 : OAI221_X1 port map( B1 => n203, B2 => n94, C1 => n205, C2 => n95, A 
                           => n156, ZN => n78);
   U116 : AOI22_X1 port map( A1 => A(20), A2 => n91, B1 => A(21), B2 => n92, ZN
                           => n156);
   U117 : OAI221_X1 port map( B1 => n230, B2 => n198, C1 => n231, C2 => n197, A
                           => n155, ZN => n117);
   U118 : AOI22_X1 port map( A1 => A(23), A2 => n232, B1 => A(22), B2 => n233, 
                           ZN => n155);
   U119 : OAI221_X1 port map( B1 => n230, B2 => n191, C1 => n231, C2 => n186, A
                           => n168, ZN => n112);
   U120 : AOI22_X1 port map( A1 => A(29), A2 => n232, B1 => A(28), B2 => n233, 
                           ZN => n168);
   U121 : OAI221_X1 port map( B1 => n94, B2 => n201, C1 => n202, C2 => n95, A 
                           => n170, ZN => n69);
   U122 : INV_X1 port map( A => A(21), ZN => n201);
   U123 : AOI22_X1 port map( A1 => A(22), A2 => n91, B1 => A(23), B2 => n92, ZN
                           => n170);
   U124 : OAI221_X1 port map( B1 => n202, B2 => n94, C1 => n203, C2 => n95, A 
                           => n150, ZN => n74);
   U125 : AOI22_X1 port map( A1 => A(21), A2 => n91, B1 => A(22), B2 => n92, ZN
                           => n150);
   U126 : OAI221_X1 port map( B1 => n230, B2 => n197, C1 => n231, C2 => n195, A
                           => n149, ZN => n115);
   U127 : AOI22_X1 port map( A1 => A(24), A2 => n232, B1 => A(23), B2 => n233, 
                           ZN => n149);
   U128 : OAI221_X1 port map( B1 => n230, B2 => n194, C1 => n231, C2 => n193, A
                           => n142, ZN => n110);
   U129 : AOI22_X1 port map( A1 => A(26), A2 => n232, B1 => A(25), B2 => n233, 
                           ZN => n142);
   U130 : OAI221_X1 port map( B1 => n230, B2 => n195, C1 => n231, C2 => n194, A
                           => n167, ZN => n113);
   U131 : AOI22_X1 port map( A1 => A(25), A2 => n232, B1 => A(24), B2 => n233, 
                           ZN => n167);
   U132 : OAI221_X1 port map( B1 => n230, B2 => n199, C1 => n231, C2 => n198, A
                           => n143, ZN => n64);
   U133 : INV_X1 port map( A => A(23), ZN => n199);
   U134 : AOI22_X1 port map( A1 => A(22), A2 => n232, B1 => A(21), B2 => n233, 
                           ZN => n143);
   U135 : OAI221_X1 port map( B1 => n230, B2 => n206, C1 => n231, C2 => n205, A
                           => n151, ZN => n73);
   U136 : INV_X1 port map( A => A(17), ZN => n206);
   U137 : AOI22_X1 port map( A1 => A(16), A2 => n232, B1 => A(15), B2 => n233, 
                           ZN => n151);
   U138 : OAI221_X1 port map( B1 => n230, B2 => n203, C1 => n231, C2 => n202, A
                           => n144, ZN => n62);
   U139 : AOI22_X1 port map( A1 => A(18), A2 => n232, B1 => A(17), B2 => n233, 
                           ZN => n144);
   U140 : OAI221_X1 port map( B1 => n230, B2 => n205, C1 => n203, C2 => n231, A
                           => n169, ZN => n68);
   U141 : AOI22_X1 port map( A1 => A(17), A2 => n232, B1 => A(16), B2 => n233, 
                           ZN => n169);
   U142 : OAI221_X1 port map( B1 => n230, B2 => n192, C1 => n231, C2 => n191, A
                           => n152, ZN => n114);
   U143 : AOI22_X1 port map( A1 => A(28), A2 => n232, B1 => A(27), B2 => n233, 
                           ZN => n152);
   U144 : OAI221_X1 port map( B1 => n230, B2 => n193, C1 => n231, C2 => n192, A
                           => n158, ZN => n116);
   U145 : AOI22_X1 port map( A1 => A(27), A2 => n232, B1 => A(26), B2 => n233, 
                           ZN => n158);
   U146 : AOI221_X1 port map( B1 => n91, B2 => A(8), C1 => n92, C2 => A(9), A 
                           => n103, ZN => n75);
   U147 : OAI22_X1 port map( A1 => n222, A2 => n94, B1 => n223, B2 => n95, ZN 
                           => n103);
   U148 : AOI221_X1 port map( B1 => n91, B2 => A(9), C1 => n92, C2 => A(10), A 
                           => n93, ZN => n70);
   U149 : OAI22_X1 port map( A1 => n221, A2 => n94, B1 => n222, B2 => n95, ZN 
                           => n93);
   U150 : AOI221_X1 port map( B1 => n91, B2 => A(7), C1 => n92, C2 => A(8), A 
                           => n130, ZN => n79);
   U151 : OAI22_X1 port map( A1 => n223, A2 => n94, B1 => n224, B2 => n95, ZN 
                           => n130);
   U152 : AOI221_X1 port map( B1 => n91, B2 => A(6), C1 => n92, C2 => A(7), A 
                           => n171, ZN => n82);
   U153 : OAI22_X1 port map( A1 => n224, A2 => n94, B1 => n225, B2 => n95, ZN 
                           => n171);
   U154 : AOI221_X1 port map( B1 => n91, B2 => A(11), C1 => n92, C2 => A(12), A
                           => n127, ZN => n57);
   U155 : OAI22_X1 port map( A1 => n219, A2 => n94, B1 => n220, B2 => n95, ZN 
                           => n127);
   U156 : AOI221_X1 port map( B1 => n91, B2 => A(12), C1 => n92, C2 => A(13), A
                           => n159, ZN => n101);
   U157 : OAI22_X1 port map( A1 => n217, A2 => n94, B1 => n219, B2 => n95, ZN 
                           => n159);
   U158 : AOI221_X1 port map( B1 => n91, B2 => A(13), C1 => n92, C2 => A(14), A
                           => n153, ZN => n89);
   U159 : OAI22_X1 port map( A1 => n215, A2 => n94, B1 => n217, B2 => n95, ZN 
                           => n153);
   U160 : INV_X1 port map( A => A(12), ZN => n215);
   U161 : AOI221_X1 port map( B1 => n91, B2 => A(16), C1 => n92, C2 => A(17), A
                           => n210, ZN => n138);
   U162 : INV_X1 port map( A => n157, ZN => n210);
   U163 : AOI22_X1 port map( A1 => A(15), A2 => n232, B1 => A(14), B2 => n233, 
                           ZN => n157);
   U164 : AOI221_X1 port map( B1 => n91, B2 => A(15), C1 => n92, C2 => A(16), A
                           => n211, ZN => n129);
   U165 : INV_X1 port map( A => n145, ZN => n211);
   U166 : AOI22_X1 port map( A1 => A(14), A2 => n232, B1 => A(13), B2 => n233, 
                           ZN => n145);
   U167 : AOI221_X1 port map( B1 => n91, B2 => A(14), C1 => n92, C2 => A(15), A
                           => n214, ZN => n146);
   U168 : INV_X1 port map( A => n165, ZN => n214);
   U169 : AOI22_X1 port map( A1 => A(13), A2 => n232, B1 => A(12), B2 => n233, 
                           ZN => n165);
   U170 : AOI221_X1 port map( B1 => n91, B2 => A(10), C1 => n92, C2 => A(11), A
                           => n162, ZN => n65);
   U171 : OAI22_X1 port map( A1 => n220, A2 => n94, B1 => n221, B2 => n95, ZN 
                           => n162);
   U172 : AOI222_X1 port map( A1 => n63, A2 => n73, B1 => n229, B2 => n88, C1 
                           => n61, C2 => n212, ZN => n87);
   U173 : OAI221_X1 port map( B1 => n230, B2 => n224, C1 => n231, C2 => n223, A
                           => n90, ZN => n88);
   U175 : AOI22_X1 port map( A1 => A(4), A2 => n232, B1 => A(3), B2 => n233, ZN
                           => n90);
   U176 : AOI222_X1 port map( A1 => n63, A2 => n208, B1 => n229, B2 => n126, C1
                           => n61, C2 => n216, ZN => n125);
   U177 : OAI221_X1 port map( B1 => n230, B2 => n226, C1 => n231, C2 => n225, A
                           => n128, ZN => n126);
   U178 : AOI22_X1 port map( A1 => A(2), A2 => n232, B1 => A(1), B2 => n233, ZN
                           => n128);
   U179 : AOI222_X1 port map( A1 => n63, A2 => n209, B1 => n229, B2 => n161, C1
                           => n61, C2 => n218, ZN => n160);
   U180 : OAI221_X1 port map( B1 => n230, B2 => n227, C1 => n231, C2 => n226, A
                           => n164, ZN => n161);
   U181 : INV_X1 port map( A => A(2), ZN => n227);
   U182 : AOI22_X1 port map( A1 => A(1), A2 => n232, B1 => A(0), B2 => n233, ZN
                           => n164);
   U183 : AOI222_X1 port map( A1 => n63, A2 => n207, B1 => n229, B2 => n100, C1
                           => n61, C2 => n213, ZN => n99);
   U184 : OAI221_X1 port map( B1 => n230, B2 => n225, C1 => n231, C2 => n224, A
                           => n102, ZN => n100);
   U185 : AOI22_X1 port map( A1 => A(3), A2 => n232, B1 => A(2), B2 => n233, ZN
                           => n102);
   U186 : OAI221_X1 port map( B1 => n82, B2 => n85, C1 => n136, C2 => n177, A 
                           => n160, ZN => B_0_port);
   U187 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n132);
   U188 : INV_X1 port map( A => A(19), ZN => n203);
   U189 : INV_X1 port map( A => A(5), ZN => n224);
   U190 : INV_X1 port map( A => A(18), ZN => n205);
   U191 : INV_X1 port map( A => A(6), ZN => n223);
   U192 : INV_X1 port map( A => A(4), ZN => n225);
   U193 : INV_X1 port map( A => A(29), ZN => n192);
   U194 : INV_X1 port map( A => A(20), ZN => n202);
   U195 : INV_X1 port map( A => A(31), ZN => n186);
   U196 : INV_X1 port map( A => A(9), ZN => n220);
   U197 : INV_X1 port map( A => A(11), ZN => n217);
   U198 : INV_X1 port map( A => A(10), ZN => n219);
   U199 : INV_X1 port map( A => A(8), ZN => n221);
   U200 : INV_X1 port map( A => A(7), ZN => n222);
   U201 : INV_X1 port map( A => A(3), ZN => n226);
   U202 : INV_X1 port map( A => A(27), ZN => n194);
   U203 : INV_X1 port map( A => A(26), ZN => n195);
   U204 : INV_X1 port map( A => A(25), ZN => n197);
   U205 : INV_X1 port map( A => A(28), ZN => n193);
   U206 : INV_X1 port map( A => A(24), ZN => n198);
   U207 : INV_X1 port map( A => A(30), ZN => n191);
   U208 : INV_X1 port map( A => SH(1), ZN => n173);
   U209 : INV_X1 port map( A => SH(2), ZN => n174);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW_rash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228 : std_logic;

begin
   
   U3 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n96);
   U5 : NOR2_X2 port map( A1 => n167, A2 => SH(1), ZN => n95);
   U141 : MUX2_X1 port map( A => n112, B => n98, S => SH(2), Z => n123);
   U4 : INV_X1 port map( A => n57, ZN => n223);
   U6 : NAND2_X1 port map( A1 => n224, A2 => n177, ZN => n57);
   U7 : INV_X1 port map( A => n174, ZN => n177);
   U8 : INV_X1 port map( A => n87, ZN => n222);
   U9 : NAND2_X1 port map( A1 => n110, A2 => n177, ZN => n87);
   U10 : NOR2_X1 port map( A1 => n177, A2 => n138, ZN => n129);
   U11 : INV_X1 port map( A => n138, ZN => n224);
   U12 : NOR2_X1 port map( A1 => n170, A2 => n171, ZN => n155);
   U13 : BUF_X1 port map( A => n176, Z => n171);
   U14 : BUF_X1 port map( A => n175, Z => n173);
   U15 : BUF_X1 port map( A => n176, Z => n172);
   U16 : BUF_X1 port map( A => n175, Z => n174);
   U17 : INV_X1 port map( A => n96, ZN => n227);
   U18 : INV_X1 port map( A => n95, ZN => n228);
   U19 : NOR2_X2 port map( A1 => n168, A2 => n169, ZN => n110);
   U20 : INV_X1 port map( A => n92, ZN => n226);
   U21 : INV_X1 port map( A => n93, ZN => n225);
   U22 : AND2_X1 port map( A1 => n155, A2 => n168, ZN => n61);
   U23 : NOR2_X1 port map( A1 => n168, A2 => n170, ZN => n125);
   U24 : INV_X1 port map( A => SH(3), ZN => n170);
   U25 : NAND2_X1 port map( A1 => n168, A2 => n170, ZN => n138);
   U26 : BUF_X1 port map( A => n93, Z => n164);
   U27 : BUF_X1 port map( A => n93, Z => n165);
   U28 : BUF_X1 port map( A => n93, Z => n166);
   U29 : INV_X1 port map( A => n123, ZN => n182);
   U30 : BUF_X1 port map( A => SH(4), Z => n175);
   U31 : BUF_X1 port map( A => SH(4), Z => n176);
   U32 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n92);
   U33 : OAI222_X1 port map( A1 => n228, A2 => n185, B1 => n164, B2 => n184, C1
                           => n227, C2 => n186, ZN => n106);
   U34 : AND2_X1 port map( A1 => SH(2), A2 => n155, ZN => n63);
   U35 : NOR2_X1 port map( A1 => n170, A2 => SH(2), ZN => n113);
   U36 : OAI22_X1 port map( A1 => n227, A2 => n185, B1 => n228, B2 => n184, ZN 
                           => n99);
   U37 : AOI222_X1 port map( A1 => n112, A2 => n110, B1 => n98, B2 => n113, C1 
                           => n114, C2 => n224, ZN => n72);
   U38 : AOI222_X1 port map( A1 => n115, A2 => n110, B1 => n99, B2 => n113, C1 
                           => n116, C2 => n224, ZN => n77);
   U39 : AOI222_X1 port map( A1 => n109, A2 => n110, B1 => n106, B2 => n113, C1
                           => n64, C2 => n224, ZN => n82);
   U40 : AOI222_X1 port map( A1 => n111, A2 => n110, B1 => n107, B2 => n113, C1
                           => n70, C2 => n224, ZN => n85);
   U41 : AOI222_X1 port map( A1 => n75, A2 => n224, B1 => n114, B2 => n110, C1 
                           => n123, C2 => n169, ZN => n88);
   U42 : AOI221_X1 port map( B1 => n116, B2 => n110, C1 => n80, C2 => n224, A 
                           => n181, ZN => n100);
   U43 : INV_X1 port map( A => n124, ZN => n181);
   U44 : AOI22_X1 port map( A1 => n125, A2 => n99, B1 => n113, B2 => n115, ZN 
                           => n124);
   U45 : AOI221_X1 port map( B1 => n64, B2 => n110, C1 => n62, C2 => n224, A =>
                           n183, ZN => n117);
   U46 : INV_X1 port map( A => n126, ZN => n183);
   U47 : AOI22_X1 port map( A1 => n125, A2 => n106, B1 => n113, B2 => n109, ZN 
                           => n126);
   U48 : AOI221_X1 port map( B1 => n70, B2 => n110, C1 => n69, C2 => n224, A =>
                           n180, ZN => n127);
   U49 : INV_X1 port map( A => n158, ZN => n180);
   U50 : AOI22_X1 port map( A1 => n125, A2 => n107, B1 => n113, B2 => n111, ZN 
                           => n158);
   U51 : AOI222_X1 port map( A1 => n63, A2 => n109, B1 => n129, B2 => n106, C1 
                           => n61, C2 => n64, ZN => n131);
   U52 : AOI222_X1 port map( A1 => n222, A2 => n79, B1 => n61, B2 => n80, C1 =>
                           n63, C2 => n116, ZN => n146);
   U53 : AOI222_X1 port map( A1 => n222, A2 => n60, B1 => n61, B2 => n62, C1 =>
                           n63, C2 => n64, ZN => n59);
   U54 : AOI222_X1 port map( A1 => n222, A2 => n68, B1 => n61, B2 => n69, C1 =>
                           n63, C2 => n70, ZN => n67);
   U55 : AOI222_X1 port map( A1 => n222, A2 => n208, B1 => n61, B2 => n79, C1 
                           => n63, C2 => n80, ZN => n78);
   U56 : AOI222_X1 port map( A1 => n222, A2 => n210, B1 => n61, B2 => n60, C1 
                           => n63, C2 => n62, ZN => n83);
   U57 : AOI222_X1 port map( A1 => n222, A2 => n212, B1 => n61, B2 => n68, C1 
                           => n63, C2 => n69, ZN => n86);
   U58 : AOI222_X1 port map( A1 => n63, A2 => n115, B1 => n129, B2 => n99, C1 
                           => n61, C2 => n116, ZN => n130);
   U59 : AOI222_X1 port map( A1 => n222, A2 => n207, B1 => n61, B2 => n74, C1 
                           => n63, C2 => n75, ZN => n73);
   U60 : AOI222_X1 port map( A1 => n63, A2 => n112, B1 => n129, B2 => n98, C1 
                           => n61, C2 => n114, ZN => n128);
   U61 : AND2_X1 port map( A1 => n99, A2 => n223, ZN => B(30));
   U62 : AND2_X1 port map( A1 => n106, A2 => n223, ZN => B(29));
   U63 : AND2_X1 port map( A1 => n107, A2 => n223, ZN => B(28));
   U64 : NOR3_X1 port map( A1 => n182, A2 => n171, A3 => n169, ZN => B(27));
   U65 : NOR2_X1 port map( A1 => n171, A2 => n108, ZN => B(26));
   U66 : NOR2_X1 port map( A1 => n172, A2 => n58, ZN => B(25));
   U67 : NOR2_X1 port map( A1 => n172, A2 => n66, ZN => B(24));
   U68 : NOR2_X1 port map( A1 => n172, A2 => n72, ZN => B(23));
   U69 : NOR2_X1 port map( A1 => n173, A2 => n77, ZN => B(22));
   U70 : NOR2_X1 port map( A1 => n173, A2 => n82, ZN => B(21));
   U71 : NOR2_X1 port map( A1 => n173, A2 => n85, ZN => B(20));
   U72 : NOR2_X1 port map( A1 => n173, A2 => n88, ZN => B(19));
   U73 : NOR2_X1 port map( A1 => n174, A2 => n100, ZN => B(18));
   U74 : NOR2_X1 port map( A1 => n172, A2 => n117, ZN => B(17));
   U75 : NOR2_X1 port map( A1 => n171, A2 => n127, ZN => B(16));
   U76 : OAI221_X1 port map( B1 => n193, B2 => n87, C1 => n199, C2 => n57, A =>
                           n128, ZN => B(15));
   U77 : OAI221_X1 port map( B1 => n194, B2 => n87, C1 => n201, C2 => n57, A =>
                           n130, ZN => B(14));
   U78 : OAI221_X1 port map( B1 => n196, B2 => n87, C1 => n203, C2 => n57, A =>
                           n131, ZN => B(13));
   U79 : INV_X1 port map( A => n136, ZN => B(12));
   U80 : OAI221_X1 port map( B1 => n199, B2 => n87, C1 => n91, C2 => n57, A => 
                           n139, ZN => B(11));
   U81 : OAI221_X1 port map( B1 => n103, B2 => n57, C1 => n108, C2 => n177, A 
                           => n146, ZN => B(10));
   U82 : OAI221_X1 port map( B1 => n76, B2 => n87, C1 => n100, C2 => n177, A =>
                           n101, ZN => B(2));
   U83 : OAI221_X1 port map( B1 => n81, B2 => n87, C1 => n117, C2 => n177, A =>
                           n118, ZN => B(1));
   U84 : OAI221_X1 port map( B1 => n56, B2 => n57, C1 => n58, C2 => n177, A => 
                           n59, ZN => B(9));
   U85 : OAI221_X1 port map( B1 => n65, B2 => n57, C1 => n66, C2 => n177, A => 
                           n67, ZN => B(8));
   U86 : OAI221_X1 port map( B1 => n71, B2 => n57, C1 => n72, C2 => n177, A => 
                           n73, ZN => B(7));
   U87 : OAI221_X1 port map( B1 => n76, B2 => n57, C1 => n77, C2 => n177, A => 
                           n78, ZN => B(6));
   U88 : OAI221_X1 port map( B1 => n81, B2 => n57, C1 => n82, C2 => n177, A => 
                           n83, ZN => B(5));
   U89 : OAI221_X1 port map( B1 => n84, B2 => n57, C1 => n85, C2 => n177, A => 
                           n86, ZN => B(4));
   U90 : OAI221_X1 port map( B1 => n71, B2 => n87, C1 => n88, C2 => n177, A => 
                           n89, ZN => B(3));
   U91 : AOI221_X1 port map( B1 => n63, B2 => n114, C1 => n61, C2 => n75, A => 
                           n140, ZN => n139);
   U92 : NOR3_X1 port map( A1 => n177, A2 => n169, A3 => n182, ZN => n140);
   U93 : AOI221_X1 port map( B1 => n69, B2 => n222, C1 => n68, C2 => n223, A =>
                           n179, ZN => n136);
   U94 : INV_X1 port map( A => n137, ZN => n179);
   U95 : AOI222_X1 port map( A1 => n63, A2 => n111, B1 => n129, B2 => n107, C1 
                           => n61, C2 => n70, ZN => n137);
   U96 : NOR2_X1 port map( A1 => n184, A2 => n227, ZN => n98);
   U97 : AOI22_X1 port map( A1 => n115, A2 => n224, B1 => n99, B2 => n110, ZN 
                           => n108);
   U98 : AOI22_X1 port map( A1 => n109, A2 => n224, B1 => n106, B2 => n110, ZN 
                           => n58);
   U99 : AOI22_X1 port map( A1 => n111, A2 => n224, B1 => n107, B2 => n110, ZN 
                           => n66);
   U100 : NAND2_X1 port map( A1 => SH(1), A2 => n167, ZN => n93);
   U101 : INV_X1 port map( A => n74, ZN => n199);
   U102 : INV_X1 port map( A => n103, ZN => n208);
   U103 : INV_X1 port map( A => n56, ZN => n210);
   U104 : INV_X1 port map( A => n65, ZN => n212);
   U105 : INV_X1 port map( A => n91, ZN => n207);
   U106 : INV_X1 port map( A => n80, ZN => n194);
   U107 : INV_X1 port map( A => n62, ZN => n196);
   U108 : INV_X1 port map( A => n75, ZN => n193);
   U109 : INV_X1 port map( A => n79, ZN => n201);
   U110 : INV_X1 port map( A => n60, ZN => n203);
   U111 : OAI221_X1 port map( B1 => n92, B2 => n184, C1 => n165, C2 => n185, A 
                           => n160, ZN => n107);
   U112 : AOI22_X1 port map( A1 => A(29), A2 => n95, B1 => A(28), B2 => n96, ZN
                           => n160);
   U113 : OAI221_X1 port map( B1 => n92, B2 => n195, C1 => n197, C2 => n165, A 
                           => n148, ZN => n80);
   U114 : AOI22_X1 port map( A1 => n95, A2 => A(19), B1 => n96, B2 => A(18), ZN
                           => n148);
   U115 : OAI221_X1 port map( B1 => n92, B2 => n197, C1 => n165, C2 => n198, A 
                           => n135, ZN => n62);
   U116 : AOI22_X1 port map( A1 => A(18), A2 => n95, B1 => A(17), B2 => n96, ZN
                           => n135);
   U117 : OAI221_X1 port map( B1 => n92, B2 => n198, C1 => n165, C2 => n200, A 
                           => n161, ZN => n69);
   U118 : AOI22_X1 port map( A1 => A(17), A2 => n95, B1 => A(16), B2 => n96, ZN
                           => n161);
   U119 : OAI221_X1 port map( B1 => n92, B2 => n202, C1 => n166, C2 => n204, A 
                           => n149, ZN => n79);
   U120 : AOI22_X1 port map( A1 => A(15), A2 => n95, B1 => A(14), B2 => n96, ZN
                           => n149);
   U121 : OAI221_X1 port map( B1 => n92, B2 => n204, C1 => n164, C2 => n205, A 
                           => n134, ZN => n60);
   U122 : AOI22_X1 port map( A1 => A(14), A2 => n95, B1 => A(13), B2 => n96, ZN
                           => n134);
   U123 : OAI221_X1 port map( B1 => n92, B2 => n205, C1 => n164, C2 => n206, A 
                           => n157, ZN => n68);
   U124 : INV_X1 port map( A => A(14), ZN => n206);
   U125 : AOI22_X1 port map( A1 => A(13), A2 => n95, B1 => A(12), B2 => n96, ZN
                           => n157);
   U126 : OAI221_X1 port map( B1 => n92, B2 => n186, C1 => n164, C2 => n187, A 
                           => n150, ZN => n115);
   U127 : AOI22_X1 port map( A1 => A(27), A2 => n95, B1 => A(26), B2 => n96, ZN
                           => n150);
   U128 : OAI221_X1 port map( B1 => n92, B2 => n187, C1 => n164, C2 => n188, A 
                           => n133, ZN => n109);
   U129 : AOI22_X1 port map( A1 => A(26), A2 => n95, B1 => A(25), B2 => n96, ZN
                           => n133);
   U130 : OAI221_X1 port map( B1 => n92, B2 => n188, C1 => n165, C2 => n189, A 
                           => n159, ZN => n111);
   U131 : AOI22_X1 port map( A1 => A(25), A2 => n95, B1 => A(24), B2 => n96, ZN
                           => n159);
   U132 : OAI221_X1 port map( B1 => n92, B2 => n190, C1 => n166, C2 => n191, A 
                           => n147, ZN => n116);
   U133 : AOI22_X1 port map( A1 => A(23), A2 => n95, B1 => A(22), B2 => n96, ZN
                           => n147);
   U134 : OAI221_X1 port map( B1 => n92, B2 => n191, C1 => n164, C2 => n192, A 
                           => n132, ZN => n64);
   U135 : INV_X1 port map( A => A(23), ZN => n192);
   U136 : AOI22_X1 port map( A1 => A(22), A2 => n95, B1 => A(21), B2 => n96, ZN
                           => n132);
   U137 : OAI221_X1 port map( B1 => n92, B2 => n189, C1 => n165, C2 => n190, A 
                           => n143, ZN => n114);
   U138 : AOI22_X1 port map( A1 => A(24), A2 => n95, B1 => A(23), B2 => n96, ZN
                           => n143);
   U139 : OAI221_X1 port map( B1 => n197, B2 => n228, C1 => n198, C2 => n227, A
                           => n142, ZN => n75);
   U140 : AOI22_X1 port map( A1 => A(22), A2 => n226, B1 => A(21), B2 => n225, 
                           ZN => n142);
   U142 : OAI221_X1 port map( B1 => n228, B2 => n195, C1 => n197, C2 => n227, A
                           => n162, ZN => n70);
   U143 : AOI22_X1 port map( A1 => A(23), A2 => n226, B1 => A(22), B2 => n225, 
                           ZN => n162);
   U144 : OAI221_X1 port map( B1 => n92, B2 => n200, C1 => n166, C2 => n202, A 
                           => n145, ZN => n74);
   U145 : AOI22_X1 port map( A1 => A(16), A2 => n95, B1 => A(15), B2 => n96, ZN
                           => n145);
   U146 : AOI221_X1 port map( B1 => n226, B2 => A(10), C1 => n225, C2 => A(9), 
                           A => n97, ZN => n71);
   U147 : OAI22_X1 port map( A1 => n215, A2 => n228, B1 => n216, B2 => n227, ZN
                           => n97);
   U148 : AOI221_X1 port map( B1 => n226, B2 => A(9), C1 => n225, C2 => A(8), A
                           => n105, ZN => n76);
   U149 : OAI22_X1 port map( A1 => n216, A2 => n228, B1 => n217, B2 => n227, ZN
                           => n105);
   U150 : AOI221_X1 port map( B1 => n226, B2 => A(8), C1 => n225, C2 => A(7), A
                           => n122, ZN => n81);
   U151 : OAI22_X1 port map( A1 => n217, A2 => n228, B1 => n218, B2 => n227, ZN
                           => n122);
   U152 : AOI221_X1 port map( B1 => n226, B2 => A(7), C1 => n225, C2 => A(6), A
                           => n163, ZN => n84);
   U153 : OAI22_X1 port map( A1 => n218, A2 => n228, B1 => n219, B2 => n227, ZN
                           => n163);
   U154 : AOI221_X1 port map( B1 => n226, B2 => A(13), C1 => n225, C2 => A(12),
                           A => n151, ZN => n103);
   U155 : OAI22_X1 port map( A1 => n211, A2 => n228, B1 => n213, B2 => n227, ZN
                           => n151);
   U156 : AOI221_X1 port map( B1 => n226, B2 => A(12), C1 => n225, C2 => A(11),
                           A => n120, ZN => n56);
   U157 : OAI22_X1 port map( A1 => n213, A2 => n228, B1 => n214, B2 => n227, ZN
                           => n120);
   U158 : AOI221_X1 port map( B1 => n226, B2 => A(11), C1 => n225, C2 => A(10),
                           A => n154, ZN => n65);
   U159 : OAI22_X1 port map( A1 => n214, A2 => n228, B1 => n215, B2 => n227, ZN
                           => n154);
   U160 : AOI221_X1 port map( B1 => n226, B2 => A(14), C1 => n225, C2 => A(13),
                           A => n144, ZN => n91);
   U161 : OAI22_X1 port map( A1 => n209, A2 => n228, B1 => n211, B2 => n227, ZN
                           => n144);
   U162 : INV_X1 port map( A => A(12), ZN => n209);
   U163 : OAI221_X1 port map( B1 => n92, B2 => n185, C1 => n165, C2 => n186, A 
                           => n141, ZN => n112);
   U164 : AOI22_X1 port map( A1 => A(28), A2 => n95, B1 => A(27), B2 => n96, ZN
                           => n141);
   U165 : AOI222_X1 port map( A1 => n63, A2 => n74, B1 => n223, B2 => n90, C1 
                           => n61, C2 => n207, ZN => n89);
   U166 : OAI221_X1 port map( B1 => n92, B2 => n217, C1 => n166, C2 => n218, A 
                           => n94, ZN => n90);
   U167 : AOI22_X1 port map( A1 => A(4), A2 => n95, B1 => A(3), B2 => n96, ZN 
                           => n94);
   U168 : AOI222_X1 port map( A1 => n63, A2 => n79, B1 => n223, B2 => n102, C1 
                           => n61, C2 => n208, ZN => n101);
   U169 : OAI221_X1 port map( B1 => n92, B2 => n218, C1 => n166, C2 => n219, A 
                           => n104, ZN => n102);
   U170 : AOI22_X1 port map( A1 => A(3), A2 => n95, B1 => A(2), B2 => n96, ZN 
                           => n104);
   U171 : AOI222_X1 port map( A1 => n63, A2 => n60, B1 => n223, B2 => n119, C1 
                           => n61, C2 => n210, ZN => n118);
   U172 : OAI221_X1 port map( B1 => n92, B2 => n219, C1 => n166, C2 => n220, A 
                           => n121, ZN => n119);
   U173 : AOI22_X1 port map( A1 => A(2), A2 => n95, B1 => A(1), B2 => n96, ZN 
                           => n121);
   U174 : OAI221_X1 port map( B1 => n84, B2 => n87, C1 => n127, C2 => n177, A 
                           => n152, ZN => B(0));
   U175 : AOI222_X1 port map( A1 => n63, A2 => n68, B1 => n223, B2 => n153, C1 
                           => n61, C2 => n212, ZN => n152);
   U176 : AND2_X1 port map( A1 => n223, A2 => n98, ZN => B(31));
   U177 : OAI221_X1 port map( B1 => n92, B2 => n220, C1 => n164, C2 => n221, A 
                           => n156, ZN => n153);
   U178 : INV_X1 port map( A => A(2), ZN => n221);
   U179 : AOI22_X1 port map( A1 => A(1), A2 => n95, B1 => A(0), B2 => n96, ZN 
                           => n156);
   U180 : INV_X1 port map( A => A(31), ZN => n184);
   U181 : INV_X1 port map( A => A(20), ZN => n197);
   U182 : INV_X1 port map( A => A(5), ZN => n218);
   U183 : INV_X1 port map( A => A(30), ZN => n185);
   U184 : INV_X1 port map( A => A(4), ZN => n219);
   U185 : INV_X1 port map( A => A(6), ZN => n217);
   U186 : INV_X1 port map( A => A(29), ZN => n186);
   U187 : INV_X1 port map( A => A(19), ZN => n198);
   U188 : INV_X1 port map( A => A(17), ZN => n202);
   U189 : INV_X1 port map( A => A(16), ZN => n204);
   U190 : INV_X1 port map( A => A(15), ZN => n205);
   U191 : INV_X1 port map( A => A(21), ZN => n195);
   U192 : INV_X1 port map( A => A(9), ZN => n214);
   U193 : INV_X1 port map( A => A(11), ZN => n211);
   U194 : INV_X1 port map( A => A(10), ZN => n213);
   U195 : INV_X1 port map( A => A(8), ZN => n215);
   U196 : INV_X1 port map( A => A(7), ZN => n216);
   U197 : INV_X1 port map( A => A(3), ZN => n220);
   U198 : INV_X1 port map( A => A(28), ZN => n187);
   U199 : INV_X1 port map( A => A(27), ZN => n188);
   U200 : INV_X1 port map( A => A(26), ZN => n189);
   U201 : INV_X1 port map( A => A(25), ZN => n190);
   U202 : INV_X1 port map( A => A(24), ZN => n191);
   U203 : INV_X1 port map( A => A(18), ZN => n200);
   U204 : INV_X1 port map( A => SH(0), ZN => n167);
   U205 : INV_X1 port map( A => SH(2), ZN => n168);
   U206 : INV_X1 port map( A => n170, ZN => n169);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_sla_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sla_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sla_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251 : std_logic;

begin
   B <= ( B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, A(0) );
   
   U10 : NOR2_X2 port map( A1 => n189, A2 => SH(3), ZN => n114);
   U12 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n116);
   U181 : MUX2_X1 port map( A => A(0), B => A(1), S => n178, Z => n119);
   U2 : NAND2_X1 port map( A1 => n196, A2 => A(0), ZN => n62);
   U3 : INV_X1 port map( A => n196, ZN => n192);
   U4 : INV_X1 port map( A => n69, ZN => n250);
   U5 : NAND2_X1 port map( A1 => n114, A2 => n192, ZN => n69);
   U6 : INV_X1 port map( A => n100, ZN => n251);
   U7 : BUF_X1 port map( A => n190, Z => n193);
   U8 : BUF_X1 port map( A => n191, Z => n195);
   U9 : BUF_X1 port map( A => n190, Z => n194);
   U11 : BUF_X1 port map( A => n191, Z => n196);
   U13 : NAND2_X1 port map( A1 => n116, A2 => n192, ZN => n100);
   U14 : AND2_X1 port map( A1 => n152, A2 => n189, ZN => n75);
   U15 : AND2_X1 port map( A1 => SH(3), A2 => n189, ZN => n118);
   U16 : BUF_X1 port map( A => n80, Z => n180);
   U17 : BUF_X1 port map( A => n80, Z => n179);
   U18 : BUF_X1 port map( A => n77, Z => n186);
   U19 : BUF_X1 port map( A => n77, Z => n185);
   U20 : BUF_X1 port map( A => n175, Z => n177);
   U21 : BUF_X1 port map( A => n175, Z => n176);
   U22 : BUF_X1 port map( A => n78, Z => n182);
   U23 : BUF_X1 port map( A => n78, Z => n183);
   U24 : BUF_X1 port map( A => n175, Z => n178);
   U25 : BUF_X1 port map( A => n80, Z => n181);
   U26 : BUF_X1 port map( A => n77, Z => n187);
   U27 : BUF_X1 port map( A => n78, Z => n184);
   U28 : AND2_X1 port map( A1 => SH(3), A2 => n192, ZN => n152);
   U29 : BUF_X1 port map( A => SH(4), Z => n191);
   U30 : BUF_X1 port map( A => SH(4), Z => n190);
   U31 : AND2_X1 port map( A1 => n152, A2 => SH(2), ZN => n72);
   U32 : AOI221_X1 port map( B1 => n125, B2 => n114, C1 => n126, C2 => n116, A 
                           => n249, ZN => n63);
   U33 : AOI221_X1 port map( B1 => n131, B2 => n114, C1 => n132, C2 => n116, A 
                           => n249, ZN => n64);
   U34 : AOI221_X1 port map( B1 => n244, B2 => n114, C1 => n136, C2 => n116, A 
                           => n249, ZN => n65);
   U35 : AOI221_X1 port map( B1 => n119, B2 => n114, C1 => n113, C2 => n116, A 
                           => n249, ZN => n66);
   U36 : AOI221_X1 port map( B1 => n130, B2 => n114, C1 => n103, C2 => n116, A 
                           => n234, ZN => n70);
   U37 : INV_X1 port map( A => n154, ZN => n234);
   U38 : AOI22_X1 port map( A1 => n155, A2 => n131, B1 => n118, B2 => n132, ZN 
                           => n154);
   U39 : AOI221_X1 port map( B1 => n135, B2 => n114, C1 => n108, C2 => n116, A 
                           => n236, ZN => n81);
   U40 : INV_X1 port map( A => n157, ZN => n236);
   U41 : AOI22_X1 port map( A1 => n155, A2 => n244, B1 => n118, B2 => n136, ZN 
                           => n157);
   U42 : AOI221_X1 port map( B1 => n119, B2 => n155, C1 => n113, C2 => n118, A 
                           => n226, ZN => n88);
   U43 : INV_X1 port map( A => n159, ZN => n226);
   U44 : AOI22_X1 port map( A1 => n114, A2 => n115, B1 => n116, B2 => n112, ZN 
                           => n159);
   U45 : AOI221_X1 port map( B1 => n126, B2 => n114, C1 => n124, C2 => n116, A 
                           => n239, ZN => n94);
   U46 : INV_X1 port map( A => n163, ZN => n239);
   U47 : AOI21_X1 port map( B1 => n118, B2 => n125, A => n120, ZN => n163);
   U48 : AOI221_X1 port map( B1 => n132, B2 => n114, C1 => n130, C2 => n116, A 
                           => n241, ZN => n101);
   U49 : INV_X1 port map( A => n167, ZN => n241);
   U50 : AOI21_X1 port map( B1 => n118, B2 => n131, A => n120, ZN => n167);
   U51 : AOI221_X1 port map( B1 => n136, B2 => n114, C1 => n135, C2 => n116, A 
                           => n243, ZN => n106);
   U52 : INV_X1 port map( A => n171, ZN => n243);
   U53 : AOI21_X1 port map( B1 => n118, B2 => n244, A => n120, ZN => n171);
   U54 : AOI221_X1 port map( B1 => n113, B2 => n114, C1 => n115, C2 => n116, A 
                           => n246, ZN => n61);
   U55 : INV_X1 port map( A => n117, ZN => n246);
   U56 : AOI21_X1 port map( B1 => n118, B2 => n119, A => n120, ZN => n117);
   U57 : AOI222_X1 port map( A1 => n250, A2 => n76, B1 => n75, B2 => n73, C1 =>
                           n72, C2 => n103, ZN => n102);
   U58 : AOI222_X1 port map( A1 => n250, A2 => n85, B1 => n75, B2 => n83, C1 =>
                           n72, C2 => n108, ZN => n107);
   U59 : AOI222_X1 port map( A1 => n250, A2 => n92, B1 => n75, B2 => n90, C1 =>
                           n72, C2 => n112, ZN => n111);
   U60 : AOI222_X1 port map( A1 => n250, A2 => n98, B1 => n75, B2 => n96, C1 =>
                           n72, C2 => n124, ZN => n123);
   U61 : AOI222_X1 port map( A1 => n250, A2 => n73, B1 => n75, B2 => n103, C1 
                           => n72, C2 => n130, ZN => n129);
   U62 : AOI222_X1 port map( A1 => n250, A2 => n83, B1 => n75, B2 => n108, C1 
                           => n72, C2 => n135, ZN => n134);
   U63 : AOI222_X1 port map( A1 => n250, A2 => n90, B1 => n75, B2 => n112, C1 
                           => n72, C2 => n115, ZN => n138);
   U64 : AOI222_X1 port map( A1 => n250, A2 => n96, B1 => n75, B2 => n124, C1 
                           => n72, C2 => n126, ZN => n141);
   U65 : AOI222_X1 port map( A1 => n250, A2 => n103, B1 => n75, B2 => n130, C1 
                           => n72, C2 => n132, ZN => n145);
   U66 : AOI222_X1 port map( A1 => n250, A2 => n108, B1 => n75, B2 => n135, C1 
                           => n72, C2 => n136, ZN => n147);
   U67 : AOI222_X1 port map( A1 => n250, A2 => n112, B1 => n75, B2 => n115, C1 
                           => n72, C2 => n113, ZN => n149);
   U68 : OAI221_X1 port map( B1 => n202, B2 => n69, C1 => n81, C2 => n192, A =>
                           n82, ZN => B_30_port);
   U69 : OAI221_X1 port map( B1 => n204, B2 => n69, C1 => n88, C2 => n192, A =>
                           n89, ZN => B_29_port);
   U70 : OAI221_X1 port map( B1 => n206, B2 => n69, C1 => n94, C2 => n192, A =>
                           n95, ZN => B_28_port);
   U71 : OAI221_X1 port map( B1 => n200, B2 => n100, C1 => n101, C2 => n192, A 
                           => n102, ZN => B_27_port);
   U72 : OAI221_X1 port map( B1 => n202, B2 => n100, C1 => n106, C2 => n192, A 
                           => n107, ZN => B_26_port);
   U73 : OAI221_X1 port map( B1 => n204, B2 => n100, C1 => n61, C2 => n192, A 
                           => n111, ZN => B_25_port);
   U74 : OAI221_X1 port map( B1 => n206, B2 => n100, C1 => n63, C2 => n192, A 
                           => n123, ZN => B_24_port);
   U75 : OAI221_X1 port map( B1 => n208, B2 => n100, C1 => n64, C2 => n192, A 
                           => n129, ZN => B_23_port);
   U76 : OAI221_X1 port map( B1 => n210, B2 => n100, C1 => n65, C2 => n192, A 
                           => n134, ZN => B_22_port);
   U77 : OAI221_X1 port map( B1 => n212, B2 => n100, C1 => n66, C2 => n192, A 
                           => n138, ZN => B_21_port);
   U78 : OAI221_X1 port map( B1 => n214, B2 => n100, C1 => n67, C2 => n192, A 
                           => n141, ZN => B_20_port);
   U79 : OAI221_X1 port map( B1 => n216, B2 => n100, C1 => n68, C2 => n192, A 
                           => n145, ZN => B_19_port);
   U80 : OAI221_X1 port map( B1 => n218, B2 => n100, C1 => n87, C2 => n192, A 
                           => n147, ZN => B_18_port);
   U81 : OAI221_X1 port map( B1 => n220, B2 => n100, C1 => n144, C2 => n192, A 
                           => n149, ZN => B_17_port);
   U82 : OAI221_X1 port map( B1 => n228, B2 => n69, C1 => n222, C2 => n100, A 
                           => n151, ZN => B_16_port);
   U83 : OAI21_X1 port map( B1 => n193, B2 => n70, A => n62, ZN => B_15_port);
   U84 : OAI21_X1 port map( B1 => n193, B2 => n81, A => n62, ZN => B_14_port);
   U85 : OAI21_X1 port map( B1 => n194, B2 => n88, A => n62, ZN => B_13_port);
   U86 : OAI21_X1 port map( B1 => n193, B2 => n94, A => n62, ZN => B_12_port);
   U87 : OAI21_X1 port map( B1 => n193, B2 => n101, A => n62, ZN => B_11_port);
   U88 : OAI21_X1 port map( B1 => n193, B2 => n106, A => n62, ZN => B_10_port);
   U89 : OAI21_X1 port map( B1 => n194, B2 => n87, A => n62, ZN => B_2_port);
   U90 : OAI21_X1 port map( B1 => n194, B2 => n144, A => n62, ZN => B_1_port);
   U91 : OAI21_X1 port map( B1 => n195, B2 => n61, A => n62, ZN => B_9_port);
   U92 : OAI21_X1 port map( B1 => n195, B2 => n63, A => n62, ZN => B_8_port);
   U93 : OAI21_X1 port map( B1 => n195, B2 => n64, A => n62, ZN => B_7_port);
   U94 : OAI21_X1 port map( B1 => n195, B2 => n65, A => n62, ZN => B_6_port);
   U95 : OAI21_X1 port map( B1 => n195, B2 => n66, A => n62, ZN => B_5_port);
   U96 : OAI21_X1 port map( B1 => n194, B2 => n67, A => n62, ZN => B_4_port);
   U97 : OAI21_X1 port map( B1 => n194, B2 => n68, A => n62, ZN => B_3_port);
   U98 : OAI21_X1 port map( B1 => n247, B2 => n189, A => n139, ZN => n142);
   U99 : AOI221_X1 port map( B1 => n72, B2 => n125, C1 => n75, C2 => n126, A =>
                           n248, ZN => n151);
   U100 : INV_X1 port map( A => n62, ZN => n248);
   U101 : NOR2_X1 port map( A1 => n189, A2 => n139, ZN => n120);
   U102 : AOI21_X1 port map( B1 => n125, B2 => n116, A => n142, ZN => n67);
   U103 : AOI21_X1 port map( B1 => n131, B2 => n116, A => n142, ZN => n68);
   U104 : AOI21_X1 port map( B1 => n244, B2 => n116, A => n142, ZN => n87);
   U105 : AOI21_X1 port map( B1 => n119, B2 => n116, A => n142, ZN => n144);
   U106 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n78);
   U107 : NAND2_X1 port map( A1 => SH(1), A2 => n188, ZN => n77);
   U108 : INV_X1 port map( A => n139, ZN => n249);
   U109 : NOR2_X1 port map( A1 => n188, A2 => SH(1), ZN => n80);
   U110 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n155);
   U111 : INV_X1 port map( A => n124, ZN => n228);
   U112 : INV_X1 port map( A => n73, ZN => n216);
   U113 : INV_X1 port map( A => n83, ZN => n218);
   U114 : INV_X1 port map( A => n90, ZN => n220);
   U115 : INV_X1 port map( A => n96, ZN => n222);
   U116 : NOR2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n175);
   U117 : INV_X1 port map( A => n76, ZN => n208);
   U118 : INV_X1 port map( A => n85, ZN => n210);
   U119 : INV_X1 port map( A => n92, ZN => n212);
   U120 : INV_X1 port map( A => n98, ZN => n214);
   U121 : OAI221_X1 port map( B1 => n185, B2 => n229, C1 => n182, C2 => n230, A
                           => n160, ZN => n112);
   U122 : AOI22_X1 port map( A1 => A(12), A2 => n179, B1 => A(13), B2 => n176, 
                           ZN => n160);
   U123 : OAI221_X1 port map( B1 => n185, B2 => n233, C1 => n182, C2 => n235, A
                           => n161, ZN => n115);
   U124 : AOI22_X1 port map( A1 => A(8), A2 => n179, B1 => A(9), B2 => n176, ZN
                           => n161);
   U125 : OAI221_X1 port map( B1 => n245, B2 => n187, C1 => n247, C2 => n182, A
                           => n168, ZN => n131);
   U126 : AOI22_X1 port map( A1 => n181, A2 => A(2), B1 => A(3), B2 => n176, ZN
                           => n168);
   U127 : OAI221_X1 port map( B1 => n187, B2 => n235, C1 => n184, C2 => n237, A
                           => n166, ZN => n126);
   U128 : AOI22_X1 port map( A1 => A(7), A2 => n179, B1 => A(8), B2 => n176, ZN
                           => n166);
   U129 : OAI221_X1 port map( B1 => n187, B2 => n237, C1 => n184, C2 => n238, A
                           => n170, ZN => n132);
   U130 : AOI22_X1 port map( A1 => A(6), A2 => n179, B1 => A(7), B2 => n176, ZN
                           => n170);
   U131 : OAI221_X1 port map( B1 => n186, B2 => n238, C1 => n240, C2 => n182, A
                           => n174, ZN => n136);
   U132 : AOI22_X1 port map( A1 => A(5), A2 => n180, B1 => A(6), B2 => n176, ZN
                           => n174);
   U133 : OAI221_X1 port map( B1 => n185, B2 => n230, C1 => n184, C2 => n231, A
                           => n165, ZN => n124);
   U134 : AOI22_X1 port map( A1 => A(11), A2 => n179, B1 => A(12), B2 => n176, 
                           ZN => n165);
   U135 : OAI221_X1 port map( B1 => n187, B2 => n231, C1 => n184, C2 => n232, A
                           => n169, ZN => n130);
   U136 : AOI22_X1 port map( A1 => A(10), A2 => n179, B1 => A(11), B2 => n176, 
                           ZN => n169);
   U137 : OAI221_X1 port map( B1 => n187, B2 => n232, C1 => n184, C2 => n233, A
                           => n173, ZN => n135);
   U138 : AOI22_X1 port map( A1 => A(9), A2 => n179, B1 => A(10), B2 => n176, 
                           ZN => n173);
   U139 : OAI221_X1 port map( B1 => n185, B2 => n219, C1 => n182, C2 => n221, A
                           => n146, ZN => n73);
   U140 : AOI22_X1 port map( A1 => A(18), A2 => n180, B1 => A(19), B2 => n177, 
                           ZN => n146);
   U141 : OAI221_X1 port map( B1 => n185, B2 => n221, C1 => n182, C2 => n223, A
                           => n148, ZN => n83);
   U142 : AOI22_X1 port map( A1 => A(17), A2 => n180, B1 => A(18), B2 => n177, 
                           ZN => n148);
   U143 : OAI221_X1 port map( B1 => n185, B2 => n223, C1 => n182, C2 => n224, A
                           => n150, ZN => n90);
   U144 : AOI22_X1 port map( A1 => A(16), A2 => n180, B1 => A(17), B2 => n177, 
                           ZN => n150);
   U145 : OAI221_X1 port map( B1 => n185, B2 => n224, C1 => n182, C2 => n225, A
                           => n153, ZN => n96);
   U146 : AOI22_X1 port map( A1 => A(15), A2 => n179, B1 => A(16), B2 => n177, 
                           ZN => n153);
   U147 : OAI221_X1 port map( B1 => n185, B2 => n225, C1 => n182, C2 => n227, A
                           => n156, ZN => n103);
   U148 : AOI22_X1 port map( A1 => A(14), A2 => n179, B1 => A(15), B2 => n177, 
                           ZN => n156);
   U149 : OAI221_X1 port map( B1 => n185, B2 => n227, C1 => n182, C2 => n229, A
                           => n158, ZN => n108);
   U150 : AOI22_X1 port map( A1 => A(13), A2 => n179, B1 => A(14), B2 => n176, 
                           ZN => n158);
   U151 : OAI221_X1 port map( B1 => n185, B2 => n242, C1 => n245, C2 => n182, A
                           => n164, ZN => n125);
   U152 : AOI22_X1 port map( A1 => n181, A2 => A(3), B1 => A(4), B2 => n176, ZN
                           => n164);
   U153 : OAI221_X1 port map( B1 => n185, B2 => n240, C1 => n182, C2 => n242, A
                           => n162, ZN => n113);
   U154 : AOI22_X1 port map( A1 => A(4), A2 => n179, B1 => A(5), B2 => n176, ZN
                           => n162);
   U155 : OAI221_X1 port map( B1 => n186, B2 => n211, C1 => n183, C2 => n213, A
                           => n133, ZN => n76);
   U156 : AOI22_X1 port map( A1 => A(22), A2 => n180, B1 => A(23), B2 => n177, 
                           ZN => n133);
   U157 : OAI221_X1 port map( B1 => n186, B2 => n213, C1 => n183, C2 => n215, A
                           => n137, ZN => n85);
   U158 : AOI22_X1 port map( A1 => A(21), A2 => n180, B1 => A(22), B2 => n177, 
                           ZN => n137);
   U159 : OAI221_X1 port map( B1 => n186, B2 => n215, C1 => n183, C2 => n217, A
                           => n140, ZN => n92);
   U160 : AOI22_X1 port map( A1 => A(20), A2 => n180, B1 => A(21), B2 => n177, 
                           ZN => n140);
   U161 : OAI221_X1 port map( B1 => n185, B2 => n217, C1 => n183, C2 => n219, A
                           => n143, ZN => n98);
   U162 : AOI22_X1 port map( A1 => A(19), A2 => n180, B1 => A(20), B2 => n177, 
                           ZN => n143);
   U163 : AOI222_X1 port map( A1 => n72, A2 => n83, B1 => n251, B2 => n84, C1 
                           => n75, C2 => n85, ZN => n82);
   U164 : OAI221_X1 port map( B1 => n186, B2 => n198, C1 => n183, C2 => n199, A
                           => n86, ZN => n84);
   U165 : AOI22_X1 port map( A1 => A(29), A2 => n181, B1 => A(30), B2 => n178, 
                           ZN => n86);
   U166 : AOI222_X1 port map( A1 => n72, A2 => n90, B1 => n251, B2 => n91, C1 
                           => n75, C2 => n92, ZN => n89);
   U167 : OAI221_X1 port map( B1 => n186, B2 => n199, C1 => n183, C2 => n201, A
                           => n93, ZN => n91);
   U168 : AOI22_X1 port map( A1 => A(28), A2 => n181, B1 => A(29), B2 => n178, 
                           ZN => n93);
   U169 : AOI222_X1 port map( A1 => n72, A2 => n96, B1 => n251, B2 => n97, C1 
                           => n75, C2 => n98, ZN => n95);
   U170 : OAI221_X1 port map( B1 => n186, B2 => n201, C1 => n183, C2 => n203, A
                           => n99, ZN => n97);
   U171 : AOI22_X1 port map( A1 => A(27), A2 => n181, B1 => A(28), B2 => n178, 
                           ZN => n99);
   U172 : OAI221_X1 port map( B1 => n200, B2 => n69, C1 => n70, C2 => n192, A 
                           => n71, ZN => B_31_port);
   U173 : AOI222_X1 port map( A1 => n72, A2 => n73, B1 => n251, B2 => n74, C1 
                           => n75, C2 => n76, ZN => n71);
   U174 : OAI221_X1 port map( B1 => n186, B2 => n197, C1 => n183, C2 => n198, A
                           => n79, ZN => n74);
   U175 : INV_X1 port map( A => A(29), ZN => n197);
   U176 : AOI22_X1 port map( A1 => A(30), A2 => n179, B1 => A(31), B2 => n177, 
                           ZN => n79);
   U177 : NAND2_X1 port map( A1 => SH(3), A2 => A(0), ZN => n139);
   U178 : INV_X1 port map( A => n172, ZN => n244);
   U179 : AOI222_X1 port map( A1 => n178, A2 => A(2), B1 => A(1), B2 => n181, 
                           C1 => A(0), C2 => SH(1), ZN => n172);
   U180 : INV_X1 port map( A => A(12), ZN => n227);
   U182 : INV_X1 port map( A => A(13), ZN => n225);
   U183 : INV_X1 port map( A => A(14), ZN => n224);
   U184 : INV_X1 port map( A => A(23), ZN => n207);
   U185 : INV_X1 port map( A => A(22), ZN => n209);
   U186 : INV_X1 port map( A => A(17), ZN => n219);
   U187 : INV_X1 port map( A => A(16), ZN => n221);
   U188 : INV_X1 port map( A => A(15), ZN => n223);
   U189 : INV_X1 port map( A => A(21), ZN => n211);
   U190 : INV_X1 port map( A => A(9), ZN => n231);
   U191 : INV_X1 port map( A => A(11), ZN => n229);
   U192 : INV_X1 port map( A => A(10), ZN => n230);
   U193 : INV_X1 port map( A => A(8), ZN => n232);
   U194 : INV_X1 port map( A => A(7), ZN => n233);
   U195 : INV_X1 port map( A => A(2), ZN => n242);
   U196 : INV_X1 port map( A => A(28), ZN => n198);
   U197 : INV_X1 port map( A => A(27), ZN => n199);
   U198 : INV_X1 port map( A => A(26), ZN => n201);
   U199 : INV_X1 port map( A => A(25), ZN => n203);
   U200 : INV_X1 port map( A => A(24), ZN => n205);
   U201 : INV_X1 port map( A => A(3), ZN => n240);
   U202 : INV_X1 port map( A => A(18), ZN => n217);
   U203 : INV_X1 port map( A => A(0), ZN => n247);
   U204 : INV_X1 port map( A => A(6), ZN => n235);
   U205 : INV_X1 port map( A => A(4), ZN => n238);
   U206 : INV_X1 port map( A => A(1), ZN => n245);
   U207 : INV_X1 port map( A => A(19), ZN => n215);
   U208 : INV_X1 port map( A => A(20), ZN => n213);
   U209 : INV_X1 port map( A => A(5), ZN => n237);
   U210 : INV_X1 port map( A => n127, ZN => n206);
   U211 : OAI221_X1 port map( B1 => n186, B2 => n209, C1 => n183, C2 => n211, A
                           => n128, ZN => n127);
   U212 : AOI22_X1 port map( A1 => A(23), A2 => n180, B1 => A(24), B2 => n177, 
                           ZN => n128);
   U213 : INV_X1 port map( A => n104, ZN => n200);
   U214 : OAI221_X1 port map( B1 => n186, B2 => n203, C1 => n183, C2 => n205, A
                           => n105, ZN => n104);
   U215 : AOI22_X1 port map( A1 => A(26), A2 => n180, B1 => A(27), B2 => n178, 
                           ZN => n105);
   U216 : INV_X1 port map( A => n109, ZN => n202);
   U217 : OAI221_X1 port map( B1 => n186, B2 => n205, C1 => n183, C2 => n207, A
                           => n110, ZN => n109);
   U218 : AOI22_X1 port map( A1 => A(25), A2 => n180, B1 => A(26), B2 => n178, 
                           ZN => n110);
   U219 : INV_X1 port map( A => n121, ZN => n204);
   U220 : OAI221_X1 port map( B1 => n186, B2 => n207, C1 => n183, C2 => n209, A
                           => n122, ZN => n121);
   U221 : AOI22_X1 port map( A1 => A(24), A2 => n180, B1 => A(25), B2 => n177, 
                           ZN => n122);
   U222 : INV_X1 port map( A => SH(0), ZN => n188);
   U223 : INV_X1 port map( A => SH(2), ZN => n189);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW01_ash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW01_ash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40
      , n41, n42, n43 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n34, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n34, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n34, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n34, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n34, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n34, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => SH(4), Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n34, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => n36, S => SH(4), Z 
                           => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => n37, S => n34, Z => 
                           B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => n38, S => SH(4), Z 
                           => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => n39, S => n34, Z => 
                           B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => n40, S => SH(4), Z 
                           => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => n41, S => SH(4), Z 
                           => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => n42, S => SH(4), Z 
                           => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => n43, S => SH(4), Z 
                           => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n32, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n32, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n32, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n32, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n32, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n32, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n32, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n32, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n32, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => SH(3), Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n32, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n32, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n32, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n32, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n32, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n32, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n32, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n32, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n32, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n32, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n32, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n32, Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => n30, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n29, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n30, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => n29, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n30, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n29, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n30, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n30, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n30, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n30, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n30, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n30, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => n30, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n30, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => n30, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n30, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n30, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n29, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n29, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n29, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => n29, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n29, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n29, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n29, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n29, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n29, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n29, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n29, Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => n27, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => n26, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => n27, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => n26, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n27, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => n26, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => n27, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => n26, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => n27, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n27, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => n27, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => n27, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n27, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n27, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => n27, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n27, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => n27, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n27, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n27, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n26, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n26, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n26, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n26, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n26, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n26, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n26, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n26, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n26, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n26, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n26, Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n24, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n23, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n24, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n23, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n24, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n23, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n24, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n23, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n24, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n24, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n24, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n24, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n24, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n24, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n24, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n24, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n24, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n24, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n24, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n24, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n23, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n23, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n23, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n23, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n23, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n23, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n23, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n23, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n23, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n23, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n23, Z => 
                           ML_int_1_1_port);
   U3 : INV_X1 port map( A => n15, ZN => n36);
   U4 : INV_X1 port map( A => n16, ZN => n37);
   U5 : INV_X1 port map( A => n17, ZN => n38);
   U6 : INV_X1 port map( A => n18, ZN => n39);
   U7 : INV_X1 port map( A => n19, ZN => n40);
   U8 : INV_X1 port map( A => n20, ZN => n41);
   U9 : INV_X1 port map( A => n21, ZN => n42);
   U10 : INV_X1 port map( A => n22, ZN => n43);
   U11 : INV_X1 port map( A => n33, ZN => n32);
   U12 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n33, ZN => n15);
   U13 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n33, ZN => n16);
   U14 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n33, ZN => n17);
   U15 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n33, ZN => n18);
   U16 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n33, ZN => n19);
   U17 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n33, ZN => n20);
   U18 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n33, ZN => n21);
   U19 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n33, ZN => n22);
   U20 : INV_X1 port map( A => n25, ZN => n24);
   U21 : INV_X1 port map( A => n25, ZN => n23);
   U22 : INV_X1 port map( A => n28, ZN => n27);
   U23 : INV_X1 port map( A => n28, ZN => n26);
   U24 : INV_X1 port map( A => n31, ZN => n30);
   U25 : INV_X1 port map( A => SH(4), ZN => n35);
   U26 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n31, ZN => 
                           ML_int_3_3_port);
   U27 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n31, ZN => 
                           ML_int_3_2_port);
   U28 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n31, ZN => 
                           ML_int_3_1_port);
   U29 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n31, ZN => 
                           ML_int_3_0_port);
   U30 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n35, ZN => B(15));
   U31 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n35, ZN => B(14));
   U32 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n35, ZN => B(13));
   U33 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n35, ZN => B(12));
   U34 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n35, ZN => B(11));
   U35 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n35, ZN => B(10));
   U36 : NOR2_X1 port map( A1 => n34, A2 => n20, ZN => B(2));
   U37 : NOR2_X1 port map( A1 => n34, A2 => n21, ZN => B(1));
   U38 : NOR2_X1 port map( A1 => n34, A2 => n22, ZN => B(0));
   U39 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n35, ZN => B(9));
   U40 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n35, ZN => B(8));
   U41 : NOR2_X1 port map( A1 => n34, A2 => n15, ZN => B(7));
   U42 : NOR2_X1 port map( A1 => n34, A2 => n16, ZN => B(6));
   U43 : NOR2_X1 port map( A1 => n34, A2 => n17, ZN => B(5));
   U44 : NOR2_X1 port map( A1 => n34, A2 => n18, ZN => B(4));
   U45 : NOR2_X1 port map( A1 => n34, A2 => n19, ZN => B(3));
   U46 : INV_X1 port map( A => SH(0), ZN => n25);
   U47 : INV_X1 port map( A => SH(1), ZN => n28);
   U48 : INV_X1 port map( A => SH(2), ZN => n31);
   U49 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n28, ZN => 
                           ML_int_2_1_port);
   U50 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n28, ZN => 
                           ML_int_2_0_port);
   U51 : AND2_X1 port map( A1 => A(0), A2 => n25, ZN => ML_int_1_0_port);
   U52 : INV_X1 port map( A => n31, ZN => n29);
   U53 : INV_X1 port map( A => SH(3), ZN => n33);
   U54 : INV_X1 port map( A => n35, ZN => n34);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_574 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_574;

architecture SYN_ARCH2 of ND2_574 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0;

architecture SYN_ARCH2 of ND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_64 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_64;

architecture SYN_STRUCTURAL of MUX21_64 is

   component ND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_64
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_64 port map( A => S, Y => SB);
   UND1 : ND2_192 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_191 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_190 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P4_ADDER_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4_ADDER_NBIT32;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32 is

   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal Cout_gen_6_port, Cout_gen_5_port, Cout_gen_4_port, Cout_gen_3_port, 
      Cout_gen_2_port, Cout_gen_1_port, Cout_gen_0_port : std_logic;

begin
   
   carry_logic : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 port map( A(31) => 
                           A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           Cin => Cin, Co(7) => Cout, Co(6) => Cout_gen_6_port,
                           Co(5) => Cout_gen_5_port, Co(4) => Cout_gen_4_port, 
                           Co(3) => Cout_gen_3_port, Co(2) => Cout_gen_2_port, 
                           Co(1) => Cout_gen_1_port, Co(0) => Cout_gen_0_port);
   sum_logic : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31),
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           Cout_gen_6_port, Ci(6) => Cout_gen_5_port, Ci(5) => 
                           Cout_gen_4_port, Ci(4) => Cout_gen_3_port, Ci(3) => 
                           Cout_gen_2_port, Ci(2) => Cout_gen_1_port, Ci(1) => 
                           Cout_gen_0_port, Ci(0) => Cin, S(31) => S(31), S(30)
                           => S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
         downto 0);  LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE : in std_logic;  
         OUTPUT : out std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32;

architecture SYN_BEHAVIORAL of SHIFTER_GENERIC_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_lbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sla_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   signal N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, 
      N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35
      , N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, 
      N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64
      , N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109, N110, N111,
      N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, 
      N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, 
      N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, 
      N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N202, N203, N204, 
      N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, 
      N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, 
      N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, 
      N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, 
      N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, 
      N265, n1, n2, n3, n4, n5, n6, n10_port, n11_port, n12_port, n19_port, 
      n20_port, n21_port, n22_port, n23_port, n24_port, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, 
      n62_port, n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, 
      n69_port, n70_port, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105_port, n106_port, 
      n107_port, n108_port : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';
   n6 <= '0';
   sll_49 : SHIFTER_GENERIC_N32_DW01_ash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n1, SH(4) => 
                           n105_port, SH(3) => n104, SH(2) => B(2), SH(1) => 
                           B(1), SH(0) => B(0), SH_TC => n1, B(31) => N265, 
                           B(30) => N264, B(29) => N263, B(28) => N262, B(27) 
                           => N261, B(26) => N260, B(25) => N259, B(24) => N258
                           , B(23) => N257, B(22) => N256, B(21) => N255, B(20)
                           => N254, B(19) => N253, B(18) => N252, B(17) => N251
                           , B(16) => N250, B(15) => N249, B(14) => N248, B(13)
                           => N247, B(12) => N246, B(11) => N245, B(10) => N244
                           , B(9) => N243, B(8) => N242, B(7) => N241, B(6) => 
                           N240, B(5) => N239, B(4) => N238, B(3) => N237, B(2)
                           => N236, B(1) => N235, B(0) => N234);
   sla_47 : SHIFTER_GENERIC_N32_DW_sla_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n105_port, SH(3) => 
                           n104, SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), 
                           SH_TC => n2, B(31) => N233, B(30) => N232, B(29) => 
                           N231, B(28) => N230, B(27) => N229, B(26) => N228, 
                           B(25) => N227, B(24) => N226, B(23) => N225, B(22) 
                           => N224, B(21) => N223, B(20) => N222, B(19) => N221
                           , B(18) => N220, B(17) => N219, B(16) => N218, B(15)
                           => N217, B(14) => N216, B(13) => N215, B(12) => N214
                           , B(11) => N213, B(10) => N212, B(9) => N211, B(8) 
                           => N210, B(7) => N209, B(6) => N208, B(5) => N207, 
                           B(4) => N206, B(3) => N205, B(2) => N204, B(1) => 
                           N203, B(0) => N202);
   srl_42 : SHIFTER_GENERIC_N32_DW_rash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n3, SH(4) => 
                           n105_port, SH(3) => n104, SH(2) => B(2), SH(1) => 
                           B(1), SH(0) => B(0), SH_TC => n3, B(31) => N168, 
                           B(30) => N167, B(29) => N166, B(28) => N165, B(27) 
                           => N164, B(26) => N163, B(25) => N162, B(24) => N161
                           , B(23) => N160, B(22) => N159, B(21) => N158, B(20)
                           => N157, B(19) => N156, B(18) => N155, B(17) => N154
                           , B(16) => N153, B(15) => N152, B(14) => N151, B(13)
                           => N150, B(12) => N149, B(11) => N148, B(10) => N147
                           , B(9) => N146, B(8) => N145, B(7) => N144, B(6) => 
                           N143, B(5) => N142, B(4) => N141, B(3) => N140, B(2)
                           => N139, B(1) => N138, B(0) => N137);
   sra_40 : SHIFTER_GENERIC_N32_DW_sra_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n105_port, SH(3) => 
                           n104, SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), 
                           SH_TC => n4, B(31) => N136, B(30) => N135, B(29) => 
                           N134, B(28) => N133, B(27) => N132, B(26) => N131, 
                           B(25) => N130, B(24) => N129, B(23) => N128, B(22) 
                           => N127, B(21) => N126, B(20) => N125, B(19) => N124
                           , B(18) => N123, B(17) => N122, B(16) => N121, B(15)
                           => N120, B(14) => N119, B(13) => N118, B(12) => N117
                           , B(11) => N116, B(10) => N115, B(9) => N114, B(8) 
                           => N113, B(7) => N112, B(6) => N111, B(5) => N110, 
                           B(4) => N109, B(3) => N108, B(2) => N107, B(1) => 
                           N106, B(0) => N105);
   rol_33 : SHIFTER_GENERIC_N32_DW_lbsh_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n105_port, SH(3) => 
                           n104, SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), 
                           SH_TC => n5, B(31) => N70, B(30) => N69, B(29) => 
                           N68, B(28) => N67, B(27) => N66, B(26) => N65, B(25)
                           => N64, B(24) => N63, B(23) => N62, B(22) => N61, 
                           B(21) => N60, B(20) => N59, B(19) => N58, B(18) => 
                           N57, B(17) => N56, B(16) => N55, B(15) => N54, B(14)
                           => N53, B(13) => N52, B(12) => N51, B(11) => N50, 
                           B(10) => N49, B(9) => N48, B(8) => N47, B(7) => N46,
                           B(6) => N45, B(5) => N44, B(4) => N43, B(3) => N42, 
                           B(2) => N41, B(1) => N40, B(0) => N39);
   ror_31 : SHIFTER_GENERIC_N32_DW_rbsh_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n105_port, SH(3) => 
                           n104, SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), 
                           SH_TC => n6, B(31) => N38, B(30) => N37, B(29) => 
                           N36, B(28) => N35, B(27) => N34, B(26) => N33, B(25)
                           => N32, B(24) => N31, B(23) => N30, B(22) => N29, 
                           B(21) => N28, B(20) => N27, B(19) => N26, B(18) => 
                           N25, B(17) => N24, B(16) => N23, B(15) => N22, B(14)
                           => N21, B(13) => N20, B(12) => N19, B(11) => N18, 
                           B(10) => N17, B(9) => N16, B(8) => N15, B(7) => N14,
                           B(6) => N13, B(5) => N12, B(4) => N11, B(3) => N10, 
                           B(2) => N9, B(1) => N8, B(0) => N7);
   U1 : BUF_X1 port map( A => B(3), Z => n104);
   U2 : AOI222_X1 port map( A1 => N232, A2 => n103, B1 => N135, B2 => n99, C1 
                           => N167, C2 => n96, ZN => n39_port);
   U3 : AOI222_X1 port map( A1 => N231, A2 => n102, B1 => N134, B2 => n99, C1 
                           => N166, C2 => n96, ZN => n43_port);
   U4 : AOI222_X1 port map( A1 => N230, A2 => n102, B1 => N133, B2 => n99, C1 
                           => N165, C2 => n96, ZN => n45_port);
   U11 : AOI222_X1 port map( A1 => N229, A2 => n102, B1 => N132, B2 => n99, C1 
                           => N164, C2 => n96, ZN => n47_port);
   U12 : AOI222_X1 port map( A1 => N228, A2 => n102, B1 => N131, B2 => n99, C1 
                           => N163, C2 => n96, ZN => n49_port);
   U13 : AOI222_X1 port map( A1 => N227, A2 => n102, B1 => N130, B2 => n99, C1 
                           => N162, C2 => n96, ZN => n51_port);
   U14 : AOI222_X1 port map( A1 => N226, A2 => n102, B1 => N129, B2 => n99, C1 
                           => N161, C2 => n96, ZN => n53_port);
   U15 : AOI222_X1 port map( A1 => N225, A2 => n102, B1 => N128, B2 => n99, C1 
                           => N160, C2 => n96, ZN => n55_port);
   U16 : AOI222_X1 port map( A1 => N224, A2 => n102, B1 => N127, B2 => n99, C1 
                           => N159, C2 => n96, ZN => n57_port);
   U17 : AOI222_X1 port map( A1 => N223, A2 => n102, B1 => N126, B2 => n99, C1 
                           => N158, C2 => n96, ZN => n59_port);
   U18 : AOI222_X1 port map( A1 => N222, A2 => n102, B1 => N125, B2 => n99, C1 
                           => N157, C2 => n96, ZN => n61_port);
   U19 : AOI222_X1 port map( A1 => N221, A2 => n101, B1 => N124, B2 => n98, C1 
                           => N156, C2 => n95, ZN => n65_port);
   U20 : AOI222_X1 port map( A1 => N220, A2 => n101, B1 => N123, B2 => n98, C1 
                           => N155, C2 => n95, ZN => n67_port);
   U21 : AOI222_X1 port map( A1 => N219, A2 => n101, B1 => N122, B2 => n98, C1 
                           => N154, C2 => n95, ZN => n69_port);
   U22 : AOI222_X1 port map( A1 => N218, A2 => n101, B1 => N121, B2 => n98, C1 
                           => N153, C2 => n95, ZN => n71);
   U23 : AOI222_X1 port map( A1 => N217, A2 => n101, B1 => N120, B2 => n98, C1 
                           => N152, C2 => n95, ZN => n73);
   U24 : AOI222_X1 port map( A1 => N216, A2 => n101, B1 => N119, B2 => n98, C1 
                           => N151, C2 => n95, ZN => n75);
   U25 : AOI222_X1 port map( A1 => N215, A2 => n101, B1 => N118, B2 => n98, C1 
                           => N150, C2 => n95, ZN => n77);
   U26 : AOI222_X1 port map( A1 => N214, A2 => n101, B1 => N117, B2 => n98, C1 
                           => N149, C2 => n95, ZN => n79);
   U27 : AOI222_X1 port map( A1 => N213, A2 => n101, B1 => N116, B2 => n98, C1 
                           => N148, C2 => n95, ZN => n81);
   U28 : AOI222_X1 port map( A1 => N212, A2 => n101, B1 => N115, B2 => n98, C1 
                           => N147, C2 => n95, ZN => n83);
   U29 : AOI222_X1 port map( A1 => N204, A2 => n103, B1 => N107, B2 => n99, C1 
                           => N139, C2 => n96, ZN => n41_port);
   U30 : AOI222_X1 port map( A1 => N203, A2 => n102, B1 => N106, B2 => n98, C1 
                           => N138, C2 => n95, ZN => n63_port);
   U31 : AOI222_X1 port map( A1 => N211, A2 => n103, B1 => N114, B2 => n100, C1
                           => N146, C2 => n97, ZN => n11_port);
   U32 : AOI222_X1 port map( A1 => N210, A2 => n103, B1 => N113, B2 => n100, C1
                           => N145, C2 => n97, ZN => n25_port);
   U33 : AOI222_X1 port map( A1 => N209, A2 => n103, B1 => N112, B2 => n100, C1
                           => N144, C2 => n97, ZN => n27_port);
   U34 : AOI222_X1 port map( A1 => N208, A2 => n103, B1 => N111, B2 => n100, C1
                           => N143, C2 => n97, ZN => n29_port);
   U35 : AOI222_X1 port map( A1 => N207, A2 => n103, B1 => N110, B2 => n100, C1
                           => N142, C2 => n97, ZN => n31_port);
   U36 : AOI222_X1 port map( A1 => N206, A2 => n103, B1 => N109, B2 => n100, C1
                           => N141, C2 => n97, ZN => n33_port);
   U37 : AOI222_X1 port map( A1 => N205, A2 => n103, B1 => N108, B2 => n100, C1
                           => N140, C2 => n97, ZN => n35_port);
   U38 : AOI222_X1 port map( A1 => N69, A2 => n94, B1 => N264, B2 => n90, C1 =>
                           N37, C2 => n87, ZN => n38_port);
   U39 : AOI222_X1 port map( A1 => N68, A2 => n93, B1 => N263, B2 => n90, C1 =>
                           N36, C2 => n87, ZN => n42_port);
   U40 : AOI222_X1 port map( A1 => N67, A2 => n93, B1 => N262, B2 => n90, C1 =>
                           N35, C2 => n87, ZN => n44_port);
   U41 : AOI222_X1 port map( A1 => N66, A2 => n93, B1 => N261, B2 => n90, C1 =>
                           N34, C2 => n87, ZN => n46_port);
   U42 : AOI222_X1 port map( A1 => N65, A2 => n93, B1 => N260, B2 => n90, C1 =>
                           N33, C2 => n87, ZN => n48_port);
   U43 : AOI222_X1 port map( A1 => N64, A2 => n93, B1 => N259, B2 => n90, C1 =>
                           N32, C2 => n87, ZN => n50_port);
   U44 : AOI222_X1 port map( A1 => N63, A2 => n93, B1 => N258, B2 => n90, C1 =>
                           N31, C2 => n87, ZN => n52_port);
   U45 : AOI222_X1 port map( A1 => N62, A2 => n93, B1 => N257, B2 => n90, C1 =>
                           N30, C2 => n87, ZN => n54_port);
   U46 : AOI222_X1 port map( A1 => N61, A2 => n93, B1 => N256, B2 => n90, C1 =>
                           N29, C2 => n87, ZN => n56_port);
   U47 : AOI222_X1 port map( A1 => N60, A2 => n93, B1 => N255, B2 => n90, C1 =>
                           N28, C2 => n87, ZN => n58_port);
   U48 : AOI222_X1 port map( A1 => N59, A2 => n93, B1 => N254, B2 => n90, C1 =>
                           N27, C2 => n87, ZN => n60_port);
   U49 : AOI222_X1 port map( A1 => N58, A2 => n92, B1 => N253, B2 => n89, C1 =>
                           N26, C2 => n86, ZN => n64_port);
   U50 : AOI222_X1 port map( A1 => N57, A2 => n92, B1 => N252, B2 => n89, C1 =>
                           N25, C2 => n86, ZN => n66_port);
   U51 : AOI222_X1 port map( A1 => N56, A2 => n92, B1 => N251, B2 => n89, C1 =>
                           N24, C2 => n86, ZN => n68_port);
   U52 : AOI222_X1 port map( A1 => N55, A2 => n92, B1 => N250, B2 => n89, C1 =>
                           N23, C2 => n86, ZN => n70_port);
   U53 : AOI222_X1 port map( A1 => N54, A2 => n92, B1 => N249, B2 => n89, C1 =>
                           N22, C2 => n86, ZN => n72);
   U54 : AOI222_X1 port map( A1 => N53, A2 => n92, B1 => N248, B2 => n89, C1 =>
                           N21, C2 => n86, ZN => n74);
   U55 : AOI222_X1 port map( A1 => N52, A2 => n92, B1 => N247, B2 => n89, C1 =>
                           N20, C2 => n86, ZN => n76);
   U56 : AOI222_X1 port map( A1 => N51, A2 => n92, B1 => N246, B2 => n89, C1 =>
                           N19, C2 => n86, ZN => n78);
   U57 : AOI222_X1 port map( A1 => N50, A2 => n92, B1 => N245, B2 => n89, C1 =>
                           N18, C2 => n86, ZN => n80);
   U58 : AOI222_X1 port map( A1 => N49, A2 => n92, B1 => N244, B2 => n89, C1 =>
                           N17, C2 => n86, ZN => n82);
   U59 : AOI222_X1 port map( A1 => N41, A2 => n94, B1 => N236, B2 => n90, C1 =>
                           N9, C2 => n87, ZN => n40_port);
   U60 : AOI222_X1 port map( A1 => N40, A2 => n93, B1 => N235, B2 => n89, C1 =>
                           N8, C2 => n86, ZN => n62_port);
   U61 : AOI222_X1 port map( A1 => N39, A2 => n92, B1 => N234, B2 => n89, C1 =>
                           N7, C2 => n86, ZN => n84);
   U62 : AOI222_X1 port map( A1 => N70, A2 => n94, B1 => N265, B2 => n91, C1 =>
                           N38, C2 => n88, ZN => n36_port);
   U63 : AOI222_X1 port map( A1 => N48, A2 => n94, B1 => N243, B2 => n91, C1 =>
                           N16, C2 => n88, ZN => n10_port);
   U64 : AOI222_X1 port map( A1 => N47, A2 => n94, B1 => N242, B2 => n91, C1 =>
                           N15, C2 => n88, ZN => n24_port);
   U65 : AOI222_X1 port map( A1 => N46, A2 => n94, B1 => N241, B2 => n91, C1 =>
                           N14, C2 => n88, ZN => n26_port);
   U66 : AOI222_X1 port map( A1 => N45, A2 => n94, B1 => N240, B2 => n91, C1 =>
                           N13, C2 => n88, ZN => n28_port);
   U67 : AOI222_X1 port map( A1 => N44, A2 => n94, B1 => N239, B2 => n91, C1 =>
                           N12, C2 => n88, ZN => n30_port);
   U68 : AOI222_X1 port map( A1 => N43, A2 => n94, B1 => N238, B2 => n91, C1 =>
                           N11, C2 => n88, ZN => n32_port);
   U69 : AOI222_X1 port map( A1 => N42, A2 => n94, B1 => N237, B2 => n91, C1 =>
                           N10, C2 => n88, ZN => n34_port);
   U70 : BUF_X1 port map( A => n22_port, Z => n90);
   U71 : BUF_X1 port map( A => n22_port, Z => n89);
   U72 : BUF_X1 port map( A => n22_port, Z => n91);
   U73 : BUF_X1 port map( A => B(4), Z => n105_port);
   U74 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => OUTPUT(31));
   U75 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => OUTPUT(30));
   U76 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => OUTPUT(29));
   U77 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => OUTPUT(28));
   U78 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => OUTPUT(27));
   U79 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => OUTPUT(26));
   U80 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => OUTPUT(25));
   U81 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => OUTPUT(24));
   U82 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => OUTPUT(23));
   U83 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => OUTPUT(22));
   U84 : NAND2_X1 port map( A1 => n58_port, A2 => n59_port, ZN => OUTPUT(21));
   U85 : NAND2_X1 port map( A1 => n60_port, A2 => n61_port, ZN => OUTPUT(20));
   U86 : NAND2_X1 port map( A1 => n64_port, A2 => n65_port, ZN => OUTPUT(19));
   U87 : NAND2_X1 port map( A1 => n66_port, A2 => n67_port, ZN => OUTPUT(18));
   U88 : NAND2_X1 port map( A1 => n68_port, A2 => n69_port, ZN => OUTPUT(17));
   U89 : NAND2_X1 port map( A1 => n70_port, A2 => n71, ZN => OUTPUT(16));
   U90 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => OUTPUT(15));
   U91 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => OUTPUT(14));
   U92 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => OUTPUT(13));
   U93 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => OUTPUT(12));
   U94 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => OUTPUT(11));
   U95 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => OUTPUT(10));
   U96 : NAND2_X1 port map( A1 => n10_port, A2 => n11_port, ZN => OUTPUT(9));
   U97 : NAND2_X1 port map( A1 => n24_port, A2 => n25_port, ZN => OUTPUT(8));
   U98 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => OUTPUT(7));
   U99 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => OUTPUT(6));
   U100 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => OUTPUT(5));
   U101 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => OUTPUT(4));
   U102 : AOI222_X1 port map( A1 => N202, A2 => n101, B1 => N105, B2 => n98, C1
                           => N137, C2 => n95, ZN => n85);
   U103 : AOI222_X1 port map( A1 => N233, A2 => n103, B1 => N136, B2 => n100, 
                           C1 => N168, C2 => n97, ZN => n37_port);
   U104 : BUF_X1 port map( A => n19_port, Z => n99);
   U105 : BUF_X1 port map( A => n19_port, Z => n98);
   U106 : BUF_X1 port map( A => n20_port, Z => n96);
   U107 : BUF_X1 port map( A => n20_port, Z => n95);
   U108 : BUF_X1 port map( A => n23_port, Z => n87);
   U109 : BUF_X1 port map( A => n23_port, Z => n86);
   U110 : BUF_X1 port map( A => n12_port, Z => n102);
   U111 : BUF_X1 port map( A => n12_port, Z => n101);
   U112 : BUF_X1 port map( A => n21_port, Z => n93);
   U113 : BUF_X1 port map( A => n21_port, Z => n92);
   U114 : NOR3_X1 port map( A1 => n106_port, A2 => n108_port, A3 => n107_port, 
                           ZN => n22_port);
   U115 : BUF_X1 port map( A => n12_port, Z => n103);
   U116 : BUF_X1 port map( A => n21_port, Z => n94);
   U117 : BUF_X1 port map( A => n19_port, Z => n100);
   U118 : BUF_X1 port map( A => n20_port, Z => n97);
   U119 : BUF_X1 port map( A => n23_port, Z => n88);
   U120 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => OUTPUT(3));
   U121 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => OUTPUT(2));
   U122 : NAND2_X1 port map( A1 => n62_port, A2 => n63_port, ZN => OUTPUT(1));
   U123 : NOR3_X1 port map( A1 => n108_port, A2 => LEFT_RIGHT, A3 => n106_port,
                           ZN => n20_port);
   U124 : NOR3_X1 port map( A1 => LEFT_RIGHT, A2 => LOGIC_ARITH, A3 => 
                           n108_port, ZN => n19_port);
   U125 : NOR3_X1 port map( A1 => n108_port, A2 => LOGIC_ARITH, A3 => n107_port
                           , ZN => n12_port);
   U126 : NOR2_X1 port map( A1 => LEFT_RIGHT, A2 => SHIFT_ROTATE, ZN => 
                           n23_port);
   U127 : NOR2_X1 port map( A1 => n107_port, A2 => SHIFT_ROTATE, ZN => n21_port
                           );
   U128 : INV_X1 port map( A => LEFT_RIGHT, ZN => n107_port);
   U129 : INV_X1 port map( A => LOGIC_ARITH, ZN => n106_port);
   U130 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => OUTPUT(0));
   U131 : INV_X1 port map( A => SHIFT_ROTATE, ZN => n108_port);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity comparator is

   port( DATA1 : in std_logic_vector (31 downto 0);  DATA2i : in std_logic;  
         tipo : in std_logic_vector (0 to 5);  OUTALU : out std_logic_vector 
         (31 downto 0));

end comparator;

architecture SYN_Architectural of comparator is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N57, N58, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
      n55, n56, n57_port, n58_port, n59, n60, n61, n62, n63 : std_logic;

begin
   
   OUTALU_reg_0_inst : DLH_X1 port map( G => N57, D => N58, Q => OUTALU(0));
   OUTALU(1) <= '0';
   OUTALU(2) <= '0';
   OUTALU(3) <= '0';
   OUTALU(4) <= '0';
   OUTALU(5) <= '0';
   OUTALU(6) <= '0';
   OUTALU(7) <= '0';
   OUTALU(8) <= '0';
   OUTALU(9) <= '0';
   OUTALU(10) <= '0';
   OUTALU(11) <= '0';
   OUTALU(12) <= '0';
   OUTALU(13) <= '0';
   OUTALU(14) <= '0';
   OUTALU(15) <= '0';
   OUTALU(16) <= '0';
   OUTALU(17) <= '0';
   OUTALU(18) <= '0';
   OUTALU(19) <= '0';
   OUTALU(20) <= '0';
   OUTALU(21) <= '0';
   OUTALU(22) <= '0';
   OUTALU(23) <= '0';
   OUTALU(24) <= '0';
   OUTALU(25) <= '0';
   OUTALU(26) <= '0';
   OUTALU(27) <= '0';
   OUTALU(28) <= '0';
   OUTALU(29) <= '0';
   OUTALU(30) <= '0';
   OUTALU(31) <= '0';
   U85 : NAND3_X1 port map( A1 => tipo(0), A2 => n44, A3 => n45, ZN => n43);
   U33 : OR4_X1 port map( A1 => tipo(1), A2 => n61, A3 => n62, A4 => n57_port, 
                           ZN => n52);
   U34 : INV_X1 port map( A => n19, ZN => n53);
   U35 : NOR4_X1 port map( A1 => DATA1(23), A2 => DATA1(22), A3 => DATA1(21), 
                           A4 => DATA1(20), ZN => n27);
   U36 : NOR4_X1 port map( A1 => DATA1(9), A2 => DATA1(8), A3 => DATA1(7), A4 
                           => DATA1(6), ZN => n31);
   U37 : NOR4_X1 port map( A1 => DATA1(16), A2 => DATA1(15), A3 => DATA1(14), 
                           A4 => DATA1(13), ZN => n25);
   U38 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n19);
   U39 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n22);
   U40 : NAND4_X1 port map( A1 => n24, A2 => n25, A3 => n26, A4 => n27, ZN => 
                           n23);
   U41 : NOR4_X1 port map( A1 => DATA1(27), A2 => DATA1(26), A3 => DATA1(25), 
                           A4 => DATA1(24), ZN => n28);
   U42 : INV_X1 port map( A => DATA2i, ZN => n54);
   U43 : NOR4_X1 port map( A1 => DATA1(1), A2 => DATA1(19), A3 => DATA1(18), A4
                           => DATA1(17), ZN => n26);
   U44 : NOR4_X1 port map( A1 => DATA1(5), A2 => DATA1(4), A3 => DATA1(3), A4 
                           => DATA1(31), ZN => n30);
   U45 : NOR4_X1 port map( A1 => DATA1(30), A2 => DATA1(2), A3 => DATA1(29), A4
                           => DATA1(28), ZN => n29);
   U46 : NOR4_X1 port map( A1 => DATA1(12), A2 => DATA1(11), A3 => DATA1(10), 
                           A4 => DATA1(0), ZN => n24);
   U47 : OAI221_X1 port map( B1 => n13, B2 => n54, C1 => n58_port, C2 => n53, A
                           => n14, ZN => N58);
   U48 : INV_X1 port map( A => n20, ZN => n58_port);
   U49 : AOI21_X1 port map( B1 => n56, B2 => n53, A => n21, ZN => n13);
   U50 : AOI22_X1 port map( A1 => n15, A2 => n55, B1 => n16, B2 => n54, ZN => 
                           n14);
   U51 : OAI21_X1 port map( B1 => n17, B2 => n63, A => n18, ZN => n16);
   U52 : INV_X1 port map( A => n34, ZN => n55);
   U53 : INV_X1 port map( A => n32, ZN => n56);
   U54 : OR3_X1 port map( A1 => n20, A2 => n21, A3 => n33, ZN => N57);
   U55 : OAI211_X1 port map( C1 => n63, C2 => n17, A => n34, B => n32, ZN => 
                           n33);
   U56 : NOR4_X1 port map( A1 => n57_port, A2 => tipo(3), A3 => tipo(2), A4 => 
                           tipo(1), ZN => n35);
   U57 : OAI221_X1 port map( B1 => tipo(0), B2 => tipo(4), C1 => tipo(1), C2 =>
                           n62, A => n51, ZN => n40);
   U58 : AOI22_X1 port map( A1 => tipo(1), A2 => n61, B1 => tipo(0), B2 => 
                           tipo(3), ZN => n51);
   U59 : OAI211_X1 port map( C1 => tipo(1), C2 => tipo(2), A => n49, B => n50, 
                           ZN => n18);
   U60 : AOI211_X1 port map( C1 => tipo(1), C2 => n63, A => tipo(0), B => n44, 
                           ZN => n50);
   U61 : AOI22_X1 port map( A1 => tipo(2), A2 => n62, B1 => tipo(4), B2 => 
                           tipo(3), ZN => n49);
   U62 : INV_X1 port map( A => tipo(4), ZN => n62);
   U63 : INV_X1 port map( A => tipo(3), ZN => n61);
   U64 : NOR2_X1 port map( A1 => n63, A2 => tipo(3), ZN => n44);
   U65 : INV_X1 port map( A => tipo(0), ZN => n57_port);
   U66 : INV_X1 port map( A => tipo(1), ZN => n59);
   U67 : INV_X1 port map( A => tipo(5), ZN => n63);
   U68 : AOI21_X1 port map( B1 => n62, B2 => n35, A => n39, ZN => n17);
   U69 : AOI21_X1 port map( B1 => n52, B2 => n40, A => n60, ZN => n39);
   U70 : INV_X1 port map( A => tipo(2), ZN => n60);
   U71 : OAI21_X1 port map( B1 => n40, B2 => n48, A => n18, ZN => n20);
   U72 : NAND2_X1 port map( A1 => tipo(2), A2 => n63, ZN => n48);
   U73 : NOR2_X1 port map( A1 => tipo(4), A2 => n19, ZN => n15);
   U74 : OAI21_X1 port map( B1 => n35, B2 => n36, A => n63, ZN => n32);
   U75 : AOI211_X1 port map( C1 => tipo(1), C2 => n37, A => n38, B => tipo(3), 
                           ZN => n36);
   U76 : OR2_X1 port map( A1 => tipo(2), A2 => tipo(4), ZN => n37);
   U77 : OAI21_X1 port map( B1 => tipo(1), B2 => tipo(4), A => tipo(0), ZN => 
                           n38);
   U78 : OAI21_X1 port map( B1 => n46, B2 => n47, A => n57_port, ZN => n34);
   U79 : AND3_X1 port map( A1 => tipo(2), A2 => n59, A3 => n44, ZN => n47);
   U80 : NOR4_X1 port map( A1 => tipo(2), A2 => tipo(5), A3 => n61, A4 => n59, 
                           ZN => n46);
   U81 : OAI21_X1 port map( B1 => n42, B2 => n62, A => n43, ZN => n21);
   U82 : AOI21_X1 port map( B1 => n35, B2 => tipo(5), A => n55, ZN => n42);
   U83 : NOR3_X1 port map( A1 => n59, A2 => tipo(2), A3 => tipo(4), ZN => n45);

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity logic_N32 is

   port( FUNC : in std_logic_vector (0 to 5);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUT_ALU : out std_logic_vector (31 
         downto 0));

end logic_N32;

architecture SYN_Architectural of logic_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258 : std_logic;

begin
   
   U172 : NAND3_X1 port map( A1 => n258, A2 => n257, A3 => FUNC(2), ZN => n139)
                           ;
   U2 : BUF_X1 port map( A => n177, Z => n180);
   U3 : BUF_X1 port map( A => n177, Z => n179);
   U4 : BUF_X1 port map( A => n178, Z => n182);
   U5 : BUF_X1 port map( A => n178, Z => n183);
   U6 : BUF_X1 port map( A => n177, Z => n181);
   U7 : AOI21_X1 port map( B1 => n191, B2 => n245, A => n183, ZN => n122);
   U8 : AOI21_X1 port map( B1 => n191, B2 => n246, A => n183, ZN => n124);
   U9 : AOI21_X1 port map( B1 => n191, B2 => n247, A => n183, ZN => n126);
   U10 : AOI21_X1 port map( B1 => n191, B2 => n248, A => n183, ZN => n128);
   U11 : AOI21_X1 port map( B1 => n191, B2 => n249, A => n184, ZN => n130);
   U12 : AOI21_X1 port map( B1 => n191, B2 => n250, A => n184, ZN => n132);
   U13 : AOI21_X1 port map( B1 => n190, B2 => n193, A => n183, ZN => n112);
   U14 : AOI21_X1 port map( B1 => n189, B2 => n194, A => n182, ZN => n90);
   U15 : AOI21_X1 port map( B1 => n189, B2 => n229, A => n182, ZN => n86);
   U16 : AOI21_X1 port map( B1 => n189, B2 => n230, A => n182, ZN => n88);
   U17 : AOI21_X1 port map( B1 => n189, B2 => n231, A => n182, ZN => n92);
   U18 : AOI21_X1 port map( B1 => n189, B2 => n232, A => n182, ZN => n94);
   U19 : AOI21_X1 port map( B1 => n189, B2 => n233, A => n182, ZN => n96);
   U20 : AOI21_X1 port map( B1 => n190, B2 => n234, A => n182, ZN => n98);
   U21 : AOI21_X1 port map( B1 => n190, B2 => n235, A => n182, ZN => n100);
   U22 : AOI21_X1 port map( B1 => n190, B2 => n236, A => n182, ZN => n102);
   U23 : AOI21_X1 port map( B1 => n190, B2 => n237, A => n183, ZN => n104);
   U24 : AOI21_X1 port map( B1 => n190, B2 => n238, A => n183, ZN => n106);
   U25 : AOI21_X1 port map( B1 => n190, B2 => n239, A => n183, ZN => n108);
   U26 : AOI21_X1 port map( B1 => n190, B2 => n240, A => n183, ZN => n110);
   U27 : AOI21_X1 port map( B1 => n190, B2 => n241, A => n183, ZN => n114);
   U28 : AOI21_X1 port map( B1 => n190, B2 => n242, A => n183, ZN => n116);
   U29 : AOI21_X1 port map( B1 => n190, B2 => n243, A => n183, ZN => n118);
   U30 : AOI21_X1 port map( B1 => n190, B2 => n244, A => n183, ZN => n120);
   U31 : AOI21_X1 port map( B1 => n189, B2 => n251, A => n182, ZN => n69);
   U32 : AOI21_X1 port map( B1 => n188, B2 => n252, A => n181, ZN => n74);
   U33 : AOI21_X1 port map( B1 => n189, B2 => n253, A => n182, ZN => n76);
   U34 : AOI21_X1 port map( B1 => n189, B2 => n254, A => n181, ZN => n78);
   U35 : AOI21_X1 port map( B1 => n189, B2 => n255, A => n181, ZN => n80);
   U36 : AOI21_X1 port map( B1 => n189, B2 => n196, A => n182, ZN => n82);
   U37 : AOI21_X1 port map( B1 => n189, B2 => n195, A => n182, ZN => n84);
   U38 : OAI22_X1 port map( A1 => n85, A2 => n229, B1 => n86, B2 => n197, ZN =>
                           OUT_ALU(31));
   U39 : OAI22_X1 port map( A1 => n87, A2 => n230, B1 => n88, B2 => n198, ZN =>
                           OUT_ALU(30));
   U40 : OAI22_X1 port map( A1 => n91, A2 => n231, B1 => n92, B2 => n199, ZN =>
                           OUT_ALU(29));
   U41 : OAI22_X1 port map( A1 => n93, A2 => n232, B1 => n94, B2 => n200, ZN =>
                           OUT_ALU(28));
   U42 : OAI22_X1 port map( A1 => n95, A2 => n233, B1 => n96, B2 => n201, ZN =>
                           OUT_ALU(27));
   U43 : OAI22_X1 port map( A1 => n97, A2 => n234, B1 => n98, B2 => n202, ZN =>
                           OUT_ALU(26));
   U44 : OAI22_X1 port map( A1 => n99, A2 => n235, B1 => n100, B2 => n203, ZN 
                           => OUT_ALU(25));
   U45 : OAI22_X1 port map( A1 => n101, A2 => n236, B1 => n102, B2 => n204, ZN 
                           => OUT_ALU(24));
   U46 : OAI22_X1 port map( A1 => n103, A2 => n237, B1 => n104, B2 => n205, ZN 
                           => OUT_ALU(23));
   U47 : OAI22_X1 port map( A1 => n105, A2 => n238, B1 => n106, B2 => n206, ZN 
                           => OUT_ALU(22));
   U48 : OAI22_X1 port map( A1 => n107, A2 => n239, B1 => n108, B2 => n207, ZN 
                           => OUT_ALU(21));
   U49 : OAI22_X1 port map( A1 => n109, A2 => n240, B1 => n110, B2 => n208, ZN 
                           => OUT_ALU(20));
   U50 : OAI22_X1 port map( A1 => n113, A2 => n241, B1 => n114, B2 => n209, ZN 
                           => OUT_ALU(19));
   U51 : OAI22_X1 port map( A1 => n115, A2 => n242, B1 => n116, B2 => n210, ZN 
                           => OUT_ALU(18));
   U52 : OAI22_X1 port map( A1 => n117, A2 => n243, B1 => n118, B2 => n211, ZN 
                           => OUT_ALU(17));
   U53 : OAI22_X1 port map( A1 => n119, A2 => n244, B1 => n120, B2 => n212, ZN 
                           => OUT_ALU(16));
   U54 : OAI22_X1 port map( A1 => n121, A2 => n245, B1 => n122, B2 => n213, ZN 
                           => OUT_ALU(15));
   U55 : OAI22_X1 port map( A1 => n123, A2 => n246, B1 => n124, B2 => n214, ZN 
                           => OUT_ALU(14));
   U56 : OAI22_X1 port map( A1 => n125, A2 => n247, B1 => n126, B2 => n215, ZN 
                           => OUT_ALU(13));
   U57 : OAI22_X1 port map( A1 => n127, A2 => n248, B1 => n128, B2 => n216, ZN 
                           => OUT_ALU(12));
   U58 : OAI22_X1 port map( A1 => n129, A2 => n249, B1 => n130, B2 => n217, ZN 
                           => OUT_ALU(11));
   U59 : OAI22_X1 port map( A1 => n131, A2 => n250, B1 => n132, B2 => n218, ZN 
                           => OUT_ALU(10));
   U60 : OAI22_X1 port map( A1 => n68, A2 => n251, B1 => n69, B2 => n219, ZN =>
                           OUT_ALU(9));
   U61 : OAI22_X1 port map( A1 => n73, A2 => n252, B1 => n74, B2 => n220, ZN =>
                           OUT_ALU(8));
   U62 : OAI22_X1 port map( A1 => n75, A2 => n253, B1 => n76, B2 => n221, ZN =>
                           OUT_ALU(7));
   U63 : OAI22_X1 port map( A1 => n77, A2 => n254, B1 => n78, B2 => n222, ZN =>
                           OUT_ALU(6));
   U64 : OAI22_X1 port map( A1 => n79, A2 => n255, B1 => n80, B2 => n223, ZN =>
                           OUT_ALU(5));
   U65 : OAI22_X1 port map( A1 => n81, A2 => n196, B1 => n82, B2 => n224, ZN =>
                           OUT_ALU(4));
   U66 : BUF_X1 port map( A => n178, Z => n184);
   U67 : AOI221_X1 port map( B1 => n186, B2 => n219, C1 => n176, C2 => DATA1(9)
                           , A => n179, ZN => n68);
   U68 : AOI221_X1 port map( B1 => n188, B2 => n200, C1 => DATA1(28), C2 => 
                           n175, A => n181, ZN => n93);
   U69 : AOI221_X1 port map( B1 => n188, B2 => n202, C1 => DATA1(26), C2 => 
                           n175, A => n180, ZN => n97);
   U70 : AOI221_X1 port map( B1 => n188, B2 => n203, C1 => DATA1(25), C2 => 
                           n175, A => n181, ZN => n99);
   U71 : AOI221_X1 port map( B1 => n188, B2 => n204, C1 => DATA1(24), C2 => 
                           n175, A => n181, ZN => n101);
   U72 : AOI221_X1 port map( B1 => n187, B2 => n205, C1 => DATA1(23), C2 => 
                           n175, A => n180, ZN => n103);
   U73 : AOI221_X1 port map( B1 => n188, B2 => n206, C1 => DATA1(22), C2 => 
                           n175, A => n180, ZN => n105);
   U74 : AOI221_X1 port map( B1 => n187, B2 => n211, C1 => DATA1(17), C2 => 
                           n174, A => n180, ZN => n117);
   U75 : AOI221_X1 port map( B1 => n187, B2 => n212, C1 => DATA1(16), C2 => 
                           n174, A => n179, ZN => n119);
   U76 : AOI221_X1 port map( B1 => n186, B2 => n213, C1 => DATA1(15), C2 => 
                           n174, A => n179, ZN => n121);
   U77 : AOI221_X1 port map( B1 => n186, B2 => n214, C1 => DATA1(14), C2 => 
                           n174, A => n179, ZN => n123);
   U78 : AOI221_X1 port map( B1 => n186, B2 => n215, C1 => DATA1(13), C2 => 
                           n174, A => n179, ZN => n125);
   U79 : AOI221_X1 port map( B1 => n186, B2 => n216, C1 => DATA1(12), C2 => 
                           n174, A => n179, ZN => n127);
   U80 : AOI221_X1 port map( B1 => n188, B2 => n197, C1 => DATA1(31), C2 => 
                           n176, A => n181, ZN => n85);
   U81 : AOI221_X1 port map( B1 => n188, B2 => n199, C1 => DATA1(29), C2 => 
                           n175, A => n181, ZN => n91);
   U82 : AOI221_X1 port map( B1 => n188, B2 => n201, C1 => DATA1(27), C2 => 
                           n175, A => n181, ZN => n95);
   U83 : AOI221_X1 port map( B1 => n187, B2 => n207, C1 => DATA1(21), C2 => 
                           n175, A => n180, ZN => n107);
   U84 : AOI221_X1 port map( B1 => n187, B2 => n208, C1 => DATA1(20), C2 => 
                           n175, A => n180, ZN => n109);
   U85 : AOI221_X1 port map( B1 => n187, B2 => n209, C1 => DATA1(19), C2 => 
                           n174, A => n180, ZN => n113);
   U86 : AOI221_X1 port map( B1 => n186, B2 => n217, C1 => DATA1(11), C2 => 
                           n174, A => n179, ZN => n129);
   U87 : AOI221_X1 port map( B1 => n186, B2 => n218, C1 => DATA1(10), C2 => 
                           n174, A => n179, ZN => n131);
   U88 : AOI221_X1 port map( B1 => n186, B2 => n220, C1 => DATA1(8), C2 => n176
                           , A => n179, ZN => n73);
   U89 : AOI221_X1 port map( B1 => n186, B2 => n221, C1 => DATA1(7), C2 => n176
                           , A => n179, ZN => n75);
   U90 : AOI221_X1 port map( B1 => n186, B2 => n222, C1 => DATA1(6), C2 => n176
                           , A => n179, ZN => n77);
   U91 : AOI221_X1 port map( B1 => n187, B2 => n223, C1 => DATA1(5), C2 => n176
                           , A => n180, ZN => n79);
   U92 : AOI221_X1 port map( B1 => n187, B2 => n224, C1 => DATA1(4), C2 => n176
                           , A => n180, ZN => n81);
   U93 : AOI221_X1 port map( B1 => n187, B2 => n225, C1 => DATA1(3), C2 => n176
                           , A => n180, ZN => n83);
   U94 : AOI221_X1 port map( B1 => n188, B2 => n226, C1 => DATA1(2), C2 => n175
                           , A => n181, ZN => n89);
   U95 : AOI221_X1 port map( B1 => n188, B2 => n198, C1 => DATA1(30), C2 => 
                           n175, A => n181, ZN => n87);
   U96 : AOI221_X1 port map( B1 => n187, B2 => n210, C1 => DATA1(18), C2 => 
                           n174, A => n180, ZN => n115);
   U97 : AOI221_X1 port map( B1 => n187, B2 => n227, C1 => DATA1(1), C2 => n174
                           , A => n180, ZN => n111);
   U98 : BUF_X1 port map( A => n72, Z => n175);
   U99 : BUF_X1 port map( A => n72, Z => n174);
   U100 : OAI22_X1 port map( A1 => n133, A2 => n192, B1 => n134, B2 => n228, ZN
                           => OUT_ALU(0));
   U101 : AOI21_X1 port map( B1 => n188, B2 => n192, A => n181, ZN => n134);
   U102 : AOI221_X1 port map( B1 => n186, B2 => n228, C1 => DATA1(0), C2 => 
                           n174, A => n179, ZN => n133);
   U103 : BUF_X1 port map( A => n185, Z => n188);
   U104 : BUF_X1 port map( A => n185, Z => n189);
   U105 : BUF_X1 port map( A => n185, Z => n190);
   U106 : BUF_X1 port map( A => n72, Z => n176);
   U107 : BUF_X1 port map( A => n185, Z => n187);
   U108 : BUF_X1 port map( A => n185, Z => n186);
   U109 : INV_X1 port map( A => DATA1(12), ZN => n216);
   U110 : INV_X1 port map( A => DATA1(13), ZN => n215);
   U111 : INV_X1 port map( A => DATA1(14), ZN => n214);
   U112 : INV_X1 port map( A => DATA1(23), ZN => n205);
   U113 : INV_X1 port map( A => DATA1(22), ZN => n206);
   U114 : INV_X1 port map( A => DATA1(17), ZN => n211);
   U115 : INV_X1 port map( A => DATA1(16), ZN => n212);
   U116 : INV_X1 port map( A => DATA1(15), ZN => n213);
   U117 : INV_X1 port map( A => DATA1(21), ZN => n207);
   U118 : INV_X1 port map( A => DATA1(9), ZN => n219);
   U119 : INV_X1 port map( A => DATA1(11), ZN => n217);
   U120 : INV_X1 port map( A => DATA1(10), ZN => n218);
   U121 : INV_X1 port map( A => DATA1(8), ZN => n220);
   U122 : INV_X1 port map( A => DATA1(7), ZN => n221);
   U123 : INV_X1 port map( A => DATA1(2), ZN => n226);
   U124 : INV_X1 port map( A => DATA1(3), ZN => n225);
   U125 : INV_X1 port map( A => DATA1(28), ZN => n200);
   U126 : INV_X1 port map( A => DATA1(27), ZN => n201);
   U127 : INV_X1 port map( A => DATA1(26), ZN => n202);
   U128 : INV_X1 port map( A => DATA1(25), ZN => n203);
   U129 : INV_X1 port map( A => DATA1(24), ZN => n204);
   U130 : INV_X1 port map( A => DATA1(18), ZN => n210);
   U131 : INV_X1 port map( A => DATA1(0), ZN => n228);
   U132 : INV_X1 port map( A => DATA1(6), ZN => n222);
   U133 : INV_X1 port map( A => DATA1(29), ZN => n199);
   U134 : INV_X1 port map( A => DATA1(4), ZN => n224);
   U135 : INV_X1 port map( A => DATA1(1), ZN => n227);
   U136 : INV_X1 port map( A => DATA1(19), ZN => n209);
   U137 : INV_X1 port map( A => DATA1(20), ZN => n208);
   U138 : INV_X1 port map( A => DATA1(31), ZN => n197);
   U139 : INV_X1 port map( A => DATA1(5), ZN => n223);
   U140 : INV_X1 port map( A => DATA1(30), ZN => n198);
   U141 : BUF_X1 port map( A => n71, Z => n177);
   U142 : BUF_X1 port map( A => n71, Z => n178);
   U143 : INV_X1 port map( A => DATA2(31), ZN => n229);
   U144 : INV_X1 port map( A => DATA2(30), ZN => n230);
   U145 : INV_X1 port map( A => DATA2(29), ZN => n231);
   U146 : INV_X1 port map( A => DATA2(28), ZN => n232);
   U147 : INV_X1 port map( A => DATA2(27), ZN => n233);
   U148 : INV_X1 port map( A => DATA2(26), ZN => n234);
   U149 : INV_X1 port map( A => DATA2(25), ZN => n235);
   U150 : INV_X1 port map( A => DATA2(24), ZN => n236);
   U151 : INV_X1 port map( A => DATA2(23), ZN => n237);
   U152 : INV_X1 port map( A => DATA2(22), ZN => n238);
   U153 : INV_X1 port map( A => DATA2(21), ZN => n239);
   U154 : INV_X1 port map( A => DATA2(20), ZN => n240);
   U155 : INV_X1 port map( A => DATA2(19), ZN => n241);
   U156 : INV_X1 port map( A => DATA2(18), ZN => n242);
   U157 : INV_X1 port map( A => DATA2(17), ZN => n243);
   U158 : INV_X1 port map( A => DATA2(16), ZN => n244);
   U159 : INV_X1 port map( A => DATA2(15), ZN => n245);
   U160 : INV_X1 port map( A => DATA2(14), ZN => n246);
   U161 : INV_X1 port map( A => DATA2(13), ZN => n247);
   U162 : INV_X1 port map( A => DATA2(12), ZN => n248);
   U163 : INV_X1 port map( A => DATA2(11), ZN => n249);
   U164 : INV_X1 port map( A => DATA2(10), ZN => n250);
   U165 : INV_X1 port map( A => DATA2(9), ZN => n251);
   U166 : INV_X1 port map( A => DATA2(8), ZN => n252);
   U167 : INV_X1 port map( A => DATA2(7), ZN => n253);
   U168 : INV_X1 port map( A => DATA2(6), ZN => n254);
   U169 : INV_X1 port map( A => DATA2(5), ZN => n255);
   U170 : OAI22_X1 port map( A1 => n83, A2 => n195, B1 => n84, B2 => n225, ZN 
                           => OUT_ALU(3));
   U171 : OAI22_X1 port map( A1 => n89, A2 => n194, B1 => n90, B2 => n226, ZN 
                           => OUT_ALU(2));
   U173 : OAI22_X1 port map( A1 => n111, A2 => n193, B1 => n112, B2 => n227, ZN
                           => OUT_ALU(1));
   U174 : AOI211_X1 port map( C1 => n135, C2 => n136, A => FUNC(2), B => 
                           FUNC(0), ZN => n71);
   U175 : OR4_X1 port map( A1 => FUNC(3), A2 => FUNC(4), A3 => FUNC(5), A4 => 
                           n257, ZN => n135);
   U176 : NAND4_X1 port map( A1 => n257, A2 => FUNC(5), A3 => FUNC(4), A4 => 
                           FUNC(3), ZN => n136);
   U177 : INV_X1 port map( A => FUNC(1), ZN => n257);
   U178 : INV_X1 port map( A => FUNC(5), ZN => n258);
   U179 : AND3_X1 port map( A1 => FUNC(3), A2 => FUNC(4), A3 => n137, ZN => n72
                           );
   U180 : AOI211_X1 port map( C1 => FUNC(2), C2 => n258, A => FUNC(0), B => 
                           FUNC(1), ZN => n137);
   U181 : BUF_X1 port map( A => n70, Z => n185);
   U182 : NOR4_X1 port map( A1 => n256, A2 => FUNC(4), A3 => FUNC(3), A4 => 
                           FUNC(0), ZN => n70);
   U183 : INV_X1 port map( A => n138, ZN => n256);
   U184 : OAI21_X1 port map( B1 => FUNC(2), B2 => n257, A => n139, ZN => n138);
   U185 : CLKBUF_X1 port map( A => n185, Z => n191);
   U186 : INV_X1 port map( A => DATA2(0), ZN => n192);
   U187 : INV_X1 port map( A => DATA2(1), ZN => n193);
   U188 : INV_X1 port map( A => DATA2(2), ZN => n194);
   U189 : INV_X1 port map( A => DATA2(3), ZN => n195);
   U190 : INV_X1 port map( A => DATA2(4), ZN => n196);

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_192;

architecture SYN_STRUCTURAL of MUX21_192 is

   component ND2_574
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_575
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_576
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_192
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_192 port map( A => S, Y => SB);
   UND1 : ND2_576 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_575 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_574 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in26_N_out32 is

   port( IR_out : in std_logic_vector (25 downto 0);  signed_val : in std_logic
         ;  Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in26_N_out32;

architecture SYN_BHV of sign_eval_N_in26_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N0, n2 : std_logic;

begin
   Immediate <= ( N0, N0, N0, N0, N0, N0, IR_out(25), IR_out(24), IR_out(23), 
      IR_out(22), IR_out(21), IR_out(20), IR_out(19), IR_out(18), IR_out(17), 
      IR_out(16), IR_out(15), IR_out(14), IR_out(13), IR_out(12), IR_out(11), 
      IR_out(10), IR_out(9), IR_out(8), IR_out(7), IR_out(6), IR_out(5), 
      IR_out(4), IR_out(3), IR_out(2), IR_out(1), IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n2, ZN => N0);
   U2 : INV_X1 port map( A => IR_out(25), ZN => n2);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in16_N_out32 is

   port( IR_out : in std_logic_vector (15 downto 0);  signed_val : in std_logic
         ;  Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in16_N_out32;

architecture SYN_BHV of sign_eval_N_in16_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N0, n2 : std_logic;

begin
   Immediate <= ( N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, 
      N0, IR_out(15), IR_out(14), IR_out(13), IR_out(12), IR_out(11), 
      IR_out(10), IR_out(9), IR_out(8), IR_out(7), IR_out(6), IR_out(5), 
      IR_out(4), IR_out(3), IR_out(2), IR_out(1), IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n2, ZN => N0);
   U2 : INV_X1 port map( A => IR_out(15), ZN => n2);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in5_N_out32 is

   port( IR_out : in std_logic_vector (4 downto 0);  signed_val : in std_logic;
         Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in5_N_out32;

architecture SYN_BHV of sign_eval_N_in5_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N0, n2 : std_logic;

begin
   Immediate <= ( N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, 
      N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, IR_out(4), IR_out(3), 
      IR_out(2), IR_out(1), IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n2, ZN => N0);
   U2 : INV_X1 port map( A => IR_out(4), ZN => n2);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0;

architecture SYN_STRUCTURAL of MUX21_0 is

   component ND2_766
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_767
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0 port map( A => S, Y => SB);
   UND1 : ND2_0 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_767 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_766 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end DATAPTH_NBIT32_REG_BIT5_DW01_inc_0;

architecture SYN_rpl of DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U2 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_1;

architecture SYN_struct of MUX21_GENERIC_NBIT32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_61
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_62
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_63
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_64
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   gen1_0 : MUX21_64 port map( A => A(0), B => B(0), S => n3, Y => Y(0));
   gen1_1 : MUX21_63 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   gen1_2 : MUX21_62 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   gen1_3 : MUX21_61 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   gen1_4 : MUX21_60 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   gen1_5 : MUX21_59 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   gen1_6 : MUX21_58 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   gen1_7 : MUX21_57 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   gen1_8 : MUX21_56 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   gen1_9 : MUX21_55 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   gen1_10 : MUX21_54 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   gen1_11 : MUX21_53 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   gen1_12 : MUX21_52 port map( A => A(12), B => B(12), S => n1, Y => Y(12));
   gen1_13 : MUX21_51 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   gen1_14 : MUX21_50 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   gen1_15 : MUX21_49 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   gen1_16 : MUX21_48 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   gen1_17 : MUX21_47 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   gen1_18 : MUX21_46 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   gen1_19 : MUX21_45 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   gen1_20 : MUX21_44 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   gen1_21 : MUX21_43 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   gen1_22 : MUX21_42 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   gen1_23 : MUX21_41 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   gen1_24 : MUX21_40 port map( A => A(24), B => B(24), S => n2, Y => Y(24));
   gen1_25 : MUX21_39 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   gen1_26 : MUX21_38 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   gen1_27 : MUX21_37 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   gen1_28 : MUX21_36 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   gen1_29 : MUX21_35 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   gen1_30 : MUX21_34 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   gen1_31 : MUX21_33 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_1 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_1;

architecture SYN_SYNC_BHV of FF_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n6, n5, n3, n7, n8, n_1076 : std_logic;

begin
   Q <= n6;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => n6, QN => n_1076);
   U3 : NOR2_X1 port map( A1 => n3, A2 => n7, ZN => n5);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => n6, B2 => n8, ZN => n3);
   U5 : INV_X1 port map( A => EN, ZN => n8);
   U6 : INV_X1 port map( A => RESET, ZN => n7);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity load_data is

   port( data_in : in std_logic_vector (31 downto 0);  signed_val, load_op : in
         std_logic;  load_type : in std_logic_vector (1 downto 0);  data_out : 
         out std_logic_vector (31 downto 0));

end load_data;

architecture SYN_bhv_load of load_data is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
      N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64
      , N65, N66, N67, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n31, n32, n33, n34 : std_logic;

begin
   
   data_out_reg_31_inst : DLH_X1 port map( G => load_op, D => N67, Q => 
                           data_out(31));
   data_out_reg_30_inst : DLH_X1 port map( G => load_op, D => N66, Q => 
                           data_out(30));
   data_out_reg_29_inst : DLH_X1 port map( G => load_op, D => N65, Q => 
                           data_out(29));
   data_out_reg_28_inst : DLH_X1 port map( G => load_op, D => N64, Q => 
                           data_out(28));
   data_out_reg_27_inst : DLH_X1 port map( G => load_op, D => N63, Q => 
                           data_out(27));
   data_out_reg_26_inst : DLH_X1 port map( G => load_op, D => N62, Q => 
                           data_out(26));
   data_out_reg_25_inst : DLH_X1 port map( G => load_op, D => N61, Q => 
                           data_out(25));
   data_out_reg_24_inst : DLH_X1 port map( G => load_op, D => N60, Q => 
                           data_out(24));
   data_out_reg_23_inst : DLH_X1 port map( G => load_op, D => N59, Q => 
                           data_out(23));
   data_out_reg_22_inst : DLH_X1 port map( G => load_op, D => N58, Q => 
                           data_out(22));
   data_out_reg_21_inst : DLH_X1 port map( G => load_op, D => N57, Q => 
                           data_out(21));
   data_out_reg_20_inst : DLH_X1 port map( G => load_op, D => N56, Q => 
                           data_out(20));
   data_out_reg_19_inst : DLH_X1 port map( G => load_op, D => N55, Q => 
                           data_out(19));
   data_out_reg_18_inst : DLH_X1 port map( G => load_op, D => N54, Q => 
                           data_out(18));
   data_out_reg_17_inst : DLH_X1 port map( G => load_op, D => N53, Q => 
                           data_out(17));
   data_out_reg_16_inst : DLH_X1 port map( G => load_op, D => N52, Q => 
                           data_out(16));
   data_out_reg_15_inst : DLH_X1 port map( G => load_op, D => N51, Q => 
                           data_out(15));
   data_out_reg_14_inst : DLH_X1 port map( G => load_op, D => N50, Q => 
                           data_out(14));
   data_out_reg_13_inst : DLH_X1 port map( G => load_op, D => N49, Q => 
                           data_out(13));
   data_out_reg_12_inst : DLH_X1 port map( G => load_op, D => N48, Q => 
                           data_out(12));
   data_out_reg_11_inst : DLH_X1 port map( G => load_op, D => N47, Q => 
                           data_out(11));
   data_out_reg_10_inst : DLH_X1 port map( G => load_op, D => N46, Q => 
                           data_out(10));
   data_out_reg_9_inst : DLH_X1 port map( G => load_op, D => N45, Q => 
                           data_out(9));
   data_out_reg_8_inst : DLH_X1 port map( G => load_op, D => N44, Q => 
                           data_out(8));
   data_out_reg_7_inst : DLH_X1 port map( G => load_op, D => N43, Q => 
                           data_out(7));
   data_out_reg_6_inst : DLH_X1 port map( G => load_op, D => N42, Q => 
                           data_out(6));
   data_out_reg_5_inst : DLH_X1 port map( G => load_op, D => N41, Q => 
                           data_out(5));
   data_out_reg_4_inst : DLH_X1 port map( G => load_op, D => N40, Q => 
                           data_out(4));
   data_out_reg_3_inst : DLH_X1 port map( G => load_op, D => N39, Q => 
                           data_out(3));
   data_out_reg_2_inst : DLH_X1 port map( G => load_op, D => N38, Q => 
                           data_out(2));
   data_out_reg_1_inst : DLH_X1 port map( G => load_op, D => N37, Q => 
                           data_out(1));
   data_out_reg_0_inst : DLH_X1 port map( G => load_op, D => N36, Q => 
                           data_out(0));
   U2 : INV_X1 port map( A => n4, ZN => n32);
   U3 : BUF_X1 port map( A => n5, Z => n30);
   U4 : BUF_X1 port map( A => n5, Z => n31);
   U5 : OAI21_X1 port map( B1 => n4, B2 => n34, A => n30, ZN => N67);
   U6 : NAND2_X1 port map( A1 => load_type(1), A2 => n33, ZN => n29);
   U7 : INV_X1 port map( A => load_type(0), ZN => n33);
   U8 : NAND2_X1 port map( A1 => load_type(1), A2 => load_type(0), ZN => n4);
   U9 : OR4_X1 port map( A1 => load_type(0), A2 => n34, A3 => signed_val, A4 =>
                           load_type(1), ZN => n5);
   U10 : INV_X1 port map( A => data_in(31), ZN => n34);
   U11 : NAND2_X1 port map( A1 => n31, A2 => n28, ZN => N44);
   U12 : NAND2_X1 port map( A1 => data_in(8), A2 => load_type(0), ZN => n28);
   U13 : NAND2_X1 port map( A1 => n31, A2 => n27, ZN => N45);
   U14 : NAND2_X1 port map( A1 => data_in(9), A2 => load_type(0), ZN => n27);
   U15 : NAND2_X1 port map( A1 => n31, A2 => n26, ZN => N46);
   U16 : NAND2_X1 port map( A1 => data_in(10), A2 => load_type(0), ZN => n26);
   U17 : NAND2_X1 port map( A1 => n31, A2 => n25, ZN => N47);
   U18 : NAND2_X1 port map( A1 => data_in(11), A2 => load_type(0), ZN => n25);
   U19 : NAND2_X1 port map( A1 => n31, A2 => n24, ZN => N48);
   U20 : NAND2_X1 port map( A1 => data_in(12), A2 => load_type(0), ZN => n24);
   U21 : NAND2_X1 port map( A1 => n31, A2 => n23, ZN => N49);
   U22 : NAND2_X1 port map( A1 => data_in(13), A2 => load_type(0), ZN => n23);
   U23 : NAND2_X1 port map( A1 => n31, A2 => n22, ZN => N50);
   U24 : NAND2_X1 port map( A1 => data_in(14), A2 => load_type(0), ZN => n22);
   U25 : NAND2_X1 port map( A1 => n31, A2 => n21, ZN => N51);
   U26 : NAND2_X1 port map( A1 => data_in(15), A2 => load_type(0), ZN => n21);
   U27 : NAND2_X1 port map( A1 => n30, A2 => n16, ZN => N56);
   U28 : NAND2_X1 port map( A1 => data_in(20), A2 => n32, ZN => n16);
   U29 : NAND2_X1 port map( A1 => n30, A2 => n15, ZN => N57);
   U30 : NAND2_X1 port map( A1 => data_in(21), A2 => n32, ZN => n15);
   U31 : NAND2_X1 port map( A1 => n30, A2 => n14, ZN => N58);
   U32 : NAND2_X1 port map( A1 => data_in(22), A2 => n32, ZN => n14);
   U33 : NAND2_X1 port map( A1 => n30, A2 => n13, ZN => N59);
   U34 : NAND2_X1 port map( A1 => data_in(23), A2 => n32, ZN => n13);
   U35 : NAND2_X1 port map( A1 => n30, A2 => n12, ZN => N60);
   U36 : NAND2_X1 port map( A1 => data_in(24), A2 => n32, ZN => n12);
   U37 : NAND2_X1 port map( A1 => n30, A2 => n11, ZN => N61);
   U38 : NAND2_X1 port map( A1 => data_in(25), A2 => n32, ZN => n11);
   U39 : NAND2_X1 port map( A1 => n30, A2 => n10, ZN => N62);
   U40 : NAND2_X1 port map( A1 => data_in(26), A2 => n32, ZN => n10);
   U41 : NAND2_X1 port map( A1 => n30, A2 => n9, ZN => N63);
   U42 : NAND2_X1 port map( A1 => data_in(27), A2 => n32, ZN => n9);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n8, ZN => N64);
   U44 : NAND2_X1 port map( A1 => data_in(28), A2 => n32, ZN => n8);
   U45 : NAND2_X1 port map( A1 => n30, A2 => n7, ZN => N65);
   U46 : NAND2_X1 port map( A1 => data_in(29), A2 => n32, ZN => n7);
   U47 : NAND2_X1 port map( A1 => n30, A2 => n6, ZN => N66);
   U48 : NAND2_X1 port map( A1 => data_in(30), A2 => n32, ZN => n6);
   U49 : NAND2_X1 port map( A1 => n31, A2 => n20, ZN => N52);
   U50 : NAND2_X1 port map( A1 => data_in(16), A2 => n32, ZN => n20);
   U51 : NAND2_X1 port map( A1 => n31, A2 => n19, ZN => N53);
   U52 : NAND2_X1 port map( A1 => data_in(17), A2 => n32, ZN => n19);
   U53 : NAND2_X1 port map( A1 => n31, A2 => n18, ZN => N54);
   U54 : NAND2_X1 port map( A1 => data_in(18), A2 => n32, ZN => n18);
   U55 : NAND2_X1 port map( A1 => n31, A2 => n17, ZN => N55);
   U56 : NAND2_X1 port map( A1 => data_in(19), A2 => n32, ZN => n17);
   U57 : AND2_X1 port map( A1 => data_in(0), A2 => n29, ZN => N36);
   U58 : AND2_X1 port map( A1 => data_in(1), A2 => n29, ZN => N37);
   U59 : AND2_X1 port map( A1 => data_in(2), A2 => n29, ZN => N38);
   U60 : AND2_X1 port map( A1 => data_in(3), A2 => n29, ZN => N39);
   U61 : AND2_X1 port map( A1 => data_in(4), A2 => n29, ZN => N40);
   U62 : AND2_X1 port map( A1 => data_in(5), A2 => n29, ZN => N41);
   U63 : AND2_X1 port map( A1 => data_in(6), A2 => n29, ZN => N42);
   U64 : AND2_X1 port map( A1 => data_in(7), A2 => n29, ZN => N43);

end SYN_bhv_load;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_3;

architecture SYN_struct of MUX21_GENERIC_NBIT32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_97
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_98
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_99
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_100
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_101
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_102
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_103
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_104
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_105
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_106
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_107
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_108
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_109
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_110
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_111
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_112
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_113
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_114
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_115
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_116
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_117
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_118
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_119
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_120
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_121
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_122
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_123
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_124
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_125
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_126
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_127
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   gen1_0 : MUX21_128 port map( A => A(0), B => B(0), S => n4, Y => Y(0));
   gen1_1 : MUX21_127 port map( A => A(1), B => B(1), S => n4, Y => Y(1));
   gen1_2 : MUX21_126 port map( A => A(2), B => B(2), S => n4, Y => Y(2));
   gen1_3 : MUX21_125 port map( A => A(3), B => B(3), S => n4, Y => Y(3));
   gen1_4 : MUX21_124 port map( A => A(4), B => B(4), S => n4, Y => Y(4));
   gen1_5 : MUX21_123 port map( A => A(5), B => B(5), S => n4, Y => Y(5));
   gen1_6 : MUX21_122 port map( A => A(6), B => B(6), S => n4, Y => Y(6));
   gen1_7 : MUX21_121 port map( A => A(7), B => B(7), S => n4, Y => Y(7));
   gen1_8 : MUX21_120 port map( A => A(8), B => B(8), S => n4, Y => Y(8));
   gen1_9 : MUX21_119 port map( A => A(9), B => B(9), S => n4, Y => Y(9));
   gen1_10 : MUX21_118 port map( A => A(10), B => B(10), S => n4, Y => Y(10));
   gen1_11 : MUX21_117 port map( A => A(11), B => B(11), S => n4, Y => Y(11));
   gen1_12 : MUX21_116 port map( A => A(12), B => B(12), S => n5, Y => Y(12));
   gen1_13 : MUX21_115 port map( A => A(13), B => B(13), S => n5, Y => Y(13));
   gen1_14 : MUX21_114 port map( A => A(14), B => B(14), S => n5, Y => Y(14));
   gen1_15 : MUX21_113 port map( A => A(15), B => B(15), S => n5, Y => Y(15));
   gen1_16 : MUX21_112 port map( A => A(16), B => B(16), S => n5, Y => Y(16));
   gen1_17 : MUX21_111 port map( A => A(17), B => B(17), S => n5, Y => Y(17));
   gen1_18 : MUX21_110 port map( A => A(18), B => B(18), S => n5, Y => Y(18));
   gen1_19 : MUX21_109 port map( A => A(19), B => B(19), S => n5, Y => Y(19));
   gen1_20 : MUX21_108 port map( A => A(20), B => B(20), S => n5, Y => Y(20));
   gen1_21 : MUX21_107 port map( A => A(21), B => B(21), S => n5, Y => Y(21));
   gen1_22 : MUX21_106 port map( A => A(22), B => B(22), S => n5, Y => Y(22));
   gen1_23 : MUX21_105 port map( A => A(23), B => B(23), S => n5, Y => Y(23));
   gen1_24 : MUX21_104 port map( A => A(24), B => B(24), S => n6, Y => Y(24));
   gen1_25 : MUX21_103 port map( A => A(25), B => B(25), S => n6, Y => Y(25));
   gen1_26 : MUX21_102 port map( A => A(26), B => B(26), S => n6, Y => Y(26));
   gen1_27 : MUX21_101 port map( A => A(27), B => B(27), S => n6, Y => Y(27));
   gen1_28 : MUX21_100 port map( A => A(28), B => B(28), S => n6, Y => Y(28));
   gen1_29 : MUX21_99 port map( A => A(29), B => B(29), S => n6, Y => Y(29));
   gen1_30 : MUX21_98 port map( A => A(30), B => B(30), S => n6, Y => Y(30));
   gen1_31 : MUX21_97 port map( A => A(31), B => B(31), S => n6, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n4);
   U2 : BUF_X1 port map( A => SEL, Z => n5);
   U3 : BUF_X1 port map( A => SEL, Z => n6);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_4 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_4;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n65);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n66);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n67);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n68);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n69);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n98, Q => Q(26), 
                           QN => n70);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n98, Q => Q(25), 
                           QN => n71);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n98, Q => Q(24), 
                           QN => n72);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n73);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n98, Q => Q(22),
                           QN => n74);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n98, Q => Q(21),
                           QN => n75);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n99, Q => Q(20),
                           QN => n76);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n97, Q => Q(19),
                           QN => n77);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n99, Q => Q(18),
                           QN => n78);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n99, Q => Q(17),
                           QN => n79);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n99, Q => Q(16),
                           QN => n80);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n97, Q => Q(15),
                           QN => n81);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n99, Q => Q(14),
                           QN => n82);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n99, Q => Q(13),
                           QN => n83);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n99, Q => Q(12),
                           QN => n84);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n85);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n86);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n98, Q => Q(9), 
                           QN => n87);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n98, Q => Q(8), 
                           QN => n88);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n97, Q => Q(7), 
                           QN => n89);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n97, Q => Q(6), 
                           QN => n90);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n91);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n92);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n98, Q => Q(3), 
                           QN => n93);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n98, Q => Q(2), 
                           QN => n94);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n95);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n97, Q => Q(0), 
                           QN => n96);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n96, B2 => ENABLE, A => n39, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n39);
   U7 : OAI21_X1 port map( B1 => n95, B2 => ENABLE, A => n40, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n40);
   U9 : OAI21_X1 port map( B1 => n94, B2 => ENABLE, A => n41, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n41);
   U11 : OAI21_X1 port map( B1 => n93, B2 => ENABLE, A => n43, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n43);
   U13 : OAI21_X1 port map( B1 => n92, B2 => ENABLE, A => n44, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n44);
   U15 : OAI21_X1 port map( B1 => n91, B2 => ENABLE, A => n45, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n45);
   U17 : OAI21_X1 port map( B1 => n90, B2 => ENABLE, A => n46, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n46);
   U19 : OAI21_X1 port map( B1 => n89, B2 => ENABLE, A => n47, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n47);
   U21 : OAI21_X1 port map( B1 => n88, B2 => ENABLE, A => n48, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n48);
   U23 : OAI21_X1 port map( B1 => n87, B2 => ENABLE, A => n49, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n49);
   U25 : OAI21_X1 port map( B1 => n86, B2 => ENABLE, A => n50, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n50);
   U27 : OAI21_X1 port map( B1 => n85, B2 => ENABLE, A => n51, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n51);
   U29 : OAI21_X1 port map( B1 => n84, B2 => ENABLE, A => n52, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n52);
   U31 : OAI21_X1 port map( B1 => n83, B2 => ENABLE, A => n54, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n54);
   U33 : OAI21_X1 port map( B1 => n82, B2 => ENABLE, A => n55, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n55);
   U35 : OAI21_X1 port map( B1 => n81, B2 => ENABLE, A => n56, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n56);
   U37 : OAI21_X1 port map( B1 => n80, B2 => ENABLE, A => n57, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n57);
   U39 : OAI21_X1 port map( B1 => n79, B2 => ENABLE, A => n58, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n58);
   U41 : OAI21_X1 port map( B1 => n78, B2 => ENABLE, A => n59, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n59);
   U43 : OAI21_X1 port map( B1 => n77, B2 => ENABLE, A => n60, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n60);
   U45 : OAI21_X1 port map( B1 => n76, B2 => ENABLE, A => n61, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n61);
   U47 : OAI21_X1 port map( B1 => n75, B2 => ENABLE, A => n62, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n62);
   U49 : OAI21_X1 port map( B1 => n74, B2 => ENABLE, A => n63, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n63);
   U51 : OAI21_X1 port map( B1 => n72, B2 => ENABLE, A => n34, ZN => n8);
   U52 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n34);
   U53 : OAI21_X1 port map( B1 => n71, B2 => ENABLE, A => n35, ZN => n7);
   U54 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n35);
   U55 : OAI21_X1 port map( B1 => n70, B2 => ENABLE, A => n36, ZN => n6);
   U56 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n36);
   U57 : OAI21_X1 port map( B1 => n69, B2 => ENABLE, A => n37, ZN => n5);
   U58 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n37);
   U59 : OAI21_X1 port map( B1 => n68, B2 => ENABLE, A => n38, ZN => n4);
   U60 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n38);
   U61 : OAI21_X1 port map( B1 => n67, B2 => ENABLE, A => n42, ZN => n3);
   U62 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n42);
   U63 : OAI21_X1 port map( B1 => n66, B2 => ENABLE, A => n53, ZN => n2);
   U64 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n53);
   U65 : OAI21_X1 port map( B1 => n65, B2 => ENABLE, A => n64, ZN => n1);
   U66 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n64);
   U67 : OAI21_X1 port map( B1 => n73, B2 => ENABLE, A => n33, ZN => n9);
   U68 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n33);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity COND_BT_NBIT32 is

   port( ZERO_BIT, OPCODE_0, branch_op : in std_logic;  con_sign : out 
         std_logic);

end COND_BT_NBIT32;

architecture SYN_BHV of COND_BT_NBIT32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ZERO_BIT, B => OPCODE_0, Z => n1);
   U2 : AND2_X1 port map( A1 => branch_op, A2 => n1, ZN => con_sign);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity zero_eval_NBIT32 is

   port( input : in std_logic_vector (31 downto 0);  res : out std_logic);

end zero_eval_NBIT32;

architecture SYN_bhv of zero_eval_NBIT32 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : NOR4_X1 port map( A1 => input(23), A2 => input(22), A3 => input(21), A4
                           => input(20), ZN => n6);
   U2 : NOR4_X1 port map( A1 => input(9), A2 => input(8), A3 => input(7), A4 =>
                           input(6), ZN => n10);
   U3 : NOR4_X1 port map( A1 => input(5), A2 => input(4), A3 => input(3), A4 =>
                           input(31), ZN => n9);
   U4 : NOR4_X1 port map( A1 => input(30), A2 => input(2), A3 => input(29), A4 
                           => input(28), ZN => n8);
   U5 : NOR4_X1 port map( A1 => input(27), A2 => input(26), A3 => input(25), A4
                           => input(24), ZN => n7);
   U6 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => n2);
   U7 : NOR4_X1 port map( A1 => input(12), A2 => input(11), A3 => input(10), A4
                           => input(0), ZN => n3);
   U8 : NOR4_X1 port map( A1 => input(16), A2 => input(15), A3 => input(14), A4
                           => input(13), ZN => n4);
   U9 : NOR4_X1 port map( A1 => input(1), A2 => input(19), A3 => input(18), A4 
                           => input(17), ZN => n5);
   U10 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => res);
   U11 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => n9, A4 => n10, ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ALU_N32 is

   port( CLK : in std_logic;  FUNC : in std_logic_vector (0 to 5);  DATA1, 
         DATA2 : in std_logic_vector (31 downto 0);  OUT_ALU : out 
         std_logic_vector (31 downto 0));

end ALU_N32;

architecture SYN_Architectural of ALU_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component P4_ADDER_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component SHIFTER_GENERIC_N32
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
            downto 0);  LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE : in std_logic;  
            OUTPUT : out std_logic_vector (31 downto 0));
   end component;
   
   component comparator
      port( DATA1 : in std_logic_vector (31 downto 0);  DATA2i : in std_logic; 
            tipo : in std_logic_vector (0 to 5);  OUTALU : out std_logic_vector
            (31 downto 0));
   end component;
   
   component logic_N32
      port( FUNC : in std_logic_vector (0 to 5);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUT_ALU : out std_logic_vector (31
            downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal OUTPUT_alu_i_31_port, OUTPUT_alu_i_30_port, OUTPUT_alu_i_29_port, 
      OUTPUT_alu_i_28_port, OUTPUT_alu_i_27_port, OUTPUT_alu_i_26_port, 
      OUTPUT_alu_i_25_port, OUTPUT_alu_i_24_port, OUTPUT_alu_i_23_port, 
      OUTPUT_alu_i_22_port, OUTPUT_alu_i_21_port, OUTPUT_alu_i_20_port, 
      OUTPUT_alu_i_19_port, OUTPUT_alu_i_18_port, OUTPUT_alu_i_17_port, 
      OUTPUT_alu_i_16_port, OUTPUT_alu_i_15_port, OUTPUT_alu_i_14_port, 
      OUTPUT_alu_i_13_port, OUTPUT_alu_i_12_port, OUTPUT_alu_i_11_port, 
      OUTPUT_alu_i_10_port, OUTPUT_alu_i_9_port, OUTPUT_alu_i_8_port, 
      OUTPUT_alu_i_7_port, OUTPUT_alu_i_6_port, OUTPUT_alu_i_5_port, 
      OUTPUT_alu_i_4_port, OUTPUT_alu_i_3_port, OUTPUT_alu_i_2_port, 
      OUTPUT_alu_i_1_port, OUTPUT_alu_i_0_port, OUTPUT4_31_port, 
      OUTPUT4_30_port, OUTPUT4_29_port, OUTPUT4_28_port, OUTPUT4_27_port, 
      OUTPUT4_26_port, OUTPUT4_25_port, OUTPUT4_24_port, OUTPUT4_23_port, 
      OUTPUT4_22_port, OUTPUT4_21_port, OUTPUT4_20_port, OUTPUT4_19_port, 
      OUTPUT4_18_port, OUTPUT4_17_port, OUTPUT4_16_port, OUTPUT4_15_port, 
      OUTPUT4_14_port, OUTPUT4_13_port, OUTPUT4_12_port, OUTPUT4_11_port, 
      OUTPUT4_10_port, OUTPUT4_9_port, OUTPUT4_8_port, OUTPUT4_7_port, 
      OUTPUT4_6_port, OUTPUT4_5_port, OUTPUT4_4_port, OUTPUT4_3_port, 
      OUTPUT4_2_port, OUTPUT4_1_port, OUTPUT4_0_port, OUTPUT2_31_port, 
      OUTPUT2_30_port, OUTPUT2_29_port, OUTPUT2_28_port, OUTPUT2_27_port, 
      OUTPUT2_26_port, OUTPUT2_25_port, OUTPUT2_24_port, OUTPUT2_23_port, 
      OUTPUT2_22_port, OUTPUT2_21_port, OUTPUT2_20_port, OUTPUT2_19_port, 
      OUTPUT2_18_port, OUTPUT2_17_port, OUTPUT2_16_port, OUTPUT2_15_port, 
      OUTPUT2_14_port, OUTPUT2_13_port, OUTPUT2_12_port, OUTPUT2_11_port, 
      OUTPUT2_10_port, OUTPUT2_9_port, OUTPUT2_8_port, OUTPUT2_7_port, 
      OUTPUT2_6_port, OUTPUT2_5_port, OUTPUT2_4_port, OUTPUT2_3_port, 
      OUTPUT2_2_port, OUTPUT2_1_port, OUTPUT2_0_port, Cout_i, OUTPUT3_0_port, 
      LOGIC_ARITH_i, LEFT_RIGHT_i, SHIFT_ROTATE_i, OUTPUT1_31_port, 
      OUTPUT1_30_port, OUTPUT1_29_port, OUTPUT1_28_port, OUTPUT1_27_port, 
      OUTPUT1_26_port, OUTPUT1_25_port, OUTPUT1_24_port, OUTPUT1_23_port, 
      OUTPUT1_22_port, OUTPUT1_21_port, OUTPUT1_20_port, OUTPUT1_19_port, 
      OUTPUT1_18_port, OUTPUT1_17_port, OUTPUT1_16_port, OUTPUT1_15_port, 
      OUTPUT1_14_port, OUTPUT1_13_port, OUTPUT1_12_port, OUTPUT1_11_port, 
      OUTPUT1_10_port, OUTPUT1_9_port, OUTPUT1_8_port, OUTPUT1_7_port, 
      OUTPUT1_6_port, OUTPUT1_5_port, OUTPUT1_4_port, OUTPUT1_3_port, 
      OUTPUT1_2_port, OUTPUT1_1_port, OUTPUT1_0_port, data1i_31_port, 
      data1i_30_port, data1i_29_port, data1i_28_port, data1i_27_port, 
      data1i_26_port, data1i_25_port, data1i_24_port, data1i_23_port, 
      data1i_22_port, data1i_21_port, data1i_20_port, data1i_19_port, 
      data1i_18_port, data1i_17_port, data1i_16_port, data1i_15_port, 
      data1i_14_port, data1i_13_port, data1i_12_port, data1i_11_port, 
      data1i_10_port, data1i_9_port, data1i_8_port, data1i_7_port, 
      data1i_6_port, data1i_5_port, data1i_4_port, data1i_3_port, data1i_2_port
      , data1i_1_port, data1i_0_port, data2i_31_port, data2i_30_port, 
      data2i_29_port, data2i_28_port, data2i_27_port, data2i_26_port, 
      data2i_25_port, data2i_24_port, data2i_23_port, data2i_22_port, 
      data2i_21_port, data2i_20_port, data2i_19_port, data2i_18_port, 
      data2i_17_port, data2i_16_port, data2i_15_port, data2i_14_port, 
      data2i_13_port, data2i_12_port, data2i_11_port, data2i_10_port, 
      data2i_9_port, data2i_8_port, data2i_7_port, data2i_6_port, data2i_5_port
      , data2i_4_port, data2i_3_port, data2i_2_port, data2i_1_port, 
      data2i_0_port, Cin_i, N139, N141, N142, N174, N175, N176, N177, N178, 
      N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, 
      N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, 
      N203, N204, N205, N206, n87, n79, n80, n81, n82, n83, n84, n85, n86, n88,
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139_port, n140, n141_port, n142_port, n143, n144, n145, n146, n147, n148
      , n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174_port, n175_port, n176_port, n177_port, n178_port, n179_port, 
      n180_port, n181_port, n182_port, n183_port, n184_port, n185_port, 
      n186_port, n187_port, n188_port, n189_port, n190_port, n191_port, 
      n192_port, n193_port, n194_port, n195_port, n196_port, n197_port, 
      n198_port, n199_port, n200_port, n201_port, n202_port, n203_port, 
      n204_port, n205_port, n206_port, n207, n208, n209, n210, n211, n212, n213
      , n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139 : std_logic;

begin
   
   Cin_i_reg : DLH_X1 port map( G => n164, D => n87, Q => Cin_i);
   data2i_reg_31_inst : DLH_X1 port map( G => n164, D => N205, Q => 
                           data2i_31_port);
   data2i_reg_30_inst : DLH_X1 port map( G => n162, D => N204, Q => 
                           data2i_30_port);
   data2i_reg_29_inst : DLH_X1 port map( G => n162, D => N203, Q => 
                           data2i_29_port);
   data2i_reg_28_inst : DLH_X1 port map( G => n164, D => N202, Q => 
                           data2i_28_port);
   data2i_reg_27_inst : DLH_X1 port map( G => n162, D => N201, Q => 
                           data2i_27_port);
   data2i_reg_26_inst : DLH_X1 port map( G => n162, D => N200, Q => 
                           data2i_26_port);
   data2i_reg_25_inst : DLH_X1 port map( G => n162, D => N199, Q => 
                           data2i_25_port);
   data2i_reg_24_inst : DLH_X1 port map( G => n162, D => N198, Q => 
                           data2i_24_port);
   data2i_reg_23_inst : DLH_X1 port map( G => n164, D => N197, Q => 
                           data2i_23_port);
   data2i_reg_22_inst : DLH_X1 port map( G => n162, D => N196, Q => 
                           data2i_22_port);
   data2i_reg_21_inst : DLH_X1 port map( G => n163, D => N195, Q => 
                           data2i_21_port);
   data2i_reg_20_inst : DLH_X1 port map( G => n162, D => N194, Q => 
                           data2i_20_port);
   data2i_reg_19_inst : DLH_X1 port map( G => n163, D => N193, Q => 
                           data2i_19_port);
   data2i_reg_18_inst : DLH_X1 port map( G => n163, D => N192, Q => 
                           data2i_18_port);
   data2i_reg_17_inst : DLH_X1 port map( G => n163, D => N191, Q => 
                           data2i_17_port);
   data2i_reg_16_inst : DLH_X1 port map( G => n163, D => N190, Q => 
                           data2i_16_port);
   data2i_reg_15_inst : DLH_X1 port map( G => n164, D => N189, Q => 
                           data2i_15_port);
   data2i_reg_14_inst : DLH_X1 port map( G => n163, D => N188, Q => 
                           data2i_14_port);
   data2i_reg_13_inst : DLH_X1 port map( G => n163, D => N187, Q => 
                           data2i_13_port);
   data2i_reg_12_inst : DLH_X1 port map( G => n163, D => N186, Q => 
                           data2i_12_port);
   data2i_reg_11_inst : DLH_X1 port map( G => n162, D => N185, Q => 
                           data2i_11_port);
   data2i_reg_10_inst : DLH_X1 port map( G => n162, D => N184, Q => 
                           data2i_10_port);
   data2i_reg_9_inst : DLH_X1 port map( G => n163, D => N183, Q => 
                           data2i_9_port);
   data2i_reg_8_inst : DLH_X1 port map( G => n162, D => N182, Q => 
                           data2i_8_port);
   data2i_reg_7_inst : DLH_X1 port map( G => n164, D => N181, Q => 
                           data2i_7_port);
   data2i_reg_6_inst : DLH_X1 port map( G => n164, D => N180, Q => 
                           data2i_6_port);
   data2i_reg_5_inst : DLH_X1 port map( G => n163, D => N179, Q => 
                           data2i_5_port);
   data2i_reg_4_inst : DLH_X1 port map( G => n163, D => N178, Q => 
                           data2i_4_port);
   data2i_reg_3_inst : DLH_X1 port map( G => n163, D => N177, Q => 
                           data2i_3_port);
   data2i_reg_2_inst : DLH_X1 port map( G => n162, D => N176, Q => 
                           data2i_2_port);
   data2i_reg_1_inst : DLH_X1 port map( G => n163, D => N175, Q => 
                           data2i_1_port);
   data2i_reg_0_inst : DLH_X1 port map( G => n164, D => N174, Q => 
                           data2i_0_port);
   data1i_reg_31_inst : DLH_X1 port map( G => n164, D => DATA1(31), Q => 
                           data1i_31_port);
   data1i_reg_30_inst : DLH_X1 port map( G => n162, D => DATA1(30), Q => 
                           data1i_30_port);
   data1i_reg_29_inst : DLH_X1 port map( G => n162, D => DATA1(29), Q => 
                           data1i_29_port);
   data1i_reg_28_inst : DLH_X1 port map( G => n164, D => DATA1(28), Q => 
                           data1i_28_port);
   data1i_reg_27_inst : DLH_X1 port map( G => n162, D => DATA1(27), Q => 
                           data1i_27_port);
   data1i_reg_26_inst : DLH_X1 port map( G => n162, D => DATA1(26), Q => 
                           data1i_26_port);
   data1i_reg_25_inst : DLH_X1 port map( G => n162, D => DATA1(25), Q => 
                           data1i_25_port);
   data1i_reg_24_inst : DLH_X1 port map( G => n162, D => DATA1(24), Q => 
                           data1i_24_port);
   data1i_reg_23_inst : DLH_X1 port map( G => n164, D => DATA1(23), Q => 
                           data1i_23_port);
   data1i_reg_22_inst : DLH_X1 port map( G => n162, D => DATA1(22), Q => 
                           data1i_22_port);
   data1i_reg_21_inst : DLH_X1 port map( G => n163, D => DATA1(21), Q => 
                           data1i_21_port);
   data1i_reg_20_inst : DLH_X1 port map( G => n162, D => DATA1(20), Q => 
                           data1i_20_port);
   data1i_reg_19_inst : DLH_X1 port map( G => n164, D => DATA1(19), Q => 
                           data1i_19_port);
   data1i_reg_18_inst : DLH_X1 port map( G => n163, D => DATA1(18), Q => 
                           data1i_18_port);
   data1i_reg_17_inst : DLH_X1 port map( G => n163, D => DATA1(17), Q => 
                           data1i_17_port);
   data1i_reg_16_inst : DLH_X1 port map( G => n163, D => DATA1(16), Q => 
                           data1i_16_port);
   data1i_reg_15_inst : DLH_X1 port map( G => n164, D => DATA1(15), Q => 
                           data1i_15_port);
   data1i_reg_14_inst : DLH_X1 port map( G => n163, D => DATA1(14), Q => 
                           data1i_14_port);
   data1i_reg_13_inst : DLH_X1 port map( G => n163, D => DATA1(13), Q => 
                           data1i_13_port);
   data1i_reg_12_inst : DLH_X1 port map( G => n163, D => DATA1(12), Q => 
                           data1i_12_port);
   data1i_reg_11_inst : DLH_X1 port map( G => n162, D => DATA1(11), Q => 
                           data1i_11_port);
   data1i_reg_10_inst : DLH_X1 port map( G => n162, D => DATA1(10), Q => 
                           data1i_10_port);
   data1i_reg_9_inst : DLH_X1 port map( G => n163, D => DATA1(9), Q => 
                           data1i_9_port);
   data1i_reg_8_inst : DLH_X1 port map( G => n162, D => DATA1(8), Q => 
                           data1i_8_port);
   data1i_reg_7_inst : DLH_X1 port map( G => n164, D => DATA1(7), Q => 
                           data1i_7_port);
   data1i_reg_6_inst : DLH_X1 port map( G => n164, D => DATA1(6), Q => 
                           data1i_6_port);
   data1i_reg_5_inst : DLH_X1 port map( G => n163, D => DATA1(5), Q => 
                           data1i_5_port);
   data1i_reg_4_inst : DLH_X1 port map( G => n163, D => DATA1(4), Q => 
                           data1i_4_port);
   data1i_reg_3_inst : DLH_X1 port map( G => n163, D => DATA1(3), Q => 
                           data1i_3_port);
   data1i_reg_2_inst : DLH_X1 port map( G => n163, D => DATA1(2), Q => 
                           data1i_2_port);
   data1i_reg_1_inst : DLH_X1 port map( G => n163, D => DATA1(1), Q => 
                           data1i_1_port);
   data1i_reg_0_inst : DLH_X1 port map( G => n164, D => DATA1(0), Q => 
                           data1i_0_port);
   LOGIC_ARITH_i_reg : DLH_X1 port map( G => n157, D => n142_port, Q => 
                           LOGIC_ARITH_i);
   LEFT_RIGHT_i_reg : DLH_X1 port map( G => n157, D => n142_port, Q => 
                           LEFT_RIGHT_i);
   OUTPUT_alu_i_reg_0_inst : DLH_X1 port map( G => n158, D => N142, Q => 
                           OUTPUT_alu_i_0_port);
   OUT_ALU_reg_0_inst : DFF_X1 port map( D => OUTPUT_alu_i_0_port, CK => CLK, Q
                           => OUT_ALU(0), QN => n_1077);
   OUTPUT_alu_i_reg_1_inst : DLH_X1 port map( G => n161, D => n197_port, Q => 
                           OUTPUT_alu_i_1_port);
   OUT_ALU_reg_1_inst : DFF_X1 port map( D => OUTPUT_alu_i_1_port, CK => CLK, Q
                           => OUT_ALU(1), QN => n_1078);
   OUTPUT_alu_i_reg_2_inst : DLH_X1 port map( G => n160, D => n195_port, Q => 
                           OUTPUT_alu_i_2_port);
   OUT_ALU_reg_2_inst : DFF_X1 port map( D => OUTPUT_alu_i_2_port, CK => CLK, Q
                           => OUT_ALU(2), QN => n_1079);
   OUTPUT_alu_i_reg_3_inst : DLH_X1 port map( G => n159, D => n199_port, Q => 
                           OUTPUT_alu_i_3_port);
   OUT_ALU_reg_3_inst : DFF_X1 port map( D => OUTPUT_alu_i_3_port, CK => CLK, Q
                           => OUT_ALU(3), QN => n_1080);
   OUTPUT_alu_i_reg_4_inst : DLH_X1 port map( G => n160, D => n194_port, Q => 
                           OUTPUT_alu_i_4_port);
   OUT_ALU_reg_4_inst : DFF_X1 port map( D => OUTPUT_alu_i_4_port, CK => CLK, Q
                           => OUT_ALU(4), QN => n_1081);
   OUTPUT_alu_i_reg_5_inst : DLH_X1 port map( G => n160, D => n198_port, Q => 
                           OUTPUT_alu_i_5_port);
   OUT_ALU_reg_5_inst : DFF_X1 port map( D => OUTPUT_alu_i_5_port, CK => CLK, Q
                           => OUT_ALU(5), QN => n_1082);
   OUTPUT_alu_i_reg_6_inst : DLH_X1 port map( G => n158, D => n196_port, Q => 
                           OUTPUT_alu_i_6_port);
   OUT_ALU_reg_6_inst : DFF_X1 port map( D => OUTPUT_alu_i_6_port, CK => CLK, Q
                           => OUT_ALU(6), QN => n_1083);
   OUTPUT_alu_i_reg_7_inst : DLH_X1 port map( G => n158, D => n200_port, Q => 
                           OUTPUT_alu_i_7_port);
   OUT_ALU_reg_7_inst : DFF_X1 port map( D => OUTPUT_alu_i_7_port, CK => CLK, Q
                           => OUT_ALU(7), QN => n_1084);
   OUTPUT_alu_i_reg_8_inst : DLH_X1 port map( G => n159, D => n173, Q => 
                           OUTPUT_alu_i_8_port);
   OUT_ALU_reg_8_inst : DFF_X1 port map( D => OUTPUT_alu_i_8_port, CK => CLK, Q
                           => OUT_ALU(8), QN => n_1085);
   OUTPUT_alu_i_reg_9_inst : DLH_X1 port map( G => n159, D => n172, Q => 
                           OUTPUT_alu_i_9_port);
   OUT_ALU_reg_9_inst : DFF_X1 port map( D => OUTPUT_alu_i_9_port, CK => CLK, Q
                           => OUT_ALU(9), QN => n_1086);
   OUTPUT_alu_i_reg_10_inst : DLH_X1 port map( G => n159, D => n171, Q => 
                           OUTPUT_alu_i_10_port);
   OUT_ALU_reg_10_inst : DFF_X1 port map( D => OUTPUT_alu_i_10_port, CK => CLK,
                           Q => OUT_ALU(10), QN => n_1087);
   OUTPUT_alu_i_reg_11_inst : DLH_X1 port map( G => n159, D => n170, Q => 
                           OUTPUT_alu_i_11_port);
   OUT_ALU_reg_11_inst : DFF_X1 port map( D => OUTPUT_alu_i_11_port, CK => CLK,
                           Q => OUT_ALU(11), QN => n_1088);
   OUTPUT_alu_i_reg_12_inst : DLH_X1 port map( G => n160, D => n177_port, Q => 
                           OUTPUT_alu_i_12_port);
   OUT_ALU_reg_12_inst : DFF_X1 port map( D => OUTPUT_alu_i_12_port, CK => CLK,
                           Q => OUT_ALU(12), QN => n_1089);
   OUTPUT_alu_i_reg_13_inst : DLH_X1 port map( G => n160, D => n176_port, Q => 
                           OUTPUT_alu_i_13_port);
   OUT_ALU_reg_13_inst : DFF_X1 port map( D => OUTPUT_alu_i_13_port, CK => CLK,
                           Q => OUT_ALU(13), QN => n_1090);
   OUTPUT_alu_i_reg_14_inst : DLH_X1 port map( G => n160, D => n175_port, Q => 
                           OUTPUT_alu_i_14_port);
   OUT_ALU_reg_14_inst : DFF_X1 port map( D => OUTPUT_alu_i_14_port, CK => CLK,
                           Q => OUT_ALU(14), QN => n_1091);
   OUTPUT_alu_i_reg_15_inst : DLH_X1 port map( G => n158, D => n174_port, Q => 
                           OUTPUT_alu_i_15_port);
   OUT_ALU_reg_15_inst : DFF_X1 port map( D => OUTPUT_alu_i_15_port, CK => CLK,
                           Q => OUT_ALU(15), QN => n_1092);
   OUTPUT_alu_i_reg_16_inst : DLH_X1 port map( G => n160, D => n181_port, Q => 
                           OUTPUT_alu_i_16_port);
   OUT_ALU_reg_16_inst : DFF_X1 port map( D => OUTPUT_alu_i_16_port, CK => CLK,
                           Q => OUT_ALU(16), QN => n_1093);
   OUTPUT_alu_i_reg_17_inst : DLH_X1 port map( G => n160, D => n180_port, Q => 
                           OUTPUT_alu_i_17_port);
   OUT_ALU_reg_17_inst : DFF_X1 port map( D => OUTPUT_alu_i_17_port, CK => CLK,
                           Q => OUT_ALU(17), QN => n_1094);
   OUTPUT_alu_i_reg_18_inst : DLH_X1 port map( G => n161, D => n179_port, Q => 
                           OUTPUT_alu_i_18_port);
   OUT_ALU_reg_18_inst : DFF_X1 port map( D => OUTPUT_alu_i_18_port, CK => CLK,
                           Q => OUT_ALU(18), QN => n_1095);
   OUTPUT_alu_i_reg_19_inst : DLH_X1 port map( G => n158, D => n178_port, Q => 
                           OUTPUT_alu_i_19_port);
   OUT_ALU_reg_19_inst : DFF_X1 port map( D => OUTPUT_alu_i_19_port, CK => CLK,
                           Q => OUT_ALU(19), QN => n_1096);
   OUTPUT_alu_i_reg_20_inst : DLH_X1 port map( G => n160, D => n185_port, Q => 
                           OUTPUT_alu_i_20_port);
   OUT_ALU_reg_20_inst : DFF_X1 port map( D => OUTPUT_alu_i_20_port, CK => CLK,
                           Q => OUT_ALU(20), QN => n_1097);
   OUTPUT_alu_i_reg_21_inst : DLH_X1 port map( G => n159, D => n184_port, Q => 
                           OUTPUT_alu_i_21_port);
   OUT_ALU_reg_21_inst : DFF_X1 port map( D => OUTPUT_alu_i_21_port, CK => CLK,
                           Q => OUT_ALU(21), QN => n_1098);
   OUTPUT_alu_i_reg_22_inst : DLH_X1 port map( G => n159, D => n183_port, Q => 
                           OUTPUT_alu_i_22_port);
   OUT_ALU_reg_22_inst : DFF_X1 port map( D => OUTPUT_alu_i_22_port, CK => CLK,
                           Q => OUT_ALU(22), QN => n_1099);
   OUTPUT_alu_i_reg_23_inst : DLH_X1 port map( G => n158, D => n182_port, Q => 
                           OUTPUT_alu_i_23_port);
   OUT_ALU_reg_23_inst : DFF_X1 port map( D => OUTPUT_alu_i_23_port, CK => CLK,
                           Q => OUT_ALU(23), QN => n_1100);
   OUTPUT_alu_i_reg_24_inst : DLH_X1 port map( G => n160, D => n189_port, Q => 
                           OUTPUT_alu_i_24_port);
   OUT_ALU_reg_24_inst : DFF_X1 port map( D => OUTPUT_alu_i_24_port, CK => CLK,
                           Q => OUT_ALU(24), QN => n_1101);
   OUTPUT_alu_i_reg_25_inst : DLH_X1 port map( G => n159, D => n188_port, Q => 
                           OUTPUT_alu_i_25_port);
   OUT_ALU_reg_25_inst : DFF_X1 port map( D => OUTPUT_alu_i_25_port, CK => CLK,
                           Q => OUT_ALU(25), QN => n_1102);
   OUTPUT_alu_i_reg_26_inst : DLH_X1 port map( G => n159, D => n187_port, Q => 
                           OUTPUT_alu_i_26_port);
   OUT_ALU_reg_26_inst : DFF_X1 port map( D => OUTPUT_alu_i_26_port, CK => CLK,
                           Q => OUT_ALU(26), QN => n_1103);
   OUTPUT_alu_i_reg_27_inst : DLH_X1 port map( G => n159, D => n186_port, Q => 
                           OUTPUT_alu_i_27_port);
   OUT_ALU_reg_27_inst : DFF_X1 port map( D => OUTPUT_alu_i_27_port, CK => CLK,
                           Q => OUT_ALU(27), QN => n_1104);
   OUTPUT_alu_i_reg_28_inst : DLH_X1 port map( G => n158, D => n193_port, Q => 
                           OUTPUT_alu_i_28_port);
   OUT_ALU_reg_28_inst : DFF_X1 port map( D => OUTPUT_alu_i_28_port, CK => CLK,
                           Q => OUT_ALU(28), QN => n_1105);
   OUTPUT_alu_i_reg_29_inst : DLH_X1 port map( G => n158, D => n192_port, Q => 
                           OUTPUT_alu_i_29_port);
   OUT_ALU_reg_29_inst : DFF_X1 port map( D => OUTPUT_alu_i_29_port, CK => CLK,
                           Q => OUT_ALU(29), QN => n_1106);
   OUTPUT_alu_i_reg_30_inst : DLH_X1 port map( G => n158, D => n191_port, Q => 
                           OUTPUT_alu_i_30_port);
   OUT_ALU_reg_30_inst : DFF_X1 port map( D => OUTPUT_alu_i_30_port, CK => CLK,
                           Q => OUT_ALU(30), QN => n_1107);
   OUTPUT_alu_i_reg_31_inst : DLH_X1 port map( G => n158, D => n190_port, Q => 
                           OUTPUT_alu_i_31_port);
   OUT_ALU_reg_31_inst : DFF_X1 port map( D => OUTPUT_alu_i_31_port, CK => CLK,
                           Q => OUT_ALU(31), QN => n_1108);
   SHIFT_ROTATE_i <= '1';
   U177 : NAND3_X1 port map( A1 => n112, A2 => n113, A3 => n229, ZN => n87);
   U178 : OAI33_X1 port map( A1 => n131, A2 => n239, A3 => n240, B1 => n132, B2
                           => FUNC(2), B3 => FUNC(3), ZN => n130);
   U179 : NAND3_X1 port map( A1 => n112, A2 => n113, A3 => n151, ZN => n80);
   U180 : NAND3_X1 port map( A1 => FUNC(2), A2 => n237, A3 => FUNC(0), ZN => 
                           n131);
   U181 : NAND3_X1 port map( A1 => n140, A2 => n126, A3 => n235, ZN => 
                           n139_port);
   log : logic_N32 port map( FUNC(0) => FUNC(0), FUNC(1) => FUNC(1), FUNC(2) =>
                           FUNC(2), FUNC(3) => FUNC(3), FUNC(4) => FUNC(4), 
                           FUNC(5) => FUNC(5), DATA1(31) => DATA1(31), 
                           DATA1(30) => DATA1(30), DATA1(29) => DATA1(29), 
                           DATA1(28) => DATA1(28), DATA1(27) => DATA1(27), 
                           DATA1(26) => DATA1(26), DATA1(25) => DATA1(25), 
                           DATA1(24) => DATA1(24), DATA1(23) => DATA1(23), 
                           DATA1(22) => DATA1(22), DATA1(21) => DATA1(21), 
                           DATA1(20) => DATA1(20), DATA1(19) => DATA1(19), 
                           DATA1(18) => DATA1(18), DATA1(17) => DATA1(17), 
                           DATA1(16) => DATA1(16), DATA1(15) => DATA1(15), 
                           DATA1(14) => DATA1(14), DATA1(13) => DATA1(13), 
                           DATA1(12) => DATA1(12), DATA1(11) => DATA1(11), 
                           DATA1(10) => DATA1(10), DATA1(9) => DATA1(9), 
                           DATA1(8) => DATA1(8), DATA1(7) => DATA1(7), DATA1(6)
                           => DATA1(6), DATA1(5) => DATA1(5), DATA1(4) => 
                           DATA1(4), DATA1(3) => DATA1(3), DATA1(2) => DATA1(2)
                           , DATA1(1) => DATA1(1), DATA1(0) => DATA1(0), 
                           DATA2(31) => DATA2(31), DATA2(30) => DATA2(30), 
                           DATA2(29) => DATA2(29), DATA2(28) => DATA2(28), 
                           DATA2(27) => DATA2(27), DATA2(26) => DATA2(26), 
                           DATA2(25) => DATA2(25), DATA2(24) => DATA2(24), 
                           DATA2(23) => DATA2(23), DATA2(22) => DATA2(22), 
                           DATA2(21) => DATA2(21), DATA2(20) => DATA2(20), 
                           DATA2(19) => DATA2(19), DATA2(18) => DATA2(18), 
                           DATA2(17) => DATA2(17), DATA2(16) => DATA2(16), 
                           DATA2(15) => DATA2(15), DATA2(14) => DATA2(14), 
                           DATA2(13) => DATA2(13), DATA2(12) => DATA2(12), 
                           DATA2(11) => DATA2(11), DATA2(10) => DATA2(10), 
                           DATA2(9) => DATA2(9), DATA2(8) => DATA2(8), DATA2(7)
                           => DATA2(7), DATA2(6) => DATA2(6), DATA2(5) => 
                           DATA2(5), DATA2(4) => DATA2(4), DATA2(3) => DATA2(3)
                           , DATA2(2) => DATA2(2), DATA2(1) => DATA2(1), 
                           DATA2(0) => DATA2(0), OUT_ALU(31) => OUTPUT4_31_port
                           , OUT_ALU(30) => OUTPUT4_30_port, OUT_ALU(29) => 
                           OUTPUT4_29_port, OUT_ALU(28) => OUTPUT4_28_port, 
                           OUT_ALU(27) => OUTPUT4_27_port, OUT_ALU(26) => 
                           OUTPUT4_26_port, OUT_ALU(25) => OUTPUT4_25_port, 
                           OUT_ALU(24) => OUTPUT4_24_port, OUT_ALU(23) => 
                           OUTPUT4_23_port, OUT_ALU(22) => OUTPUT4_22_port, 
                           OUT_ALU(21) => OUTPUT4_21_port, OUT_ALU(20) => 
                           OUTPUT4_20_port, OUT_ALU(19) => OUTPUT4_19_port, 
                           OUT_ALU(18) => OUTPUT4_18_port, OUT_ALU(17) => 
                           OUTPUT4_17_port, OUT_ALU(16) => OUTPUT4_16_port, 
                           OUT_ALU(15) => OUTPUT4_15_port, OUT_ALU(14) => 
                           OUTPUT4_14_port, OUT_ALU(13) => OUTPUT4_13_port, 
                           OUT_ALU(12) => OUTPUT4_12_port, OUT_ALU(11) => 
                           OUTPUT4_11_port, OUT_ALU(10) => OUTPUT4_10_port, 
                           OUT_ALU(9) => OUTPUT4_9_port, OUT_ALU(8) => 
                           OUTPUT4_8_port, OUT_ALU(7) => OUTPUT4_7_port, 
                           OUT_ALU(6) => OUTPUT4_6_port, OUT_ALU(5) => 
                           OUTPUT4_5_port, OUT_ALU(4) => OUTPUT4_4_port, 
                           OUT_ALU(3) => OUTPUT4_3_port, OUT_ALU(2) => 
                           OUTPUT4_2_port, OUT_ALU(1) => OUTPUT4_1_port, 
                           OUT_ALU(0) => OUTPUT4_0_port);
   comp : comparator port map( DATA1(31) => OUTPUT2_31_port, DATA1(30) => 
                           OUTPUT2_30_port, DATA1(29) => OUTPUT2_29_port, 
                           DATA1(28) => OUTPUT2_28_port, DATA1(27) => 
                           OUTPUT2_27_port, DATA1(26) => OUTPUT2_26_port, 
                           DATA1(25) => OUTPUT2_25_port, DATA1(24) => 
                           OUTPUT2_24_port, DATA1(23) => OUTPUT2_23_port, 
                           DATA1(22) => OUTPUT2_22_port, DATA1(21) => 
                           OUTPUT2_21_port, DATA1(20) => OUTPUT2_20_port, 
                           DATA1(19) => OUTPUT2_19_port, DATA1(18) => 
                           OUTPUT2_18_port, DATA1(17) => OUTPUT2_17_port, 
                           DATA1(16) => OUTPUT2_16_port, DATA1(15) => 
                           OUTPUT2_15_port, DATA1(14) => OUTPUT2_14_port, 
                           DATA1(13) => OUTPUT2_13_port, DATA1(12) => 
                           OUTPUT2_12_port, DATA1(11) => OUTPUT2_11_port, 
                           DATA1(10) => OUTPUT2_10_port, DATA1(9) => 
                           OUTPUT2_9_port, DATA1(8) => OUTPUT2_8_port, DATA1(7)
                           => OUTPUT2_7_port, DATA1(6) => OUTPUT2_6_port, 
                           DATA1(5) => OUTPUT2_5_port, DATA1(4) => 
                           OUTPUT2_4_port, DATA1(3) => OUTPUT2_3_port, DATA1(2)
                           => OUTPUT2_2_port, DATA1(1) => OUTPUT2_1_port, 
                           DATA1(0) => OUTPUT2_0_port, DATA2i => Cout_i, 
                           tipo(0) => FUNC(0), tipo(1) => FUNC(1), tipo(2) => 
                           FUNC(2), tipo(3) => FUNC(3), tipo(4) => FUNC(4), 
                           tipo(5) => FUNC(5), OUTALU(31) => n_1109, OUTALU(30)
                           => n_1110, OUTALU(29) => n_1111, OUTALU(28) => 
                           n_1112, OUTALU(27) => n_1113, OUTALU(26) => n_1114, 
                           OUTALU(25) => n_1115, OUTALU(24) => n_1116, 
                           OUTALU(23) => n_1117, OUTALU(22) => n_1118, 
                           OUTALU(21) => n_1119, OUTALU(20) => n_1120, 
                           OUTALU(19) => n_1121, OUTALU(18) => n_1122, 
                           OUTALU(17) => n_1123, OUTALU(16) => n_1124, 
                           OUTALU(15) => n_1125, OUTALU(14) => n_1126, 
                           OUTALU(13) => n_1127, OUTALU(12) => n_1128, 
                           OUTALU(11) => n_1129, OUTALU(10) => n_1130, 
                           OUTALU(9) => n_1131, OUTALU(8) => n_1132, OUTALU(7) 
                           => n_1133, OUTALU(6) => n_1134, OUTALU(5) => n_1135,
                           OUTALU(4) => n_1136, OUTALU(3) => n_1137, OUTALU(2) 
                           => n_1138, OUTALU(1) => n_1139, OUTALU(0) => 
                           OUTPUT3_0_port);
   shifter : SHIFTER_GENERIC_N32 port map( A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28), 
                           A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), B(4) => 
                           DATA2(4), B(3) => DATA2(3), B(2) => DATA2(2), B(1) 
                           => DATA2(1), B(0) => DATA2(0), LOGIC_ARITH => 
                           LOGIC_ARITH_i, LEFT_RIGHT => LEFT_RIGHT_i, 
                           SHIFT_ROTATE => SHIFT_ROTATE_i, OUTPUT(31) => 
                           OUTPUT1_31_port, OUTPUT(30) => OUTPUT1_30_port, 
                           OUTPUT(29) => OUTPUT1_29_port, OUTPUT(28) => 
                           OUTPUT1_28_port, OUTPUT(27) => OUTPUT1_27_port, 
                           OUTPUT(26) => OUTPUT1_26_port, OUTPUT(25) => 
                           OUTPUT1_25_port, OUTPUT(24) => OUTPUT1_24_port, 
                           OUTPUT(23) => OUTPUT1_23_port, OUTPUT(22) => 
                           OUTPUT1_22_port, OUTPUT(21) => OUTPUT1_21_port, 
                           OUTPUT(20) => OUTPUT1_20_port, OUTPUT(19) => 
                           OUTPUT1_19_port, OUTPUT(18) => OUTPUT1_18_port, 
                           OUTPUT(17) => OUTPUT1_17_port, OUTPUT(16) => 
                           OUTPUT1_16_port, OUTPUT(15) => OUTPUT1_15_port, 
                           OUTPUT(14) => OUTPUT1_14_port, OUTPUT(13) => 
                           OUTPUT1_13_port, OUTPUT(12) => OUTPUT1_12_port, 
                           OUTPUT(11) => OUTPUT1_11_port, OUTPUT(10) => 
                           OUTPUT1_10_port, OUTPUT(9) => OUTPUT1_9_port, 
                           OUTPUT(8) => OUTPUT1_8_port, OUTPUT(7) => 
                           OUTPUT1_7_port, OUTPUT(6) => OUTPUT1_6_port, 
                           OUTPUT(5) => OUTPUT1_5_port, OUTPUT(4) => 
                           OUTPUT1_4_port, OUTPUT(3) => OUTPUT1_3_port, 
                           OUTPUT(2) => OUTPUT1_2_port, OUTPUT(1) => 
                           OUTPUT1_1_port, OUTPUT(0) => OUTPUT1_0_port);
   adder : P4_ADDER_NBIT32 port map( A(31) => data1i_31_port, A(30) => 
                           data1i_30_port, A(29) => data1i_29_port, A(28) => 
                           data1i_28_port, A(27) => data1i_27_port, A(26) => 
                           data1i_26_port, A(25) => data1i_25_port, A(24) => 
                           data1i_24_port, A(23) => data1i_23_port, A(22) => 
                           data1i_22_port, A(21) => data1i_21_port, A(20) => 
                           data1i_20_port, A(19) => data1i_19_port, A(18) => 
                           data1i_18_port, A(17) => data1i_17_port, A(16) => 
                           data1i_16_port, A(15) => data1i_15_port, A(14) => 
                           data1i_14_port, A(13) => data1i_13_port, A(12) => 
                           data1i_12_port, A(11) => data1i_11_port, A(10) => 
                           data1i_10_port, A(9) => data1i_9_port, A(8) => 
                           data1i_8_port, A(7) => data1i_7_port, A(6) => 
                           data1i_6_port, A(5) => data1i_5_port, A(4) => 
                           data1i_4_port, A(3) => data1i_3_port, A(2) => 
                           data1i_2_port, A(1) => data1i_1_port, A(0) => 
                           data1i_0_port, B(31) => data2i_31_port, B(30) => 
                           data2i_30_port, B(29) => data2i_29_port, B(28) => 
                           data2i_28_port, B(27) => data2i_27_port, B(26) => 
                           data2i_26_port, B(25) => data2i_25_port, B(24) => 
                           data2i_24_port, B(23) => data2i_23_port, B(22) => 
                           data2i_22_port, B(21) => data2i_21_port, B(20) => 
                           data2i_20_port, B(19) => data2i_19_port, B(18) => 
                           data2i_18_port, B(17) => data2i_17_port, B(16) => 
                           data2i_16_port, B(15) => data2i_15_port, B(14) => 
                           data2i_14_port, B(13) => data2i_13_port, B(12) => 
                           data2i_12_port, B(11) => data2i_11_port, B(10) => 
                           data2i_10_port, B(9) => data2i_9_port, B(8) => 
                           data2i_8_port, B(7) => data2i_7_port, B(6) => 
                           data2i_6_port, B(5) => data2i_5_port, B(4) => 
                           data2i_4_port, B(3) => data2i_3_port, B(2) => 
                           data2i_2_port, B(1) => data2i_1_port, B(0) => 
                           data2i_0_port, Cin => Cin_i, S(31) => 
                           OUTPUT2_31_port, S(30) => OUTPUT2_30_port, S(29) => 
                           OUTPUT2_29_port, S(28) => OUTPUT2_28_port, S(27) => 
                           OUTPUT2_27_port, S(26) => OUTPUT2_26_port, S(25) => 
                           OUTPUT2_25_port, S(24) => OUTPUT2_24_port, S(23) => 
                           OUTPUT2_23_port, S(22) => OUTPUT2_22_port, S(21) => 
                           OUTPUT2_21_port, S(20) => OUTPUT2_20_port, S(19) => 
                           OUTPUT2_19_port, S(18) => OUTPUT2_18_port, S(17) => 
                           OUTPUT2_17_port, S(16) => OUTPUT2_16_port, S(15) => 
                           OUTPUT2_15_port, S(14) => OUTPUT2_14_port, S(13) => 
                           OUTPUT2_13_port, S(12) => OUTPUT2_12_port, S(11) => 
                           OUTPUT2_11_port, S(10) => OUTPUT2_10_port, S(9) => 
                           OUTPUT2_9_port, S(8) => OUTPUT2_8_port, S(7) => 
                           OUTPUT2_7_port, S(6) => OUTPUT2_6_port, S(5) => 
                           OUTPUT2_5_port, S(4) => OUTPUT2_4_port, S(3) => 
                           OUTPUT2_3_port, S(2) => OUTPUT2_2_port, S(1) => 
                           OUTPUT2_1_port, S(0) => OUTPUT2_0_port, Cout => 
                           Cout_i);
   U4 : BUF_X1 port map( A => N139, Z => n163);
   U5 : BUF_X1 port map( A => n228, Z => n143);
   U6 : BUF_X1 port map( A => n228, Z => n144);
   U7 : BUF_X1 port map( A => N139, Z => n162);
   U8 : BUF_X1 port map( A => n228, Z => n145);
   U9 : BUF_X1 port map( A => N139, Z => n164);
   U10 : BUF_X1 port map( A => n80, Z => n152);
   U11 : BUF_X1 port map( A => n80, Z => n153);
   U12 : BUF_X1 port map( A => n80, Z => n154);
   U13 : INV_X1 port map( A => n140, ZN => n234);
   U14 : INV_X1 port map( A => n87, ZN => n228);
   U15 : INV_X1 port map( A => n118, ZN => n240);
   U16 : OR2_X1 port map( A1 => n154, A2 => n114, ZN => N139);
   U17 : OR3_X1 port map( A1 => n162, A2 => n155, A3 => n148, ZN => N141);
   U18 : INV_X1 port map( A => n111, ZN => n190_port);
   U19 : AOI222_X1 port map( A1 => OUTPUT1_31_port, A2 => n155, B1 => 
                           OUTPUT4_31_port, B2 => n148, C1 => OUTPUT2_31_port, 
                           C2 => n154, ZN => n111);
   U20 : INV_X1 port map( A => n110, ZN => n191_port);
   U21 : AOI222_X1 port map( A1 => OUTPUT1_30_port, A2 => n157, B1 => 
                           OUTPUT4_30_port, B2 => n148, C1 => OUTPUT2_30_port, 
                           C2 => n154, ZN => n110);
   U22 : INV_X1 port map( A => n109, ZN => n192_port);
   U23 : AOI222_X1 port map( A1 => OUTPUT1_29_port, A2 => n157, B1 => 
                           OUTPUT4_29_port, B2 => n148, C1 => OUTPUT2_29_port, 
                           C2 => n154, ZN => n109);
   U24 : INV_X1 port map( A => n108, ZN => n193_port);
   U25 : AOI222_X1 port map( A1 => OUTPUT1_28_port, A2 => n157, B1 => 
                           OUTPUT4_28_port, B2 => n148, C1 => OUTPUT2_28_port, 
                           C2 => n154, ZN => n108);
   U26 : INV_X1 port map( A => n107, ZN => n186_port);
   U27 : AOI222_X1 port map( A1 => OUTPUT1_27_port, A2 => n157, B1 => 
                           OUTPUT4_27_port, B2 => n148, C1 => OUTPUT2_27_port, 
                           C2 => n154, ZN => n107);
   U28 : INV_X1 port map( A => n106, ZN => n187_port);
   U29 : AOI222_X1 port map( A1 => OUTPUT1_26_port, A2 => n157, B1 => 
                           OUTPUT4_26_port, B2 => n148, C1 => OUTPUT2_26_port, 
                           C2 => n154, ZN => n106);
   U30 : INV_X1 port map( A => n105, ZN => n188_port);
   U31 : AOI222_X1 port map( A1 => OUTPUT1_25_port, A2 => n157, B1 => 
                           OUTPUT4_25_port, B2 => n148, C1 => OUTPUT2_25_port, 
                           C2 => n154, ZN => n105);
   U32 : INV_X1 port map( A => n104, ZN => n189_port);
   U33 : AOI222_X1 port map( A1 => OUTPUT1_24_port, A2 => n157, B1 => 
                           OUTPUT4_24_port, B2 => n148, C1 => OUTPUT2_24_port, 
                           C2 => n154, ZN => n104);
   U34 : INV_X1 port map( A => n103, ZN => n182_port);
   U35 : AOI222_X1 port map( A1 => OUTPUT1_23_port, A2 => n157, B1 => 
                           OUTPUT4_23_port, B2 => n147, C1 => OUTPUT2_23_port, 
                           C2 => n153, ZN => n103);
   U36 : INV_X1 port map( A => n102, ZN => n183_port);
   U37 : AOI222_X1 port map( A1 => OUTPUT1_22_port, A2 => n157, B1 => 
                           OUTPUT4_22_port, B2 => n147, C1 => OUTPUT2_22_port, 
                           C2 => n153, ZN => n102);
   U38 : INV_X1 port map( A => n101, ZN => n184_port);
   U39 : AOI222_X1 port map( A1 => OUTPUT1_21_port, A2 => n156, B1 => 
                           OUTPUT4_21_port, B2 => n147, C1 => OUTPUT2_21_port, 
                           C2 => n153, ZN => n101);
   U40 : INV_X1 port map( A => n100, ZN => n185_port);
   U41 : AOI222_X1 port map( A1 => OUTPUT1_20_port, A2 => n156, B1 => 
                           OUTPUT4_20_port, B2 => n147, C1 => OUTPUT2_20_port, 
                           C2 => n153, ZN => n100);
   U42 : INV_X1 port map( A => n99, ZN => n178_port);
   U43 : AOI222_X1 port map( A1 => OUTPUT1_19_port, A2 => n156, B1 => 
                           OUTPUT4_19_port, B2 => n147, C1 => OUTPUT2_19_port, 
                           C2 => n153, ZN => n99);
   U44 : INV_X1 port map( A => n98, ZN => n179_port);
   U45 : AOI222_X1 port map( A1 => OUTPUT1_18_port, A2 => n156, B1 => 
                           OUTPUT4_18_port, B2 => n147, C1 => OUTPUT2_18_port, 
                           C2 => n153, ZN => n98);
   U46 : INV_X1 port map( A => n97, ZN => n180_port);
   U47 : AOI222_X1 port map( A1 => OUTPUT1_17_port, A2 => n156, B1 => 
                           OUTPUT4_17_port, B2 => n147, C1 => OUTPUT2_17_port, 
                           C2 => n153, ZN => n97);
   U48 : INV_X1 port map( A => n96, ZN => n181_port);
   U49 : AOI222_X1 port map( A1 => OUTPUT1_16_port, A2 => n156, B1 => 
                           OUTPUT4_16_port, B2 => n147, C1 => OUTPUT2_16_port, 
                           C2 => n153, ZN => n96);
   U50 : INV_X1 port map( A => n95, ZN => n174_port);
   U51 : AOI222_X1 port map( A1 => OUTPUT1_15_port, A2 => n156, B1 => 
                           OUTPUT4_15_port, B2 => n147, C1 => OUTPUT2_15_port, 
                           C2 => n153, ZN => n95);
   U52 : INV_X1 port map( A => n94, ZN => n175_port);
   U53 : AOI222_X1 port map( A1 => OUTPUT1_14_port, A2 => n156, B1 => 
                           OUTPUT4_14_port, B2 => n147, C1 => OUTPUT2_14_port, 
                           C2 => n153, ZN => n94);
   U54 : INV_X1 port map( A => n93, ZN => n176_port);
   U55 : AOI222_X1 port map( A1 => OUTPUT1_13_port, A2 => n156, B1 => 
                           OUTPUT4_13_port, B2 => n147, C1 => OUTPUT2_13_port, 
                           C2 => n153, ZN => n93);
   U56 : INV_X1 port map( A => n92, ZN => n177_port);
   U57 : AOI222_X1 port map( A1 => OUTPUT1_12_port, A2 => n156, B1 => 
                           OUTPUT4_12_port, B2 => n146, C1 => OUTPUT2_12_port, 
                           C2 => n152, ZN => n92);
   U58 : INV_X1 port map( A => n91, ZN => n170);
   U59 : AOI222_X1 port map( A1 => OUTPUT1_11_port, A2 => n156, B1 => 
                           OUTPUT4_11_port, B2 => n146, C1 => OUTPUT2_11_port, 
                           C2 => n152, ZN => n91);
   U60 : INV_X1 port map( A => n90, ZN => n171);
   U61 : AOI222_X1 port map( A1 => OUTPUT1_10_port, A2 => n155, B1 => 
                           OUTPUT4_10_port, B2 => n146, C1 => OUTPUT2_10_port, 
                           C2 => n152, ZN => n90);
   U62 : INV_X1 port map( A => n89, ZN => n172);
   U63 : AOI222_X1 port map( A1 => OUTPUT1_9_port, A2 => n155, B1 => 
                           OUTPUT4_9_port, B2 => n146, C1 => OUTPUT2_9_port, C2
                           => n152, ZN => n89);
   U64 : INV_X1 port map( A => n88, ZN => n173);
   U65 : AOI222_X1 port map( A1 => OUTPUT1_8_port, A2 => n155, B1 => 
                           OUTPUT4_8_port, B2 => n146, C1 => OUTPUT2_8_port, C2
                           => n152, ZN => n88);
   U66 : INV_X1 port map( A => n86, ZN => n200_port);
   U67 : AOI222_X1 port map( A1 => OUTPUT1_7_port, A2 => n156, B1 => 
                           OUTPUT4_7_port, B2 => n146, C1 => OUTPUT2_7_port, C2
                           => n152, ZN => n86);
   U68 : INV_X1 port map( A => n85, ZN => n196_port);
   U69 : AOI222_X1 port map( A1 => OUTPUT1_6_port, A2 => n155, B1 => 
                           OUTPUT4_6_port, B2 => n146, C1 => OUTPUT2_6_port, C2
                           => n152, ZN => n85);
   U70 : INV_X1 port map( A => n84, ZN => n198_port);
   U71 : AOI222_X1 port map( A1 => OUTPUT1_5_port, A2 => n155, B1 => 
                           OUTPUT4_5_port, B2 => n146, C1 => OUTPUT2_5_port, C2
                           => n152, ZN => n84);
   U72 : INV_X1 port map( A => n83, ZN => n194_port);
   U73 : AOI222_X1 port map( A1 => OUTPUT1_4_port, A2 => n155, B1 => 
                           OUTPUT4_4_port, B2 => n146, C1 => OUTPUT2_4_port, C2
                           => n152, ZN => n83);
   U74 : OAI221_X1 port map( B1 => n241, B2 => n126, C1 => n118, C2 => n231, A 
                           => n128, ZN => n114);
   U75 : INV_X1 port map( A => n133, ZN => n231);
   U76 : NOR2_X1 port map( A1 => n129, A2 => n130, ZN => n128);
   U77 : AOI21_X1 port map( B1 => n242, B2 => n241, A => n122, ZN => n129);
   U78 : NOR2_X1 port map( A1 => n241, A2 => n242, ZN => n118);
   U79 : AOI221_X1 port map( B1 => n127, B2 => n237, C1 => n139_port, C2 => 
                           n242, A => n119, ZN => n135);
   U80 : INV_X1 port map( A => n121, ZN => n235);
   U81 : BUF_X1 port map( A => n232, Z => n149);
   U82 : BUF_X1 port map( A => n232, Z => n150);
   U83 : BUF_X1 port map( A => n232, Z => n151);
   U84 : BUF_X1 port map( A => N206, Z => n157);
   U85 : BUF_X1 port map( A => n230, Z => n148);
   U86 : BUF_X1 port map( A => n230, Z => n146);
   U87 : BUF_X1 port map( A => n230, Z => n147);
   U88 : BUF_X1 port map( A => N206, Z => n155);
   U89 : BUF_X1 port map( A => N206, Z => n156);
   U90 : OAI22_X1 port map( A1 => DATA2(0), A2 => n143, B1 => n149, B2 => n165,
                           ZN => N174);
   U91 : OAI22_X1 port map( A1 => DATA2(1), A2 => n143, B1 => n149, B2 => n166,
                           ZN => N175);
   U92 : OAI22_X1 port map( A1 => DATA2(2), A2 => n143, B1 => n149, B2 => n167,
                           ZN => N176);
   U93 : OAI22_X1 port map( A1 => DATA2(3), A2 => n143, B1 => n149, B2 => n168,
                           ZN => N177);
   U94 : OAI22_X1 port map( A1 => DATA2(4), A2 => n143, B1 => n149, B2 => n169,
                           ZN => N178);
   U95 : OAI22_X1 port map( A1 => DATA2(5), A2 => n143, B1 => n149, B2 => n227,
                           ZN => N179);
   U96 : INV_X1 port map( A => DATA2(5), ZN => n227);
   U97 : OAI22_X1 port map( A1 => DATA2(6), A2 => n143, B1 => n149, B2 => n226,
                           ZN => N180);
   U98 : INV_X1 port map( A => DATA2(6), ZN => n226);
   U99 : OAI22_X1 port map( A1 => DATA2(7), A2 => n143, B1 => n149, B2 => n225,
                           ZN => N181);
   U100 : INV_X1 port map( A => DATA2(7), ZN => n225);
   U101 : OAI22_X1 port map( A1 => DATA2(8), A2 => n143, B1 => n149, B2 => n224
                           , ZN => N182);
   U102 : INV_X1 port map( A => DATA2(8), ZN => n224);
   U103 : OAI22_X1 port map( A1 => DATA2(9), A2 => n143, B1 => n149, B2 => n223
                           , ZN => N183);
   U104 : INV_X1 port map( A => DATA2(9), ZN => n223);
   U105 : OAI22_X1 port map( A1 => DATA2(10), A2 => n143, B1 => n149, B2 => 
                           n222, ZN => N184);
   U106 : INV_X1 port map( A => DATA2(10), ZN => n222);
   U107 : OAI22_X1 port map( A1 => DATA2(11), A2 => n143, B1 => n150, B2 => 
                           n221, ZN => N185);
   U108 : INV_X1 port map( A => DATA2(11), ZN => n221);
   U109 : OAI22_X1 port map( A1 => DATA2(12), A2 => n144, B1 => n150, B2 => 
                           n220, ZN => N186);
   U110 : INV_X1 port map( A => DATA2(12), ZN => n220);
   U111 : OAI22_X1 port map( A1 => DATA2(13), A2 => n144, B1 => n150, B2 => 
                           n219, ZN => N187);
   U112 : INV_X1 port map( A => DATA2(13), ZN => n219);
   U113 : OAI22_X1 port map( A1 => DATA2(14), A2 => n144, B1 => n150, B2 => 
                           n218, ZN => N188);
   U114 : INV_X1 port map( A => DATA2(14), ZN => n218);
   U115 : OAI22_X1 port map( A1 => DATA2(15), A2 => n144, B1 => n150, B2 => 
                           n217, ZN => N189);
   U116 : INV_X1 port map( A => DATA2(15), ZN => n217);
   U117 : OAI22_X1 port map( A1 => DATA2(16), A2 => n144, B1 => n150, B2 => 
                           n216, ZN => N190);
   U118 : INV_X1 port map( A => DATA2(16), ZN => n216);
   U119 : OAI22_X1 port map( A1 => DATA2(17), A2 => n144, B1 => n150, B2 => 
                           n215, ZN => N191);
   U120 : INV_X1 port map( A => DATA2(17), ZN => n215);
   U121 : OAI22_X1 port map( A1 => DATA2(18), A2 => n144, B1 => n150, B2 => 
                           n214, ZN => N192);
   U122 : INV_X1 port map( A => DATA2(18), ZN => n214);
   U123 : OAI22_X1 port map( A1 => DATA2(19), A2 => n144, B1 => n150, B2 => 
                           n213, ZN => N193);
   U124 : INV_X1 port map( A => DATA2(19), ZN => n213);
   U125 : OAI22_X1 port map( A1 => DATA2(20), A2 => n144, B1 => n150, B2 => 
                           n212, ZN => N194);
   U126 : INV_X1 port map( A => DATA2(20), ZN => n212);
   U127 : OAI22_X1 port map( A1 => DATA2(21), A2 => n144, B1 => n150, B2 => 
                           n211, ZN => N195);
   U128 : INV_X1 port map( A => DATA2(21), ZN => n211);
   U129 : OAI22_X1 port map( A1 => DATA2(22), A2 => n144, B1 => n151, B2 => 
                           n210, ZN => N196);
   U130 : INV_X1 port map( A => DATA2(22), ZN => n210);
   U131 : OAI22_X1 port map( A1 => DATA2(23), A2 => n144, B1 => n151, B2 => 
                           n209, ZN => N197);
   U132 : INV_X1 port map( A => DATA2(23), ZN => n209);
   U133 : OAI22_X1 port map( A1 => DATA2(24), A2 => n145, B1 => n151, B2 => 
                           n208, ZN => N198);
   U134 : INV_X1 port map( A => DATA2(24), ZN => n208);
   U135 : OAI22_X1 port map( A1 => DATA2(25), A2 => n145, B1 => n151, B2 => 
                           n207, ZN => N199);
   U136 : INV_X1 port map( A => DATA2(25), ZN => n207);
   U137 : OAI22_X1 port map( A1 => DATA2(26), A2 => n145, B1 => n151, B2 => 
                           n206_port, ZN => N200);
   U138 : INV_X1 port map( A => DATA2(26), ZN => n206_port);
   U139 : OAI22_X1 port map( A1 => DATA2(27), A2 => n145, B1 => n151, B2 => 
                           n205_port, ZN => N201);
   U140 : INV_X1 port map( A => DATA2(27), ZN => n205_port);
   U141 : OAI22_X1 port map( A1 => DATA2(28), A2 => n145, B1 => n151, B2 => 
                           n204_port, ZN => N202);
   U142 : INV_X1 port map( A => DATA2(28), ZN => n204_port);
   U143 : OAI22_X1 port map( A1 => DATA2(29), A2 => n145, B1 => n151, B2 => 
                           n203_port, ZN => N203);
   U144 : INV_X1 port map( A => DATA2(29), ZN => n203_port);
   U145 : OAI22_X1 port map( A1 => DATA2(30), A2 => n145, B1 => n151, B2 => 
                           n202_port, ZN => N204);
   U146 : INV_X1 port map( A => DATA2(30), ZN => n202_port);
   U147 : OAI22_X1 port map( A1 => DATA2(31), A2 => n145, B1 => n151, B2 => 
                           n201_port, ZN => N205);
   U148 : INV_X1 port map( A => DATA2(31), ZN => n201_port);
   U149 : INV_X1 port map( A => n127, ZN => n236);
   U150 : INV_X1 port map( A => n114, ZN => n229);
   U151 : NAND2_X1 port map( A1 => n141_port, A2 => n239, ZN => n140);
   U152 : INV_X1 port map( A => n82, ZN => n199_port);
   U153 : AOI222_X1 port map( A1 => OUTPUT1_3_port, A2 => n155, B1 => 
                           OUTPUT4_3_port, B2 => n146, C1 => OUTPUT2_3_port, C2
                           => n152, ZN => n82);
   U154 : INV_X1 port map( A => n81, ZN => n195_port);
   U155 : AOI222_X1 port map( A1 => OUTPUT1_2_port, A2 => n155, B1 => 
                           OUTPUT4_2_port, B2 => n146, C1 => OUTPUT2_2_port, C2
                           => n152, ZN => n81);
   U156 : INV_X1 port map( A => n79, ZN => n197_port);
   U157 : AOI222_X1 port map( A1 => OUTPUT1_1_port, A2 => n155, B1 => 
                           OUTPUT4_1_port, B2 => n147, C1 => OUTPUT2_1_port, C2
                           => n153, ZN => n79);
   U158 : NOR4_X1 port map( A1 => n239, A2 => FUNC(2), A3 => FUNC(1), A4 => 
                           FUNC(0), ZN => n121);
   U159 : NOR4_X1 port map( A1 => n239, A2 => n238, A3 => FUNC(1), A4 => 
                           FUNC(0), ZN => n119);
   U160 : OAI21_X1 port map( B1 => n237, B2 => n241, A => FUNC(0), ZN => n132);
   U161 : NAND4_X1 port map( A1 => FUNC(2), A2 => n239, A3 => n237, A4 => n233,
                           ZN => n122);
   U162 : INV_X1 port map( A => FUNC(4), ZN => n241);
   U163 : NOR3_X1 port map( A1 => FUNC(2), A2 => FUNC(0), A3 => FUNC(3), ZN => 
                           n127);
   U164 : INV_X1 port map( A => FUNC(3), ZN => n239);
   U165 : NOR3_X1 port map( A1 => n237, A2 => FUNC(0), A3 => n238, ZN => 
                           n141_port);
   U166 : INV_X1 port map( A => FUNC(1), ZN => n237);
   U167 : OAI21_X1 port map( B1 => FUNC(3), B2 => n131, A => n138, ZN => n133);
   U168 : NAND4_X1 port map( A1 => FUNC(3), A2 => FUNC(1), A3 => n238, A4 => 
                           n233, ZN => n138);
   U169 : INV_X1 port map( A => FUNC(2), ZN => n238);
   U170 : OAI211_X1 port map( C1 => n241, C2 => n236, A => n123, B => n124, ZN 
                           => N206);
   U171 : OR3_X1 port map( A1 => n242, A2 => FUNC(4), A3 => n126, ZN => n123);
   U172 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => FUNC(3), A4 => n125,
                           ZN => n124);
   U173 : NOR2_X1 port map( A1 => n240, A2 => n233, ZN => n125);
   U174 : INV_X1 port map( A => FUNC(0), ZN => n233);
   U175 : NAND2_X1 port map( A1 => n141_port, A2 => FUNC(3), ZN => n126);
   U176 : INV_X1 port map( A => FUNC(5), ZN => n242);
   U182 : OAI211_X1 port map( C1 => n119, C2 => n234, A => n242, B => FUNC(4), 
                           ZN => n113);
   U183 : NOR3_X1 port map( A1 => n241, A2 => FUNC(5), A3 => n236, ZN => 
                           n142_port);
   U184 : OAI211_X1 port map( C1 => n234, C2 => n121, A => n241, B => FUNC(5), 
                           ZN => n112);
   U185 : INV_X1 port map( A => n117, ZN => n230);
   U186 : AOI222_X1 port map( A1 => n118, A2 => n119, B1 => n241, B2 => n120, 
                           C1 => FUNC(4), C2 => n121, ZN => n117);
   U187 : OAI22_X1 port map( A1 => n236, A2 => n237, B1 => n122, B2 => FUNC(5),
                           ZN => n120);
   U188 : INV_X1 port map( A => n134, ZN => n232);
   U189 : OAI211_X1 port map( C1 => FUNC(4), C2 => n135, A => n136, B => n137, 
                           ZN => n134);
   U190 : OR3_X1 port map( A1 => n239, A2 => n118, A3 => n131, ZN => n137);
   U191 : OAI21_X1 port map( B1 => n234, B2 => n133, A => n118, ZN => n136);
   U192 : INV_X1 port map( A => DATA2(2), ZN => n167);
   U193 : INV_X1 port map( A => DATA2(1), ZN => n166);
   U194 : NAND2_X1 port map( A1 => n115, A2 => n116, ZN => N142);
   U195 : AOI22_X1 port map( A1 => OUTPUT2_0_port, A2 => n152, B1 => 
                           OUTPUT1_0_port, B2 => n155, ZN => n115);
   U196 : AOI22_X1 port map( A1 => OUTPUT4_0_port, A2 => n146, B1 => 
                           OUTPUT3_0_port, B2 => n114, ZN => n116);
   U197 : CLKBUF_X1 port map( A => N141, Z => n158);
   U198 : CLKBUF_X1 port map( A => N141, Z => n159);
   U199 : CLKBUF_X1 port map( A => N141, Z => n160);
   U200 : CLKBUF_X1 port map( A => N141, Z => n161);
   U201 : INV_X1 port map( A => DATA2(0), ZN => n165);
   U202 : INV_X1 port map( A => DATA2(3), ZN => n168);
   U203 : INV_X1 port map( A => DATA2(4), ZN => n169);

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_5;

architecture SYN_struct of MUX21_GENERIC_NBIT32_5 is

   component MUX21_161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_192 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_191 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_190 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_189 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_188 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_187 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_186 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_185 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_184 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_183 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_182 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_181 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_180 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_179 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_178 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_177 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_176 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_175 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_174 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_173 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_172 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_171 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_170 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_169 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_168 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_167 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_166 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_165 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_164 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_163 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_162 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_161 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_6;

architecture SYN_struct of MUX21_GENERIC_NBIT32_6 is

   component MUX21_193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_218
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_219
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_220
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_221
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_222
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_223
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_224
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_224 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_223 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_222 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_221 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_220 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_219 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_218 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_217 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_216 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_215 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_214 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_213 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_212 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_211 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_210 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_209 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_208 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_207 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_206 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_205 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_204 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_203 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_202 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_201 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_200 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_199 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_198 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_197 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_196 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_195 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_194 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_193 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT6_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 downto 
         0);  Q : out std_logic_vector (5 downto 0));

end regFFD_NBIT6_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT6_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   Q_reg_5_inst : DFFR_X1 port map( D => n1, CK => CK, RN => RESET, Q => Q(5), 
                           QN => n13);
   Q_reg_4_inst : DFFR_X1 port map( D => n2, CK => CK, RN => RESET, Q => Q(4), 
                           QN => n14);
   Q_reg_3_inst : DFFR_X1 port map( D => n3, CK => CK, RN => RESET, Q => Q(3), 
                           QN => n15);
   Q_reg_2_inst : DFFR_X1 port map( D => n4, CK => CK, RN => RESET, Q => Q(2), 
                           QN => n16);
   Q_reg_1_inst : DFFR_X1 port map( D => n5, CK => CK, RN => RESET, Q => Q(1), 
                           QN => n17);
   Q_reg_0_inst : DFFR_X1 port map( D => n6, CK => CK, RN => RESET, Q => Q(0), 
                           QN => n18);
   U2 : OAI21_X1 port map( B1 => n13, B2 => ENABLE, A => n12, ZN => n1);
   U3 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n12);
   U4 : OAI21_X1 port map( B1 => n16, B2 => ENABLE, A => n9, ZN => n4);
   U5 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n9);
   U6 : OAI21_X1 port map( B1 => n14, B2 => ENABLE, A => n11, ZN => n2);
   U7 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n11);
   U8 : OAI21_X1 port map( B1 => n15, B2 => ENABLE, A => n10, ZN => n3);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n10);
   U10 : OAI21_X1 port map( B1 => n17, B2 => ENABLE, A => n8, ZN => n5);
   U11 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n8);
   U12 : OAI21_X1 port map( B1 => n18, B2 => ENABLE, A => n7, ZN => n6);
   U13 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n7);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15 : 
      std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n1, CK => CK, RN => RESET, Q => Q(4), 
                           QN => n11);
   Q_reg_3_inst : DFFR_X1 port map( D => n2, CK => CK, RN => RESET, Q => Q(3), 
                           QN => n12);
   Q_reg_2_inst : DFFR_X1 port map( D => n3, CK => CK, RN => RESET, Q => Q(2), 
                           QN => n13);
   Q_reg_1_inst : DFFR_X1 port map( D => n4, CK => CK, RN => RESET, Q => Q(1), 
                           QN => n14);
   Q_reg_0_inst : DFFR_X1 port map( D => n5, CK => CK, RN => RESET, Q => Q(0), 
                           QN => n15);
   U2 : OAI21_X1 port map( B1 => n14, B2 => ENABLE, A => n7, ZN => n4);
   U3 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n7);
   U4 : OAI21_X1 port map( B1 => n13, B2 => ENABLE, A => n8, ZN => n3);
   U5 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n8);
   U6 : OAI21_X1 port map( B1 => n12, B2 => ENABLE, A => n9, ZN => n2);
   U7 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n9);
   U8 : OAI21_X1 port map( B1 => n11, B2 => ENABLE, A => n10, ZN => n1);
   U9 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n10);
   U10 : OAI21_X1 port map( B1 => n15, B2 => ENABLE, A => n6, ZN => n5);
   U11 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n6);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_8 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_8;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n65);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n66);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n67);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n68);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n69);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n70);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n71);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n98, Q => Q(24), 
                           QN => n72);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n73);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n98, Q => Q(22),
                           QN => n74);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n75);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n76);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n97, Q => Q(19),
                           QN => n77);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n78);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n97, Q => Q(17),
                           QN => n79);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n80);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n81);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n82);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n83);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n84);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n85);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n86);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n87);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n88);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n89);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n90);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n91);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n92);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n93);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n94);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n95);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n96);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n96, B2 => ENABLE, A => n39, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n39);
   U7 : OAI21_X1 port map( B1 => n95, B2 => ENABLE, A => n40, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n40);
   U9 : OAI21_X1 port map( B1 => n94, B2 => ENABLE, A => n41, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n41);
   U11 : OAI21_X1 port map( B1 => n93, B2 => ENABLE, A => n43, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n43);
   U13 : OAI21_X1 port map( B1 => n92, B2 => ENABLE, A => n44, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n44);
   U15 : OAI21_X1 port map( B1 => n91, B2 => ENABLE, A => n45, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n45);
   U17 : OAI21_X1 port map( B1 => n90, B2 => ENABLE, A => n46, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n46);
   U19 : OAI21_X1 port map( B1 => n89, B2 => ENABLE, A => n47, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n47);
   U21 : OAI21_X1 port map( B1 => n88, B2 => ENABLE, A => n48, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n48);
   U23 : OAI21_X1 port map( B1 => n87, B2 => ENABLE, A => n49, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n49);
   U25 : OAI21_X1 port map( B1 => n86, B2 => ENABLE, A => n50, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n50);
   U27 : OAI21_X1 port map( B1 => n85, B2 => ENABLE, A => n51, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n51);
   U29 : OAI21_X1 port map( B1 => n84, B2 => ENABLE, A => n52, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n52);
   U31 : OAI21_X1 port map( B1 => n83, B2 => ENABLE, A => n54, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n54);
   U33 : OAI21_X1 port map( B1 => n82, B2 => ENABLE, A => n55, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n55);
   U35 : OAI21_X1 port map( B1 => n81, B2 => ENABLE, A => n56, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n56);
   U37 : OAI21_X1 port map( B1 => n80, B2 => ENABLE, A => n57, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n57);
   U39 : OAI21_X1 port map( B1 => n79, B2 => ENABLE, A => n58, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n58);
   U41 : OAI21_X1 port map( B1 => n78, B2 => ENABLE, A => n59, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n59);
   U43 : OAI21_X1 port map( B1 => n77, B2 => ENABLE, A => n60, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n60);
   U45 : OAI21_X1 port map( B1 => n76, B2 => ENABLE, A => n61, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n61);
   U47 : OAI21_X1 port map( B1 => n75, B2 => ENABLE, A => n62, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n62);
   U49 : OAI21_X1 port map( B1 => n74, B2 => ENABLE, A => n63, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n63);
   U51 : OAI21_X1 port map( B1 => n73, B2 => ENABLE, A => n33, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n33);
   U53 : OAI21_X1 port map( B1 => n72, B2 => ENABLE, A => n34, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n34);
   U55 : OAI21_X1 port map( B1 => n71, B2 => ENABLE, A => n35, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n35);
   U57 : OAI21_X1 port map( B1 => n70, B2 => ENABLE, A => n36, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n36);
   U59 : OAI21_X1 port map( B1 => n69, B2 => ENABLE, A => n37, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n37);
   U61 : OAI21_X1 port map( B1 => n68, B2 => ENABLE, A => n38, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n38);
   U63 : OAI21_X1 port map( B1 => n67, B2 => ENABLE, A => n42, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n42);
   U65 : OAI21_X1 port map( B1 => n66, B2 => ENABLE, A => n53, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n53);
   U67 : OAI21_X1 port map( B1 => n65, B2 => ENABLE, A => n64, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n64);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_9 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_9;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n99, Q => Q(31), 
                           QN => n65);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n66);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n67);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n99, Q => Q(28), 
                           QN => n68);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n69);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n70);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n71);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n72);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n99, Q => Q(23), 
                           QN => n73);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n74);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n98, Q => Q(21),
                           QN => n75);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n97, Q => Q(20),
                           QN => n76);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n99, Q => Q(19),
                           QN => n77);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n78);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n79);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n80);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n99, Q => Q(15),
                           QN => n81);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n82);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n83);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n84);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n97, Q => Q(11),
                           QN => n85);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n97, Q => Q(10),
                           QN => n86);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n87);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n97, Q => Q(8), 
                           QN => n88);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n89);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n90);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n98, Q => Q(5), 
                           QN => n91);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n98, Q => Q(4), 
                           QN => n92);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n93);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n98, Q => Q(2), 
                           QN => n94);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n98, Q => Q(1), 
                           QN => n95);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n96);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n96, B2 => ENABLE, A => n39, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n39);
   U7 : OAI21_X1 port map( B1 => n95, B2 => ENABLE, A => n40, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n40);
   U9 : OAI21_X1 port map( B1 => n94, B2 => ENABLE, A => n41, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n41);
   U11 : OAI21_X1 port map( B1 => n93, B2 => ENABLE, A => n43, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n43);
   U13 : OAI21_X1 port map( B1 => n92, B2 => ENABLE, A => n44, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n44);
   U15 : OAI21_X1 port map( B1 => n91, B2 => ENABLE, A => n45, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n45);
   U17 : OAI21_X1 port map( B1 => n90, B2 => ENABLE, A => n46, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n46);
   U19 : OAI21_X1 port map( B1 => n89, B2 => ENABLE, A => n47, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n47);
   U21 : OAI21_X1 port map( B1 => n88, B2 => ENABLE, A => n48, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n48);
   U23 : OAI21_X1 port map( B1 => n87, B2 => ENABLE, A => n49, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n49);
   U25 : OAI21_X1 port map( B1 => n86, B2 => ENABLE, A => n50, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n50);
   U27 : OAI21_X1 port map( B1 => n85, B2 => ENABLE, A => n51, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n51);
   U29 : OAI21_X1 port map( B1 => n84, B2 => ENABLE, A => n52, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n52);
   U31 : OAI21_X1 port map( B1 => n83, B2 => ENABLE, A => n54, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n54);
   U33 : OAI21_X1 port map( B1 => n82, B2 => ENABLE, A => n55, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n55);
   U35 : OAI21_X1 port map( B1 => n81, B2 => ENABLE, A => n56, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n56);
   U37 : OAI21_X1 port map( B1 => n80, B2 => ENABLE, A => n57, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n57);
   U39 : OAI21_X1 port map( B1 => n79, B2 => ENABLE, A => n58, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n58);
   U41 : OAI21_X1 port map( B1 => n78, B2 => ENABLE, A => n59, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n59);
   U43 : OAI21_X1 port map( B1 => n77, B2 => ENABLE, A => n60, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n60);
   U45 : OAI21_X1 port map( B1 => n76, B2 => ENABLE, A => n61, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n61);
   U47 : OAI21_X1 port map( B1 => n75, B2 => ENABLE, A => n62, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n62);
   U49 : OAI21_X1 port map( B1 => n74, B2 => ENABLE, A => n63, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n63);
   U51 : OAI21_X1 port map( B1 => n73, B2 => ENABLE, A => n33, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n33);
   U53 : OAI21_X1 port map( B1 => n72, B2 => ENABLE, A => n34, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n34);
   U55 : OAI21_X1 port map( B1 => n71, B2 => ENABLE, A => n35, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n35);
   U57 : OAI21_X1 port map( B1 => n70, B2 => ENABLE, A => n36, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n36);
   U59 : OAI21_X1 port map( B1 => n69, B2 => ENABLE, A => n37, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n37);
   U61 : OAI21_X1 port map( B1 => n68, B2 => ENABLE, A => n38, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n38);
   U63 : OAI21_X1 port map( B1 => n67, B2 => ENABLE, A => n42, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n42);
   U65 : OAI21_X1 port map( B1 => n66, B2 => ENABLE, A => n53, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n53);
   U67 : OAI21_X1 port map( B1 => n65, B2 => ENABLE, A => n64, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n64);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_10 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_10;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n99, Q => Q(31), 
                           QN => n65);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n99, Q => Q(30), 
                           QN => n66);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n99, Q => Q(29), 
                           QN => n67);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n99, Q => Q(28), 
                           QN => n68);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n98, Q => Q(27), 
                           QN => n69);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n98, Q => Q(26), 
                           QN => n70);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n98, Q => Q(25), 
                           QN => n71);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n98, Q => Q(24), 
                           QN => n72);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n99, Q => Q(23), 
                           QN => n73);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n98, Q => Q(22),
                           QN => n74);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n98, Q => Q(21),
                           QN => n75);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n97, Q => Q(20),
                           QN => n76);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n99, Q => Q(19),
                           QN => n77);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n97, Q => Q(18),
                           QN => n78);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n97, Q => Q(17),
                           QN => n79);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n97, Q => Q(16),
                           QN => n80);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n99, Q => Q(15),
                           QN => n81);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n97, Q => Q(14),
                           QN => n82);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n97, Q => Q(13),
                           QN => n83);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n97, Q => Q(12),
                           QN => n84);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n85);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n86);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n98, Q => Q(9), 
                           QN => n87);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n98, Q => Q(8), 
                           QN => n88);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n89);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n90);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n97, Q => Q(5), 
                           QN => n91);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n97, Q => Q(4), 
                           QN => n92);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n98, Q => Q(3), 
                           QN => n93);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n97, Q => Q(2), 
                           QN => n94);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n97, Q => Q(1), 
                           QN => n95);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n96);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n96, B2 => ENABLE, A => n39, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n39);
   U7 : OAI21_X1 port map( B1 => n95, B2 => ENABLE, A => n40, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n40);
   U9 : OAI21_X1 port map( B1 => n94, B2 => ENABLE, A => n41, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n41);
   U11 : OAI21_X1 port map( B1 => n93, B2 => ENABLE, A => n43, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n43);
   U13 : OAI21_X1 port map( B1 => n92, B2 => ENABLE, A => n44, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n44);
   U15 : OAI21_X1 port map( B1 => n91, B2 => ENABLE, A => n45, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n45);
   U17 : OAI21_X1 port map( B1 => n90, B2 => ENABLE, A => n46, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n46);
   U19 : OAI21_X1 port map( B1 => n89, B2 => ENABLE, A => n47, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n47);
   U21 : OAI21_X1 port map( B1 => n88, B2 => ENABLE, A => n48, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n48);
   U23 : OAI21_X1 port map( B1 => n87, B2 => ENABLE, A => n49, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n49);
   U25 : OAI21_X1 port map( B1 => n86, B2 => ENABLE, A => n50, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n50);
   U27 : OAI21_X1 port map( B1 => n85, B2 => ENABLE, A => n51, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n51);
   U29 : OAI21_X1 port map( B1 => n84, B2 => ENABLE, A => n52, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n52);
   U31 : OAI21_X1 port map( B1 => n83, B2 => ENABLE, A => n54, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n54);
   U33 : OAI21_X1 port map( B1 => n82, B2 => ENABLE, A => n55, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n55);
   U35 : OAI21_X1 port map( B1 => n81, B2 => ENABLE, A => n56, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n56);
   U37 : OAI21_X1 port map( B1 => n80, B2 => ENABLE, A => n57, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n57);
   U39 : OAI21_X1 port map( B1 => n79, B2 => ENABLE, A => n58, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n58);
   U41 : OAI21_X1 port map( B1 => n78, B2 => ENABLE, A => n59, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n59);
   U43 : OAI21_X1 port map( B1 => n77, B2 => ENABLE, A => n60, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n60);
   U45 : OAI21_X1 port map( B1 => n76, B2 => ENABLE, A => n61, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n61);
   U47 : OAI21_X1 port map( B1 => n75, B2 => ENABLE, A => n62, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n62);
   U49 : OAI21_X1 port map( B1 => n74, B2 => ENABLE, A => n63, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n63);
   U51 : OAI21_X1 port map( B1 => n73, B2 => ENABLE, A => n33, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n33);
   U53 : OAI21_X1 port map( B1 => n72, B2 => ENABLE, A => n34, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n34);
   U55 : OAI21_X1 port map( B1 => n71, B2 => ENABLE, A => n35, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n35);
   U57 : OAI21_X1 port map( B1 => n70, B2 => ENABLE, A => n36, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n36);
   U59 : OAI21_X1 port map( B1 => n69, B2 => ENABLE, A => n37, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n37);
   U61 : OAI21_X1 port map( B1 => n68, B2 => ENABLE, A => n38, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n38);
   U63 : OAI21_X1 port map( B1 => n67, B2 => ENABLE, A => n42, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n42);
   U65 : OAI21_X1 port map( B1 => n66, B2 => ENABLE, A => n53, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n53);
   U67 : OAI21_X1 port map( B1 => n65, B2 => ENABLE, A => n64, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n64);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_0 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_0;

architecture SYN_SYNC_BHV of FF_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n2, n4, n3, n5, n_1140 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n2, CK => CLK, Q => Q_port, QN => n_1140);
   U3 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => n2);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => n5, B2 => Q_port, ZN => n4)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n5);
   U6 : INV_X1 port map( A => RESET, ZN => n3);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity windRF_M8_N8_F5_NBIT32 is

   port( CLK, RESET, ENABLE, CALL, RETRN : in std_logic;  FILL, SPILL : out 
         std_logic;  BUSin : in std_logic_vector (31 downto 0);  BUSout : out 
         std_logic_vector (31 downto 0);  RD1, RD2, WR : in std_logic;  ADD_WR,
         ADD_RD1, ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0);  wr_signal : in std_logic);

end windRF_M8_N8_F5_NBIT32;

architecture SYN_bhv of windRF_M8_N8_F5_NBIT32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N2170, N2171, N2172, N2173, N8434, N8435, N8436, N8437, N8578, N8579,
      N8580, N8581, N8702, N8703, N8704, N8705, N8706, N8707, N8708, N8709, 
      N8710, N8711, N8712, N8713, N8714, N8715, N8716, N8717, N8718, N8719, 
      N8720, N8721, N8722, N8723, N8724, N8725, N8726, N8727, N8728, N8729, 
      N8730, N8731, N8732, N8733, N8734, N8735, N8736, N8737, N8738, N8739, 
      N8740, N8741, N8742, N8743, N8744, N8745, N8746, N8747, N8748, N8749, 
      N8750, N8751, N8752, N8753, N8754, N8755, N8756, N8757, N8758, N8759, 
      N8760, N8761, N8762, N8763, N8764, N8765, N8766, N8767, U3_U97_Z_4, 
      U3_U97_Z_5, U3_U97_Z_6, U3_U98_Z_4, U3_U98_Z_5, U3_U98_Z_6, U3_U99_Z_4, 
      U3_U99_Z_5, U3_U99_Z_6, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
      n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, 
      n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
      n730, n731, n732, n733, n734, n735, n736, n737, n770, n771, n772, n773, 
      n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, 
      n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, 
      n798, n799, n800, n801, n2754, n2755, n2756, n2757, n2758, n2759, n2760, 
      n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, 
      n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, 
      n2781, n2782, n2783, n2784, n2785, n2818, n2819, n2820, n2821, n2822, 
      n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
      n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, 
      n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2882, n2883, n2884, 
      n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, 
      n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, 
      n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2935, 
      n2936, n2937, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
      n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, 
      n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, 
      n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
      n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, 
      n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, 
      n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, 
      n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, 
      n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, 
      n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, 
      n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, 
      n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, 
      n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
      n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, 
      n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, 
      n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
      n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, 
      n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, 
      n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, 
      n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
      n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, 
      n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, 
      n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, 
      n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
      n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, 
      n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
      n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, 
      n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, 
      n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, 
      n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, 
      n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, 
      n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, 
      n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, 
      n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, 
      n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, 
      n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, 
      n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, 
      n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, 
      n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, 
      n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, 
      n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
      n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, 
      n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, 
      n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, 
      n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, 
      n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, 
      n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, 
      n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, 
      n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, 
      n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, 
      n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, 
      n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, 
      n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, 
      n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, 
      n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
      n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
      n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
      n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, 
      n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, 
      n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, 
      n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, 
      n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, 
      n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, 
      n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, 
      n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, 
      n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, 
      n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, 
      n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, 
      n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
      n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, 
      n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, 
      n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, 
      n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, 
      n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, 
      n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, 
      n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, 
      n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, 
      n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, 
      n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, 
      n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, 
      n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, 
      n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, 
      n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
      n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, 
      n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, 
      n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, 
      n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
      n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, 
      n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
      n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, 
      n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, 
      n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, 
      n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, 
      n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, 
      n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, 
      n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, 
      n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, 
      n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, 
      n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
      n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434_port, n8435_port, n8436_port, n8437_port, n8438, n8439, n8440, 
      n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, 
      n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, 
      n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, 
      n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, 
      n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, 
      n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, 
      n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, 
      n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, 
      n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, 
      n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, 
      n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, 
      n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, 
      n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, 
      n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578_port, n8579_port, 
      n8580_port, n8581_port, n8582, n8583, n8584, n8585, n8586, n8587, n8588, 
      n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, 
      n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, 
      n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, 
      n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, 
      n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, 
      n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, 
      n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, 
      n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, 
      n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, 
      n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, 
      n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, 
      n8699, n8700, n8701, n8702_port, n8703_port, n8704_port, n8705_port, 
      n8706_port, n8707_port, n8708_port, n8709_port, n8710_port, n8711_port, 
      n8712_port, n8713_port, n8714_port, n8715_port, n8716_port, n8717_port, 
      n8718_port, n8719_port, n8720_port, n8721_port, n8722_port, n8723_port, 
      n8724_port, n8725_port, n8726_port, n8727_port, n8728_port, n8729_port, 
      n8730_port, n8731_port, n8732_port, n8733_port, n8734_port, n8735_port, 
      n8736_port, n8737_port, n8738_port, n8739_port, n8740_port, n8741_port, 
      n8742_port, n8743_port, n8744_port, n8745_port, n8746_port, n8747_port, 
      n8748_port, n8749_port, n8750_port, n8751_port, n8752_port, n8753_port, 
      n8754_port, n8755_port, n8756_port, n8757_port, n8758_port, n8759_port, 
      n8760_port, n8761_port, n8762_port, n8763_port, n8764_port, n8765_port, 
      n8766_port, n8767_port, n8768, n8769, n8770, n8771, n8772, n8773, n8774, 
      n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, 
      n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, 
      n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, 
      n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, 
      n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, 
      n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, 
      n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, 
      n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, 
      n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, 
      n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, 
      n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, 
      n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, 
      n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, 
      n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, 
      n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, 
      n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, 
      n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, 
      n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, 
      n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, 
      n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, 
      n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, 
      n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, 
      n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, 
      n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, 
      n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, 
      n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, 
      n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, 
      n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, 
      n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, 
      n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, 
      n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, 
      n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, 
      n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, 
      n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, 
      n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, 
      n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n141, n142
      , n143, n153, n154, n155, n165, n166, n167, n177, n178, n179, n189, n190,
      n191, n201, n202, n203, n213, n214, n215, n225, n226, n227, n237, n238, 
      n239, n249, n250, n251, n261, n262, n263, n273, n274, n275, n285, n286, 
      n287, n297, n298, n299, n309, n310, n311, n321, n322, n323, n333, n334, 
      n335, n345, n346, n347, n357, n358, n359, n369, n370, n371, n381, n382, 
      n383, n393, n394, n395, n405, n406, n407, n417, n418, n419, n429, n430, 
      n431, n441, n442, n443, n453, n454, n455, n465, n466, n467, n477, n478, 
      n479, n489, n490, n491, n501, n502, n503, n513, n514, n515, n868, n871, 
      n872, n875, n876, n879, n880, n883, n884, n887, n888, n891, n892, n895, 
      n896, n899, n900, n903, n904, n907, n908, n911, n912, n915, n916, n919, 
      n920, n923, n924, n927, n928, n929, n931, n932, n933, n935, n936, n937, 
      n939, n940, n941, n943, n944, n945, n947, n948, n949, n951, n952, n953, 
      n955, n956, n957, n959, n960, n961, n963, n964, n965, n967, n968, n969, 
      n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, 
      n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, 
      n995, n996, n997, n998, n999, n1029, n1041, n1042, n1043, n1053, n1054, 
      n1055, n1065, n1066, n1067, n1077, n1078, n1079, n1089, n1090, n1091, 
      n1101, n1102, n1103, n1113, n1114, n1115, n1125, n1126, n1127, n1137, 
      n1138, n1139, n1149, n1150, n1151, n1161, n1162, n1163, n1173, n1174, 
      n1175, n1185, n1186, n1187, n1197, n1198, n1199, n1209, n1210, n1211, 
      n1221, n1222, n1223, n1233, n1234, n1235, n1245, n1246, n1247, n1257, 
      n1258, n1259, n1269, n1270, n1271, n1281, n1282, n1283, n1293, n1294, 
      n1295, n1305, n1306, n1307, n1317, n1318, n1319, n1329, n1330, n1331, 
      n1341, n1342, n1343, n1385, n1386, n1387, n1397, n1398, n1399, n1409, 
      n1442, n1443, n1735, n1739, n1743, n1747, n1751, n1755, n1759, n1763, 
      n1767, n1771, n1775, n1779, n1783, n1787, n1791, n1795, n1799, n1803, 
      n1807, n1811, n1815, n1819, n1823, n1827, n1831, n1835, n1839, n1843, 
      n1847, n1851, n1855, n1859, n1868, n1869, n1870, n1871, n1880, n1881, 
      n1882, n1883, n1892, n1893, n1894, n1895, n1904, n1905, n1906, n1907, 
      n1916, n1917, n1918, n1919, n1928, n1929, n1930, n1931, n1940, n1941, 
      n1942, n1943, n1952, n1953, n1954, n1955, n1964, n1965, n1966, n1967, 
      n1976, n1977, n1978, n1979, n1988, n1989, n1990, n1991, n2000, n2001, 
      n2002, n2003, n2012, n2013, n2014, n2015, n2024, n2025, n2026, n2027, 
      n2036, n2037, n2038, n2039, n2048, n2049, n2082, n2083, n2093, n2094, 
      n2095, n2105, n2106, n2107, n2149, n2150, n2151, n2161, n2162, n2163, 
      n2173_port, n2174, n2175, n2217, n2218, n2219, n2229, n2230, n2231, n2241
      , n2242, n2243, n2253, n2254, n2255, n2265, n2266, n2267, n2277, n2278, 
      n2279, n2289, n2290, n2291, n2301, n2302, n2303, n2313, n2314, n2315, 
      n2325, n2326, n2327, n2337, n2338, n2339, n9216, n9217, n9218, n9219, 
      n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, 
      n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, 
      n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9265, n9266, 
      n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, 
      n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, 
      n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, 
      n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, 
      n9307, n9308, n9309, n9310, n9312, n9313, n9314, n9315, n9316, n9317, 
      n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, 
      n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, 
      n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, 
      n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, 
      n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, 
      n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, 
      n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, 
      n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, 
      n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, 
      n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, 
      n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, 
      n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, 
      n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, 
      n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, 
      n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, 
      n9564, n9565, n9566, n9567, n9664, n9665, n9666, n9667, n9668, n9669, 
      n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, 
      n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, 
      n9690, n9691, n9692, n9693, n9694, n9695, n9702, n9703, n9704, n9705, 
      n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, 
      n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, 
      n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, 
      n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, 
      n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, 
      n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, 
      n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, 
      n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, 
      n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, 
      n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, 
      n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, 
      n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, 
      n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, 
      n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, 
      n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, 
      n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, 
      n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, 
      n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, 
      n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, 
      n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n2477, n2478, 
      n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, 
      n2489, n2490, n2491, n2492, n2494, n2496, n2498, n2500, n2566, n2568, 
      n2570, n2571, n2573, n2574, n2576, n2578, n2580, n2582, n2584, n2586, 
      n2588, n2597, n2599, n2615, n2617, n2698, n2715, n2716, n2717, n2719, 
      n2721, n2723, n2725, n2730, n2735, n2739, n2740, n2741, n2742, n2743, 
      n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
      n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, 
      n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, 
      n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
      n2816, n2817, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, 
      n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, 
      n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, 
      n2878, n2879, n2880, n2881, n2914, n2915, n2916, n2917, n2918, n2919, 
      n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
      n2930, n2931, n2932, n2933, n2934, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, 
      n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, 
      n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
      n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, 
      n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
      n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, 
      n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
      n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, 
      n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
      n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
      n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
      n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, 
      n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
      n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, 
      n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
      n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, 
      n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
      n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, 
      n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, 
      n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
      n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, 
      n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
      n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, 
      n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
      n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, 
      n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
      n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, 
      n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
      n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, 
      n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
      n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, 
      n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
      n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, 
      n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
      n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, 
      n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, 
      n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
      n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, 
      n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, 
      n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, 
      n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
      n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, 
      n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, 
      n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, 
      n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
      n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, 
      n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, 
      n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, 
      n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
      n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
      n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
      n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, 
      n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
      n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
      n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, 
      n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, 
      n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
      n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
      n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, 
      n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, 
      n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, 
      n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
      n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, 
      n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, 
      n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, 
      n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
      n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, 
      n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, 
      n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, 
      n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, 
      n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, 
      n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, 
      n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, 
      n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, 
      n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, 
      n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, 
      n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, 
      n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, 
      n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, 
      n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, 
      n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, 
      n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, 
      n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
      n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, 
      n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, 
      n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, 
      n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, 
      n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, 
      n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, 
      n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, 
      n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, 
      n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, 
      n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, 
      n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, 
      n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, 
      n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, 
      n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, 
      n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, 
      n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, 
      n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, 
      n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, 
      n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, 
      n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, 
      n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, 
      n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
      n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, 
      n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, 
      n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, 
      n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, 
      n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, 
      n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, 
      n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, 
      n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, 
      n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, 
      n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, 
      n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, 
      n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, 
      n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, 
      n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, 
      n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, 
      n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, 
      n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, 
      n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, 
      n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, 
      n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, 
      n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, 
      n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, 
      n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, 
      n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, 
      n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, 
      n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, 
      n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, 
      n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, 
      n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, 
      n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, 
      n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, 
      n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, 
      n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, 
      n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, 
      n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, 
      n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, 
      n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, 
      n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, 
      n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, 
      n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, 
      n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, 
      n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, 
      n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, 
      n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, 
      n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, 
      n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, 
      n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, 
      n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, 
      n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, 
      n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, 
      n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, 
      n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, 
      n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, 
      n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, 
      n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, 
      n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, 
      n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, 
      n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, 
      n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, 
      n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, 
      n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, 
      n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, 
      n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, 
      n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, 
      n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, 
      n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, 
      n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, 
      n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, 
      n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, 
      n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, 
      n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, 
      n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, 
      n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
      n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, 
      n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
      n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, 
      n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, 
      n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, 
      n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, 
      n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, 
      n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, 
      n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, 
      n5943, n5944, n5945, n5946, n5947, n5948, n5981, n5982, n5983, n5984, 
      n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, 
      n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, 
      n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6044, n6140, 
      n6236, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, 
      n6310, n6311, n6312, n6313, n6314, n6315, n9134, n9135, n9136, n9137, 
      n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, 
      n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, 
      n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, 
      n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, 
      n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, 
      n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, 
      n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, 
      n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9248, n9249, 
      n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, 
      n9260, n9261, n9262, n9263, n9264, n9311, n9568, n9569, n9570, n9571, 
      n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, 
      n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, 
      n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, 
      n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, 
      n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, 
      n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, 
      n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, 
      n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, 
      n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, 
      n9662, n9663, n9696, n9697, n9698, n9699, n9700, n9701, n10000, n10001, 
      n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, 
      n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, 
      n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, 
      n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, 
      n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, 
      n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, 
      n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, 
      n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, 
      n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, 
      n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, 
      n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, 
      n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, 
      n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, 
      n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, 
      n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, 
      n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, 
      n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, 
      n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, 
      n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, 
      n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, 
      n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, 
      n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, 
      n10200, n10201, n10202, n10203, n10204, n10205, n10208, n10209, n10210, 
      n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, 
      n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, 
      n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, 
      n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, 
      n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, 
      n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, 
      n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, 
      n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, 
      n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, 
      n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, 
      n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, 
      n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, 
      n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, 
      n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, 
      n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, 
      n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, 
      n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, 
      n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, 
      n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, 
      n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, 
      n10394, n10395, n10396, n10400, n10401, n10402, n10403, n10404, n10405, 
      n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, 
      n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, 
      n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, 
      n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, 
      n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, 
      n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, 
      n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, 
      n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, 
      n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, 
      n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, 
      n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, 
      n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, 
      n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, 
      n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, 
      n10532, n10533, n10534, n10535, n10536, n10537, r486_n4, 
      r486_carry_4_port, r486_carry_5_port, r486_A_3_port, r480_n4, 
      r480_carry_4_port, r480_carry_5_port, r480_A_3_port, r472_n4, 
      r472_carry_4_port, r472_carry_5_port, r472_B_3_port, n10538, n10539, 
      n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, 
      n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, 
      n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, 
      n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, 
      n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, 
      n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, 
      n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, 
      n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, 
      n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, 
      n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, 
      n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, 
      n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, 
      n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, 
      n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, 
      n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, 
      n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, 
      n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, 
      n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, 
      n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, 
      n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, 
      n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, 
      n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, 
      n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, 
      n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, 
      n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, 
      n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, 
      n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, 
      n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, 
      n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, 
      n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, 
      n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, 
      n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, 
      n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, 
      n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, 
      n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, 
      n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, 
      n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, 
      n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, 
      n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, 
      n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, 
      n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, 
      n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, 
      n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, 
      n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, 
      n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, 
      n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, 
      n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, 
      n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, 
      n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, 
      n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, 
      n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, 
      n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, 
      n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, 
      n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, 
      n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, 
      n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, 
      n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, 
      n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, 
      n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, 
      n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, 
      n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, 
      n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, 
      n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, 
      n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, 
      n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, 
      n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, 
      n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, 
      n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, 
      n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, 
      n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, 
      n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, 
      n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, 
      n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, 
      n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, 
      n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, 
      n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, 
      n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, 
      n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, 
      n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, 
      n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, 
      n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, 
      n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, 
      n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, 
      n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, 
      n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, 
      n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, 
      n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, 
      n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, 
      n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, 
      n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, 
      n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, 
      n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, 
      n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, 
      n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, 
      n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, 
      n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, 
      n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, 
      n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, 
      n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, 
      n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, 
      n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, 
      n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, 
      n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, 
      n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, 
      n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, 
      n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, 
      n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, 
      n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, 
      n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, 
      n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, 
      n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, 
      n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, 
      n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, 
      n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, 
      n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, 
      n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, 
      n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, 
      n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, 
      n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, 
      n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, 
      n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, 
      n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, 
      n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, 
      n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, 
      n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, 
      n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, 
      n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, 
      n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, 
      n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, 
      n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, 
      n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, 
      n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, 
      n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, 
      n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, 
      n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, 
      n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, 
      n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, 
      n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, 
      n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, 
      n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, 
      n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, 
      n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, 
      n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, 
      n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, 
      n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, 
      n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, 
      n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, 
      n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, 
      n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, 
      n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, 
      n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, 
      n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, 
      n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, 
      n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, 
      n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, 
      n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, 
      n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, 
      n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, 
      n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, 
      n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, 
      n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, 
      n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, 
      n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, 
      n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, 
      n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, 
      n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, 
      n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, 
      n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, 
      n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, 
      n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, 
      n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, 
      n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, 
      n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, 
      n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, 
      n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, 
      n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, 
      n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, 
      n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, 
      n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, 
      n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, 
      n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, 
      n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, 
      n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, 
      n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, 
      n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, 
      n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, 
      n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, 
      n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, 
      n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, 
      n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, 
      n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, 
      n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, 
      n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, 
      n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, 
      n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, 
      n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, 
      n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, 
      n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, 
      n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, 
      n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, 
      n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, 
      n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, 
      n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, 
      n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, 
      n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, 
      n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, 
      n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, 
      n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, 
      n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, 
      n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, 
      n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, 
      n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, 
      n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, 
      n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, 
      n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, 
      n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, 
      n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, 
      n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, 
      n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, 
      n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, 
      n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, 
      n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, 
      n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, 
      n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, 
      n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, 
      n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, 
      n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, 
      n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, 
      n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, 
      n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, 
      n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, 
      n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, 
      n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, 
      n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, 
      n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, 
      n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, 
      n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, 
      n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, 
      n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, 
      n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, 
      n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, 
      n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, 
      n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, 
      n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, 
      n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, 
      n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, 
      n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, 
      n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, 
      n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, 
      n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, 
      n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, 
      n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, 
      n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, 
      n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, 
      n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, 
      n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, 
      n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, 
      n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, 
      n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, 
      n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, 
      n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, 
      n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, 
      n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, 
      n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, 
      n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, 
      n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, 
      n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, 
      n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, 
      n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, 
      n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, 
      n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, 
      n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, 
      n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, 
      n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, 
      n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, 
      n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, 
      n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, 
      n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, 
      n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, 
      n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, 
      n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, 
      n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, 
      n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, 
      n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, 
      n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, 
      n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, 
      n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, 
      n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, 
      n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, 
      n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, 
      n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, 
      n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, 
      n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, 
      n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, 
      n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, 
      n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, 
      n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, 
      n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, 
      n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, 
      n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, 
      n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, 
      n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, 
      n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, 
      n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, 
      n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, 
      n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, 
      n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, 
      n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, 
      n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, 
      n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, 
      n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, 
      n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, 
      n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, 
      n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, 
      n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, 
      n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, 
      n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, 
      n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, 
      n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, 
      n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, 
      n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, 
      n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, 
      n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, 
      n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, 
      n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, 
      n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, 
      n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, 
      n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, 
      n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, 
      n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, 
      n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, 
      n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, 
      n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, 
      n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, 
      n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, 
      n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, 
      n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, 
      n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, 
      n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, 
      n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, 
      n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, 
      n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, 
      n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, 
      n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, 
      n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, 
      n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, 
      n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, 
      n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, 
      n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, 
      n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, 
      n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, 
      n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, 
      n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, 
      n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, 
      n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, 
      n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, 
      n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, 
      n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, 
      n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, 
      n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, 
      n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, 
      n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, 
      n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, 
      n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, 
      n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, 
      n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, 
      n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, 
      n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, 
      n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, 
      n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, 
      n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, 
      n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, 
      n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, 
      n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, 
      n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, 
      n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, 
      n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, 
      n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, 
      n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, 
      n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, 
      n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, 
      n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, 
      n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, 
      n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, 
      n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, 
      n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, 
      n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, 
      n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, 
      n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, 
      n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, 
      n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, 
      n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, 
      n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, 
      n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, 
      n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, 
      n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, 
      n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, 
      n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, 
      n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, 
      n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, 
      n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, 
      n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, 
      n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, 
      n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, 
      n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, 
      n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, 
      n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, 
      n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, 
      n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, 
      n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, 
      n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, 
      n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, 
      n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, 
      n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, 
      n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, 
      n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, 
      n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, 
      n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, 
      n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, 
      n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, 
      n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, 
      n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, 
      n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, 
      n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, 
      n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, 
      n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, 
      n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, 
      n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, 
      n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, 
      n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, 
      n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, 
      n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, 
      n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, 
      n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, 
      n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, 
      n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, 
      n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, 
      n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, 
      n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, 
      n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, 
      n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, 
      n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, 
      n14518, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, 
      n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, 
      n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, 
      n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, 
      n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, 
      n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, 
      n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, 
      n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, 
      n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, 
      n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, 
      n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, 
      n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, 
      n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, 
      n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, 
      n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, 
      n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, 
      n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, 
      n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, 
      n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, 
      n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, 
      n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, 
      n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, 
      n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, 
      n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, 
      n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, 
      n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, 
      n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, 
      n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, 
      n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, 
      n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, 
      n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, 
      n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, 
      n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, 
      n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, 
      n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, 
      n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, 
      n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, 
      n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, 
      n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, 
      n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, 
      n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, 
      n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, 
      n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, 
      n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, 
      n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, 
      n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, 
      n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, 
      n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, 
      n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, 
      n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, 
      n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, 
      n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, 
      n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, 
      n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, 
      n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, 
      n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, 
      n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, 
      n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, 
      n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, 
      n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, 
      n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, 
      n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, 
      n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, 
      n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, 
      n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, 
      n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, 
      n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, 
      n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, 
      n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, 
      n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, 
      n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, 
      n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, 
      n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, 
      n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, 
      n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, 
      n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, 
      n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, 
      n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, 
      n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, 
      n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, 
      n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, 
      n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, 
      n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, 
      n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, 
      n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, 
      n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, 
      n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, 
      n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, 
      n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, 
      n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, 
      n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, 
      n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, 
      n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, 
      n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, 
      n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, 
      n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, 
      n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, 
      n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, 
      n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, 
      n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, 
      n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, 
      n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, 
      n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, 
      n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, 
      n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, 
      n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, 
      n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, 
      n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, 
      n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, 
      n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, 
      n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, 
      n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, 
      n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, 
      n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, 
      n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, 
      n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, 
      n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, 
      n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, 
      n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, 
      n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, 
      n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, 
      n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, 
      n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, 
      n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, 
      n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, 
      n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, 
      n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, 
      n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, 
      n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, 
      n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, 
      n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, 
      n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, 
      n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, 
      n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, 
      n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, 
      n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, 
      n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, 
      n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, 
      n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, 
      n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, 
      n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, 
      n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, 
      n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, 
      n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, 
      n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, 
      n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, 
      n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, 
      n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, 
      n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, 
      n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, 
      n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, 
      n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, 
      n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, 
      n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, 
      n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, 
      n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, 
      n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, 
      n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, 
      n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, 
      n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, 
      n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, 
      n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, 
      n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, 
      n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, 
      n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, 
      n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, 
      n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, 
      n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, 
      n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, 
      n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, 
      n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, 
      n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, 
      n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, 
      n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, 
      n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, 
      n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, 
      n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, 
      n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, 
      n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, 
      n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, 
      n_2963, n_2964, n_2965 : std_logic;

begin
   
   CWP_reg_6_inst : DFFR_X1 port map( D => n9132, CK => CLK, RN => n12662, Q =>
                           n_1173, QN => n2935);
   CWP_reg_4_inst : DFFR_X1 port map( D => n12778, CK => CLK, RN => n12662, Q 
                           => n10625, QN => n2937);
   CWP_reg_5_inst : DFFR_X1 port map( D => n9133, CK => CLK, RN => n12662, Q =>
                           n10626, QN => n2936);
   REGISTERS_reg_0_31_inst : DFFR_X1 port map( D => n6316, CK => CLK, RN => 
                           n12655, Q => n_1174, QN => n1871);
   REGISTERS_reg_0_30_inst : DFFR_X1 port map( D => n6317, CK => CLK, RN => 
                           n12618, Q => n_1175, QN => n1883);
   REGISTERS_reg_0_29_inst : DFFR_X1 port map( D => n6318, CK => CLK, RN => 
                           n12604, Q => n_1176, QN => n1895);
   REGISTERS_reg_0_28_inst : DFFR_X1 port map( D => n6319, CK => CLK, RN => 
                           n12611, Q => n_1177, QN => n1907);
   REGISTERS_reg_0_27_inst : DFFR_X1 port map( D => n6320, CK => CLK, RN => 
                           n12582, Q => n_1178, QN => n1919);
   REGISTERS_reg_0_26_inst : DFFR_X1 port map( D => n6321, CK => CLK, RN => 
                           n12560, Q => n_1179, QN => n1931);
   REGISTERS_reg_0_25_inst : DFFR_X1 port map( D => n6322, CK => CLK, RN => 
                           n12538, Q => n_1180, QN => n1943);
   REGISTERS_reg_0_24_inst : DFFR_X1 port map( D => n6323, CK => CLK, RN => 
                           n12512, Q => n_1181, QN => n1955);
   REGISTERS_reg_0_23_inst : DFFR_X1 port map( D => n6324, CK => CLK, RN => 
                           n12626, Q => n_1182, QN => n1967);
   REGISTERS_reg_0_22_inst : DFFR_X1 port map( D => n6325, CK => CLK, RN => 
                           n12485, Q => n_1183, QN => n1979);
   REGISTERS_reg_0_21_inst : DFFR_X1 port map( D => n6326, CK => CLK, RN => 
                           n12523, Q => n_1184, QN => n1991);
   REGISTERS_reg_0_20_inst : DFFR_X1 port map( D => n6327, CK => CLK, RN => 
                           n12498, Q => n_1185, QN => n2003);
   REGISTERS_reg_0_19_inst : DFFR_X1 port map( D => n6328, CK => CLK, RN => 
                           n12589, Q => n_1186, QN => n2015);
   REGISTERS_reg_0_18_inst : DFFR_X1 port map( D => n6329, CK => CLK, RN => 
                           n12440, Q => n_1187, QN => n2027);
   REGISTERS_reg_0_17_inst : DFFR_X1 port map( D => n6330, CK => CLK, RN => 
                           n12447, Q => n_1188, QN => n2039);
   REGISTERS_reg_0_16_inst : DFFR_X1 port map( D => n6331, CK => CLK, RN => 
                           n12499, Q => n_1189, QN => n2083);
   REGISTERS_reg_0_15_inst : DFFR_X1 port map( D => n6332, CK => CLK, RN => 
                           n12633, Q => n_1190, QN => n2095);
   REGISTERS_reg_0_14_inst : DFFR_X1 port map( D => n6333, CK => CLK, RN => 
                           n12461, Q => n_1191, QN => n2107);
   REGISTERS_reg_0_13_inst : DFFR_X1 port map( D => n6334, CK => CLK, RN => 
                           n12468, Q => n_1192, QN => n2151);
   REGISTERS_reg_0_12_inst : DFFR_X1 port map( D => n6335, CK => CLK, RN => 
                           n12476, Q => n_1193, QN => n2163);
   REGISTERS_reg_0_11_inst : DFFR_X1 port map( D => n6336, CK => CLK, RN => 
                           n12567, Q => n_1194, QN => n2175);
   REGISTERS_reg_0_10_inst : DFFR_X1 port map( D => n6337, CK => CLK, RN => 
                           n12545, Q => n_1195, QN => n2219);
   REGISTERS_reg_0_9_inst : DFFR_X1 port map( D => n6338, CK => CLK, RN => 
                           n12552, Q => n_1196, QN => n2231);
   REGISTERS_reg_0_8_inst : DFFR_X1 port map( D => n6339, CK => CLK, RN => 
                           n12530, Q => n_1197, QN => n2243);
   REGISTERS_reg_0_7_inst : DFFR_X1 port map( D => n6340, CK => CLK, RN => 
                           n12640, Q => n_1198, QN => n2255);
   REGISTERS_reg_0_6_inst : DFFR_X1 port map( D => n6341, CK => CLK, RN => 
                           n12596, Q => n_1199, QN => n2267);
   REGISTERS_reg_0_5_inst : DFFR_X1 port map( D => n6342, CK => CLK, RN => 
                           n12483, Q => n_1200, QN => n2279);
   REGISTERS_reg_0_4_inst : DFFR_X1 port map( D => n6343, CK => CLK, RN => 
                           n12490, Q => n_1201, QN => n2291);
   REGISTERS_reg_0_3_inst : DFFR_X1 port map( D => n6344, CK => CLK, RN => 
                           n12574, Q => n_1202, QN => n2303);
   REGISTERS_reg_0_2_inst : DFFR_X1 port map( D => n6345, CK => CLK, RN => 
                           n12505, Q => n_1203, QN => n2315);
   REGISTERS_reg_0_1_inst : DFFR_X1 port map( D => n6346, CK => CLK, RN => 
                           n12433, Q => n_1204, QN => n2327);
   REGISTERS_reg_0_0_inst : DFFR_X1 port map( D => n6347, CK => CLK, RN => 
                           n12648, Q => n_1205, QN => n2339);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n6348, CK => CLK, RN => 
                           n12655, Q => n_1206, QN => n143);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n6349, CK => CLK, RN => 
                           n12618, Q => n_1207, QN => n155);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n6350, CK => CLK, RN => 
                           n12604, Q => n_1208, QN => n167);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n6351, CK => CLK, RN => 
                           n12611, Q => n_1209, QN => n179);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n6352, CK => CLK, RN => 
                           n12582, Q => n_1210, QN => n191);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n6353, CK => CLK, RN => 
                           n12560, Q => n_1211, QN => n203);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n6354, CK => CLK, RN => 
                           n12538, Q => n_1212, QN => n215);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n6355, CK => CLK, RN => 
                           n12512, Q => n_1213, QN => n227);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n6356, CK => CLK, RN => 
                           n12626, Q => n_1214, QN => n239);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n6357, CK => CLK, RN => 
                           n12484, Q => n_1215, QN => n251);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n6358, CK => CLK, RN => 
                           n12523, Q => n_1216, QN => n263);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n6359, CK => CLK, RN => 
                           n12498, Q => n_1217, QN => n275);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n6360, CK => CLK, RN => 
                           n12589, Q => n_1218, QN => n287);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n6361, CK => CLK, RN => 
                           n12440, Q => n_1219, QN => n299);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n6362, CK => CLK, RN => 
                           n12447, Q => n_1220, QN => n311);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n6363, CK => CLK, RN => 
                           n12498, Q => n_1221, QN => n323);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n6364, CK => CLK, RN => 
                           n12633, Q => n_1222, QN => n335);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n6365, CK => CLK, RN => 
                           n12461, Q => n_1223, QN => n347);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n6366, CK => CLK, RN => 
                           n12468, Q => n_1224, QN => n359);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n6367, CK => CLK, RN => 
                           n12476, Q => n_1225, QN => n371);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n6368, CK => CLK, RN => 
                           n12567, Q => n_1226, QN => n383);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n6369, CK => CLK, RN => 
                           n12545, Q => n_1227, QN => n395);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n6370, CK => CLK, RN => 
                           n12552, Q => n_1228, QN => n407);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n6371, CK => CLK, RN => 
                           n12530, Q => n_1229, QN => n419);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n6372, CK => CLK, RN => 
                           n12640, Q => n_1230, QN => n431);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n6373, CK => CLK, RN => 
                           n12596, Q => n_1231, QN => n443);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n6374, CK => CLK, RN => 
                           n12483, Q => n_1232, QN => n455);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n6375, CK => CLK, RN => 
                           n12490, Q => n_1233, QN => n467);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n6376, CK => CLK, RN => 
                           n12574, Q => n_1234, QN => n479);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n6377, CK => CLK, RN => 
                           n12505, Q => n_1235, QN => n491);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n6378, CK => CLK, RN => 
                           n12433, Q => n_1236, QN => n503);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n6379, CK => CLK, RN => 
                           n12648, Q => n_1237, QN => n515);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n6380, CK => CLK, RN => 
                           n12655, Q => n_1238, QN => n12780);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n6381, CK => CLK, RN => 
                           n12618, Q => n_1239, QN => n12781);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n6382, CK => CLK, RN => 
                           n12604, Q => n_1240, QN => n12782);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n6383, CK => CLK, RN => 
                           n12611, Q => n_1241, QN => n1043);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n6384, CK => CLK, RN => 
                           n12582, Q => n_1242, QN => n1055);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n6385, CK => CLK, RN => 
                           n12560, Q => n_1243, QN => n1067);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n6386, CK => CLK, RN => 
                           n12538, Q => n_1244, QN => n1079);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n6387, CK => CLK, RN => 
                           n12512, Q => n_1245, QN => n1091);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n6388, CK => CLK, RN => 
                           n12626, Q => n_1246, QN => n1103);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n6389, CK => CLK, RN => 
                           n12483, Q => n_1247, QN => n1115);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n6390, CK => CLK, RN => 
                           n12523, Q => n_1248, QN => n1127);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n6391, CK => CLK, RN => 
                           n12498, Q => n_1249, QN => n1139);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n6392, CK => CLK, RN => 
                           n12589, Q => n_1250, QN => n1151);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n6393, CK => CLK, RN => 
                           n12440, Q => n_1251, QN => n1163);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n6394, CK => CLK, RN => 
                           n12447, Q => n_1252, QN => n1175);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n6395, CK => CLK, RN => 
                           n12497, Q => n_1253, QN => n1187);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n6396, CK => CLK, RN => 
                           n12633, Q => n_1254, QN => n1199);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n6397, CK => CLK, RN => 
                           n12461, Q => n_1255, QN => n1211);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n6398, CK => CLK, RN => 
                           n12468, Q => n_1256, QN => n1223);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n6399, CK => CLK, RN => 
                           n12476, Q => n_1257, QN => n1235);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n6400, CK => CLK, RN => 
                           n12567, Q => n_1258, QN => n1247);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n6401, CK => CLK, RN => 
                           n12545, Q => n_1259, QN => n1259);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n6402, CK => CLK, RN => 
                           n12552, Q => n_1260, QN => n1271);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n6403, CK => CLK, RN => 
                           n12530, Q => n_1261, QN => n1283);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n6404, CK => CLK, RN => 
                           n12640, Q => n_1262, QN => n1295);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n6405, CK => CLK, RN => 
                           n12596, Q => n_1263, QN => n1307);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n6406, CK => CLK, RN => 
                           n12483, Q => n_1264, QN => n1319);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n6407, CK => CLK, RN => 
                           n12490, Q => n_1265, QN => n1331);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n6408, CK => CLK, RN => 
                           n12574, Q => n_1266, QN => n1343);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n6409, CK => CLK, RN => 
                           n12505, Q => n_1267, QN => n1387);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n6410, CK => CLK, RN => 
                           n12433, Q => n_1268, QN => n1399);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n6411, CK => CLK, RN => 
                           n12648, Q => n_1269, QN => n1443);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n6412, CK => CLK, RN => 
                           n12655, Q => n_1270, QN => n1870);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n6413, CK => CLK, RN => 
                           n12618, Q => n_1271, QN => n1882);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n6414, CK => CLK, RN => 
                           n12604, Q => n_1272, QN => n1894);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n6415, CK => CLK, RN => 
                           n12611, Q => n_1273, QN => n1906);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n6416, CK => CLK, RN => 
                           n12582, Q => n_1274, QN => n1918);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n6417, CK => CLK, RN => 
                           n12560, Q => n_1275, QN => n1930);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n6418, CK => CLK, RN => 
                           n12538, Q => n_1276, QN => n1942);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n6419, CK => CLK, RN => 
                           n12512, Q => n_1277, QN => n1954);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n6420, CK => CLK, RN => 
                           n12626, Q => n_1278, QN => n1966);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n6421, CK => CLK, RN => 
                           n12482, Q => n_1279, QN => n1978);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n6422, CK => CLK, RN => 
                           n12523, Q => n_1280, QN => n1990);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n6423, CK => CLK, RN => 
                           n12498, Q => n_1281, QN => n2002);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n6424, CK => CLK, RN => 
                           n12589, Q => n_1282, QN => n2014);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n6425, CK => CLK, RN => 
                           n12440, Q => n_1283, QN => n2026);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n6426, CK => CLK, RN => 
                           n12447, Q => n_1284, QN => n2038);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n6427, CK => CLK, RN => 
                           n12496, Q => n_1285, QN => n2082);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n6428, CK => CLK, RN => 
                           n12633, Q => n_1286, QN => n2094);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n6429, CK => CLK, RN => 
                           n12461, Q => n_1287, QN => n2106);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n6430, CK => CLK, RN => 
                           n12468, Q => n_1288, QN => n2150);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n6431, CK => CLK, RN => 
                           n12476, Q => n_1289, QN => n2162);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n6432, CK => CLK, RN => 
                           n12567, Q => n_1290, QN => n2174);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n6433, CK => CLK, RN => 
                           n12545, Q => n_1291, QN => n2218);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n6434, CK => CLK, RN => 
                           n12552, Q => n_1292, QN => n2230);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n6435, CK => CLK, RN => 
                           n12530, Q => n_1293, QN => n2242);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n6436, CK => CLK, RN => 
                           n12640, Q => n_1294, QN => n2254);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n6437, CK => CLK, RN => 
                           n12596, Q => n_1295, QN => n2266);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n6438, CK => CLK, RN => 
                           n12483, Q => n_1296, QN => n2278);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n6439, CK => CLK, RN => 
                           n12490, Q => n_1297, QN => n2290);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n6440, CK => CLK, RN => 
                           n12574, Q => n_1298, QN => n2302);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n6441, CK => CLK, RN => 
                           n12505, Q => n_1299, QN => n2314);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n6442, CK => CLK, RN => 
                           n12433, Q => n_1300, QN => n2326);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n6443, CK => CLK, RN => 
                           n12648, Q => n_1301, QN => n2338);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n6444, CK => CLK, RN => 
                           n12655, Q => n_1302, QN => n142);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n6445, CK => CLK, RN => 
                           n12619, Q => n_1303, QN => n154);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n6446, CK => CLK, RN => 
                           n12604, Q => n_1304, QN => n166);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n6447, CK => CLK, RN => 
                           n12611, Q => n_1305, QN => n178);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n6448, CK => CLK, RN => 
                           n12582, Q => n_1306, QN => n190);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n6449, CK => CLK, RN => 
                           n12560, Q => n_1307, QN => n202);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n6450, CK => CLK, RN => 
                           n12538, Q => n_1308, QN => n214);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n6451, CK => CLK, RN => 
                           n12513, Q => n_1309, QN => n226);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n6452, CK => CLK, RN => 
                           n12626, Q => n_1310, QN => n238);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n6453, CK => CLK, RN => 
                           n12474, Q => n_1311, QN => n250);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n6454, CK => CLK, RN => 
                           n12523, Q => n_1312, QN => n262);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n6455, CK => CLK, RN => 
                           n12498, Q => n_1313, QN => n274);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n6456, CK => CLK, RN => 
                           n12589, Q => n_1314, QN => n286);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n6457, CK => CLK, RN => 
                           n12440, Q => n_1315, QN => n298);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n6458, CK => CLK, RN => 
                           n12448, Q => n_1316, QN => n310);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n6459, CK => CLK, RN => 
                           n12495, Q => n_1317, QN => n322);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n6460, CK => CLK, RN => 
                           n12633, Q => n_1318, QN => n334);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n6461, CK => CLK, RN => 
                           n12461, Q => n_1319, QN => n346);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n6462, CK => CLK, RN => 
                           n12469, Q => n_1320, QN => n358);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n6463, CK => CLK, RN => 
                           n12476, Q => n_1321, QN => n370);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n6464, CK => CLK, RN => 
                           n12567, Q => n_1322, QN => n382);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n6465, CK => CLK, RN => 
                           n12545, Q => n_1323, QN => n394);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n6466, CK => CLK, RN => 
                           n12553, Q => n_1324, QN => n406);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n6467, CK => CLK, RN => 
                           n12531, Q => n_1325, QN => n418);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n6468, CK => CLK, RN => 
                           n12641, Q => n_1326, QN => n430);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n6469, CK => CLK, RN => 
                           n12597, Q => n_1327, QN => n442);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n6470, CK => CLK, RN => 
                           n12483, Q => n_1328, QN => n454);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n6471, CK => CLK, RN => 
                           n12491, Q => n_1329, QN => n466);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n6472, CK => CLK, RN => 
                           n12575, Q => n_1330, QN => n478);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n6473, CK => CLK, RN => 
                           n12505, Q => n_1331, QN => n490);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n6474, CK => CLK, RN => 
                           n12433, Q => n_1332, QN => n502);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n6475, CK => CLK, RN => 
                           n12648, Q => n_1333, QN => n514);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n6476, CK => CLK, RN => 
                           n12655, Q => n_1334, QN => n12783);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n6477, CK => CLK, RN => 
                           n12619, Q => n_1335, QN => n12784);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n6478, CK => CLK, RN => 
                           n12604, Q => n_1336, QN => n12785);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n6479, CK => CLK, RN => 
                           n12611, Q => n_1337, QN => n1042);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n6480, CK => CLK, RN => 
                           n12582, Q => n_1338, QN => n1054);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n6481, CK => CLK, RN => 
                           n12560, Q => n_1339, QN => n1066);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n6482, CK => CLK, RN => 
                           n12538, Q => n_1340, QN => n1078);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n6483, CK => CLK, RN => 
                           n12513, Q => n_1341, QN => n1090);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n6484, CK => CLK, RN => 
                           n12626, Q => n_1342, QN => n1102);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n6485, CK => CLK, RN => 
                           n12516, Q => n_1343, QN => n1114);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n6486, CK => CLK, RN => 
                           n12523, Q => n_1344, QN => n1126);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n6487, CK => CLK, RN => 
                           n12498, Q => n_1345, QN => n1138);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n6488, CK => CLK, RN => 
                           n12589, Q => n_1346, QN => n1150);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n6489, CK => CLK, RN => 
                           n12440, Q => n_1347, QN => n1162);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n6490, CK => CLK, RN => 
                           n12448, Q => n_1348, QN => n1174);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n6491, CK => CLK, RN => 
                           n12494, Q => n_1349, QN => n1186);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n6492, CK => CLK, RN => 
                           n12633, Q => n_1350, QN => n1198);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n6493, CK => CLK, RN => 
                           n12461, Q => n_1351, QN => n1210);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n6494, CK => CLK, RN => 
                           n12469, Q => n_1352, QN => n1222);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n6495, CK => CLK, RN => 
                           n12476, Q => n_1353, QN => n1234);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n6496, CK => CLK, RN => 
                           n12567, Q => n_1354, QN => n1246);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n6497, CK => CLK, RN => 
                           n12545, Q => n_1355, QN => n1258);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n6498, CK => CLK, RN => 
                           n12553, Q => n_1356, QN => n1270);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n6499, CK => CLK, RN => 
                           n12531, Q => n_1357, QN => n1282);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n6500, CK => CLK, RN => 
                           n12641, Q => n_1358, QN => n1294);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n6501, CK => CLK, RN => 
                           n12597, Q => n_1359, QN => n1306);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n6502, CK => CLK, RN => 
                           n12483, Q => n_1360, QN => n1318);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n6503, CK => CLK, RN => 
                           n12491, Q => n_1361, QN => n1330);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n6504, CK => CLK, RN => 
                           n12575, Q => n_1362, QN => n1342);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n6505, CK => CLK, RN => 
                           n12505, Q => n_1363, QN => n1386);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n6506, CK => CLK, RN => 
                           n12433, Q => n_1364, QN => n1398);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n6507, CK => CLK, RN => 
                           n12648, Q => n_1365, QN => n1442);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n6508, CK => CLK, RN => 
                           n12655, Q => n_1366, QN => n1869);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n6509, CK => CLK, RN => 
                           n12619, Q => n_1367, QN => n1881);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n6510, CK => CLK, RN => 
                           n12604, Q => n_1368, QN => n1893);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n6511, CK => CLK, RN => 
                           n12611, Q => n_1369, QN => n1905);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n6512, CK => CLK, RN => 
                           n12582, Q => n_1370, QN => n1917);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n6513, CK => CLK, RN => 
                           n12560, Q => n_1371, QN => n1929);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n6514, CK => CLK, RN => 
                           n12538, Q => n_1372, QN => n1941);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n6515, CK => CLK, RN => 
                           n12513, Q => n_1373, QN => n1953);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n6516, CK => CLK, RN => 
                           n12626, Q => n_1374, QN => n1965);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n6517, CK => CLK, RN => 
                           n12473, Q => n_1375, QN => n1977);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n6518, CK => CLK, RN => 
                           n12523, Q => n_1376, QN => n1989);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n6519, CK => CLK, RN => 
                           n12498, Q => n_1377, QN => n2001);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n6520, CK => CLK, RN => 
                           n12589, Q => n_1378, QN => n2013);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n6521, CK => CLK, RN => 
                           n12440, Q => n_1379, QN => n2025);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n6522, CK => CLK, RN => 
                           n12448, Q => n_1380, QN => n2037);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n6523, CK => CLK, RN => 
                           n12493, Q => n_1381, QN => n2049);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n6524, CK => CLK, RN => 
                           n12633, Q => n_1382, QN => n2093);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n6525, CK => CLK, RN => 
                           n12461, Q => n_1383, QN => n2105);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n6526, CK => CLK, RN => 
                           n12469, Q => n_1384, QN => n2149);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n6527, CK => CLK, RN => 
                           n12476, Q => n_1385, QN => n2161);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n6528, CK => CLK, RN => 
                           n12567, Q => n_1386, QN => n2173_port);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n6529, CK => CLK, RN => 
                           n12545, Q => n_1387, QN => n2217);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n6530, CK => CLK, RN => 
                           n12553, Q => n_1388, QN => n2229);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n6531, CK => CLK, RN => 
                           n12531, Q => n_1389, QN => n2241);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n6532, CK => CLK, RN => 
                           n12641, Q => n_1390, QN => n2253);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n6533, CK => CLK, RN => 
                           n12597, Q => n_1391, QN => n2265);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n6534, CK => CLK, RN => 
                           n12483, Q => n_1392, QN => n2277);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n6535, CK => CLK, RN => 
                           n12491, Q => n_1393, QN => n2289);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n6536, CK => CLK, RN => 
                           n12575, Q => n_1394, QN => n2301);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n6537, CK => CLK, RN => 
                           n12505, Q => n_1395, QN => n2313);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n6538, CK => CLK, RN => 
                           n12433, Q => n_1396, QN => n2325);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n6539, CK => CLK, RN => 
                           n12648, Q => n_1397, QN => n2337);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n6540, CK => CLK, RN => 
                           n12655, Q => n_1398, QN => n141);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n6541, CK => CLK, RN => 
                           n12619, Q => n_1399, QN => n153);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n6542, CK => CLK, RN => 
                           n12604, Q => n_1400, QN => n165);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n6543, CK => CLK, RN => 
                           n12611, Q => n_1401, QN => n177);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n6544, CK => CLK, RN => 
                           n12582, Q => n_1402, QN => n189);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n6545, CK => CLK, RN => 
                           n12560, Q => n_1403, QN => n201);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n6546, CK => CLK, RN => 
                           n12538, Q => n_1404, QN => n213);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n6547, CK => CLK, RN => 
                           n12513, Q => n_1405, QN => n225);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n6548, CK => CLK, RN => 
                           n12626, Q => n_1406, QN => n237);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n6549, CK => CLK, RN => 
                           n12472, Q => n_1407, QN => n249);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n6550, CK => CLK, RN => 
                           n12523, Q => n_1408, QN => n261);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n6551, CK => CLK, RN => 
                           n12498, Q => n_1409, QN => n273);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n6552, CK => CLK, RN => 
                           n12589, Q => n_1410, QN => n285);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n6553, CK => CLK, RN => 
                           n12440, Q => n_1411, QN => n297);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n6554, CK => CLK, RN => 
                           n12448, Q => n_1412, QN => n309);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n6555, CK => CLK, RN => 
                           n12492, Q => n_1413, QN => n321);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n6556, CK => CLK, RN => 
                           n12633, Q => n_1414, QN => n333);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n6557, CK => CLK, RN => 
                           n12461, Q => n_1415, QN => n345);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n6558, CK => CLK, RN => 
                           n12469, Q => n_1416, QN => n357);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n6559, CK => CLK, RN => 
                           n12476, Q => n_1417, QN => n369);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n6560, CK => CLK, RN => 
                           n12567, Q => n_1418, QN => n381);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n6561, CK => CLK, RN => 
                           n12545, Q => n_1419, QN => n393);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n6562, CK => CLK, RN => 
                           n12553, Q => n_1420, QN => n405);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n6563, CK => CLK, RN => 
                           n12531, Q => n_1421, QN => n417);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n6564, CK => CLK, RN => 
                           n12641, Q => n_1422, QN => n429);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n6565, CK => CLK, RN => 
                           n12597, Q => n_1423, QN => n441);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n6566, CK => CLK, RN => 
                           n12483, Q => n_1424, QN => n453);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n6567, CK => CLK, RN => 
                           n12491, Q => n_1425, QN => n465);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n6568, CK => CLK, RN => 
                           n12575, Q => n_1426, QN => n477);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n6569, CK => CLK, RN => 
                           n12505, Q => n_1427, QN => n489);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n6570, CK => CLK, RN => 
                           n12433, Q => n_1428, QN => n501);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n6571, CK => CLK, RN => 
                           n12648, Q => n_1429, QN => n513);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n6572, CK => CLK, RN => 
                           n12656, Q => n_1430, QN => n12786);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n6573, CK => CLK, RN => 
                           n12619, Q => n_1431, QN => n12787);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n6574, CK => CLK, RN => 
                           n12604, Q => n_1432, QN => n1029);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n6575, CK => CLK, RN => 
                           n12612, Q => n_1433, QN => n1041);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n6576, CK => CLK, RN => 
                           n12582, Q => n_1434, QN => n1053);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n6577, CK => CLK, RN => 
                           n12560, Q => n_1435, QN => n1065);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n6578, CK => CLK, RN => 
                           n12538, Q => n_1436, QN => n1077);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n6579, CK => CLK, RN => 
                           n12513, Q => n_1437, QN => n1089);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n6580, CK => CLK, RN => 
                           n12626, Q => n_1438, QN => n1101);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n6581, CK => CLK, RN => 
                           n12471, Q => n_1439, QN => n1113);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n6582, CK => CLK, RN => 
                           n12524, Q => n_1440, QN => n1125);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n6583, CK => CLK, RN => 
                           n12498, Q => n_1441, QN => n1137);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n6584, CK => CLK, RN => 
                           n12590, Q => n_1442, QN => n1149);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n6585, CK => CLK, RN => 
                           n12441, Q => n_1443, QN => n1161);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n6586, CK => CLK, RN => 
                           n12448, Q => n_1444, QN => n1173);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n6587, CK => CLK, RN => 
                           n12491, Q => n_1445, QN => n1185);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n6588, CK => CLK, RN => 
                           n12634, Q => n_1446, QN => n1197);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n6589, CK => CLK, RN => 
                           n12462, Q => n_1447, QN => n1209);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n6590, CK => CLK, RN => 
                           n12469, Q => n_1448, QN => n1221);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n6591, CK => CLK, RN => 
                           n12476, Q => n_1449, QN => n1233);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n6592, CK => CLK, RN => 
                           n12568, Q => n_1450, QN => n1245);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n6593, CK => CLK, RN => 
                           n12546, Q => n_1451, QN => n1257);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n6594, CK => CLK, RN => 
                           n12553, Q => n_1452, QN => n1269);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n6595, CK => CLK, RN => 
                           n12531, Q => n_1453, QN => n1281);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n6596, CK => CLK, RN => 
                           n12641, Q => n_1454, QN => n1293);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n6597, CK => CLK, RN => 
                           n12597, Q => n_1455, QN => n1305);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n6598, CK => CLK, RN => 
                           n12484, Q => n_1456, QN => n1317);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n6599, CK => CLK, RN => 
                           n12491, Q => n_1457, QN => n1329);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n6600, CK => CLK, RN => 
                           n12575, Q => n_1458, QN => n1341);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n6601, CK => CLK, RN => 
                           n12506, Q => n_1459, QN => n1385);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n6602, CK => CLK, RN => 
                           n12433, Q => n_1460, QN => n1397);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n6603, CK => CLK, RN => 
                           n12648, Q => n_1461, QN => n1409);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n6604, CK => CLK, RN => 
                           n12656, Q => n_1462, QN => n871);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n6605, CK => CLK, RN => 
                           n12619, Q => n_1463, QN => n875);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n6606, CK => CLK, RN => 
                           n12604, Q => n_1464, QN => n879);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n6607, CK => CLK, RN => 
                           n12612, Q => n_1465, QN => n883);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n6608, CK => CLK, RN => 
                           n12582, Q => n_1466, QN => n887);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n6609, CK => CLK, RN => 
                           n12560, Q => n_1467, QN => n891);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n6610, CK => CLK, RN => 
                           n12538, Q => n_1468, QN => n895);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n6611, CK => CLK, RN => 
                           n12513, Q => n_1469, QN => n899);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n6612, CK => CLK, RN => 
                           n12626, Q => n_1470, QN => n903);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n6613, CK => CLK, RN => 
                           n12470, Q => n_1471, QN => n907);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n6614, CK => CLK, RN => 
                           n12524, Q => n_1472, QN => n911);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n6615, CK => CLK, RN => 
                           n12498, Q => n_1473, QN => n915);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n6616, CK => CLK, RN => 
                           n12590, Q => n_1474, QN => n919);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n6617, CK => CLK, RN => 
                           n12441, Q => n_1475, QN => n923);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n6618, CK => CLK, RN => 
                           n12448, Q => n_1476, QN => n927);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n6619, CK => CLK, RN => 
                           n12490, Q => n_1477, QN => n931);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n6620, CK => CLK, RN => 
                           n12634, Q => n_1478, QN => n935);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n6621, CK => CLK, RN => 
                           n12462, Q => n_1479, QN => n939);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n6622, CK => CLK, RN => 
                           n12469, Q => n_1480, QN => n943);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n6623, CK => CLK, RN => 
                           n12476, Q => n_1481, QN => n947);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n6624, CK => CLK, RN => 
                           n12568, Q => n_1482, QN => n951);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n6625, CK => CLK, RN => 
                           n12546, Q => n_1483, QN => n955);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n6626, CK => CLK, RN => 
                           n12553, Q => n_1484, QN => n959);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n6627, CK => CLK, RN => 
                           n12531, Q => n_1485, QN => n963);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n6628, CK => CLK, RN => 
                           n12641, Q => n_1486, QN => n967);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n6629, CK => CLK, RN => 
                           n12597, Q => n_1487, QN => n971);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n6630, CK => CLK, RN => 
                           n12484, Q => n_1488, QN => n975);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n6631, CK => CLK, RN => 
                           n12491, Q => n_1489, QN => n979);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n6632, CK => CLK, RN => 
                           n12575, Q => n_1490, QN => n983);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n6633, CK => CLK, RN => 
                           n12506, Q => n_1491, QN => n987);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n6634, CK => CLK, RN => 
                           n12433, Q => n_1492, QN => n991);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n6635, CK => CLK, RN => 
                           n12648, Q => n_1493, QN => n995);
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n6636, CK => CLK, RN => 
                           n12656, Q => n_1494, QN => n1735);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n6637, CK => CLK, RN => 
                           n12619, Q => n_1495, QN => n1739);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n6638, CK => CLK, RN => 
                           n12604, Q => n_1496, QN => n1743);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n6639, CK => CLK, RN => 
                           n12612, Q => n_1497, QN => n1747);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n6640, CK => CLK, RN => 
                           n12582, Q => n_1498, QN => n1751);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n6641, CK => CLK, RN => 
                           n12560, Q => n_1499, QN => n1755);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n6642, CK => CLK, RN => 
                           n12538, Q => n_1500, QN => n1759);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n6643, CK => CLK, RN => 
                           n12513, Q => n_1501, QN => n1763);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n6644, CK => CLK, RN => 
                           n12626, Q => n_1502, QN => n1767);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n6645, CK => CLK, RN => 
                           n12486, Q => n_1503, QN => n1771);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n6646, CK => CLK, RN => 
                           n12524, Q => n_1504, QN => n1775);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n6647, CK => CLK, RN => 
                           n12498, Q => n_1505, QN => n1779);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n6648, CK => CLK, RN => 
                           n12590, Q => n_1506, QN => n1783);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n6649, CK => CLK, RN => 
                           n12441, Q => n_1507, QN => n1787);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n6650, CK => CLK, RN => 
                           n12448, Q => n_1508, QN => n1791);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n6651, CK => CLK, RN => 
                           n12500, Q => n_1509, QN => n1795);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n6652, CK => CLK, RN => 
                           n12634, Q => n_1510, QN => n1799);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n6653, CK => CLK, RN => 
                           n12462, Q => n_1511, QN => n1803);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n6654, CK => CLK, RN => 
                           n12469, Q => n_1512, QN => n1807);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n6655, CK => CLK, RN => 
                           n12476, Q => n_1513, QN => n1811);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n6656, CK => CLK, RN => 
                           n12568, Q => n_1514, QN => n1815);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n6657, CK => CLK, RN => 
                           n12546, Q => n_1515, QN => n1819);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n6658, CK => CLK, RN => 
                           n12553, Q => n_1516, QN => n1823);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n6659, CK => CLK, RN => 
                           n12531, Q => n_1517, QN => n1827);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n6660, CK => CLK, RN => 
                           n12641, Q => n_1518, QN => n1831);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n6661, CK => CLK, RN => 
                           n12597, Q => n_1519, QN => n1835);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n6662, CK => CLK, RN => 
                           n12484, Q => n_1520, QN => n1839);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n6663, CK => CLK, RN => 
                           n12491, Q => n_1521, QN => n1843);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n6664, CK => CLK, RN => 
                           n12575, Q => n_1522, QN => n1847);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n6665, CK => CLK, RN => 
                           n12506, Q => n_1523, QN => n1851);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n6666, CK => CLK, RN => 
                           n12433, Q => n_1524, QN => n1855);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n6667, CK => CLK, RN => 
                           n12648, Q => n_1525, QN => n1859);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n6700, CK => CLK, RN => 
                           n12656, Q => n_1526, QN => n5736);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n6701, CK => CLK, RN => 
                           n12619, Q => n_1527, QN => n5768);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n6702, CK => CLK, RN => 
                           n12605, Q => n_1528, QN => n5800);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n6703, CK => CLK, RN => 
                           n12612, Q => n_1529, QN => n5832);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n6704, CK => CLK, RN => 
                           n12583, Q => n_1530, QN => n5864);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n6705, CK => CLK, RN => 
                           n12561, Q => n_1531, QN => n5896);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n6706, CK => CLK, RN => 
                           n12539, Q => n_1532, QN => n5928);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n6707, CK => CLK, RN => 
                           n12513, Q => n_1533, QN => n5992);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n6708, CK => CLK, RN => 
                           n12627, Q => n_1534, QN => n6309);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n6709, CK => CLK, RN => 
                           n12517, Q => n_1535, QN => n9159);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n6710, CK => CLK, RN => 
                           n12524, Q => n_1536, QN => n9191);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n6711, CK => CLK, RN => 
                           n12499, Q => n_1537, QN => n9255);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n6712, CK => CLK, RN => 
                           n12590, Q => n_1538, QN => n9589);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n6713, CK => CLK, RN => 
                           n12441, Q => n_1539, QN => n9621);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n6714, CK => CLK, RN => 
                           n12448, Q => n_1540, QN => n9653);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n6715, CK => CLK, RN => 
                           n12455, Q => n_1541, QN => n10015);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n6716, CK => CLK, RN => 
                           n12634, Q => n_1542, QN => n10047);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n6717, CK => CLK, RN => 
                           n12462, Q => n_1543, QN => n10079);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n6718, CK => CLK, RN => 
                           n12469, Q => n_1544, QN => n10111);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n6719, CK => CLK, RN => 
                           n12477, Q => n_1545, QN => n10143);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n6720, CK => CLK, RN => 
                           n12568, Q => n_1546, QN => n10175);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n6721, CK => CLK, RN => 
                           n12546, Q => n_1547, QN => n10209);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n6722, CK => CLK, RN => 
                           n12553, Q => n_1548, QN => n10241);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n6723, CK => CLK, RN => 
                           n12531, Q => n_1549, QN => n10273);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n6724, CK => CLK, RN => 
                           n12641, Q => n_1550, QN => n10308);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n6725, CK => CLK, RN => 
                           n12597, Q => n_1551, QN => n10340);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n6726, CK => CLK, RN => 
                           n12484, Q => n_1552, QN => n10372);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n6727, CK => CLK, RN => 
                           n12491, Q => n_1553, QN => n10407);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n6728, CK => CLK, RN => 
                           n12575, Q => n_1554, QN => n10439);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n6729, CK => CLK, RN => 
                           n12506, Q => n_1555, QN => n10471);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n6730, CK => CLK, RN => 
                           n12434, Q => n_1556, QN => n10503);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n6731, CK => CLK, RN => 
                           n12649, Q => n_1557, QN => n10535);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n6732, CK => CLK, RN => 
                           n12656, Q => n_1558, QN => n5734);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n6733, CK => CLK, RN => 
                           n12619, Q => n_1559, QN => n5766);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n6734, CK => CLK, RN => 
                           n12605, Q => n_1560, QN => n5798);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n6735, CK => CLK, RN => 
                           n12612, Q => n_1561, QN => n5830);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n6736, CK => CLK, RN => 
                           n12583, Q => n_1562, QN => n5862);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n6737, CK => CLK, RN => 
                           n12561, Q => n_1563, QN => n5894);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n6738, CK => CLK, RN => 
                           n12539, Q => n_1564, QN => n5926);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n6739, CK => CLK, RN => 
                           n12513, Q => n_1565, QN => n5990);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n6740, CK => CLK, RN => 
                           n12627, Q => n_1566, QN => n6307);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n6741, CK => CLK, RN => 
                           n12517, Q => n_1567, QN => n9157);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n6742, CK => CLK, RN => 
                           n12524, Q => n_1568, QN => n9189);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n6743, CK => CLK, RN => 
                           n12499, Q => n_1569, QN => n9253);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n6744, CK => CLK, RN => 
                           n12590, Q => n_1570, QN => n9587);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n6745, CK => CLK, RN => 
                           n12441, Q => n_1571, QN => n9619);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n6746, CK => CLK, RN => 
                           n12448, Q => n_1572, QN => n9651);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n6747, CK => CLK, RN => 
                           n12455, Q => n_1573, QN => n10013);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n6748, CK => CLK, RN => 
                           n12634, Q => n_1574, QN => n10045);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n6749, CK => CLK, RN => 
                           n12462, Q => n_1575, QN => n10077);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n6750, CK => CLK, RN => 
                           n12469, Q => n_1576, QN => n10109);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n6751, CK => CLK, RN => 
                           n12477, Q => n_1577, QN => n10141);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n6752, CK => CLK, RN => 
                           n12568, Q => n_1578, QN => n10173);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n6753, CK => CLK, RN => 
                           n12546, Q => n_1579, QN => n10205);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n6754, CK => CLK, RN => 
                           n12553, Q => n_1580, QN => n10239);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n6755, CK => CLK, RN => 
                           n12531, Q => n_1581, QN => n10271);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n6756, CK => CLK, RN => 
                           n12641, Q => n_1582, QN => n10306);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n6757, CK => CLK, RN => 
                           n12597, Q => n_1583, QN => n10338);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n6758, CK => CLK, RN => 
                           n12484, Q => n_1584, QN => n10370);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n6759, CK => CLK, RN => 
                           n12491, Q => n_1585, QN => n10405);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n6760, CK => CLK, RN => 
                           n12575, Q => n_1586, QN => n10437);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n6761, CK => CLK, RN => 
                           n12506, Q => n_1587, QN => n10469);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n6762, CK => CLK, RN => 
                           n12434, Q => n_1588, QN => n10501);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n6763, CK => CLK, RN => 
                           n12649, Q => n_1589, QN => n10533);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n6764, CK => CLK, RN => 
                           n12656, Q => n_1590, QN => n5735);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n6765, CK => CLK, RN => 
                           n12619, Q => n_1591, QN => n5767);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n6766, CK => CLK, RN => 
                           n12605, Q => n_1592, QN => n5799);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n6767, CK => CLK, RN => 
                           n12612, Q => n_1593, QN => n5831);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n6768, CK => CLK, RN => 
                           n12583, Q => n_1594, QN => n5863);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n6769, CK => CLK, RN => 
                           n12561, Q => n_1595, QN => n5895);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n6770, CK => CLK, RN => 
                           n12539, Q => n_1596, QN => n5927);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n6771, CK => CLK, RN => 
                           n12513, Q => n_1597, QN => n5991);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n6772, CK => CLK, RN => 
                           n12627, Q => n_1598, QN => n6308);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n6773, CK => CLK, RN => 
                           n12517, Q => n_1599, QN => n9158);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n6774, CK => CLK, RN => 
                           n12524, Q => n_1600, QN => n9190);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n6775, CK => CLK, RN => 
                           n12499, Q => n_1601, QN => n9254);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n6776, CK => CLK, RN => 
                           n12590, Q => n_1602, QN => n9588);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n6777, CK => CLK, RN => 
                           n12441, Q => n_1603, QN => n9620);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n6778, CK => CLK, RN => 
                           n12448, Q => n_1604, QN => n9652);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n6779, CK => CLK, RN => 
                           n12455, Q => n_1605, QN => n10014);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n6780, CK => CLK, RN => 
                           n12634, Q => n_1606, QN => n10046);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n6781, CK => CLK, RN => 
                           n12462, Q => n_1607, QN => n10078);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n6782, CK => CLK, RN => 
                           n12469, Q => n_1608, QN => n10110);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n6783, CK => CLK, RN => 
                           n12477, Q => n_1609, QN => n10142);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n6784, CK => CLK, RN => 
                           n12568, Q => n_1610, QN => n10174);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n6785, CK => CLK, RN => 
                           n12546, Q => n_1611, QN => n10208);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n6786, CK => CLK, RN => 
                           n12553, Q => n_1612, QN => n10240);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n6787, CK => CLK, RN => 
                           n12531, Q => n_1613, QN => n10272);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n6788, CK => CLK, RN => 
                           n12641, Q => n_1614, QN => n10307);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n6789, CK => CLK, RN => 
                           n12597, Q => n_1615, QN => n10339);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n6790, CK => CLK, RN => 
                           n12484, Q => n_1616, QN => n10371);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n6791, CK => CLK, RN => 
                           n12491, Q => n_1617, QN => n10406);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n6792, CK => CLK, RN => 
                           n12575, Q => n_1618, QN => n10438);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n6793, CK => CLK, RN => 
                           n12506, Q => n_1619, QN => n10470);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n6794, CK => CLK, RN => 
                           n12434, Q => n_1620, QN => n10502);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n6795, CK => CLK, RN => 
                           n12649, Q => n_1621, QN => n10534);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n7036, CK => CLK, RN => 
                           n12635, Q => n9999, QN => n13060);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n7037, CK => CLK, RN => 
                           n12463, Q => n9998, QN => n13061);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n7038, CK => CLK, RN => 
                           n12470, Q => n9997, QN => n13062);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n7039, CK => CLK, RN => 
                           n12477, Q => n9996, QN => n13063);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n7040, CK => CLK, RN => 
                           n12569, Q => n9995, QN => n13064);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n7041, CK => CLK, RN => 
                           n12547, Q => n9994, QN => n13065);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n7042, CK => CLK, RN => 
                           n12554, Q => n9993, QN => n13066);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n7043, CK => CLK, RN => 
                           n12532, Q => n9992, QN => n13067);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n7044, CK => CLK, RN => 
                           n12642, Q => n9991, QN => n13068);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n7045, CK => CLK, RN => 
                           n12598, Q => n9990, QN => n13069);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n7046, CK => CLK, RN => 
                           n12485, Q => n9989, QN => n13070);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n7047, CK => CLK, RN => 
                           n12492, Q => n9988, QN => n13071);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n7048, CK => CLK, RN => 
                           n12576, Q => n9987, QN => n13072);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n7049, CK => CLK, RN => 
                           n12507, Q => n9986, QN => n13073);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n7050, CK => CLK, RN => 
                           n12434, Q => n9985, QN => n13074);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n7051, CK => CLK, RN => 
                           n12649, Q => n9984, QN => n13075);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n7052, CK => CLK, RN => 
                           n12657, Q => n9983, QN => n13076);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n7053, CK => CLK, RN => 
                           n12620, Q => n9982, QN => n13077);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n7054, CK => CLK, RN => 
                           n12605, Q => n9981, QN => n13078);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n7055, CK => CLK, RN => 
                           n12613, Q => n9980, QN => n13079);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n7056, CK => CLK, RN => 
                           n12583, Q => n9979, QN => n13080);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n7057, CK => CLK, RN => 
                           n12561, Q => n9978, QN => n13081);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n7058, CK => CLK, RN => 
                           n12539, Q => n9977, QN => n13082);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n7059, CK => CLK, RN => 
                           n12514, Q => n9976, QN => n13083);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n7060, CK => CLK, RN => 
                           n12627, Q => n9975, QN => n13084);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n7061, CK => CLK, RN => 
                           n12517, Q => n9974, QN => n13085);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n7062, CK => CLK, RN => 
                           n12525, Q => n9973, QN => n13086);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n7063, CK => CLK, RN => 
                           n12499, Q => n9972, QN => n13087);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n7064, CK => CLK, RN => 
                           n12591, Q => n9971, QN => n13088);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n7065, CK => CLK, RN => 
                           n12442, Q => n9970, QN => n13089);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n7066, CK => CLK, RN => 
                           n12449, Q => n9969, QN => n13090);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n7067, CK => CLK, RN => 
                           n12455, Q => n9968, QN => n13091);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n7068, CK => CLK, RN => 
                           n12635, Q => n9967, QN => n13092);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n7069, CK => CLK, RN => 
                           n12463, Q => n9966, QN => n13093);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n7070, CK => CLK, RN => 
                           n12470, Q => n9965, QN => n13094);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n7071, CK => CLK, RN => 
                           n12477, Q => n9964, QN => n13095);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n7072, CK => CLK, RN => 
                           n12569, Q => n9963, QN => n13096);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n7073, CK => CLK, RN => 
                           n12547, Q => n9962, QN => n13097);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n7074, CK => CLK, RN => 
                           n12554, Q => n9961, QN => n13098);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n7075, CK => CLK, RN => 
                           n12532, Q => n9960, QN => n13099);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n7076, CK => CLK, RN => 
                           n12642, Q => n9959, QN => n13100);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n7077, CK => CLK, RN => 
                           n12598, Q => n9958, QN => n13101);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n7078, CK => CLK, RN => 
                           n12485, Q => n9957, QN => n13102);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n7079, CK => CLK, RN => 
                           n12492, Q => n9956, QN => n13103);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n7080, CK => CLK, RN => 
                           n12576, Q => n9955, QN => n13104);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n7081, CK => CLK, RN => 
                           n12507, Q => n9954, QN => n13105);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n7082, CK => CLK, RN => 
                           n12434, Q => n9953, QN => n13106);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n7083, CK => CLK, RN => 
                           n12649, Q => n9952, QN => n13107);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n7084, CK => CLK, RN => 
                           n12657, Q => n_1622, QN => n13108);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n7085, CK => CLK, RN => 
                           n12620, Q => n_1623, QN => n13109);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n7086, CK => CLK, RN => 
                           n12606, Q => n_1624, QN => n13110);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n7087, CK => CLK, RN => 
                           n12613, Q => n_1625, QN => n13111);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n7088, CK => CLK, RN => 
                           n12584, Q => n_1626, QN => n13112);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n7089, CK => CLK, RN => 
                           n12562, Q => n_1627, QN => n13113);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n7090, CK => CLK, RN => 
                           n12540, Q => n_1628, QN => n13114);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n7091, CK => CLK, RN => 
                           n12514, Q => n_1629, QN => n13115);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n7092, CK => CLK, RN => 
                           n12628, Q => n_1630, QN => n13116);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n7093, CK => CLK, RN => 
                           n12518, Q => n_1631, QN => n13117);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n7094, CK => CLK, RN => 
                           n12525, Q => n_1632, QN => n13118);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n7095, CK => CLK, RN => 
                           n12500, Q => n_1633, QN => n13119);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n7096, CK => CLK, RN => 
                           n12591, Q => n_1634, QN => n13120);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n7097, CK => CLK, RN => 
                           n12442, Q => n_1635, QN => n13121);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n7098, CK => CLK, RN => 
                           n12449, Q => n_1636, QN => n13122);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n7099, CK => CLK, RN => 
                           n12456, Q => n_1637, QN => n13123);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n7100, CK => CLK, RN => 
                           n12635, Q => n_1638, QN => n13124);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n7101, CK => CLK, RN => 
                           n12463, Q => n_1639, QN => n13125);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n7102, CK => CLK, RN => 
                           n12470, Q => n_1640, QN => n13126);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n7103, CK => CLK, RN => 
                           n12478, Q => n_1641, QN => n13127);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n7104, CK => CLK, RN => 
                           n12569, Q => n_1642, QN => n13128);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n7105, CK => CLK, RN => 
                           n12547, Q => n_1643, QN => n13129);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n7106, CK => CLK, RN => 
                           n12554, Q => n_1644, QN => n13130);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n7107, CK => CLK, RN => 
                           n12532, Q => n_1645, QN => n13131);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n7108, CK => CLK, RN => 
                           n12642, Q => n_1646, QN => n13132);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n7109, CK => CLK, RN => 
                           n12598, Q => n_1647, QN => n13133);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n7110, CK => CLK, RN => 
                           n12485, Q => n_1648, QN => n13134);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n7111, CK => CLK, RN => 
                           n12492, Q => n_1649, QN => n13135);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n7112, CK => CLK, RN => 
                           n12576, Q => n_1650, QN => n13136);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n7113, CK => CLK, RN => 
                           n12507, Q => n_1651, QN => n13137);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n7114, CK => CLK, RN => 
                           n12435, Q => n_1652, QN => n13138);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n7115, CK => CLK, RN => 
                           n12650, Q => n_1653, QN => n13139);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n7116, CK => CLK, RN => 
                           n12657, Q => n_1654, QN => n13140);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n7117, CK => CLK, RN => 
                           n12620, Q => n_1655, QN => n13141);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n7118, CK => CLK, RN => 
                           n12606, Q => n_1656, QN => n13142);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n7119, CK => CLK, RN => 
                           n12613, Q => n_1657, QN => n13143);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n7120, CK => CLK, RN => 
                           n12584, Q => n_1658, QN => n13144);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n7121, CK => CLK, RN => 
                           n12562, Q => n_1659, QN => n13145);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n7122, CK => CLK, RN => 
                           n12540, Q => n_1660, QN => n13146);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n7123, CK => CLK, RN => 
                           n12514, Q => n_1661, QN => n13147);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n7124, CK => CLK, RN => 
                           n12628, Q => n_1662, QN => n13148);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n7125, CK => CLK, RN => 
                           n12518, Q => n_1663, QN => n13149);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n7126, CK => CLK, RN => 
                           n12525, Q => n_1664, QN => n13150);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n7127, CK => CLK, RN => 
                           n12500, Q => n_1665, QN => n13151);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n7128, CK => CLK, RN => 
                           n12591, Q => n_1666, QN => n13152);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n7129, CK => CLK, RN => 
                           n12442, Q => n_1667, QN => n13153);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n7130, CK => CLK, RN => 
                           n12449, Q => n_1668, QN => n13154);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n7131, CK => CLK, RN => 
                           n12456, Q => n_1669, QN => n13155);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n7132, CK => CLK, RN => 
                           n12635, Q => n_1670, QN => n13156);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n7133, CK => CLK, RN => 
                           n12463, Q => n_1671, QN => n13157);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n7134, CK => CLK, RN => 
                           n12470, Q => n_1672, QN => n13158);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n7135, CK => CLK, RN => 
                           n12478, Q => n_1673, QN => n13159);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n7136, CK => CLK, RN => 
                           n12569, Q => n_1674, QN => n13160);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n7137, CK => CLK, RN => 
                           n12547, Q => n_1675, QN => n13161);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n7138, CK => CLK, RN => 
                           n12554, Q => n_1676, QN => n13162);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n7139, CK => CLK, RN => 
                           n12532, Q => n_1677, QN => n13163);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n7140, CK => CLK, RN => 
                           n12642, Q => n_1678, QN => n13164);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n7141, CK => CLK, RN => 
                           n12598, Q => n_1679, QN => n13165);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n7142, CK => CLK, RN => 
                           n12485, Q => n_1680, QN => n13166);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n7143, CK => CLK, RN => 
                           n12492, Q => n_1681, QN => n13167);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n7144, CK => CLK, RN => 
                           n12576, Q => n_1682, QN => n13168);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n7145, CK => CLK, RN => 
                           n12507, Q => n_1683, QN => n13169);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n7146, CK => CLK, RN => 
                           n12435, Q => n_1684, QN => n13170);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n7147, CK => CLK, RN => 
                           n12650, Q => n_1685, QN => n13171);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n7148, CK => CLK, RN => 
                           n12657, Q => n_1686, QN => n13172);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n7149, CK => CLK, RN => 
                           n12620, Q => n_1687, QN => n13173);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n7150, CK => CLK, RN => 
                           n12606, Q => n_1688, QN => n13174);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n7151, CK => CLK, RN => 
                           n12613, Q => n_1689, QN => n13175);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n7152, CK => CLK, RN => 
                           n12584, Q => n_1690, QN => n13176);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n7153, CK => CLK, RN => 
                           n12562, Q => n_1691, QN => n13177);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n7154, CK => CLK, RN => 
                           n12540, Q => n_1692, QN => n13178);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n7155, CK => CLK, RN => 
                           n12514, Q => n_1693, QN => n13179);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n7156, CK => CLK, RN => 
                           n12628, Q => n_1694, QN => n13180);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n7157, CK => CLK, RN => 
                           n12518, Q => n_1695, QN => n13181);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n7158, CK => CLK, RN => 
                           n12525, Q => n_1696, QN => n13182);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n7159, CK => CLK, RN => 
                           n12500, Q => n_1697, QN => n13183);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n7160, CK => CLK, RN => 
                           n12591, Q => n_1698, QN => n13184);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n7161, CK => CLK, RN => 
                           n12442, Q => n_1699, QN => n13185);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n7162, CK => CLK, RN => 
                           n12449, Q => n_1700, QN => n13186);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n7163, CK => CLK, RN => 
                           n12456, Q => n_1701, QN => n13187);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n7164, CK => CLK, RN => 
                           n12635, Q => n_1702, QN => n13188);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n7165, CK => CLK, RN => 
                           n12463, Q => n_1703, QN => n13189);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n7166, CK => CLK, RN => 
                           n12470, Q => n_1704, QN => n13190);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n7167, CK => CLK, RN => 
                           n12478, Q => n_1705, QN => n13191);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n7168, CK => CLK, RN => 
                           n12569, Q => n_1706, QN => n13192);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n7169, CK => CLK, RN => 
                           n12547, Q => n_1707, QN => n13193);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n7170, CK => CLK, RN => 
                           n12554, Q => n_1708, QN => n13194);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n7171, CK => CLK, RN => 
                           n12532, Q => n_1709, QN => n13195);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n7172, CK => CLK, RN => 
                           n12642, Q => n_1710, QN => n13196);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n7173, CK => CLK, RN => 
                           n12598, Q => n_1711, QN => n13197);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n7174, CK => CLK, RN => 
                           n12485, Q => n_1712, QN => n13198);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n7175, CK => CLK, RN => 
                           n12492, Q => n_1713, QN => n13199);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n7176, CK => CLK, RN => 
                           n12576, Q => n_1714, QN => n13200);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n7177, CK => CLK, RN => 
                           n12507, Q => n_1715, QN => n13201);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n7178, CK => CLK, RN => 
                           n12435, Q => n_1716, QN => n13202);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n7179, CK => CLK, RN => 
                           n12650, Q => n_1717, QN => n13203);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n7180, CK => CLK, RN => 
                           n12657, Q => n9855, QN => n13204);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n7181, CK => CLK, RN => 
                           n12620, Q => n9854, QN => n13205);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n7182, CK => CLK, RN => 
                           n12606, Q => n9853, QN => n13206);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n7183, CK => CLK, RN => 
                           n12613, Q => n9852, QN => n13207);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n7184, CK => CLK, RN => 
                           n12584, Q => n9851, QN => n13208);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n7185, CK => CLK, RN => 
                           n12562, Q => n9850, QN => n13209);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n7186, CK => CLK, RN => 
                           n12540, Q => n9849, QN => n13210);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n7187, CK => CLK, RN => 
                           n12514, Q => n9848, QN => n13211);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n7188, CK => CLK, RN => 
                           n12628, Q => n9847, QN => n13212);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n7189, CK => CLK, RN => 
                           n12518, Q => n9846, QN => n13213);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n7190, CK => CLK, RN => 
                           n12525, Q => n9845, QN => n13214);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n7191, CK => CLK, RN => 
                           n12500, Q => n9844, QN => n13215);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n7192, CK => CLK, RN => 
                           n12591, Q => n9843, QN => n13216);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n7193, CK => CLK, RN => 
                           n12442, Q => n9842, QN => n13217);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n7194, CK => CLK, RN => 
                           n12449, Q => n9841, QN => n13218);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n7195, CK => CLK, RN => 
                           n12456, Q => n9840, QN => n13219);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n7196, CK => CLK, RN => 
                           n12635, Q => n9839, QN => n13220);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n7197, CK => CLK, RN => 
                           n12463, Q => n9838, QN => n13221);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n7198, CK => CLK, RN => 
                           n12470, Q => n9837, QN => n13222);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n7199, CK => CLK, RN => 
                           n12478, Q => n9836, QN => n13223);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n7200, CK => CLK, RN => 
                           n12569, Q => n9835, QN => n13224);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n7201, CK => CLK, RN => 
                           n12547, Q => n9834, QN => n13225);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n7202, CK => CLK, RN => 
                           n12554, Q => n9833, QN => n13226);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n7203, CK => CLK, RN => 
                           n12532, Q => n9832, QN => n13227);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n7204, CK => CLK, RN => 
                           n12642, Q => n9831, QN => n13228);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n7205, CK => CLK, RN => 
                           n12598, Q => n9830, QN => n13229);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n7206, CK => CLK, RN => 
                           n12485, Q => n9829, QN => n13230);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n7207, CK => CLK, RN => 
                           n12492, Q => n9828, QN => n13231);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n7208, CK => CLK, RN => 
                           n12576, Q => n9827, QN => n13232);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n7209, CK => CLK, RN => 
                           n12507, Q => n9826, QN => n13233);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n7210, CK => CLK, RN => 
                           n12435, Q => n9825, QN => n13234);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n7211, CK => CLK, RN => 
                           n12650, Q => n9824, QN => n13235);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n7212, CK => CLK, RN => 
                           n12657, Q => n9823, QN => n13236);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n7213, CK => CLK, RN => 
                           n12621, Q => n9822, QN => n13237);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n7214, CK => CLK, RN => 
                           n12606, Q => n9821, QN => n13238);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n7215, CK => CLK, RN => 
                           n12613, Q => n9820, QN => n13239);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n7216, CK => CLK, RN => 
                           n12584, Q => n9819, QN => n13240);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n7217, CK => CLK, RN => 
                           n12562, Q => n9818, QN => n13241);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n7218, CK => CLK, RN => 
                           n12540, Q => n9817, QN => n13242);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n7219, CK => CLK, RN => 
                           n12515, Q => n9816, QN => n13243);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n7220, CK => CLK, RN => 
                           n12628, Q => n9815, QN => n13244);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n7221, CK => CLK, RN => 
                           n12518, Q => n9814, QN => n13245);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n7222, CK => CLK, RN => 
                           n12525, Q => n9813, QN => n13246);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n7223, CK => CLK, RN => 
                           n12500, Q => n9812, QN => n13247);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n7224, CK => CLK, RN => 
                           n12591, Q => n9811, QN => n13248);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n7225, CK => CLK, RN => 
                           n12442, Q => n9810, QN => n13249);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n7226, CK => CLK, RN => 
                           n12450, Q => n9809, QN => n13250);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n7227, CK => CLK, RN => 
                           n12456, Q => n9808, QN => n13251);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n7228, CK => CLK, RN => 
                           n12635, Q => n9807, QN => n13252);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n7229, CK => CLK, RN => 
                           n12463, Q => n9806, QN => n13253);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n7230, CK => CLK, RN => 
                           n12471, Q => n9805, QN => n13254);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n7231, CK => CLK, RN => 
                           n12478, Q => n9804, QN => n13255);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n7232, CK => CLK, RN => 
                           n12569, Q => n9803, QN => n13256);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n7233, CK => CLK, RN => 
                           n12547, Q => n9802, QN => n13257);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n7234, CK => CLK, RN => 
                           n12555, Q => n9801, QN => n13258);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n7235, CK => CLK, RN => 
                           n12533, Q => n9800, QN => n13259);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n7236, CK => CLK, RN => 
                           n12643, Q => n9799, QN => n13260);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n7237, CK => CLK, RN => 
                           n12599, Q => n9798, QN => n13261);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n7238, CK => CLK, RN => 
                           n12485, Q => n9797, QN => n13262);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n7239, CK => CLK, RN => 
                           n12493, Q => n9796, QN => n13263);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n7240, CK => CLK, RN => 
                           n12577, Q => n9795, QN => n13264);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n7241, CK => CLK, RN => 
                           n12507, Q => n9794, QN => n13265);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n7242, CK => CLK, RN => 
                           n12435, Q => n9793, QN => n13266);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n7243, CK => CLK, RN => 
                           n12650, Q => n9792, QN => n13267);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n7244, CK => CLK, RN => 
                           n12657, Q => n9791, QN => n13268);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n7245, CK => CLK, RN => 
                           n12621, Q => n9790, QN => n13269);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n7246, CK => CLK, RN => 
                           n12606, Q => n9789, QN => n13270);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n7247, CK => CLK, RN => 
                           n12613, Q => n9788, QN => n13271);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n7248, CK => CLK, RN => 
                           n12584, Q => n9787, QN => n13272);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n7249, CK => CLK, RN => 
                           n12562, Q => n9786, QN => n13273);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n7250, CK => CLK, RN => 
                           n12540, Q => n9785, QN => n13274);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n7251, CK => CLK, RN => 
                           n12515, Q => n9784, QN => n13275);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n7252, CK => CLK, RN => 
                           n12628, Q => n9783, QN => n13276);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n7253, CK => CLK, RN => 
                           n12518, Q => n9782, QN => n13277);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n7254, CK => CLK, RN => 
                           n12525, Q => n9781, QN => n13278);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n7255, CK => CLK, RN => 
                           n12500, Q => n9780, QN => n13279);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n7256, CK => CLK, RN => 
                           n12591, Q => n9779, QN => n13280);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n7257, CK => CLK, RN => 
                           n12442, Q => n9778, QN => n13281);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n7258, CK => CLK, RN => 
                           n12450, Q => n9777, QN => n13282);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n7259, CK => CLK, RN => 
                           n12456, Q => n9776, QN => n13283);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n7260, CK => CLK, RN => 
                           n12635, Q => n9775, QN => n13284);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n7261, CK => CLK, RN => 
                           n12463, Q => n9774, QN => n13285);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n7262, CK => CLK, RN => 
                           n12471, Q => n9773, QN => n13286);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n7263, CK => CLK, RN => 
                           n12478, Q => n9772, QN => n13287);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n7264, CK => CLK, RN => 
                           n12569, Q => n9771, QN => n13288);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n7265, CK => CLK, RN => 
                           n12547, Q => n9770, QN => n13289);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n7266, CK => CLK, RN => 
                           n12555, Q => n9769, QN => n13290);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n7267, CK => CLK, RN => 
                           n12533, Q => n9768, QN => n13291);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n7268, CK => CLK, RN => 
                           n12643, Q => n9767, QN => n13292);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n7269, CK => CLK, RN => 
                           n12599, Q => n9766, QN => n13293);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n7270, CK => CLK, RN => 
                           n12485, Q => n9765, QN => n13294);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n7271, CK => CLK, RN => 
                           n12493, Q => n9764, QN => n13295);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n7272, CK => CLK, RN => 
                           n12577, Q => n9763, QN => n13296);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n7273, CK => CLK, RN => 
                           n12507, Q => n9762, QN => n13297);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n7274, CK => CLK, RN => 
                           n12435, Q => n9761, QN => n13298);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n7275, CK => CLK, RN => 
                           n12650, Q => n9760, QN => n13299);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n7276, CK => CLK, RN => 
                           n12657, Q => n9759, QN => n13300);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n7277, CK => CLK, RN => 
                           n12621, Q => n9758, QN => n13301);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n7278, CK => CLK, RN => 
                           n12606, Q => n9757, QN => n13302);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n7279, CK => CLK, RN => 
                           n12613, Q => n9756, QN => n13303);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n7280, CK => CLK, RN => 
                           n12584, Q => n9755, QN => n13304);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n7281, CK => CLK, RN => 
                           n12562, Q => n9754, QN => n13305);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n7282, CK => CLK, RN => 
                           n12540, Q => n9753, QN => n13306);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n7283, CK => CLK, RN => 
                           n12515, Q => n9752, QN => n13307);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n7284, CK => CLK, RN => 
                           n12628, Q => n9751, QN => n13308);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n7285, CK => CLK, RN => 
                           n12518, Q => n9750, QN => n13309);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n7286, CK => CLK, RN => 
                           n12525, Q => n9749, QN => n13310);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n7287, CK => CLK, RN => 
                           n12500, Q => n9748, QN => n13311);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n7288, CK => CLK, RN => 
                           n12591, Q => n9747, QN => n13312);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n7289, CK => CLK, RN => 
                           n12442, Q => n9746, QN => n13313);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n7290, CK => CLK, RN => 
                           n12450, Q => n9745, QN => n13314);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n7291, CK => CLK, RN => 
                           n12456, Q => n9744, QN => n13315);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n7292, CK => CLK, RN => 
                           n12635, Q => n9743, QN => n13316);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n7293, CK => CLK, RN => 
                           n12463, Q => n9742, QN => n13317);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n7294, CK => CLK, RN => 
                           n12471, Q => n9741, QN => n13318);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n7295, CK => CLK, RN => 
                           n12478, Q => n9740, QN => n13319);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n7296, CK => CLK, RN => 
                           n12569, Q => n9739, QN => n13320);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n7297, CK => CLK, RN => 
                           n12547, Q => n9738, QN => n13321);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n7298, CK => CLK, RN => 
                           n12555, Q => n9737, QN => n13322);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n7299, CK => CLK, RN => 
                           n12533, Q => n9736, QN => n13323);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n7300, CK => CLK, RN => 
                           n12643, Q => n9735, QN => n13324);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n7301, CK => CLK, RN => 
                           n12599, Q => n9734, QN => n13325);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n7302, CK => CLK, RN => 
                           n12485, Q => n9733, QN => n13326);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n7303, CK => CLK, RN => 
                           n12493, Q => n9732, QN => n13327);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n7304, CK => CLK, RN => 
                           n12577, Q => n9731, QN => n13328);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n7305, CK => CLK, RN => 
                           n12507, Q => n9730, QN => n13329);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n7306, CK => CLK, RN => 
                           n12435, Q => n9729, QN => n13330);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n7307, CK => CLK, RN => 
                           n12650, Q => n9728, QN => n13331);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n7308, CK => CLK, RN => 
                           n12657, Q => n9727, QN => n13332);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n7309, CK => CLK, RN => 
                           n12621, Q => n9726, QN => n13333);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n7310, CK => CLK, RN => 
                           n12606, Q => n9725, QN => n13334);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n7311, CK => CLK, RN => 
                           n12613, Q => n9724, QN => n13335);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n7312, CK => CLK, RN => 
                           n12584, Q => n9723, QN => n13336);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n7313, CK => CLK, RN => 
                           n12562, Q => n9722, QN => n13337);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n7314, CK => CLK, RN => 
                           n12540, Q => n9721, QN => n13338);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n7315, CK => CLK, RN => 
                           n12515, Q => n9720, QN => n13339);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n7316, CK => CLK, RN => 
                           n12628, Q => n9719, QN => n13340);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n7317, CK => CLK, RN => 
                           n12518, Q => n9718, QN => n13341);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n7318, CK => CLK, RN => 
                           n12525, Q => n9717, QN => n13342);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n7319, CK => CLK, RN => 
                           n12500, Q => n9716, QN => n13343);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n7320, CK => CLK, RN => 
                           n12591, Q => n9715, QN => n13344);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n7321, CK => CLK, RN => 
                           n12442, Q => n9714, QN => n13345);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n7322, CK => CLK, RN => 
                           n12450, Q => n9713, QN => n13346);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n7323, CK => CLK, RN => 
                           n12456, Q => n9712, QN => n13347);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n7324, CK => CLK, RN => 
                           n12635, Q => n9711, QN => n13348);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n7325, CK => CLK, RN => 
                           n12463, Q => n9710, QN => n13349);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n7326, CK => CLK, RN => 
                           n12471, Q => n9709, QN => n13350);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n7327, CK => CLK, RN => 
                           n12478, Q => n9708, QN => n13351);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n7328, CK => CLK, RN => 
                           n12569, Q => n9707, QN => n13352);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n7329, CK => CLK, RN => 
                           n12547, Q => n9706, QN => n13353);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n7330, CK => CLK, RN => 
                           n12555, Q => n9705, QN => n13354);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n7331, CK => CLK, RN => 
                           n12533, Q => n9704, QN => n13355);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n7332, CK => CLK, RN => 
                           n12643, Q => n9703, QN => n13356);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n7333, CK => CLK, RN => 
                           n12599, Q => n9702, QN => n13357);
   REGISTERS_reg_32_31_inst : DFFR_X1 port map( D => n7340, CK => CLK, RN => 
                           n12658, Q => n9695, QN => n13364);
   REGISTERS_reg_32_30_inst : DFFR_X1 port map( D => n7341, CK => CLK, RN => 
                           n12621, Q => n9694, QN => n13365);
   REGISTERS_reg_32_29_inst : DFFR_X1 port map( D => n7342, CK => CLK, RN => 
                           n12606, Q => n9693, QN => n13366);
   REGISTERS_reg_32_28_inst : DFFR_X1 port map( D => n7343, CK => CLK, RN => 
                           n12614, Q => n9692, QN => n13367);
   REGISTERS_reg_32_27_inst : DFFR_X1 port map( D => n7344, CK => CLK, RN => 
                           n12584, Q => n9691, QN => n13368);
   REGISTERS_reg_32_26_inst : DFFR_X1 port map( D => n7345, CK => CLK, RN => 
                           n12562, Q => n9690, QN => n13369);
   REGISTERS_reg_32_25_inst : DFFR_X1 port map( D => n7346, CK => CLK, RN => 
                           n12540, Q => n9689, QN => n13370);
   REGISTERS_reg_32_24_inst : DFFR_X1 port map( D => n7347, CK => CLK, RN => 
                           n12515, Q => n9688, QN => n13371);
   REGISTERS_reg_32_23_inst : DFFR_X1 port map( D => n7348, CK => CLK, RN => 
                           n12628, Q => n9687, QN => n13372);
   REGISTERS_reg_32_22_inst : DFFR_X1 port map( D => n7349, CK => CLK, RN => 
                           n12518, Q => n9686, QN => n13373);
   REGISTERS_reg_32_21_inst : DFFR_X1 port map( D => n7350, CK => CLK, RN => 
                           n12526, Q => n9685, QN => n13374);
   REGISTERS_reg_32_20_inst : DFFR_X1 port map( D => n7351, CK => CLK, RN => 
                           n12500, Q => n9684, QN => n13375);
   REGISTERS_reg_32_19_inst : DFFR_X1 port map( D => n7352, CK => CLK, RN => 
                           n12592, Q => n9683, QN => n13376);
   REGISTERS_reg_32_18_inst : DFFR_X1 port map( D => n7353, CK => CLK, RN => 
                           n12443, Q => n9682, QN => n13377);
   REGISTERS_reg_32_17_inst : DFFR_X1 port map( D => n7354, CK => CLK, RN => 
                           n12450, Q => n9681, QN => n13378);
   REGISTERS_reg_32_16_inst : DFFR_X1 port map( D => n7355, CK => CLK, RN => 
                           n12456, Q => n9680, QN => n13379);
   REGISTERS_reg_32_15_inst : DFFR_X1 port map( D => n7356, CK => CLK, RN => 
                           n12636, Q => n9679, QN => n13380);
   REGISTERS_reg_32_14_inst : DFFR_X1 port map( D => n7357, CK => CLK, RN => 
                           n12464, Q => n9678, QN => n13381);
   REGISTERS_reg_32_13_inst : DFFR_X1 port map( D => n7358, CK => CLK, RN => 
                           n12471, Q => n9677, QN => n13382);
   REGISTERS_reg_32_12_inst : DFFR_X1 port map( D => n7359, CK => CLK, RN => 
                           n12478, Q => n9676, QN => n13383);
   REGISTERS_reg_32_11_inst : DFFR_X1 port map( D => n7360, CK => CLK, RN => 
                           n12570, Q => n9675, QN => n13384);
   REGISTERS_reg_32_10_inst : DFFR_X1 port map( D => n7361, CK => CLK, RN => 
                           n12548, Q => n9674, QN => n13385);
   REGISTERS_reg_32_9_inst : DFFR_X1 port map( D => n7362, CK => CLK, RN => 
                           n12555, Q => n9673, QN => n13386);
   REGISTERS_reg_32_8_inst : DFFR_X1 port map( D => n7363, CK => CLK, RN => 
                           n12533, Q => n9672, QN => n13387);
   REGISTERS_reg_32_7_inst : DFFR_X1 port map( D => n7364, CK => CLK, RN => 
                           n12643, Q => n9671, QN => n13388);
   REGISTERS_reg_32_6_inst : DFFR_X1 port map( D => n7365, CK => CLK, RN => 
                           n12599, Q => n9670, QN => n13389);
   REGISTERS_reg_32_5_inst : DFFR_X1 port map( D => n7366, CK => CLK, RN => 
                           n12486, Q => n9669, QN => n13390);
   REGISTERS_reg_32_4_inst : DFFR_X1 port map( D => n7367, CK => CLK, RN => 
                           n12493, Q => n9668, QN => n13391);
   REGISTERS_reg_32_3_inst : DFFR_X1 port map( D => n7368, CK => CLK, RN => 
                           n12577, Q => n9667, QN => n13392);
   REGISTERS_reg_32_2_inst : DFFR_X1 port map( D => n7369, CK => CLK, RN => 
                           n12508, Q => n9666, QN => n13393);
   REGISTERS_reg_32_1_inst : DFFR_X1 port map( D => n7370, CK => CLK, RN => 
                           n12435, Q => n9665, QN => n13394);
   REGISTERS_reg_32_0_inst : DFFR_X1 port map( D => n7371, CK => CLK, RN => 
                           n12650, Q => n9664, QN => n13395);
   REGISTERS_reg_33_31_inst : DFFR_X1 port map( D => n7372, CK => CLK, RN => 
                           n12658, Q => n_1718, QN => n5729);
   REGISTERS_reg_33_30_inst : DFFR_X1 port map( D => n7373, CK => CLK, RN => 
                           n12621, Q => n_1719, QN => n5761);
   REGISTERS_reg_33_29_inst : DFFR_X1 port map( D => n7374, CK => CLK, RN => 
                           n12606, Q => n_1720, QN => n5793);
   REGISTERS_reg_33_28_inst : DFFR_X1 port map( D => n7375, CK => CLK, RN => 
                           n12614, Q => n_1721, QN => n5825);
   REGISTERS_reg_33_27_inst : DFFR_X1 port map( D => n7376, CK => CLK, RN => 
                           n12584, Q => n_1722, QN => n5857);
   REGISTERS_reg_33_26_inst : DFFR_X1 port map( D => n7377, CK => CLK, RN => 
                           n12562, Q => n_1723, QN => n5889);
   REGISTERS_reg_33_25_inst : DFFR_X1 port map( D => n7378, CK => CLK, RN => 
                           n12540, Q => n_1724, QN => n5921);
   REGISTERS_reg_33_24_inst : DFFR_X1 port map( D => n7379, CK => CLK, RN => 
                           n12515, Q => n_1725, QN => n5985);
   REGISTERS_reg_33_23_inst : DFFR_X1 port map( D => n7380, CK => CLK, RN => 
                           n12628, Q => n_1726, QN => n6302);
   REGISTERS_reg_33_22_inst : DFFR_X1 port map( D => n7381, CK => CLK, RN => 
                           n12518, Q => n_1727, QN => n9152);
   REGISTERS_reg_33_21_inst : DFFR_X1 port map( D => n7382, CK => CLK, RN => 
                           n12526, Q => n_1728, QN => n9184);
   REGISTERS_reg_33_20_inst : DFFR_X1 port map( D => n7383, CK => CLK, RN => 
                           n12500, Q => n_1729, QN => n9248);
   REGISTERS_reg_33_19_inst : DFFR_X1 port map( D => n7384, CK => CLK, RN => 
                           n12592, Q => n_1730, QN => n9582);
   REGISTERS_reg_33_18_inst : DFFR_X1 port map( D => n7385, CK => CLK, RN => 
                           n12443, Q => n_1731, QN => n9614);
   REGISTERS_reg_33_17_inst : DFFR_X1 port map( D => n7386, CK => CLK, RN => 
                           n12450, Q => n_1732, QN => n9646);
   REGISTERS_reg_33_16_inst : DFFR_X1 port map( D => n7387, CK => CLK, RN => 
                           n12456, Q => n_1733, QN => n10008);
   REGISTERS_reg_33_15_inst : DFFR_X1 port map( D => n7388, CK => CLK, RN => 
                           n12636, Q => n_1734, QN => n10040);
   REGISTERS_reg_33_14_inst : DFFR_X1 port map( D => n7389, CK => CLK, RN => 
                           n12464, Q => n_1735, QN => n10072);
   REGISTERS_reg_33_13_inst : DFFR_X1 port map( D => n7390, CK => CLK, RN => 
                           n12471, Q => n_1736, QN => n10104);
   REGISTERS_reg_33_12_inst : DFFR_X1 port map( D => n7391, CK => CLK, RN => 
                           n12478, Q => n_1737, QN => n10136);
   REGISTERS_reg_33_11_inst : DFFR_X1 port map( D => n7392, CK => CLK, RN => 
                           n12570, Q => n_1738, QN => n10168);
   REGISTERS_reg_33_10_inst : DFFR_X1 port map( D => n7393, CK => CLK, RN => 
                           n12548, Q => n_1739, QN => n10200);
   REGISTERS_reg_33_9_inst : DFFR_X1 port map( D => n7394, CK => CLK, RN => 
                           n12555, Q => n_1740, QN => n10234);
   REGISTERS_reg_33_8_inst : DFFR_X1 port map( D => n7395, CK => CLK, RN => 
                           n12533, Q => n_1741, QN => n10266);
   REGISTERS_reg_33_7_inst : DFFR_X1 port map( D => n7396, CK => CLK, RN => 
                           n12643, Q => n_1742, QN => n10298);
   REGISTERS_reg_33_6_inst : DFFR_X1 port map( D => n7397, CK => CLK, RN => 
                           n12599, Q => n_1743, QN => n10333);
   REGISTERS_reg_33_5_inst : DFFR_X1 port map( D => n7398, CK => CLK, RN => 
                           n12486, Q => n_1744, QN => n10365);
   REGISTERS_reg_33_4_inst : DFFR_X1 port map( D => n7399, CK => CLK, RN => 
                           n12493, Q => n_1745, QN => n10400);
   REGISTERS_reg_33_3_inst : DFFR_X1 port map( D => n7400, CK => CLK, RN => 
                           n12577, Q => n_1746, QN => n10432);
   REGISTERS_reg_33_2_inst : DFFR_X1 port map( D => n7401, CK => CLK, RN => 
                           n12508, Q => n_1747, QN => n10464);
   REGISTERS_reg_33_1_inst : DFFR_X1 port map( D => n7402, CK => CLK, RN => 
                           n12435, Q => n_1748, QN => n10496);
   REGISTERS_reg_33_0_inst : DFFR_X1 port map( D => n7403, CK => CLK, RN => 
                           n12650, Q => n_1749, QN => n10528);
   REGISTERS_reg_34_31_inst : DFFR_X1 port map( D => n7404, CK => CLK, RN => 
                           n12658, Q => n_1750, QN => n5728);
   REGISTERS_reg_34_30_inst : DFFR_X1 port map( D => n7405, CK => CLK, RN => 
                           n12621, Q => n_1751, QN => n5760);
   REGISTERS_reg_34_29_inst : DFFR_X1 port map( D => n7406, CK => CLK, RN => 
                           n12606, Q => n_1752, QN => n5792);
   REGISTERS_reg_34_28_inst : DFFR_X1 port map( D => n7407, CK => CLK, RN => 
                           n12614, Q => n_1753, QN => n5824);
   REGISTERS_reg_34_27_inst : DFFR_X1 port map( D => n7408, CK => CLK, RN => 
                           n12584, Q => n_1754, QN => n5856);
   REGISTERS_reg_34_26_inst : DFFR_X1 port map( D => n7409, CK => CLK, RN => 
                           n12562, Q => n_1755, QN => n5888);
   REGISTERS_reg_34_25_inst : DFFR_X1 port map( D => n7410, CK => CLK, RN => 
                           n12540, Q => n_1756, QN => n5920);
   REGISTERS_reg_34_24_inst : DFFR_X1 port map( D => n7411, CK => CLK, RN => 
                           n12515, Q => n_1757, QN => n5984);
   REGISTERS_reg_34_23_inst : DFFR_X1 port map( D => n7412, CK => CLK, RN => 
                           n12628, Q => n_1758, QN => n6301);
   REGISTERS_reg_34_22_inst : DFFR_X1 port map( D => n7413, CK => CLK, RN => 
                           n12518, Q => n_1759, QN => n9151);
   REGISTERS_reg_34_21_inst : DFFR_X1 port map( D => n7414, CK => CLK, RN => 
                           n12526, Q => n_1760, QN => n9183);
   REGISTERS_reg_34_20_inst : DFFR_X1 port map( D => n7415, CK => CLK, RN => 
                           n12500, Q => n_1761, QN => n9215);
   REGISTERS_reg_34_19_inst : DFFR_X1 port map( D => n7416, CK => CLK, RN => 
                           n12592, Q => n_1762, QN => n9581);
   REGISTERS_reg_34_18_inst : DFFR_X1 port map( D => n7417, CK => CLK, RN => 
                           n12443, Q => n_1763, QN => n9613);
   REGISTERS_reg_34_17_inst : DFFR_X1 port map( D => n7418, CK => CLK, RN => 
                           n12450, Q => n_1764, QN => n9645);
   REGISTERS_reg_34_16_inst : DFFR_X1 port map( D => n7419, CK => CLK, RN => 
                           n12456, Q => n_1765, QN => n10007);
   REGISTERS_reg_34_15_inst : DFFR_X1 port map( D => n7420, CK => CLK, RN => 
                           n12636, Q => n_1766, QN => n10039);
   REGISTERS_reg_34_14_inst : DFFR_X1 port map( D => n7421, CK => CLK, RN => 
                           n12464, Q => n_1767, QN => n10071);
   REGISTERS_reg_34_13_inst : DFFR_X1 port map( D => n7422, CK => CLK, RN => 
                           n12471, Q => n_1768, QN => n10103);
   REGISTERS_reg_34_12_inst : DFFR_X1 port map( D => n7423, CK => CLK, RN => 
                           n12478, Q => n_1769, QN => n10135);
   REGISTERS_reg_34_11_inst : DFFR_X1 port map( D => n7424, CK => CLK, RN => 
                           n12570, Q => n_1770, QN => n10167);
   REGISTERS_reg_34_10_inst : DFFR_X1 port map( D => n7425, CK => CLK, RN => 
                           n12548, Q => n_1771, QN => n10199);
   REGISTERS_reg_34_9_inst : DFFR_X1 port map( D => n7426, CK => CLK, RN => 
                           n12555, Q => n_1772, QN => n10233);
   REGISTERS_reg_34_8_inst : DFFR_X1 port map( D => n7427, CK => CLK, RN => 
                           n12533, Q => n_1773, QN => n10265);
   REGISTERS_reg_34_7_inst : DFFR_X1 port map( D => n7428, CK => CLK, RN => 
                           n12643, Q => n_1774, QN => n10297);
   REGISTERS_reg_34_6_inst : DFFR_X1 port map( D => n7429, CK => CLK, RN => 
                           n12599, Q => n_1775, QN => n10332);
   REGISTERS_reg_34_5_inst : DFFR_X1 port map( D => n7430, CK => CLK, RN => 
                           n12486, Q => n_1776, QN => n10364);
   REGISTERS_reg_34_4_inst : DFFR_X1 port map( D => n7431, CK => CLK, RN => 
                           n12493, Q => n_1777, QN => n10396);
   REGISTERS_reg_34_3_inst : DFFR_X1 port map( D => n7432, CK => CLK, RN => 
                           n12577, Q => n_1778, QN => n10431);
   REGISTERS_reg_34_2_inst : DFFR_X1 port map( D => n7433, CK => CLK, RN => 
                           n12508, Q => n_1779, QN => n10463);
   REGISTERS_reg_34_1_inst : DFFR_X1 port map( D => n7434, CK => CLK, RN => 
                           n12435, Q => n_1780, QN => n10495);
   REGISTERS_reg_34_0_inst : DFFR_X1 port map( D => n7435, CK => CLK, RN => 
                           n12650, Q => n_1781, QN => n10527);
   REGISTERS_reg_35_31_inst : DFFR_X1 port map( D => n7436, CK => CLK, RN => 
                           n12658, Q => n_1782, QN => n5726);
   REGISTERS_reg_35_30_inst : DFFR_X1 port map( D => n7437, CK => CLK, RN => 
                           n12621, Q => n_1783, QN => n5758);
   REGISTERS_reg_35_29_inst : DFFR_X1 port map( D => n7438, CK => CLK, RN => 
                           n12606, Q => n_1784, QN => n5790);
   REGISTERS_reg_35_28_inst : DFFR_X1 port map( D => n7439, CK => CLK, RN => 
                           n12614, Q => n_1785, QN => n5822);
   REGISTERS_reg_35_27_inst : DFFR_X1 port map( D => n7440, CK => CLK, RN => 
                           n12584, Q => n_1786, QN => n5854);
   REGISTERS_reg_35_26_inst : DFFR_X1 port map( D => n7441, CK => CLK, RN => 
                           n12562, Q => n_1787, QN => n5886);
   REGISTERS_reg_35_25_inst : DFFR_X1 port map( D => n7442, CK => CLK, RN => 
                           n12540, Q => n_1788, QN => n5918);
   REGISTERS_reg_35_24_inst : DFFR_X1 port map( D => n7443, CK => CLK, RN => 
                           n12515, Q => n_1789, QN => n5982);
   REGISTERS_reg_35_23_inst : DFFR_X1 port map( D => n7444, CK => CLK, RN => 
                           n12628, Q => n_1790, QN => n6140);
   REGISTERS_reg_35_22_inst : DFFR_X1 port map( D => n7445, CK => CLK, RN => 
                           n12518, Q => n_1791, QN => n9149);
   REGISTERS_reg_35_21_inst : DFFR_X1 port map( D => n7446, CK => CLK, RN => 
                           n12526, Q => n_1792, QN => n9181);
   REGISTERS_reg_35_20_inst : DFFR_X1 port map( D => n7447, CK => CLK, RN => 
                           n12500, Q => n_1793, QN => n9213);
   REGISTERS_reg_35_19_inst : DFFR_X1 port map( D => n7448, CK => CLK, RN => 
                           n12592, Q => n_1794, QN => n9579);
   REGISTERS_reg_35_18_inst : DFFR_X1 port map( D => n7449, CK => CLK, RN => 
                           n12443, Q => n_1795, QN => n9611);
   REGISTERS_reg_35_17_inst : DFFR_X1 port map( D => n7450, CK => CLK, RN => 
                           n12450, Q => n_1796, QN => n9643);
   REGISTERS_reg_35_16_inst : DFFR_X1 port map( D => n7451, CK => CLK, RN => 
                           n12456, Q => n_1797, QN => n10005);
   REGISTERS_reg_35_15_inst : DFFR_X1 port map( D => n7452, CK => CLK, RN => 
                           n12636, Q => n_1798, QN => n10037);
   REGISTERS_reg_35_14_inst : DFFR_X1 port map( D => n7453, CK => CLK, RN => 
                           n12464, Q => n_1799, QN => n10069);
   REGISTERS_reg_35_13_inst : DFFR_X1 port map( D => n7454, CK => CLK, RN => 
                           n12471, Q => n_1800, QN => n10101);
   REGISTERS_reg_35_12_inst : DFFR_X1 port map( D => n7455, CK => CLK, RN => 
                           n12478, Q => n_1801, QN => n10133);
   REGISTERS_reg_35_11_inst : DFFR_X1 port map( D => n7456, CK => CLK, RN => 
                           n12570, Q => n_1802, QN => n10165);
   REGISTERS_reg_35_10_inst : DFFR_X1 port map( D => n7457, CK => CLK, RN => 
                           n12548, Q => n_1803, QN => n10197);
   REGISTERS_reg_35_9_inst : DFFR_X1 port map( D => n7458, CK => CLK, RN => 
                           n12555, Q => n_1804, QN => n10231);
   REGISTERS_reg_35_8_inst : DFFR_X1 port map( D => n7459, CK => CLK, RN => 
                           n12533, Q => n_1805, QN => n10263);
   REGISTERS_reg_35_7_inst : DFFR_X1 port map( D => n7460, CK => CLK, RN => 
                           n12643, Q => n_1806, QN => n10295);
   REGISTERS_reg_35_6_inst : DFFR_X1 port map( D => n7461, CK => CLK, RN => 
                           n12599, Q => n_1807, QN => n10330);
   REGISTERS_reg_35_5_inst : DFFR_X1 port map( D => n7462, CK => CLK, RN => 
                           n12486, Q => n_1808, QN => n10362);
   REGISTERS_reg_35_4_inst : DFFR_X1 port map( D => n7463, CK => CLK, RN => 
                           n12493, Q => n_1809, QN => n10394);
   REGISTERS_reg_35_3_inst : DFFR_X1 port map( D => n7464, CK => CLK, RN => 
                           n12577, Q => n_1810, QN => n10429);
   REGISTERS_reg_35_2_inst : DFFR_X1 port map( D => n7465, CK => CLK, RN => 
                           n12508, Q => n_1811, QN => n10461);
   REGISTERS_reg_35_1_inst : DFFR_X1 port map( D => n7466, CK => CLK, RN => 
                           n12435, Q => n_1812, QN => n10493);
   REGISTERS_reg_35_0_inst : DFFR_X1 port map( D => n7467, CK => CLK, RN => 
                           n12650, Q => n_1813, QN => n10525);
   REGISTERS_reg_36_31_inst : DFFR_X1 port map( D => n7468, CK => CLK, RN => 
                           n12658, Q => n_1814, QN => n5727);
   REGISTERS_reg_36_30_inst : DFFR_X1 port map( D => n7469, CK => CLK, RN => 
                           n12621, Q => n_1815, QN => n5759);
   REGISTERS_reg_36_29_inst : DFFR_X1 port map( D => n7470, CK => CLK, RN => 
                           n12607, Q => n_1816, QN => n5791);
   REGISTERS_reg_36_28_inst : DFFR_X1 port map( D => n7471, CK => CLK, RN => 
                           n12614, Q => n_1817, QN => n5823);
   REGISTERS_reg_36_27_inst : DFFR_X1 port map( D => n7472, CK => CLK, RN => 
                           n12585, Q => n_1818, QN => n5855);
   REGISTERS_reg_36_26_inst : DFFR_X1 port map( D => n7473, CK => CLK, RN => 
                           n12563, Q => n_1819, QN => n5887);
   REGISTERS_reg_36_25_inst : DFFR_X1 port map( D => n7474, CK => CLK, RN => 
                           n12541, Q => n_1820, QN => n5919);
   REGISTERS_reg_36_24_inst : DFFR_X1 port map( D => n7475, CK => CLK, RN => 
                           n12515, Q => n_1821, QN => n5983);
   REGISTERS_reg_36_23_inst : DFFR_X1 port map( D => n7476, CK => CLK, RN => 
                           n12629, Q => n_1822, QN => n6236);
   REGISTERS_reg_36_22_inst : DFFR_X1 port map( D => n7477, CK => CLK, RN => 
                           n12519, Q => n_1823, QN => n9150);
   REGISTERS_reg_36_21_inst : DFFR_X1 port map( D => n7478, CK => CLK, RN => 
                           n12526, Q => n_1824, QN => n9182);
   REGISTERS_reg_36_20_inst : DFFR_X1 port map( D => n7479, CK => CLK, RN => 
                           n12501, Q => n_1825, QN => n9214);
   REGISTERS_reg_36_19_inst : DFFR_X1 port map( D => n7480, CK => CLK, RN => 
                           n12592, Q => n_1826, QN => n9580);
   REGISTERS_reg_36_18_inst : DFFR_X1 port map( D => n7481, CK => CLK, RN => 
                           n12443, Q => n_1827, QN => n9612);
   REGISTERS_reg_36_17_inst : DFFR_X1 port map( D => n7482, CK => CLK, RN => 
                           n12450, Q => n_1828, QN => n9644);
   REGISTERS_reg_36_16_inst : DFFR_X1 port map( D => n7483, CK => CLK, RN => 
                           n12457, Q => n_1829, QN => n10006);
   REGISTERS_reg_36_15_inst : DFFR_X1 port map( D => n7484, CK => CLK, RN => 
                           n12636, Q => n_1830, QN => n10038);
   REGISTERS_reg_36_14_inst : DFFR_X1 port map( D => n7485, CK => CLK, RN => 
                           n12464, Q => n_1831, QN => n10070);
   REGISTERS_reg_36_13_inst : DFFR_X1 port map( D => n7486, CK => CLK, RN => 
                           n12471, Q => n_1832, QN => n10102);
   REGISTERS_reg_36_12_inst : DFFR_X1 port map( D => n7487, CK => CLK, RN => 
                           n12479, Q => n_1833, QN => n10134);
   REGISTERS_reg_36_11_inst : DFFR_X1 port map( D => n7488, CK => CLK, RN => 
                           n12570, Q => n_1834, QN => n10166);
   REGISTERS_reg_36_10_inst : DFFR_X1 port map( D => n7489, CK => CLK, RN => 
                           n12548, Q => n_1835, QN => n10198);
   REGISTERS_reg_36_9_inst : DFFR_X1 port map( D => n7490, CK => CLK, RN => 
                           n12555, Q => n_1836, QN => n10232);
   REGISTERS_reg_36_8_inst : DFFR_X1 port map( D => n7491, CK => CLK, RN => 
                           n12533, Q => n_1837, QN => n10264);
   REGISTERS_reg_36_7_inst : DFFR_X1 port map( D => n7492, CK => CLK, RN => 
                           n12643, Q => n_1838, QN => n10296);
   REGISTERS_reg_36_6_inst : DFFR_X1 port map( D => n7493, CK => CLK, RN => 
                           n12599, Q => n_1839, QN => n10331);
   REGISTERS_reg_36_5_inst : DFFR_X1 port map( D => n7494, CK => CLK, RN => 
                           n12486, Q => n_1840, QN => n10363);
   REGISTERS_reg_36_4_inst : DFFR_X1 port map( D => n7495, CK => CLK, RN => 
                           n12493, Q => n_1841, QN => n10395);
   REGISTERS_reg_36_3_inst : DFFR_X1 port map( D => n7496, CK => CLK, RN => 
                           n12577, Q => n_1842, QN => n10430);
   REGISTERS_reg_36_2_inst : DFFR_X1 port map( D => n7497, CK => CLK, RN => 
                           n12508, Q => n_1843, QN => n10462);
   REGISTERS_reg_36_1_inst : DFFR_X1 port map( D => n7498, CK => CLK, RN => 
                           n12436, Q => n_1844, QN => n10494);
   REGISTERS_reg_36_0_inst : DFFR_X1 port map( D => n7499, CK => CLK, RN => 
                           n12651, Q => n_1845, QN => n10526);
   REGISTERS_reg_37_31_inst : DFFR_X1 port map( D => n7500, CK => CLK, RN => 
                           n12658, Q => n_1846, QN => n5725);
   REGISTERS_reg_37_30_inst : DFFR_X1 port map( D => n7501, CK => CLK, RN => 
                           n12621, Q => n_1847, QN => n5757);
   REGISTERS_reg_37_29_inst : DFFR_X1 port map( D => n7502, CK => CLK, RN => 
                           n12607, Q => n_1848, QN => n5789);
   REGISTERS_reg_37_28_inst : DFFR_X1 port map( D => n7503, CK => CLK, RN => 
                           n12614, Q => n_1849, QN => n5821);
   REGISTERS_reg_37_27_inst : DFFR_X1 port map( D => n7504, CK => CLK, RN => 
                           n12585, Q => n_1850, QN => n5853);
   REGISTERS_reg_37_26_inst : DFFR_X1 port map( D => n7505, CK => CLK, RN => 
                           n12563, Q => n_1851, QN => n5885);
   REGISTERS_reg_37_25_inst : DFFR_X1 port map( D => n7506, CK => CLK, RN => 
                           n12541, Q => n_1852, QN => n5917);
   REGISTERS_reg_37_24_inst : DFFR_X1 port map( D => n7507, CK => CLK, RN => 
                           n12515, Q => n_1853, QN => n5981);
   REGISTERS_reg_37_23_inst : DFFR_X1 port map( D => n7508, CK => CLK, RN => 
                           n12629, Q => n_1854, QN => n6044);
   REGISTERS_reg_37_22_inst : DFFR_X1 port map( D => n7509, CK => CLK, RN => 
                           n12519, Q => n_1855, QN => n9148);
   REGISTERS_reg_37_21_inst : DFFR_X1 port map( D => n7510, CK => CLK, RN => 
                           n12526, Q => n_1856, QN => n9180);
   REGISTERS_reg_37_20_inst : DFFR_X1 port map( D => n7511, CK => CLK, RN => 
                           n12501, Q => n_1857, QN => n9212);
   REGISTERS_reg_37_19_inst : DFFR_X1 port map( D => n7512, CK => CLK, RN => 
                           n12592, Q => n_1858, QN => n9578);
   REGISTERS_reg_37_18_inst : DFFR_X1 port map( D => n7513, CK => CLK, RN => 
                           n12443, Q => n_1859, QN => n9610);
   REGISTERS_reg_37_17_inst : DFFR_X1 port map( D => n7514, CK => CLK, RN => 
                           n12450, Q => n_1860, QN => n9642);
   REGISTERS_reg_37_16_inst : DFFR_X1 port map( D => n7515, CK => CLK, RN => 
                           n12457, Q => n_1861, QN => n10004);
   REGISTERS_reg_37_15_inst : DFFR_X1 port map( D => n7516, CK => CLK, RN => 
                           n12636, Q => n_1862, QN => n10036);
   REGISTERS_reg_37_14_inst : DFFR_X1 port map( D => n7517, CK => CLK, RN => 
                           n12464, Q => n_1863, QN => n10068);
   REGISTERS_reg_37_13_inst : DFFR_X1 port map( D => n7518, CK => CLK, RN => 
                           n12471, Q => n_1864, QN => n10100);
   REGISTERS_reg_37_12_inst : DFFR_X1 port map( D => n7519, CK => CLK, RN => 
                           n12479, Q => n_1865, QN => n10132);
   REGISTERS_reg_37_11_inst : DFFR_X1 port map( D => n7520, CK => CLK, RN => 
                           n12570, Q => n_1866, QN => n10164);
   REGISTERS_reg_37_10_inst : DFFR_X1 port map( D => n7521, CK => CLK, RN => 
                           n12548, Q => n_1867, QN => n10196);
   REGISTERS_reg_37_9_inst : DFFR_X1 port map( D => n7522, CK => CLK, RN => 
                           n12555, Q => n_1868, QN => n10230);
   REGISTERS_reg_37_8_inst : DFFR_X1 port map( D => n7523, CK => CLK, RN => 
                           n12533, Q => n_1869, QN => n10262);
   REGISTERS_reg_37_7_inst : DFFR_X1 port map( D => n7524, CK => CLK, RN => 
                           n12643, Q => n_1870, QN => n10294);
   REGISTERS_reg_37_6_inst : DFFR_X1 port map( D => n7525, CK => CLK, RN => 
                           n12599, Q => n_1871, QN => n10329);
   REGISTERS_reg_37_5_inst : DFFR_X1 port map( D => n7526, CK => CLK, RN => 
                           n12486, Q => n_1872, QN => n10361);
   REGISTERS_reg_37_4_inst : DFFR_X1 port map( D => n7527, CK => CLK, RN => 
                           n12493, Q => n_1873, QN => n10393);
   REGISTERS_reg_37_3_inst : DFFR_X1 port map( D => n7528, CK => CLK, RN => 
                           n12577, Q => n_1874, QN => n10428);
   REGISTERS_reg_37_2_inst : DFFR_X1 port map( D => n7529, CK => CLK, RN => 
                           n12508, Q => n_1875, QN => n10460);
   REGISTERS_reg_37_1_inst : DFFR_X1 port map( D => n7530, CK => CLK, RN => 
                           n12436, Q => n_1876, QN => n10492);
   REGISTERS_reg_37_0_inst : DFFR_X1 port map( D => n7531, CK => CLK, RN => 
                           n12651, Q => n_1877, QN => n10524);
   REGISTERS_reg_38_31_inst : DFFR_X1 port map( D => n7532, CK => CLK, RN => 
                           n12658, Q => n_1878, QN => n5723);
   REGISTERS_reg_38_30_inst : DFFR_X1 port map( D => n7533, CK => CLK, RN => 
                           n12621, Q => n_1879, QN => n5755);
   REGISTERS_reg_38_29_inst : DFFR_X1 port map( D => n7534, CK => CLK, RN => 
                           n12607, Q => n_1880, QN => n5787);
   REGISTERS_reg_38_28_inst : DFFR_X1 port map( D => n7535, CK => CLK, RN => 
                           n12614, Q => n_1881, QN => n5819);
   REGISTERS_reg_38_27_inst : DFFR_X1 port map( D => n7536, CK => CLK, RN => 
                           n12585, Q => n_1882, QN => n5851);
   REGISTERS_reg_38_26_inst : DFFR_X1 port map( D => n7537, CK => CLK, RN => 
                           n12563, Q => n_1883, QN => n5883);
   REGISTERS_reg_38_25_inst : DFFR_X1 port map( D => n7538, CK => CLK, RN => 
                           n12541, Q => n_1884, QN => n5915);
   REGISTERS_reg_38_24_inst : DFFR_X1 port map( D => n7539, CK => CLK, RN => 
                           n12515, Q => n_1885, QN => n5947);
   REGISTERS_reg_38_23_inst : DFFR_X1 port map( D => n7540, CK => CLK, RN => 
                           n12629, Q => n_1886, QN => n6011);
   REGISTERS_reg_38_22_inst : DFFR_X1 port map( D => n7541, CK => CLK, RN => 
                           n12519, Q => n_1887, QN => n9146);
   REGISTERS_reg_38_21_inst : DFFR_X1 port map( D => n7542, CK => CLK, RN => 
                           n12526, Q => n_1888, QN => n9178);
   REGISTERS_reg_38_20_inst : DFFR_X1 port map( D => n7543, CK => CLK, RN => 
                           n12501, Q => n_1889, QN => n9210);
   REGISTERS_reg_38_19_inst : DFFR_X1 port map( D => n7544, CK => CLK, RN => 
                           n12592, Q => n_1890, QN => n9576);
   REGISTERS_reg_38_18_inst : DFFR_X1 port map( D => n7545, CK => CLK, RN => 
                           n12443, Q => n_1891, QN => n9608);
   REGISTERS_reg_38_17_inst : DFFR_X1 port map( D => n7546, CK => CLK, RN => 
                           n12450, Q => n_1892, QN => n9640);
   REGISTERS_reg_38_16_inst : DFFR_X1 port map( D => n7547, CK => CLK, RN => 
                           n12457, Q => n_1893, QN => n10002);
   REGISTERS_reg_38_15_inst : DFFR_X1 port map( D => n7548, CK => CLK, RN => 
                           n12636, Q => n_1894, QN => n10034);
   REGISTERS_reg_38_14_inst : DFFR_X1 port map( D => n7549, CK => CLK, RN => 
                           n12464, Q => n_1895, QN => n10066);
   REGISTERS_reg_38_13_inst : DFFR_X1 port map( D => n7550, CK => CLK, RN => 
                           n12471, Q => n_1896, QN => n10098);
   REGISTERS_reg_38_12_inst : DFFR_X1 port map( D => n7551, CK => CLK, RN => 
                           n12479, Q => n_1897, QN => n10130);
   REGISTERS_reg_38_11_inst : DFFR_X1 port map( D => n7552, CK => CLK, RN => 
                           n12570, Q => n_1898, QN => n10162);
   REGISTERS_reg_38_10_inst : DFFR_X1 port map( D => n7553, CK => CLK, RN => 
                           n12548, Q => n_1899, QN => n10194);
   REGISTERS_reg_38_9_inst : DFFR_X1 port map( D => n7554, CK => CLK, RN => 
                           n12555, Q => n_1900, QN => n10228);
   REGISTERS_reg_38_8_inst : DFFR_X1 port map( D => n7555, CK => CLK, RN => 
                           n12533, Q => n_1901, QN => n10260);
   REGISTERS_reg_38_7_inst : DFFR_X1 port map( D => n7556, CK => CLK, RN => 
                           n12643, Q => n_1902, QN => n10292);
   REGISTERS_reg_38_6_inst : DFFR_X1 port map( D => n7557, CK => CLK, RN => 
                           n12599, Q => n_1903, QN => n10327);
   REGISTERS_reg_38_5_inst : DFFR_X1 port map( D => n7558, CK => CLK, RN => 
                           n12486, Q => n_1904, QN => n10359);
   REGISTERS_reg_38_4_inst : DFFR_X1 port map( D => n7559, CK => CLK, RN => 
                           n12493, Q => n_1905, QN => n10391);
   REGISTERS_reg_38_3_inst : DFFR_X1 port map( D => n7560, CK => CLK, RN => 
                           n12577, Q => n_1906, QN => n10426);
   REGISTERS_reg_38_2_inst : DFFR_X1 port map( D => n7561, CK => CLK, RN => 
                           n12508, Q => n_1907, QN => n10458);
   REGISTERS_reg_38_1_inst : DFFR_X1 port map( D => n7562, CK => CLK, RN => 
                           n12436, Q => n_1908, QN => n10490);
   REGISTERS_reg_38_0_inst : DFFR_X1 port map( D => n7563, CK => CLK, RN => 
                           n12651, Q => n_1909, QN => n10522);
   REGISTERS_reg_39_31_inst : DFFR_X1 port map( D => n7564, CK => CLK, RN => 
                           n12658, Q => n_1910, QN => n13396);
   REGISTERS_reg_39_30_inst : DFFR_X1 port map( D => n7565, CK => CLK, RN => 
                           n12621, Q => n_1911, QN => n13397);
   REGISTERS_reg_39_29_inst : DFFR_X1 port map( D => n7566, CK => CLK, RN => 
                           n12607, Q => n_1912, QN => n13398);
   REGISTERS_reg_39_28_inst : DFFR_X1 port map( D => n7567, CK => CLK, RN => 
                           n12614, Q => n_1913, QN => n13399);
   REGISTERS_reg_39_27_inst : DFFR_X1 port map( D => n7568, CK => CLK, RN => 
                           n12585, Q => n_1914, QN => n13400);
   REGISTERS_reg_39_26_inst : DFFR_X1 port map( D => n7569, CK => CLK, RN => 
                           n12563, Q => n_1915, QN => n13401);
   REGISTERS_reg_39_25_inst : DFFR_X1 port map( D => n7570, CK => CLK, RN => 
                           n12541, Q => n_1916, QN => n13402);
   REGISTERS_reg_39_24_inst : DFFR_X1 port map( D => n7571, CK => CLK, RN => 
                           n12515, Q => n_1917, QN => n13403);
   REGISTERS_reg_39_23_inst : DFFR_X1 port map( D => n7572, CK => CLK, RN => 
                           n12629, Q => n_1918, QN => n13404);
   REGISTERS_reg_39_22_inst : DFFR_X1 port map( D => n7573, CK => CLK, RN => 
                           n12519, Q => n_1919, QN => n13405);
   REGISTERS_reg_39_21_inst : DFFR_X1 port map( D => n7574, CK => CLK, RN => 
                           n12526, Q => n_1920, QN => n13406);
   REGISTERS_reg_39_20_inst : DFFR_X1 port map( D => n7575, CK => CLK, RN => 
                           n12501, Q => n_1921, QN => n13407);
   REGISTERS_reg_39_19_inst : DFFR_X1 port map( D => n7576, CK => CLK, RN => 
                           n12592, Q => n_1922, QN => n13408);
   REGISTERS_reg_39_18_inst : DFFR_X1 port map( D => n7577, CK => CLK, RN => 
                           n12443, Q => n_1923, QN => n13409);
   REGISTERS_reg_39_17_inst : DFFR_X1 port map( D => n7578, CK => CLK, RN => 
                           n12450, Q => n_1924, QN => n13410);
   REGISTERS_reg_39_16_inst : DFFR_X1 port map( D => n7579, CK => CLK, RN => 
                           n12457, Q => n_1925, QN => n13411);
   REGISTERS_reg_39_15_inst : DFFR_X1 port map( D => n7580, CK => CLK, RN => 
                           n12636, Q => n_1926, QN => n13412);
   REGISTERS_reg_39_14_inst : DFFR_X1 port map( D => n7581, CK => CLK, RN => 
                           n12464, Q => n_1927, QN => n13413);
   REGISTERS_reg_39_13_inst : DFFR_X1 port map( D => n7582, CK => CLK, RN => 
                           n12471, Q => n_1928, QN => n13414);
   REGISTERS_reg_39_12_inst : DFFR_X1 port map( D => n7583, CK => CLK, RN => 
                           n12479, Q => n_1929, QN => n13415);
   REGISTERS_reg_39_11_inst : DFFR_X1 port map( D => n7584, CK => CLK, RN => 
                           n12570, Q => n_1930, QN => n13416);
   REGISTERS_reg_39_10_inst : DFFR_X1 port map( D => n7585, CK => CLK, RN => 
                           n12548, Q => n_1931, QN => n13417);
   REGISTERS_reg_39_9_inst : DFFR_X1 port map( D => n7586, CK => CLK, RN => 
                           n12555, Q => n_1932, QN => n13418);
   REGISTERS_reg_39_8_inst : DFFR_X1 port map( D => n7587, CK => CLK, RN => 
                           n12533, Q => n_1933, QN => n13419);
   REGISTERS_reg_39_7_inst : DFFR_X1 port map( D => n7588, CK => CLK, RN => 
                           n12643, Q => n_1934, QN => n13420);
   REGISTERS_reg_39_6_inst : DFFR_X1 port map( D => n7589, CK => CLK, RN => 
                           n12599, Q => n_1935, QN => n13421);
   REGISTERS_reg_39_5_inst : DFFR_X1 port map( D => n7590, CK => CLK, RN => 
                           n12486, Q => n_1936, QN => n13422);
   REGISTERS_reg_39_4_inst : DFFR_X1 port map( D => n7591, CK => CLK, RN => 
                           n12493, Q => n_1937, QN => n13423);
   REGISTERS_reg_39_3_inst : DFFR_X1 port map( D => n7592, CK => CLK, RN => 
                           n12577, Q => n_1938, QN => n13424);
   REGISTERS_reg_39_2_inst : DFFR_X1 port map( D => n7593, CK => CLK, RN => 
                           n12508, Q => n_1939, QN => n13425);
   REGISTERS_reg_39_1_inst : DFFR_X1 port map( D => n7594, CK => CLK, RN => 
                           n12436, Q => n_1940, QN => n13426);
   REGISTERS_reg_39_0_inst : DFFR_X1 port map( D => n7595, CK => CLK, RN => 
                           n12651, Q => n_1941, QN => n13427);
   REGISTERS_reg_40_31_inst : DFFR_X1 port map( D => n7596, CK => CLK, RN => 
                           n12658, Q => n_1942, QN => n5724);
   REGISTERS_reg_40_30_inst : DFFR_X1 port map( D => n7597, CK => CLK, RN => 
                           n12622, Q => n_1943, QN => n5756);
   REGISTERS_reg_40_29_inst : DFFR_X1 port map( D => n7598, CK => CLK, RN => 
                           n12607, Q => n_1944, QN => n5788);
   REGISTERS_reg_40_28_inst : DFFR_X1 port map( D => n7599, CK => CLK, RN => 
                           n12614, Q => n_1945, QN => n5820);
   REGISTERS_reg_40_27_inst : DFFR_X1 port map( D => n7600, CK => CLK, RN => 
                           n12585, Q => n_1946, QN => n5852);
   REGISTERS_reg_40_26_inst : DFFR_X1 port map( D => n7601, CK => CLK, RN => 
                           n12563, Q => n_1947, QN => n5884);
   REGISTERS_reg_40_25_inst : DFFR_X1 port map( D => n7602, CK => CLK, RN => 
                           n12541, Q => n_1948, QN => n5916);
   REGISTERS_reg_40_24_inst : DFFR_X1 port map( D => n7603, CK => CLK, RN => 
                           n12516, Q => n_1949, QN => n5948);
   REGISTERS_reg_40_23_inst : DFFR_X1 port map( D => n7604, CK => CLK, RN => 
                           n12629, Q => n_1950, QN => n6012);
   REGISTERS_reg_40_22_inst : DFFR_X1 port map( D => n7605, CK => CLK, RN => 
                           n12519, Q => n_1951, QN => n9147);
   REGISTERS_reg_40_21_inst : DFFR_X1 port map( D => n7606, CK => CLK, RN => 
                           n12526, Q => n_1952, QN => n9179);
   REGISTERS_reg_40_20_inst : DFFR_X1 port map( D => n7607, CK => CLK, RN => 
                           n12501, Q => n_1953, QN => n9211);
   REGISTERS_reg_40_19_inst : DFFR_X1 port map( D => n7608, CK => CLK, RN => 
                           n12592, Q => n_1954, QN => n9577);
   REGISTERS_reg_40_18_inst : DFFR_X1 port map( D => n7609, CK => CLK, RN => 
                           n12443, Q => n_1955, QN => n9609);
   REGISTERS_reg_40_17_inst : DFFR_X1 port map( D => n7610, CK => CLK, RN => 
                           n12451, Q => n_1956, QN => n9641);
   REGISTERS_reg_40_16_inst : DFFR_X1 port map( D => n7611, CK => CLK, RN => 
                           n12457, Q => n_1957, QN => n10003);
   REGISTERS_reg_40_15_inst : DFFR_X1 port map( D => n7612, CK => CLK, RN => 
                           n12636, Q => n_1958, QN => n10035);
   REGISTERS_reg_40_14_inst : DFFR_X1 port map( D => n7613, CK => CLK, RN => 
                           n12464, Q => n_1959, QN => n10067);
   REGISTERS_reg_40_13_inst : DFFR_X1 port map( D => n7614, CK => CLK, RN => 
                           n12472, Q => n_1960, QN => n10099);
   REGISTERS_reg_40_12_inst : DFFR_X1 port map( D => n7615, CK => CLK, RN => 
                           n12479, Q => n_1961, QN => n10131);
   REGISTERS_reg_40_11_inst : DFFR_X1 port map( D => n7616, CK => CLK, RN => 
                           n12570, Q => n_1962, QN => n10163);
   REGISTERS_reg_40_10_inst : DFFR_X1 port map( D => n7617, CK => CLK, RN => 
                           n12548, Q => n_1963, QN => n10195);
   REGISTERS_reg_40_9_inst : DFFR_X1 port map( D => n7618, CK => CLK, RN => 
                           n12556, Q => n_1964, QN => n10229);
   REGISTERS_reg_40_8_inst : DFFR_X1 port map( D => n7619, CK => CLK, RN => 
                           n12534, Q => n_1965, QN => n10261);
   REGISTERS_reg_40_7_inst : DFFR_X1 port map( D => n7620, CK => CLK, RN => 
                           n12644, Q => n_1966, QN => n10293);
   REGISTERS_reg_40_6_inst : DFFR_X1 port map( D => n7621, CK => CLK, RN => 
                           n12600, Q => n_1967, QN => n10328);
   REGISTERS_reg_40_5_inst : DFFR_X1 port map( D => n7622, CK => CLK, RN => 
                           n12486, Q => n_1968, QN => n10360);
   REGISTERS_reg_40_4_inst : DFFR_X1 port map( D => n7623, CK => CLK, RN => 
                           n12494, Q => n_1969, QN => n10392);
   REGISTERS_reg_40_3_inst : DFFR_X1 port map( D => n7624, CK => CLK, RN => 
                           n12578, Q => n_1970, QN => n10427);
   REGISTERS_reg_40_2_inst : DFFR_X1 port map( D => n7625, CK => CLK, RN => 
                           n12508, Q => n_1971, QN => n10459);
   REGISTERS_reg_40_1_inst : DFFR_X1 port map( D => n7626, CK => CLK, RN => 
                           n12436, Q => n_1972, QN => n10491);
   REGISTERS_reg_40_0_inst : DFFR_X1 port map( D => n7627, CK => CLK, RN => 
                           n12651, Q => n_1973, QN => n10523);
   REGISTERS_reg_41_31_inst : DFFR_X1 port map( D => n7628, CK => CLK, RN => 
                           n12658, Q => n_1974, QN => n13428);
   REGISTERS_reg_41_30_inst : DFFR_X1 port map( D => n7629, CK => CLK, RN => 
                           n12622, Q => n_1975, QN => n13429);
   REGISTERS_reg_41_29_inst : DFFR_X1 port map( D => n7630, CK => CLK, RN => 
                           n12607, Q => n_1976, QN => n13430);
   REGISTERS_reg_41_28_inst : DFFR_X1 port map( D => n7631, CK => CLK, RN => 
                           n12614, Q => n_1977, QN => n13431);
   REGISTERS_reg_41_27_inst : DFFR_X1 port map( D => n7632, CK => CLK, RN => 
                           n12585, Q => n_1978, QN => n13432);
   REGISTERS_reg_41_26_inst : DFFR_X1 port map( D => n7633, CK => CLK, RN => 
                           n12563, Q => n_1979, QN => n13433);
   REGISTERS_reg_41_25_inst : DFFR_X1 port map( D => n7634, CK => CLK, RN => 
                           n12541, Q => n_1980, QN => n13434);
   REGISTERS_reg_41_24_inst : DFFR_X1 port map( D => n7635, CK => CLK, RN => 
                           n12516, Q => n_1981, QN => n13435);
   REGISTERS_reg_41_23_inst : DFFR_X1 port map( D => n7636, CK => CLK, RN => 
                           n12629, Q => n_1982, QN => n13436);
   REGISTERS_reg_41_22_inst : DFFR_X1 port map( D => n7637, CK => CLK, RN => 
                           n12519, Q => n_1983, QN => n13437);
   REGISTERS_reg_41_21_inst : DFFR_X1 port map( D => n7638, CK => CLK, RN => 
                           n12526, Q => n_1984, QN => n13438);
   REGISTERS_reg_41_20_inst : DFFR_X1 port map( D => n7639, CK => CLK, RN => 
                           n12501, Q => n_1985, QN => n13439);
   REGISTERS_reg_41_19_inst : DFFR_X1 port map( D => n7640, CK => CLK, RN => 
                           n12592, Q => n_1986, QN => n13440);
   REGISTERS_reg_41_18_inst : DFFR_X1 port map( D => n7641, CK => CLK, RN => 
                           n12443, Q => n_1987, QN => n13441);
   REGISTERS_reg_41_17_inst : DFFR_X1 port map( D => n7642, CK => CLK, RN => 
                           n12451, Q => n_1988, QN => n13442);
   REGISTERS_reg_41_16_inst : DFFR_X1 port map( D => n7643, CK => CLK, RN => 
                           n12457, Q => n_1989, QN => n13443);
   REGISTERS_reg_41_15_inst : DFFR_X1 port map( D => n7644, CK => CLK, RN => 
                           n12636, Q => n_1990, QN => n13444);
   REGISTERS_reg_41_14_inst : DFFR_X1 port map( D => n7645, CK => CLK, RN => 
                           n12464, Q => n_1991, QN => n13445);
   REGISTERS_reg_41_13_inst : DFFR_X1 port map( D => n7646, CK => CLK, RN => 
                           n12472, Q => n_1992, QN => n13446);
   REGISTERS_reg_41_12_inst : DFFR_X1 port map( D => n7647, CK => CLK, RN => 
                           n12479, Q => n_1993, QN => n13447);
   REGISTERS_reg_41_11_inst : DFFR_X1 port map( D => n7648, CK => CLK, RN => 
                           n12570, Q => n_1994, QN => n13448);
   REGISTERS_reg_41_10_inst : DFFR_X1 port map( D => n7649, CK => CLK, RN => 
                           n12548, Q => n_1995, QN => n13449);
   REGISTERS_reg_41_9_inst : DFFR_X1 port map( D => n7650, CK => CLK, RN => 
                           n12556, Q => n_1996, QN => n13450);
   REGISTERS_reg_41_8_inst : DFFR_X1 port map( D => n7651, CK => CLK, RN => 
                           n12534, Q => n_1997, QN => n13451);
   REGISTERS_reg_41_7_inst : DFFR_X1 port map( D => n7652, CK => CLK, RN => 
                           n12644, Q => n_1998, QN => n13452);
   REGISTERS_reg_41_6_inst : DFFR_X1 port map( D => n7653, CK => CLK, RN => 
                           n12600, Q => n_1999, QN => n13453);
   REGISTERS_reg_41_5_inst : DFFR_X1 port map( D => n7654, CK => CLK, RN => 
                           n12486, Q => n_2000, QN => n13454);
   REGISTERS_reg_41_4_inst : DFFR_X1 port map( D => n7655, CK => CLK, RN => 
                           n12494, Q => n_2001, QN => n13455);
   REGISTERS_reg_41_3_inst : DFFR_X1 port map( D => n7656, CK => CLK, RN => 
                           n12578, Q => n_2002, QN => n13456);
   REGISTERS_reg_41_2_inst : DFFR_X1 port map( D => n7657, CK => CLK, RN => 
                           n12508, Q => n_2003, QN => n13457);
   REGISTERS_reg_41_1_inst : DFFR_X1 port map( D => n7658, CK => CLK, RN => 
                           n12436, Q => n_2004, QN => n13458);
   REGISTERS_reg_41_0_inst : DFFR_X1 port map( D => n7659, CK => CLK, RN => 
                           n12651, Q => n_2005, QN => n13459);
   REGISTERS_reg_42_31_inst : DFFR_X1 port map( D => n7660, CK => CLK, RN => 
                           n12658, Q => n_2006, QN => n5730);
   REGISTERS_reg_42_30_inst : DFFR_X1 port map( D => n7661, CK => CLK, RN => 
                           n12622, Q => n_2007, QN => n5762);
   REGISTERS_reg_42_29_inst : DFFR_X1 port map( D => n7662, CK => CLK, RN => 
                           n12607, Q => n_2008, QN => n5794);
   REGISTERS_reg_42_28_inst : DFFR_X1 port map( D => n7663, CK => CLK, RN => 
                           n12614, Q => n_2009, QN => n5826);
   REGISTERS_reg_42_27_inst : DFFR_X1 port map( D => n7664, CK => CLK, RN => 
                           n12585, Q => n_2010, QN => n5858);
   REGISTERS_reg_42_26_inst : DFFR_X1 port map( D => n7665, CK => CLK, RN => 
                           n12563, Q => n_2011, QN => n5890);
   REGISTERS_reg_42_25_inst : DFFR_X1 port map( D => n7666, CK => CLK, RN => 
                           n12541, Q => n_2012, QN => n5922);
   REGISTERS_reg_42_24_inst : DFFR_X1 port map( D => n7667, CK => CLK, RN => 
                           n12516, Q => n_2013, QN => n5986);
   REGISTERS_reg_42_23_inst : DFFR_X1 port map( D => n7668, CK => CLK, RN => 
                           n12629, Q => n_2014, QN => n6303);
   REGISTERS_reg_42_22_inst : DFFR_X1 port map( D => n7669, CK => CLK, RN => 
                           n12519, Q => n_2015, QN => n9153);
   REGISTERS_reg_42_21_inst : DFFR_X1 port map( D => n7670, CK => CLK, RN => 
                           n12526, Q => n_2016, QN => n9185);
   REGISTERS_reg_42_20_inst : DFFR_X1 port map( D => n7671, CK => CLK, RN => 
                           n12501, Q => n_2017, QN => n9249);
   REGISTERS_reg_42_19_inst : DFFR_X1 port map( D => n7672, CK => CLK, RN => 
                           n12592, Q => n_2018, QN => n9583);
   REGISTERS_reg_42_18_inst : DFFR_X1 port map( D => n7673, CK => CLK, RN => 
                           n12443, Q => n_2019, QN => n9615);
   REGISTERS_reg_42_17_inst : DFFR_X1 port map( D => n7674, CK => CLK, RN => 
                           n12451, Q => n_2020, QN => n9647);
   REGISTERS_reg_42_16_inst : DFFR_X1 port map( D => n7675, CK => CLK, RN => 
                           n12457, Q => n_2021, QN => n10009);
   REGISTERS_reg_42_15_inst : DFFR_X1 port map( D => n7676, CK => CLK, RN => 
                           n12636, Q => n_2022, QN => n10041);
   REGISTERS_reg_42_14_inst : DFFR_X1 port map( D => n7677, CK => CLK, RN => 
                           n12464, Q => n_2023, QN => n10073);
   REGISTERS_reg_42_13_inst : DFFR_X1 port map( D => n7678, CK => CLK, RN => 
                           n12472, Q => n_2024, QN => n10105);
   REGISTERS_reg_42_12_inst : DFFR_X1 port map( D => n7679, CK => CLK, RN => 
                           n12479, Q => n_2025, QN => n10137);
   REGISTERS_reg_42_11_inst : DFFR_X1 port map( D => n7680, CK => CLK, RN => 
                           n12570, Q => n_2026, QN => n10169);
   REGISTERS_reg_42_10_inst : DFFR_X1 port map( D => n7681, CK => CLK, RN => 
                           n12548, Q => n_2027, QN => n10201);
   REGISTERS_reg_42_9_inst : DFFR_X1 port map( D => n7682, CK => CLK, RN => 
                           n12556, Q => n_2028, QN => n10235);
   REGISTERS_reg_42_8_inst : DFFR_X1 port map( D => n7683, CK => CLK, RN => 
                           n12534, Q => n_2029, QN => n10267);
   REGISTERS_reg_42_7_inst : DFFR_X1 port map( D => n7684, CK => CLK, RN => 
                           n12644, Q => n_2030, QN => n10299);
   REGISTERS_reg_42_6_inst : DFFR_X1 port map( D => n7685, CK => CLK, RN => 
                           n12600, Q => n_2031, QN => n10334);
   REGISTERS_reg_42_5_inst : DFFR_X1 port map( D => n7686, CK => CLK, RN => 
                           n12486, Q => n_2032, QN => n10366);
   REGISTERS_reg_42_4_inst : DFFR_X1 port map( D => n7687, CK => CLK, RN => 
                           n12494, Q => n_2033, QN => n10401);
   REGISTERS_reg_42_3_inst : DFFR_X1 port map( D => n7688, CK => CLK, RN => 
                           n12578, Q => n_2034, QN => n10433);
   REGISTERS_reg_42_2_inst : DFFR_X1 port map( D => n7689, CK => CLK, RN => 
                           n12508, Q => n_2035, QN => n10465);
   REGISTERS_reg_42_1_inst : DFFR_X1 port map( D => n7690, CK => CLK, RN => 
                           n12436, Q => n_2036, QN => n10497);
   REGISTERS_reg_42_0_inst : DFFR_X1 port map( D => n7691, CK => CLK, RN => 
                           n12651, Q => n_2037, QN => n10529);
   REGISTERS_reg_43_31_inst : DFFR_X1 port map( D => n7692, CK => CLK, RN => 
                           n12658, Q => n_2038, QN => n13460);
   REGISTERS_reg_43_30_inst : DFFR_X1 port map( D => n7693, CK => CLK, RN => 
                           n12622, Q => n_2039, QN => n13461);
   REGISTERS_reg_43_29_inst : DFFR_X1 port map( D => n7694, CK => CLK, RN => 
                           n12607, Q => n_2040, QN => n13462);
   REGISTERS_reg_43_28_inst : DFFR_X1 port map( D => n7695, CK => CLK, RN => 
                           n12614, Q => n_2041, QN => n13463);
   REGISTERS_reg_43_27_inst : DFFR_X1 port map( D => n7696, CK => CLK, RN => 
                           n12585, Q => n_2042, QN => n13464);
   REGISTERS_reg_43_26_inst : DFFR_X1 port map( D => n7697, CK => CLK, RN => 
                           n12563, Q => n_2043, QN => n13465);
   REGISTERS_reg_43_25_inst : DFFR_X1 port map( D => n7698, CK => CLK, RN => 
                           n12541, Q => n_2044, QN => n13466);
   REGISTERS_reg_43_24_inst : DFFR_X1 port map( D => n7699, CK => CLK, RN => 
                           n12516, Q => n_2045, QN => n13467);
   REGISTERS_reg_43_23_inst : DFFR_X1 port map( D => n7700, CK => CLK, RN => 
                           n12629, Q => n_2046, QN => n13468);
   REGISTERS_reg_43_22_inst : DFFR_X1 port map( D => n7701, CK => CLK, RN => 
                           n12519, Q => n_2047, QN => n13469);
   REGISTERS_reg_43_21_inst : DFFR_X1 port map( D => n7702, CK => CLK, RN => 
                           n12526, Q => n_2048, QN => n13470);
   REGISTERS_reg_43_20_inst : DFFR_X1 port map( D => n7703, CK => CLK, RN => 
                           n12501, Q => n_2049, QN => n13471);
   REGISTERS_reg_43_19_inst : DFFR_X1 port map( D => n7704, CK => CLK, RN => 
                           n12592, Q => n_2050, QN => n13472);
   REGISTERS_reg_43_18_inst : DFFR_X1 port map( D => n7705, CK => CLK, RN => 
                           n12443, Q => n_2051, QN => n13473);
   REGISTERS_reg_43_17_inst : DFFR_X1 port map( D => n7706, CK => CLK, RN => 
                           n12451, Q => n_2052, QN => n13474);
   REGISTERS_reg_43_16_inst : DFFR_X1 port map( D => n7707, CK => CLK, RN => 
                           n12457, Q => n_2053, QN => n13475);
   REGISTERS_reg_43_15_inst : DFFR_X1 port map( D => n7708, CK => CLK, RN => 
                           n12636, Q => n_2054, QN => n13476);
   REGISTERS_reg_43_14_inst : DFFR_X1 port map( D => n7709, CK => CLK, RN => 
                           n12464, Q => n_2055, QN => n13477);
   REGISTERS_reg_43_13_inst : DFFR_X1 port map( D => n7710, CK => CLK, RN => 
                           n12472, Q => n_2056, QN => n13478);
   REGISTERS_reg_43_12_inst : DFFR_X1 port map( D => n7711, CK => CLK, RN => 
                           n12479, Q => n_2057, QN => n13479);
   REGISTERS_reg_43_11_inst : DFFR_X1 port map( D => n7712, CK => CLK, RN => 
                           n12570, Q => n_2058, QN => n13480);
   REGISTERS_reg_43_10_inst : DFFR_X1 port map( D => n7713, CK => CLK, RN => 
                           n12548, Q => n_2059, QN => n13481);
   REGISTERS_reg_43_9_inst : DFFR_X1 port map( D => n7714, CK => CLK, RN => 
                           n12556, Q => n_2060, QN => n13482);
   REGISTERS_reg_43_8_inst : DFFR_X1 port map( D => n7715, CK => CLK, RN => 
                           n12534, Q => n_2061, QN => n13483);
   REGISTERS_reg_43_7_inst : DFFR_X1 port map( D => n7716, CK => CLK, RN => 
                           n12644, Q => n_2062, QN => n13484);
   REGISTERS_reg_43_6_inst : DFFR_X1 port map( D => n7717, CK => CLK, RN => 
                           n12600, Q => n_2063, QN => n13485);
   REGISTERS_reg_43_5_inst : DFFR_X1 port map( D => n7718, CK => CLK, RN => 
                           n12486, Q => n_2064, QN => n13486);
   REGISTERS_reg_43_4_inst : DFFR_X1 port map( D => n7719, CK => CLK, RN => 
                           n12494, Q => n_2065, QN => n13487);
   REGISTERS_reg_43_3_inst : DFFR_X1 port map( D => n7720, CK => CLK, RN => 
                           n12578, Q => n_2066, QN => n13488);
   REGISTERS_reg_43_2_inst : DFFR_X1 port map( D => n7721, CK => CLK, RN => 
                           n12508, Q => n_2067, QN => n13489);
   REGISTERS_reg_43_1_inst : DFFR_X1 port map( D => n7722, CK => CLK, RN => 
                           n12436, Q => n_2068, QN => n13490);
   REGISTERS_reg_43_0_inst : DFFR_X1 port map( D => n7723, CK => CLK, RN => 
                           n12651, Q => n_2069, QN => n13491);
   REGISTERS_reg_44_31_inst : DFFR_X1 port map( D => n7724, CK => CLK, RN => 
                           n12659, Q => n9567, QN => n13492);
   REGISTERS_reg_44_30_inst : DFFR_X1 port map( D => n7725, CK => CLK, RN => 
                           n12622, Q => n9566, QN => n13493);
   REGISTERS_reg_44_29_inst : DFFR_X1 port map( D => n7726, CK => CLK, RN => 
                           n12607, Q => n9565, QN => n13494);
   REGISTERS_reg_44_28_inst : DFFR_X1 port map( D => n7727, CK => CLK, RN => 
                           n12615, Q => n9564, QN => n13495);
   REGISTERS_reg_44_27_inst : DFFR_X1 port map( D => n7728, CK => CLK, RN => 
                           n12585, Q => n9563, QN => n13496);
   REGISTERS_reg_44_26_inst : DFFR_X1 port map( D => n7729, CK => CLK, RN => 
                           n12563, Q => n9562, QN => n13497);
   REGISTERS_reg_44_25_inst : DFFR_X1 port map( D => n7730, CK => CLK, RN => 
                           n12541, Q => n9561, QN => n13498);
   REGISTERS_reg_44_24_inst : DFFR_X1 port map( D => n7731, CK => CLK, RN => 
                           n12516, Q => n9560, QN => n13499);
   REGISTERS_reg_44_23_inst : DFFR_X1 port map( D => n7732, CK => CLK, RN => 
                           n12629, Q => n9559, QN => n13500);
   REGISTERS_reg_44_22_inst : DFFR_X1 port map( D => n7733, CK => CLK, RN => 
                           n12519, Q => n9558, QN => n13501);
   REGISTERS_reg_44_21_inst : DFFR_X1 port map( D => n7734, CK => CLK, RN => 
                           n12527, Q => n9557, QN => n13502);
   REGISTERS_reg_44_20_inst : DFFR_X1 port map( D => n7735, CK => CLK, RN => 
                           n12501, Q => n9556, QN => n13503);
   REGISTERS_reg_44_19_inst : DFFR_X1 port map( D => n7736, CK => CLK, RN => 
                           n12593, Q => n9555, QN => n13504);
   REGISTERS_reg_44_18_inst : DFFR_X1 port map( D => n7737, CK => CLK, RN => 
                           n12444, Q => n9554, QN => n13505);
   REGISTERS_reg_44_17_inst : DFFR_X1 port map( D => n7738, CK => CLK, RN => 
                           n12451, Q => n9553, QN => n13506);
   REGISTERS_reg_44_16_inst : DFFR_X1 port map( D => n7739, CK => CLK, RN => 
                           n12457, Q => n9552, QN => n13507);
   REGISTERS_reg_44_15_inst : DFFR_X1 port map( D => n7740, CK => CLK, RN => 
                           n12637, Q => n9551, QN => n13508);
   REGISTERS_reg_44_14_inst : DFFR_X1 port map( D => n7741, CK => CLK, RN => 
                           n12465, Q => n9550, QN => n13509);
   REGISTERS_reg_44_13_inst : DFFR_X1 port map( D => n7742, CK => CLK, RN => 
                           n12472, Q => n9549, QN => n13510);
   REGISTERS_reg_44_12_inst : DFFR_X1 port map( D => n7743, CK => CLK, RN => 
                           n12479, Q => n9548, QN => n13511);
   REGISTERS_reg_44_11_inst : DFFR_X1 port map( D => n7744, CK => CLK, RN => 
                           n12571, Q => n9547, QN => n13512);
   REGISTERS_reg_44_10_inst : DFFR_X1 port map( D => n7745, CK => CLK, RN => 
                           n12549, Q => n9546, QN => n13513);
   REGISTERS_reg_44_9_inst : DFFR_X1 port map( D => n7746, CK => CLK, RN => 
                           n12556, Q => n9545, QN => n13514);
   REGISTERS_reg_44_8_inst : DFFR_X1 port map( D => n7747, CK => CLK, RN => 
                           n12534, Q => n9544, QN => n13515);
   REGISTERS_reg_44_7_inst : DFFR_X1 port map( D => n7748, CK => CLK, RN => 
                           n12644, Q => n9543, QN => n13516);
   REGISTERS_reg_44_6_inst : DFFR_X1 port map( D => n7749, CK => CLK, RN => 
                           n12600, Q => n9542, QN => n13517);
   REGISTERS_reg_44_5_inst : DFFR_X1 port map( D => n7750, CK => CLK, RN => 
                           n12487, Q => n9541, QN => n13518);
   REGISTERS_reg_44_4_inst : DFFR_X1 port map( D => n7751, CK => CLK, RN => 
                           n12494, Q => n9540, QN => n13519);
   REGISTERS_reg_44_3_inst : DFFR_X1 port map( D => n7752, CK => CLK, RN => 
                           n12578, Q => n9539, QN => n13520);
   REGISTERS_reg_44_2_inst : DFFR_X1 port map( D => n7753, CK => CLK, RN => 
                           n12509, Q => n9538, QN => n13521);
   REGISTERS_reg_44_1_inst : DFFR_X1 port map( D => n7754, CK => CLK, RN => 
                           n12436, Q => n9537, QN => n13522);
   REGISTERS_reg_44_0_inst : DFFR_X1 port map( D => n7755, CK => CLK, RN => 
                           n12651, Q => n9536, QN => n13523);
   REGISTERS_reg_45_31_inst : DFFR_X1 port map( D => n7756, CK => CLK, RN => 
                           n12659, Q => n9535, QN => n13524);
   REGISTERS_reg_45_30_inst : DFFR_X1 port map( D => n7757, CK => CLK, RN => 
                           n12622, Q => n9534, QN => n13525);
   REGISTERS_reg_45_29_inst : DFFR_X1 port map( D => n7758, CK => CLK, RN => 
                           n12607, Q => n9533, QN => n13526);
   REGISTERS_reg_45_28_inst : DFFR_X1 port map( D => n7759, CK => CLK, RN => 
                           n12615, Q => n9532, QN => n13527);
   REGISTERS_reg_45_27_inst : DFFR_X1 port map( D => n7760, CK => CLK, RN => 
                           n12585, Q => n9531, QN => n13528);
   REGISTERS_reg_45_26_inst : DFFR_X1 port map( D => n7761, CK => CLK, RN => 
                           n12563, Q => n9530, QN => n13529);
   REGISTERS_reg_45_25_inst : DFFR_X1 port map( D => n7762, CK => CLK, RN => 
                           n12541, Q => n9529, QN => n13530);
   REGISTERS_reg_45_24_inst : DFFR_X1 port map( D => n7763, CK => CLK, RN => 
                           n12516, Q => n9528, QN => n13531);
   REGISTERS_reg_45_23_inst : DFFR_X1 port map( D => n7764, CK => CLK, RN => 
                           n12629, Q => n9527, QN => n13532);
   REGISTERS_reg_45_22_inst : DFFR_X1 port map( D => n7765, CK => CLK, RN => 
                           n12519, Q => n9526, QN => n13533);
   REGISTERS_reg_45_21_inst : DFFR_X1 port map( D => n7766, CK => CLK, RN => 
                           n12527, Q => n9525, QN => n13534);
   REGISTERS_reg_45_20_inst : DFFR_X1 port map( D => n7767, CK => CLK, RN => 
                           n12501, Q => n9524, QN => n13535);
   REGISTERS_reg_45_19_inst : DFFR_X1 port map( D => n7768, CK => CLK, RN => 
                           n12593, Q => n9523, QN => n13536);
   REGISTERS_reg_45_18_inst : DFFR_X1 port map( D => n7769, CK => CLK, RN => 
                           n12444, Q => n9522, QN => n13537);
   REGISTERS_reg_45_17_inst : DFFR_X1 port map( D => n7770, CK => CLK, RN => 
                           n12451, Q => n9521, QN => n13538);
   REGISTERS_reg_45_16_inst : DFFR_X1 port map( D => n7771, CK => CLK, RN => 
                           n12457, Q => n9520, QN => n13539);
   REGISTERS_reg_45_15_inst : DFFR_X1 port map( D => n7772, CK => CLK, RN => 
                           n12637, Q => n9519, QN => n13540);
   REGISTERS_reg_45_14_inst : DFFR_X1 port map( D => n7773, CK => CLK, RN => 
                           n12465, Q => n9518, QN => n13541);
   REGISTERS_reg_45_13_inst : DFFR_X1 port map( D => n7774, CK => CLK, RN => 
                           n12472, Q => n9517, QN => n13542);
   REGISTERS_reg_45_12_inst : DFFR_X1 port map( D => n7775, CK => CLK, RN => 
                           n12479, Q => n9516, QN => n13543);
   REGISTERS_reg_45_11_inst : DFFR_X1 port map( D => n7776, CK => CLK, RN => 
                           n12571, Q => n9515, QN => n13544);
   REGISTERS_reg_45_10_inst : DFFR_X1 port map( D => n7777, CK => CLK, RN => 
                           n12549, Q => n9514, QN => n13545);
   REGISTERS_reg_45_9_inst : DFFR_X1 port map( D => n7778, CK => CLK, RN => 
                           n12556, Q => n9513, QN => n13546);
   REGISTERS_reg_45_8_inst : DFFR_X1 port map( D => n7779, CK => CLK, RN => 
                           n12534, Q => n9512, QN => n13547);
   REGISTERS_reg_45_7_inst : DFFR_X1 port map( D => n7780, CK => CLK, RN => 
                           n12644, Q => n9511, QN => n13548);
   REGISTERS_reg_45_6_inst : DFFR_X1 port map( D => n7781, CK => CLK, RN => 
                           n12600, Q => n9510, QN => n13549);
   REGISTERS_reg_45_5_inst : DFFR_X1 port map( D => n7782, CK => CLK, RN => 
                           n12487, Q => n9509, QN => n13550);
   REGISTERS_reg_45_4_inst : DFFR_X1 port map( D => n7783, CK => CLK, RN => 
                           n12494, Q => n9508, QN => n13551);
   REGISTERS_reg_45_3_inst : DFFR_X1 port map( D => n7784, CK => CLK, RN => 
                           n12578, Q => n9507, QN => n13552);
   REGISTERS_reg_45_2_inst : DFFR_X1 port map( D => n7785, CK => CLK, RN => 
                           n12509, Q => n9506, QN => n13553);
   REGISTERS_reg_45_1_inst : DFFR_X1 port map( D => n7786, CK => CLK, RN => 
                           n12436, Q => n9505, QN => n13554);
   REGISTERS_reg_45_0_inst : DFFR_X1 port map( D => n7787, CK => CLK, RN => 
                           n12651, Q => n9504, QN => n13555);
   REGISTERS_reg_46_31_inst : DFFR_X1 port map( D => n7788, CK => CLK, RN => 
                           n12659, Q => n_2070, QN => n13556);
   REGISTERS_reg_46_30_inst : DFFR_X1 port map( D => n7789, CK => CLK, RN => 
                           n12622, Q => n_2071, QN => n13557);
   REGISTERS_reg_46_29_inst : DFFR_X1 port map( D => n7790, CK => CLK, RN => 
                           n12607, Q => n_2072, QN => n13558);
   REGISTERS_reg_46_28_inst : DFFR_X1 port map( D => n7791, CK => CLK, RN => 
                           n12615, Q => n_2073, QN => n13559);
   REGISTERS_reg_46_27_inst : DFFR_X1 port map( D => n7792, CK => CLK, RN => 
                           n12585, Q => n_2074, QN => n13560);
   REGISTERS_reg_46_26_inst : DFFR_X1 port map( D => n7793, CK => CLK, RN => 
                           n12563, Q => n_2075, QN => n13561);
   REGISTERS_reg_46_25_inst : DFFR_X1 port map( D => n7794, CK => CLK, RN => 
                           n12541, Q => n_2076, QN => n13562);
   REGISTERS_reg_46_24_inst : DFFR_X1 port map( D => n7795, CK => CLK, RN => 
                           n12516, Q => n_2077, QN => n13563);
   REGISTERS_reg_46_23_inst : DFFR_X1 port map( D => n7796, CK => CLK, RN => 
                           n12629, Q => n_2078, QN => n13564);
   REGISTERS_reg_46_22_inst : DFFR_X1 port map( D => n7797, CK => CLK, RN => 
                           n12519, Q => n_2079, QN => n13565);
   REGISTERS_reg_46_21_inst : DFFR_X1 port map( D => n7798, CK => CLK, RN => 
                           n12527, Q => n_2080, QN => n13566);
   REGISTERS_reg_46_20_inst : DFFR_X1 port map( D => n7799, CK => CLK, RN => 
                           n12501, Q => n_2081, QN => n13567);
   REGISTERS_reg_46_19_inst : DFFR_X1 port map( D => n7800, CK => CLK, RN => 
                           n12593, Q => n_2082, QN => n13568);
   REGISTERS_reg_46_18_inst : DFFR_X1 port map( D => n7801, CK => CLK, RN => 
                           n12444, Q => n_2083, QN => n13569);
   REGISTERS_reg_46_17_inst : DFFR_X1 port map( D => n7802, CK => CLK, RN => 
                           n12451, Q => n_2084, QN => n13570);
   REGISTERS_reg_46_16_inst : DFFR_X1 port map( D => n7803, CK => CLK, RN => 
                           n12457, Q => n_2085, QN => n13571);
   REGISTERS_reg_46_15_inst : DFFR_X1 port map( D => n7804, CK => CLK, RN => 
                           n12637, Q => n_2086, QN => n13572);
   REGISTERS_reg_46_14_inst : DFFR_X1 port map( D => n7805, CK => CLK, RN => 
                           n12465, Q => n_2087, QN => n13573);
   REGISTERS_reg_46_13_inst : DFFR_X1 port map( D => n7806, CK => CLK, RN => 
                           n12472, Q => n_2088, QN => n13574);
   REGISTERS_reg_46_12_inst : DFFR_X1 port map( D => n7807, CK => CLK, RN => 
                           n12479, Q => n_2089, QN => n13575);
   REGISTERS_reg_46_11_inst : DFFR_X1 port map( D => n7808, CK => CLK, RN => 
                           n12571, Q => n_2090, QN => n13576);
   REGISTERS_reg_46_10_inst : DFFR_X1 port map( D => n7809, CK => CLK, RN => 
                           n12549, Q => n_2091, QN => n13577);
   REGISTERS_reg_46_9_inst : DFFR_X1 port map( D => n7810, CK => CLK, RN => 
                           n12556, Q => n_2092, QN => n13578);
   REGISTERS_reg_46_8_inst : DFFR_X1 port map( D => n7811, CK => CLK, RN => 
                           n12534, Q => n_2093, QN => n13579);
   REGISTERS_reg_46_7_inst : DFFR_X1 port map( D => n7812, CK => CLK, RN => 
                           n12644, Q => n_2094, QN => n13580);
   REGISTERS_reg_46_6_inst : DFFR_X1 port map( D => n7813, CK => CLK, RN => 
                           n12600, Q => n_2095, QN => n13581);
   REGISTERS_reg_46_5_inst : DFFR_X1 port map( D => n7814, CK => CLK, RN => 
                           n12487, Q => n_2096, QN => n13582);
   REGISTERS_reg_46_4_inst : DFFR_X1 port map( D => n7815, CK => CLK, RN => 
                           n12494, Q => n_2097, QN => n13583);
   REGISTERS_reg_46_3_inst : DFFR_X1 port map( D => n7816, CK => CLK, RN => 
                           n12578, Q => n_2098, QN => n13584);
   REGISTERS_reg_46_2_inst : DFFR_X1 port map( D => n7817, CK => CLK, RN => 
                           n12509, Q => n_2099, QN => n13585);
   REGISTERS_reg_46_1_inst : DFFR_X1 port map( D => n7818, CK => CLK, RN => 
                           n12436, Q => n_2100, QN => n13586);
   REGISTERS_reg_46_0_inst : DFFR_X1 port map( D => n7819, CK => CLK, RN => 
                           n12651, Q => n_2101, QN => n13587);
   REGISTERS_reg_47_31_inst : DFFR_X1 port map( D => n7820, CK => CLK, RN => 
                           n12659, Q => n_2102, QN => n13588);
   REGISTERS_reg_47_30_inst : DFFR_X1 port map( D => n7821, CK => CLK, RN => 
                           n12622, Q => n_2103, QN => n13589);
   REGISTERS_reg_47_29_inst : DFFR_X1 port map( D => n7822, CK => CLK, RN => 
                           n12607, Q => n_2104, QN => n13590);
   REGISTERS_reg_47_28_inst : DFFR_X1 port map( D => n7823, CK => CLK, RN => 
                           n12615, Q => n_2105, QN => n13591);
   REGISTERS_reg_47_27_inst : DFFR_X1 port map( D => n7824, CK => CLK, RN => 
                           n12585, Q => n_2106, QN => n13592);
   REGISTERS_reg_47_26_inst : DFFR_X1 port map( D => n7825, CK => CLK, RN => 
                           n12563, Q => n_2107, QN => n13593);
   REGISTERS_reg_47_25_inst : DFFR_X1 port map( D => n7826, CK => CLK, RN => 
                           n12541, Q => n_2108, QN => n13594);
   REGISTERS_reg_47_24_inst : DFFR_X1 port map( D => n7827, CK => CLK, RN => 
                           n12516, Q => n_2109, QN => n13595);
   REGISTERS_reg_47_23_inst : DFFR_X1 port map( D => n7828, CK => CLK, RN => 
                           n12629, Q => n_2110, QN => n13596);
   REGISTERS_reg_47_22_inst : DFFR_X1 port map( D => n7829, CK => CLK, RN => 
                           n12519, Q => n_2111, QN => n13597);
   REGISTERS_reg_47_21_inst : DFFR_X1 port map( D => n7830, CK => CLK, RN => 
                           n12527, Q => n_2112, QN => n13598);
   REGISTERS_reg_47_20_inst : DFFR_X1 port map( D => n7831, CK => CLK, RN => 
                           n12501, Q => n_2113, QN => n13599);
   REGISTERS_reg_47_19_inst : DFFR_X1 port map( D => n7832, CK => CLK, RN => 
                           n12593, Q => n_2114, QN => n13600);
   REGISTERS_reg_47_18_inst : DFFR_X1 port map( D => n7833, CK => CLK, RN => 
                           n12444, Q => n_2115, QN => n13601);
   REGISTERS_reg_47_17_inst : DFFR_X1 port map( D => n7834, CK => CLK, RN => 
                           n12451, Q => n_2116, QN => n13602);
   REGISTERS_reg_47_16_inst : DFFR_X1 port map( D => n7835, CK => CLK, RN => 
                           n12457, Q => n_2117, QN => n13603);
   REGISTERS_reg_47_15_inst : DFFR_X1 port map( D => n7836, CK => CLK, RN => 
                           n12637, Q => n_2118, QN => n13604);
   REGISTERS_reg_47_14_inst : DFFR_X1 port map( D => n7837, CK => CLK, RN => 
                           n12465, Q => n_2119, QN => n13605);
   REGISTERS_reg_47_13_inst : DFFR_X1 port map( D => n7838, CK => CLK, RN => 
                           n12472, Q => n_2120, QN => n13606);
   REGISTERS_reg_47_12_inst : DFFR_X1 port map( D => n7839, CK => CLK, RN => 
                           n12479, Q => n_2121, QN => n13607);
   REGISTERS_reg_47_11_inst : DFFR_X1 port map( D => n7840, CK => CLK, RN => 
                           n12571, Q => n_2122, QN => n13608);
   REGISTERS_reg_47_10_inst : DFFR_X1 port map( D => n7841, CK => CLK, RN => 
                           n12549, Q => n_2123, QN => n13609);
   REGISTERS_reg_47_9_inst : DFFR_X1 port map( D => n7842, CK => CLK, RN => 
                           n12556, Q => n_2124, QN => n13610);
   REGISTERS_reg_47_8_inst : DFFR_X1 port map( D => n7843, CK => CLK, RN => 
                           n12534, Q => n_2125, QN => n13611);
   REGISTERS_reg_47_7_inst : DFFR_X1 port map( D => n7844, CK => CLK, RN => 
                           n12644, Q => n_2126, QN => n13612);
   REGISTERS_reg_47_6_inst : DFFR_X1 port map( D => n7845, CK => CLK, RN => 
                           n12600, Q => n_2127, QN => n13613);
   REGISTERS_reg_47_5_inst : DFFR_X1 port map( D => n7846, CK => CLK, RN => 
                           n12487, Q => n_2128, QN => n13614);
   REGISTERS_reg_47_4_inst : DFFR_X1 port map( D => n7847, CK => CLK, RN => 
                           n12494, Q => n_2129, QN => n13615);
   REGISTERS_reg_47_3_inst : DFFR_X1 port map( D => n7848, CK => CLK, RN => 
                           n12578, Q => n_2130, QN => n13616);
   REGISTERS_reg_47_2_inst : DFFR_X1 port map( D => n7849, CK => CLK, RN => 
                           n12509, Q => n_2131, QN => n13617);
   REGISTERS_reg_47_1_inst : DFFR_X1 port map( D => n7850, CK => CLK, RN => 
                           n12436, Q => n_2132, QN => n13618);
   REGISTERS_reg_47_0_inst : DFFR_X1 port map( D => n7851, CK => CLK, RN => 
                           n12651, Q => n_2133, QN => n13619);
   REGISTERS_reg_48_31_inst : DFFR_X1 port map( D => n7852, CK => CLK, RN => 
                           n12659, Q => n_2134, QN => n13620);
   REGISTERS_reg_48_30_inst : DFFR_X1 port map( D => n7853, CK => CLK, RN => 
                           n12622, Q => n_2135, QN => n13621);
   REGISTERS_reg_48_29_inst : DFFR_X1 port map( D => n7854, CK => CLK, RN => 
                           n12608, Q => n_2136, QN => n13622);
   REGISTERS_reg_48_28_inst : DFFR_X1 port map( D => n7855, CK => CLK, RN => 
                           n12615, Q => n_2137, QN => n13623);
   REGISTERS_reg_48_27_inst : DFFR_X1 port map( D => n7856, CK => CLK, RN => 
                           n12586, Q => n_2138, QN => n13624);
   REGISTERS_reg_48_26_inst : DFFR_X1 port map( D => n7857, CK => CLK, RN => 
                           n12564, Q => n_2139, QN => n13625);
   REGISTERS_reg_48_25_inst : DFFR_X1 port map( D => n7858, CK => CLK, RN => 
                           n12542, Q => n_2140, QN => n13626);
   REGISTERS_reg_48_24_inst : DFFR_X1 port map( D => n7859, CK => CLK, RN => 
                           n12516, Q => n_2141, QN => n13627);
   REGISTERS_reg_48_23_inst : DFFR_X1 port map( D => n7860, CK => CLK, RN => 
                           n12630, Q => n_2142, QN => n13628);
   REGISTERS_reg_48_22_inst : DFFR_X1 port map( D => n7861, CK => CLK, RN => 
                           n12520, Q => n_2143, QN => n13629);
   REGISTERS_reg_48_21_inst : DFFR_X1 port map( D => n7862, CK => CLK, RN => 
                           n12527, Q => n_2144, QN => n13630);
   REGISTERS_reg_48_20_inst : DFFR_X1 port map( D => n7863, CK => CLK, RN => 
                           n12502, Q => n_2145, QN => n13631);
   REGISTERS_reg_48_19_inst : DFFR_X1 port map( D => n7864, CK => CLK, RN => 
                           n12593, Q => n_2146, QN => n13632);
   REGISTERS_reg_48_18_inst : DFFR_X1 port map( D => n7865, CK => CLK, RN => 
                           n12444, Q => n_2147, QN => n13633);
   REGISTERS_reg_48_17_inst : DFFR_X1 port map( D => n7866, CK => CLK, RN => 
                           n12451, Q => n_2148, QN => n13634);
   REGISTERS_reg_48_16_inst : DFFR_X1 port map( D => n7867, CK => CLK, RN => 
                           n12458, Q => n_2149, QN => n13635);
   REGISTERS_reg_48_15_inst : DFFR_X1 port map( D => n7868, CK => CLK, RN => 
                           n12637, Q => n_2150, QN => n13636);
   REGISTERS_reg_48_14_inst : DFFR_X1 port map( D => n7869, CK => CLK, RN => 
                           n12465, Q => n_2151, QN => n13637);
   REGISTERS_reg_48_13_inst : DFFR_X1 port map( D => n7870, CK => CLK, RN => 
                           n12472, Q => n_2152, QN => n13638);
   REGISTERS_reg_48_12_inst : DFFR_X1 port map( D => n7871, CK => CLK, RN => 
                           n12480, Q => n_2153, QN => n13639);
   REGISTERS_reg_48_11_inst : DFFR_X1 port map( D => n7872, CK => CLK, RN => 
                           n12571, Q => n_2154, QN => n13640);
   REGISTERS_reg_48_10_inst : DFFR_X1 port map( D => n7873, CK => CLK, RN => 
                           n12549, Q => n_2155, QN => n13641);
   REGISTERS_reg_48_9_inst : DFFR_X1 port map( D => n7874, CK => CLK, RN => 
                           n12556, Q => n_2156, QN => n13642);
   REGISTERS_reg_48_8_inst : DFFR_X1 port map( D => n7875, CK => CLK, RN => 
                           n12534, Q => n_2157, QN => n13643);
   REGISTERS_reg_48_7_inst : DFFR_X1 port map( D => n7876, CK => CLK, RN => 
                           n12644, Q => n_2158, QN => n13644);
   REGISTERS_reg_48_6_inst : DFFR_X1 port map( D => n7877, CK => CLK, RN => 
                           n12600, Q => n_2159, QN => n13645);
   REGISTERS_reg_48_5_inst : DFFR_X1 port map( D => n7878, CK => CLK, RN => 
                           n12487, Q => n_2160, QN => n13646);
   REGISTERS_reg_48_4_inst : DFFR_X1 port map( D => n7879, CK => CLK, RN => 
                           n12494, Q => n_2161, QN => n13647);
   REGISTERS_reg_48_3_inst : DFFR_X1 port map( D => n7880, CK => CLK, RN => 
                           n12578, Q => n_2162, QN => n13648);
   REGISTERS_reg_48_2_inst : DFFR_X1 port map( D => n7881, CK => CLK, RN => 
                           n12509, Q => n_2163, QN => n13649);
   REGISTERS_reg_48_1_inst : DFFR_X1 port map( D => n7882, CK => CLK, RN => 
                           n12437, Q => n_2164, QN => n13650);
   REGISTERS_reg_48_0_inst : DFFR_X1 port map( D => n7883, CK => CLK, RN => 
                           n12652, Q => n_2165, QN => n13651);
   REGISTERS_reg_49_31_inst : DFFR_X1 port map( D => n7884, CK => CLK, RN => 
                           n12659, Q => n9407, QN => n13652);
   REGISTERS_reg_49_30_inst : DFFR_X1 port map( D => n7885, CK => CLK, RN => 
                           n12622, Q => n9406, QN => n13653);
   REGISTERS_reg_49_29_inst : DFFR_X1 port map( D => n7886, CK => CLK, RN => 
                           n12608, Q => n9405, QN => n13654);
   REGISTERS_reg_49_28_inst : DFFR_X1 port map( D => n7887, CK => CLK, RN => 
                           n12615, Q => n9404, QN => n13655);
   REGISTERS_reg_49_27_inst : DFFR_X1 port map( D => n7888, CK => CLK, RN => 
                           n12586, Q => n9403, QN => n13656);
   REGISTERS_reg_49_26_inst : DFFR_X1 port map( D => n7889, CK => CLK, RN => 
                           n12564, Q => n9402, QN => n13657);
   REGISTERS_reg_49_25_inst : DFFR_X1 port map( D => n7890, CK => CLK, RN => 
                           n12542, Q => n9401, QN => n13658);
   REGISTERS_reg_49_24_inst : DFFR_X1 port map( D => n7891, CK => CLK, RN => 
                           n12516, Q => n9400, QN => n13659);
   REGISTERS_reg_49_23_inst : DFFR_X1 port map( D => n7892, CK => CLK, RN => 
                           n12630, Q => n9399, QN => n13660);
   REGISTERS_reg_49_22_inst : DFFR_X1 port map( D => n7893, CK => CLK, RN => 
                           n12520, Q => n9398, QN => n13661);
   REGISTERS_reg_49_21_inst : DFFR_X1 port map( D => n7894, CK => CLK, RN => 
                           n12527, Q => n9397, QN => n13662);
   REGISTERS_reg_49_20_inst : DFFR_X1 port map( D => n7895, CK => CLK, RN => 
                           n12502, Q => n9396, QN => n13663);
   REGISTERS_reg_49_19_inst : DFFR_X1 port map( D => n7896, CK => CLK, RN => 
                           n12593, Q => n9395, QN => n13664);
   REGISTERS_reg_49_18_inst : DFFR_X1 port map( D => n7897, CK => CLK, RN => 
                           n12444, Q => n9394, QN => n13665);
   REGISTERS_reg_49_17_inst : DFFR_X1 port map( D => n7898, CK => CLK, RN => 
                           n12451, Q => n9393, QN => n13666);
   REGISTERS_reg_49_16_inst : DFFR_X1 port map( D => n7899, CK => CLK, RN => 
                           n12458, Q => n9392, QN => n13667);
   REGISTERS_reg_49_15_inst : DFFR_X1 port map( D => n7900, CK => CLK, RN => 
                           n12637, Q => n9391, QN => n13668);
   REGISTERS_reg_49_14_inst : DFFR_X1 port map( D => n7901, CK => CLK, RN => 
                           n12465, Q => n9390, QN => n13669);
   REGISTERS_reg_49_13_inst : DFFR_X1 port map( D => n7902, CK => CLK, RN => 
                           n12472, Q => n9389, QN => n13670);
   REGISTERS_reg_49_12_inst : DFFR_X1 port map( D => n7903, CK => CLK, RN => 
                           n12480, Q => n9388, QN => n13671);
   REGISTERS_reg_49_11_inst : DFFR_X1 port map( D => n7904, CK => CLK, RN => 
                           n12571, Q => n9387, QN => n13672);
   REGISTERS_reg_49_10_inst : DFFR_X1 port map( D => n7905, CK => CLK, RN => 
                           n12549, Q => n9386, QN => n13673);
   REGISTERS_reg_49_9_inst : DFFR_X1 port map( D => n7906, CK => CLK, RN => 
                           n12556, Q => n9385, QN => n13674);
   REGISTERS_reg_49_8_inst : DFFR_X1 port map( D => n7907, CK => CLK, RN => 
                           n12534, Q => n9384, QN => n13675);
   REGISTERS_reg_49_7_inst : DFFR_X1 port map( D => n7908, CK => CLK, RN => 
                           n12644, Q => n9383, QN => n13676);
   REGISTERS_reg_49_6_inst : DFFR_X1 port map( D => n7909, CK => CLK, RN => 
                           n12600, Q => n9382, QN => n13677);
   REGISTERS_reg_49_5_inst : DFFR_X1 port map( D => n7910, CK => CLK, RN => 
                           n12487, Q => n9381, QN => n13678);
   REGISTERS_reg_49_4_inst : DFFR_X1 port map( D => n7911, CK => CLK, RN => 
                           n12494, Q => n9380, QN => n13679);
   REGISTERS_reg_49_3_inst : DFFR_X1 port map( D => n7912, CK => CLK, RN => 
                           n12578, Q => n9379, QN => n13680);
   REGISTERS_reg_49_2_inst : DFFR_X1 port map( D => n7913, CK => CLK, RN => 
                           n12509, Q => n9378, QN => n13681);
   REGISTERS_reg_49_1_inst : DFFR_X1 port map( D => n7914, CK => CLK, RN => 
                           n12437, Q => n9377, QN => n13682);
   REGISTERS_reg_49_0_inst : DFFR_X1 port map( D => n7915, CK => CLK, RN => 
                           n12652, Q => n9376, QN => n13683);
   REGISTERS_reg_50_31_inst : DFFR_X1 port map( D => n7916, CK => CLK, RN => 
                           n12659, Q => n9375, QN => n13684);
   REGISTERS_reg_50_30_inst : DFFR_X1 port map( D => n7917, CK => CLK, RN => 
                           n12622, Q => n9374, QN => n13685);
   REGISTERS_reg_50_29_inst : DFFR_X1 port map( D => n7918, CK => CLK, RN => 
                           n12608, Q => n9373, QN => n13686);
   REGISTERS_reg_50_28_inst : DFFR_X1 port map( D => n7919, CK => CLK, RN => 
                           n12615, Q => n9372, QN => n13687);
   REGISTERS_reg_50_27_inst : DFFR_X1 port map( D => n7920, CK => CLK, RN => 
                           n12586, Q => n9371, QN => n13688);
   REGISTERS_reg_50_26_inst : DFFR_X1 port map( D => n7921, CK => CLK, RN => 
                           n12564, Q => n9370, QN => n13689);
   REGISTERS_reg_50_25_inst : DFFR_X1 port map( D => n7922, CK => CLK, RN => 
                           n12542, Q => n9369, QN => n13690);
   REGISTERS_reg_50_24_inst : DFFR_X1 port map( D => n7923, CK => CLK, RN => 
                           n12516, Q => n9368, QN => n13691);
   REGISTERS_reg_50_23_inst : DFFR_X1 port map( D => n7924, CK => CLK, RN => 
                           n12630, Q => n9367, QN => n13692);
   REGISTERS_reg_50_22_inst : DFFR_X1 port map( D => n7925, CK => CLK, RN => 
                           n12520, Q => n9366, QN => n13693);
   REGISTERS_reg_50_21_inst : DFFR_X1 port map( D => n7926, CK => CLK, RN => 
                           n12527, Q => n9365, QN => n13694);
   REGISTERS_reg_50_20_inst : DFFR_X1 port map( D => n7927, CK => CLK, RN => 
                           n12502, Q => n9364, QN => n13695);
   REGISTERS_reg_50_19_inst : DFFR_X1 port map( D => n7928, CK => CLK, RN => 
                           n12593, Q => n9363, QN => n13696);
   REGISTERS_reg_50_18_inst : DFFR_X1 port map( D => n7929, CK => CLK, RN => 
                           n12444, Q => n9362, QN => n13697);
   REGISTERS_reg_50_17_inst : DFFR_X1 port map( D => n7930, CK => CLK, RN => 
                           n12451, Q => n9361, QN => n13698);
   REGISTERS_reg_50_16_inst : DFFR_X1 port map( D => n7931, CK => CLK, RN => 
                           n12458, Q => n9360, QN => n13699);
   REGISTERS_reg_50_15_inst : DFFR_X1 port map( D => n7932, CK => CLK, RN => 
                           n12637, Q => n9359, QN => n13700);
   REGISTERS_reg_50_14_inst : DFFR_X1 port map( D => n7933, CK => CLK, RN => 
                           n12465, Q => n9358, QN => n13701);
   REGISTERS_reg_50_13_inst : DFFR_X1 port map( D => n7934, CK => CLK, RN => 
                           n12472, Q => n9357, QN => n13702);
   REGISTERS_reg_50_12_inst : DFFR_X1 port map( D => n7935, CK => CLK, RN => 
                           n12480, Q => n9356, QN => n13703);
   REGISTERS_reg_50_11_inst : DFFR_X1 port map( D => n7936, CK => CLK, RN => 
                           n12571, Q => n9355, QN => n13704);
   REGISTERS_reg_50_10_inst : DFFR_X1 port map( D => n7937, CK => CLK, RN => 
                           n12549, Q => n9354, QN => n13705);
   REGISTERS_reg_50_9_inst : DFFR_X1 port map( D => n7938, CK => CLK, RN => 
                           n12556, Q => n9353, QN => n13706);
   REGISTERS_reg_50_8_inst : DFFR_X1 port map( D => n7939, CK => CLK, RN => 
                           n12534, Q => n9352, QN => n13707);
   REGISTERS_reg_50_7_inst : DFFR_X1 port map( D => n7940, CK => CLK, RN => 
                           n12644, Q => n9351, QN => n13708);
   REGISTERS_reg_50_6_inst : DFFR_X1 port map( D => n7941, CK => CLK, RN => 
                           n12600, Q => n9350, QN => n13709);
   REGISTERS_reg_50_5_inst : DFFR_X1 port map( D => n7942, CK => CLK, RN => 
                           n12487, Q => n9349, QN => n13710);
   REGISTERS_reg_50_4_inst : DFFR_X1 port map( D => n7943, CK => CLK, RN => 
                           n12494, Q => n9348, QN => n13711);
   REGISTERS_reg_50_3_inst : DFFR_X1 port map( D => n7944, CK => CLK, RN => 
                           n12578, Q => n9347, QN => n13712);
   REGISTERS_reg_50_2_inst : DFFR_X1 port map( D => n7945, CK => CLK, RN => 
                           n12509, Q => n9346, QN => n13713);
   REGISTERS_reg_50_1_inst : DFFR_X1 port map( D => n7946, CK => CLK, RN => 
                           n12437, Q => n9345, QN => n13714);
   REGISTERS_reg_50_0_inst : DFFR_X1 port map( D => n7947, CK => CLK, RN => 
                           n12652, Q => n9344, QN => n13715);
   REGISTERS_reg_51_31_inst : DFFR_X1 port map( D => n7948, CK => CLK, RN => 
                           n12659, Q => n9343, QN => n13716);
   REGISTERS_reg_51_30_inst : DFFR_X1 port map( D => n7949, CK => CLK, RN => 
                           n12622, Q => n9342, QN => n13717);
   REGISTERS_reg_51_29_inst : DFFR_X1 port map( D => n7950, CK => CLK, RN => 
                           n12608, Q => n9341, QN => n13718);
   REGISTERS_reg_51_28_inst : DFFR_X1 port map( D => n7951, CK => CLK, RN => 
                           n12615, Q => n9340, QN => n13719);
   REGISTERS_reg_51_27_inst : DFFR_X1 port map( D => n7952, CK => CLK, RN => 
                           n12586, Q => n9339, QN => n13720);
   REGISTERS_reg_51_26_inst : DFFR_X1 port map( D => n7953, CK => CLK, RN => 
                           n12564, Q => n9338, QN => n13721);
   REGISTERS_reg_51_25_inst : DFFR_X1 port map( D => n7954, CK => CLK, RN => 
                           n12542, Q => n9337, QN => n13722);
   REGISTERS_reg_51_24_inst : DFFR_X1 port map( D => n7955, CK => CLK, RN => 
                           n12516, Q => n9336, QN => n13723);
   REGISTERS_reg_51_23_inst : DFFR_X1 port map( D => n7956, CK => CLK, RN => 
                           n12630, Q => n9335, QN => n13724);
   REGISTERS_reg_51_22_inst : DFFR_X1 port map( D => n7957, CK => CLK, RN => 
                           n12520, Q => n9334, QN => n13725);
   REGISTERS_reg_51_21_inst : DFFR_X1 port map( D => n7958, CK => CLK, RN => 
                           n12527, Q => n9333, QN => n13726);
   REGISTERS_reg_51_20_inst : DFFR_X1 port map( D => n7959, CK => CLK, RN => 
                           n12502, Q => n9332, QN => n13727);
   REGISTERS_reg_51_19_inst : DFFR_X1 port map( D => n7960, CK => CLK, RN => 
                           n12593, Q => n9331, QN => n13728);
   REGISTERS_reg_51_18_inst : DFFR_X1 port map( D => n7961, CK => CLK, RN => 
                           n12444, Q => n9330, QN => n13729);
   REGISTERS_reg_51_17_inst : DFFR_X1 port map( D => n7962, CK => CLK, RN => 
                           n12451, Q => n9329, QN => n13730);
   REGISTERS_reg_51_16_inst : DFFR_X1 port map( D => n7963, CK => CLK, RN => 
                           n12458, Q => n9328, QN => n13731);
   REGISTERS_reg_51_15_inst : DFFR_X1 port map( D => n7964, CK => CLK, RN => 
                           n12637, Q => n9327, QN => n13732);
   REGISTERS_reg_51_14_inst : DFFR_X1 port map( D => n7965, CK => CLK, RN => 
                           n12465, Q => n9326, QN => n13733);
   REGISTERS_reg_51_13_inst : DFFR_X1 port map( D => n7966, CK => CLK, RN => 
                           n12472, Q => n9325, QN => n13734);
   REGISTERS_reg_51_12_inst : DFFR_X1 port map( D => n7967, CK => CLK, RN => 
                           n12480, Q => n9324, QN => n13735);
   REGISTERS_reg_51_11_inst : DFFR_X1 port map( D => n7968, CK => CLK, RN => 
                           n12571, Q => n9323, QN => n13736);
   REGISTERS_reg_51_10_inst : DFFR_X1 port map( D => n7969, CK => CLK, RN => 
                           n12549, Q => n9322, QN => n13737);
   REGISTERS_reg_51_9_inst : DFFR_X1 port map( D => n7970, CK => CLK, RN => 
                           n12556, Q => n9321, QN => n13738);
   REGISTERS_reg_51_8_inst : DFFR_X1 port map( D => n7971, CK => CLK, RN => 
                           n12534, Q => n9320, QN => n13739);
   REGISTERS_reg_51_7_inst : DFFR_X1 port map( D => n7972, CK => CLK, RN => 
                           n12644, Q => n9319, QN => n13740);
   REGISTERS_reg_51_6_inst : DFFR_X1 port map( D => n7973, CK => CLK, RN => 
                           n12600, Q => n9318, QN => n13741);
   REGISTERS_reg_51_5_inst : DFFR_X1 port map( D => n7974, CK => CLK, RN => 
                           n12487, Q => n9317, QN => n13742);
   REGISTERS_reg_51_4_inst : DFFR_X1 port map( D => n7975, CK => CLK, RN => 
                           n12494, Q => n9316, QN => n13743);
   REGISTERS_reg_51_3_inst : DFFR_X1 port map( D => n7976, CK => CLK, RN => 
                           n12578, Q => n9315, QN => n13744);
   REGISTERS_reg_51_2_inst : DFFR_X1 port map( D => n7977, CK => CLK, RN => 
                           n12509, Q => n9314, QN => n13745);
   REGISTERS_reg_51_1_inst : DFFR_X1 port map( D => n7978, CK => CLK, RN => 
                           n12437, Q => n9313, QN => n13746);
   REGISTERS_reg_51_0_inst : DFFR_X1 port map( D => n7979, CK => CLK, RN => 
                           n12652, Q => n9312, QN => n13747);
   REGISTERS_reg_52_30_inst : DFFR_X1 port map( D => n7981, CK => CLK, RN => 
                           n12623, Q => n9310, QN => n13749);
   REGISTERS_reg_52_29_inst : DFFR_X1 port map( D => n7982, CK => CLK, RN => 
                           n12608, Q => n9309, QN => n13750);
   REGISTERS_reg_52_28_inst : DFFR_X1 port map( D => n7983, CK => CLK, RN => 
                           n12615, Q => n9308, QN => n13751);
   REGISTERS_reg_52_27_inst : DFFR_X1 port map( D => n7984, CK => CLK, RN => 
                           n12586, Q => n9307, QN => n13752);
   REGISTERS_reg_52_26_inst : DFFR_X1 port map( D => n7985, CK => CLK, RN => 
                           n12564, Q => n9306, QN => n13753);
   REGISTERS_reg_52_25_inst : DFFR_X1 port map( D => n7986, CK => CLK, RN => 
                           n12542, Q => n9305, QN => n13754);
   REGISTERS_reg_52_24_inst : DFFR_X1 port map( D => n7987, CK => CLK, RN => 
                           n12463, Q => n9304, QN => n13755);
   REGISTERS_reg_52_23_inst : DFFR_X1 port map( D => n7988, CK => CLK, RN => 
                           n12630, Q => n9303, QN => n13756);
   REGISTERS_reg_52_22_inst : DFFR_X1 port map( D => n7989, CK => CLK, RN => 
                           n12520, Q => n9302, QN => n13757);
   REGISTERS_reg_52_21_inst : DFFR_X1 port map( D => n7990, CK => CLK, RN => 
                           n12527, Q => n9301, QN => n13758);
   REGISTERS_reg_52_20_inst : DFFR_X1 port map( D => n7991, CK => CLK, RN => 
                           n12502, Q => n9300, QN => n13759);
   REGISTERS_reg_52_19_inst : DFFR_X1 port map( D => n7992, CK => CLK, RN => 
                           n12593, Q => n9299, QN => n13760);
   REGISTERS_reg_52_18_inst : DFFR_X1 port map( D => n7993, CK => CLK, RN => 
                           n12444, Q => n9298, QN => n13761);
   REGISTERS_reg_52_17_inst : DFFR_X1 port map( D => n7994, CK => CLK, RN => 
                           n12452, Q => n9297, QN => n13762);
   REGISTERS_reg_52_16_inst : DFFR_X1 port map( D => n7995, CK => CLK, RN => 
                           n12458, Q => n9296, QN => n13763);
   REGISTERS_reg_52_15_inst : DFFR_X1 port map( D => n7996, CK => CLK, RN => 
                           n12637, Q => n9295, QN => n13764);
   REGISTERS_reg_52_14_inst : DFFR_X1 port map( D => n7997, CK => CLK, RN => 
                           n12465, Q => n9294, QN => n13765);
   REGISTERS_reg_52_13_inst : DFFR_X1 port map( D => n7998, CK => CLK, RN => 
                           n12473, Q => n9293, QN => n13766);
   REGISTERS_reg_52_12_inst : DFFR_X1 port map( D => n7999, CK => CLK, RN => 
                           n12480, Q => n9292, QN => n13767);
   REGISTERS_reg_52_11_inst : DFFR_X1 port map( D => n8000, CK => CLK, RN => 
                           n12571, Q => n9291, QN => n13768);
   REGISTERS_reg_52_10_inst : DFFR_X1 port map( D => n8001, CK => CLK, RN => 
                           n12549, Q => n9290, QN => n13769);
   REGISTERS_reg_52_9_inst : DFFR_X1 port map( D => n8002, CK => CLK, RN => 
                           n12557, Q => n9289, QN => n13770);
   REGISTERS_reg_52_8_inst : DFFR_X1 port map( D => n8003, CK => CLK, RN => 
                           n12535, Q => n9288, QN => n13771);
   REGISTERS_reg_52_7_inst : DFFR_X1 port map( D => n8004, CK => CLK, RN => 
                           n12645, Q => n9287, QN => n13772);
   REGISTERS_reg_52_6_inst : DFFR_X1 port map( D => n8005, CK => CLK, RN => 
                           n12601, Q => n9286, QN => n13773);
   REGISTERS_reg_52_5_inst : DFFR_X1 port map( D => n8006, CK => CLK, RN => 
                           n12487, Q => n9285, QN => n13774);
   REGISTERS_reg_52_4_inst : DFFR_X1 port map( D => n8007, CK => CLK, RN => 
                           n12495, Q => n9284, QN => n13775);
   REGISTERS_reg_52_3_inst : DFFR_X1 port map( D => n8008, CK => CLK, RN => 
                           n12579, Q => n9283, QN => n13776);
   REGISTERS_reg_52_2_inst : DFFR_X1 port map( D => n8009, CK => CLK, RN => 
                           n12509, Q => n9282, QN => n13777);
   REGISTERS_reg_52_1_inst : DFFR_X1 port map( D => n8010, CK => CLK, RN => 
                           n12437, Q => n9281, QN => n13778);
   REGISTERS_reg_52_0_inst : DFFR_X1 port map( D => n8011, CK => CLK, RN => 
                           n12652, Q => n9280, QN => n13779);
   REGISTERS_reg_53_31_inst : DFFR_X1 port map( D => n8012, CK => CLK, RN => 
                           n12659, Q => n9279, QN => n13780);
   REGISTERS_reg_53_30_inst : DFFR_X1 port map( D => n8013, CK => CLK, RN => 
                           n12623, Q => n9278, QN => n13781);
   REGISTERS_reg_53_29_inst : DFFR_X1 port map( D => n8014, CK => CLK, RN => 
                           n12608, Q => n9277, QN => n13782);
   REGISTERS_reg_53_28_inst : DFFR_X1 port map( D => n8015, CK => CLK, RN => 
                           n12615, Q => n9276, QN => n13783);
   REGISTERS_reg_53_27_inst : DFFR_X1 port map( D => n8016, CK => CLK, RN => 
                           n12586, Q => n9275, QN => n13784);
   REGISTERS_reg_53_26_inst : DFFR_X1 port map( D => n8017, CK => CLK, RN => 
                           n12564, Q => n9274, QN => n13785);
   REGISTERS_reg_53_25_inst : DFFR_X1 port map( D => n8018, CK => CLK, RN => 
                           n12542, Q => n9273, QN => n13786);
   REGISTERS_reg_53_24_inst : DFFR_X1 port map( D => n8019, CK => CLK, RN => 
                           n12462, Q => n9272, QN => n13787);
   REGISTERS_reg_53_23_inst : DFFR_X1 port map( D => n8020, CK => CLK, RN => 
                           n12630, Q => n9271, QN => n13788);
   REGISTERS_reg_53_22_inst : DFFR_X1 port map( D => n8021, CK => CLK, RN => 
                           n12520, Q => n9270, QN => n13789);
   REGISTERS_reg_53_21_inst : DFFR_X1 port map( D => n8022, CK => CLK, RN => 
                           n12527, Q => n9269, QN => n13790);
   REGISTERS_reg_53_20_inst : DFFR_X1 port map( D => n8023, CK => CLK, RN => 
                           n12502, Q => n9268, QN => n13791);
   REGISTERS_reg_53_19_inst : DFFR_X1 port map( D => n8024, CK => CLK, RN => 
                           n12593, Q => n9267, QN => n13792);
   REGISTERS_reg_53_18_inst : DFFR_X1 port map( D => n8025, CK => CLK, RN => 
                           n12444, Q => n9266, QN => n13793);
   REGISTERS_reg_53_17_inst : DFFR_X1 port map( D => n8026, CK => CLK, RN => 
                           n12452, Q => n9265, QN => n13794);
   REGISTERS_reg_54_31_inst : DFFR_X1 port map( D => n8044, CK => CLK, RN => 
                           n12659, Q => n9247, QN => n13812);
   REGISTERS_reg_54_30_inst : DFFR_X1 port map( D => n8045, CK => CLK, RN => 
                           n12623, Q => n9246, QN => n13813);
   REGISTERS_reg_54_29_inst : DFFR_X1 port map( D => n8046, CK => CLK, RN => 
                           n12608, Q => n9245, QN => n13814);
   REGISTERS_reg_54_28_inst : DFFR_X1 port map( D => n8047, CK => CLK, RN => 
                           n12615, Q => n9244, QN => n13815);
   REGISTERS_reg_54_27_inst : DFFR_X1 port map( D => n8048, CK => CLK, RN => 
                           n12586, Q => n9243, QN => n13816);
   REGISTERS_reg_54_26_inst : DFFR_X1 port map( D => n8049, CK => CLK, RN => 
                           n12564, Q => n9242, QN => n13817);
   REGISTERS_reg_54_25_inst : DFFR_X1 port map( D => n8050, CK => CLK, RN => 
                           n12542, Q => n9241, QN => n13818);
   REGISTERS_reg_54_24_inst : DFFR_X1 port map( D => n8051, CK => CLK, RN => 
                           n12481, Q => n9240, QN => n13819);
   REGISTERS_reg_54_23_inst : DFFR_X1 port map( D => n8052, CK => CLK, RN => 
                           n12630, Q => n9239, QN => n13820);
   REGISTERS_reg_54_22_inst : DFFR_X1 port map( D => n8053, CK => CLK, RN => 
                           n12520, Q => n9238, QN => n13821);
   REGISTERS_reg_54_21_inst : DFFR_X1 port map( D => n8054, CK => CLK, RN => 
                           n12527, Q => n9237, QN => n13822);
   REGISTERS_reg_54_20_inst : DFFR_X1 port map( D => n8055, CK => CLK, RN => 
                           n12502, Q => n9236, QN => n13823);
   REGISTERS_reg_54_19_inst : DFFR_X1 port map( D => n8056, CK => CLK, RN => 
                           n12593, Q => n9235, QN => n13824);
   REGISTERS_reg_54_18_inst : DFFR_X1 port map( D => n8057, CK => CLK, RN => 
                           n12444, Q => n9234, QN => n13825);
   REGISTERS_reg_54_17_inst : DFFR_X1 port map( D => n8058, CK => CLK, RN => 
                           n12452, Q => n9233, QN => n13826);
   REGISTERS_reg_54_16_inst : DFFR_X1 port map( D => n8059, CK => CLK, RN => 
                           n12458, Q => n9232, QN => n13827);
   REGISTERS_reg_54_15_inst : DFFR_X1 port map( D => n8060, CK => CLK, RN => 
                           n12637, Q => n9231, QN => n13828);
   REGISTERS_reg_54_14_inst : DFFR_X1 port map( D => n8061, CK => CLK, RN => 
                           n12465, Q => n9230, QN => n13829);
   REGISTERS_reg_54_13_inst : DFFR_X1 port map( D => n8062, CK => CLK, RN => 
                           n12473, Q => n9229, QN => n13830);
   REGISTERS_reg_54_12_inst : DFFR_X1 port map( D => n8063, CK => CLK, RN => 
                           n12480, Q => n9228, QN => n13831);
   REGISTERS_reg_54_11_inst : DFFR_X1 port map( D => n8064, CK => CLK, RN => 
                           n12571, Q => n9227, QN => n13832);
   REGISTERS_reg_54_10_inst : DFFR_X1 port map( D => n8065, CK => CLK, RN => 
                           n12549, Q => n9226, QN => n13833);
   REGISTERS_reg_54_9_inst : DFFR_X1 port map( D => n8066, CK => CLK, RN => 
                           n12557, Q => n9225, QN => n13834);
   REGISTERS_reg_54_8_inst : DFFR_X1 port map( D => n8067, CK => CLK, RN => 
                           n12535, Q => n9224, QN => n13835);
   REGISTERS_reg_54_7_inst : DFFR_X1 port map( D => n8068, CK => CLK, RN => 
                           n12645, Q => n9223, QN => n13836);
   REGISTERS_reg_54_6_inst : DFFR_X1 port map( D => n8069, CK => CLK, RN => 
                           n12601, Q => n9222, QN => n13837);
   REGISTERS_reg_54_5_inst : DFFR_X1 port map( D => n8070, CK => CLK, RN => 
                           n12487, Q => n9221, QN => n13838);
   REGISTERS_reg_54_4_inst : DFFR_X1 port map( D => n8071, CK => CLK, RN => 
                           n12495, Q => n9220, QN => n13839);
   REGISTERS_reg_54_3_inst : DFFR_X1 port map( D => n8072, CK => CLK, RN => 
                           n12579, Q => n9219, QN => n13840);
   REGISTERS_reg_54_2_inst : DFFR_X1 port map( D => n8073, CK => CLK, RN => 
                           n12509, Q => n9218, QN => n13841);
   REGISTERS_reg_54_1_inst : DFFR_X1 port map( D => n8074, CK => CLK, RN => 
                           n12437, Q => n9217, QN => n13842);
   REGISTERS_reg_54_0_inst : DFFR_X1 port map( D => n8075, CK => CLK, RN => 
                           n12652, Q => n9216, QN => n13843);
   REGISTERS_reg_55_31_inst : DFFR_X1 port map( D => n8076, CK => CLK, RN => 
                           n12659, Q => n_2166, QN => n5721);
   REGISTERS_reg_55_30_inst : DFFR_X1 port map( D => n8077, CK => CLK, RN => 
                           n12623, Q => n_2167, QN => n5753);
   REGISTERS_reg_55_29_inst : DFFR_X1 port map( D => n8078, CK => CLK, RN => 
                           n12608, Q => n_2168, QN => n5785);
   REGISTERS_reg_55_28_inst : DFFR_X1 port map( D => n8079, CK => CLK, RN => 
                           n12615, Q => n_2169, QN => n5817);
   REGISTERS_reg_55_27_inst : DFFR_X1 port map( D => n8080, CK => CLK, RN => 
                           n12586, Q => n_2170, QN => n5849);
   REGISTERS_reg_55_26_inst : DFFR_X1 port map( D => n8081, CK => CLK, RN => 
                           n12564, Q => n_2171, QN => n5881);
   REGISTERS_reg_55_25_inst : DFFR_X1 port map( D => n8082, CK => CLK, RN => 
                           n12542, Q => n_2172, QN => n5913);
   REGISTERS_reg_55_24_inst : DFFR_X1 port map( D => n8083, CK => CLK, RN => 
                           n12480, Q => n_2173, QN => n5945);
   REGISTERS_reg_55_23_inst : DFFR_X1 port map( D => n8084, CK => CLK, RN => 
                           n12630, Q => n_2174, QN => n6009);
   REGISTERS_reg_55_22_inst : DFFR_X1 port map( D => n8085, CK => CLK, RN => 
                           n12520, Q => n_2175, QN => n9144);
   REGISTERS_reg_55_21_inst : DFFR_X1 port map( D => n8086, CK => CLK, RN => 
                           n12527, Q => n_2176, QN => n9176);
   REGISTERS_reg_55_20_inst : DFFR_X1 port map( D => n8087, CK => CLK, RN => 
                           n12502, Q => n_2177, QN => n9208);
   REGISTERS_reg_55_19_inst : DFFR_X1 port map( D => n8088, CK => CLK, RN => 
                           n12593, Q => n_2178, QN => n9574);
   REGISTERS_reg_55_18_inst : DFFR_X1 port map( D => n8089, CK => CLK, RN => 
                           n12444, Q => n_2179, QN => n9606);
   REGISTERS_reg_55_17_inst : DFFR_X1 port map( D => n8090, CK => CLK, RN => 
                           n12452, Q => n_2180, QN => n9638);
   REGISTERS_reg_55_16_inst : DFFR_X1 port map( D => n8091, CK => CLK, RN => 
                           n12458, Q => n_2181, QN => n10000);
   REGISTERS_reg_55_15_inst : DFFR_X1 port map( D => n8092, CK => CLK, RN => 
                           n12637, Q => n_2182, QN => n10032);
   REGISTERS_reg_55_14_inst : DFFR_X1 port map( D => n8093, CK => CLK, RN => 
                           n12465, Q => n_2183, QN => n10064);
   REGISTERS_reg_55_13_inst : DFFR_X1 port map( D => n8094, CK => CLK, RN => 
                           n12473, Q => n_2184, QN => n10096);
   REGISTERS_reg_55_12_inst : DFFR_X1 port map( D => n8095, CK => CLK, RN => 
                           n12480, Q => n_2185, QN => n10128);
   REGISTERS_reg_55_11_inst : DFFR_X1 port map( D => n8096, CK => CLK, RN => 
                           n12571, Q => n_2186, QN => n10160);
   REGISTERS_reg_55_10_inst : DFFR_X1 port map( D => n8097, CK => CLK, RN => 
                           n12549, Q => n_2187, QN => n10192);
   REGISTERS_reg_55_9_inst : DFFR_X1 port map( D => n8098, CK => CLK, RN => 
                           n12557, Q => n_2188, QN => n10226);
   REGISTERS_reg_55_8_inst : DFFR_X1 port map( D => n8099, CK => CLK, RN => 
                           n12535, Q => n_2189, QN => n10258);
   REGISTERS_reg_55_7_inst : DFFR_X1 port map( D => n8100, CK => CLK, RN => 
                           n12645, Q => n_2190, QN => n10290);
   REGISTERS_reg_55_6_inst : DFFR_X1 port map( D => n8101, CK => CLK, RN => 
                           n12601, Q => n_2191, QN => n10325);
   REGISTERS_reg_55_5_inst : DFFR_X1 port map( D => n8102, CK => CLK, RN => 
                           n12487, Q => n_2192, QN => n10357);
   REGISTERS_reg_55_4_inst : DFFR_X1 port map( D => n8103, CK => CLK, RN => 
                           n12495, Q => n_2193, QN => n10389);
   REGISTERS_reg_55_3_inst : DFFR_X1 port map( D => n8104, CK => CLK, RN => 
                           n12579, Q => n_2194, QN => n10424);
   REGISTERS_reg_55_2_inst : DFFR_X1 port map( D => n8105, CK => CLK, RN => 
                           n12509, Q => n_2195, QN => n10456);
   REGISTERS_reg_55_1_inst : DFFR_X1 port map( D => n8106, CK => CLK, RN => 
                           n12437, Q => n_2196, QN => n10488);
   REGISTERS_reg_55_0_inst : DFFR_X1 port map( D => n8107, CK => CLK, RN => 
                           n12652, Q => n_2197, QN => n10520);
   REGISTERS_reg_56_31_inst : DFFR_X1 port map( D => n8108, CK => CLK, RN => 
                           n12660, Q => n_2198, QN => n5720);
   REGISTERS_reg_56_30_inst : DFFR_X1 port map( D => n8109, CK => CLK, RN => 
                           n12623, Q => n_2199, QN => n5752);
   REGISTERS_reg_56_29_inst : DFFR_X1 port map( D => n8110, CK => CLK, RN => 
                           n12608, Q => n_2200, QN => n5784);
   REGISTERS_reg_56_28_inst : DFFR_X1 port map( D => n8111, CK => CLK, RN => 
                           n12616, Q => n_2201, QN => n5816);
   REGISTERS_reg_56_27_inst : DFFR_X1 port map( D => n8112, CK => CLK, RN => 
                           n12586, Q => n_2202, QN => n5848);
   REGISTERS_reg_56_26_inst : DFFR_X1 port map( D => n8113, CK => CLK, RN => 
                           n12564, Q => n_2203, QN => n5880);
   REGISTERS_reg_56_25_inst : DFFR_X1 port map( D => n8114, CK => CLK, RN => 
                           n12542, Q => n_2204, QN => n5912);
   REGISTERS_reg_56_24_inst : DFFR_X1 port map( D => n8115, CK => CLK, RN => 
                           n12479, Q => n_2205, QN => n5944);
   REGISTERS_reg_56_23_inst : DFFR_X1 port map( D => n8116, CK => CLK, RN => 
                           n12630, Q => n_2206, QN => n6008);
   REGISTERS_reg_56_22_inst : DFFR_X1 port map( D => n8117, CK => CLK, RN => 
                           n12520, Q => n_2207, QN => n9143);
   REGISTERS_reg_56_21_inst : DFFR_X1 port map( D => n8118, CK => CLK, RN => 
                           n12528, Q => n_2208, QN => n9175);
   REGISTERS_reg_56_20_inst : DFFR_X1 port map( D => n8119, CK => CLK, RN => 
                           n12502, Q => n_2209, QN => n9207);
   REGISTERS_reg_56_19_inst : DFFR_X1 port map( D => n8120, CK => CLK, RN => 
                           n12594, Q => n_2210, QN => n9573);
   REGISTERS_reg_56_18_inst : DFFR_X1 port map( D => n8121, CK => CLK, RN => 
                           n12445, Q => n_2211, QN => n9605);
   REGISTERS_reg_56_17_inst : DFFR_X1 port map( D => n8122, CK => CLK, RN => 
                           n12452, Q => n_2212, QN => n9637);
   REGISTERS_reg_56_16_inst : DFFR_X1 port map( D => n8123, CK => CLK, RN => 
                           n12458, Q => n_2213, QN => n9701);
   REGISTERS_reg_56_15_inst : DFFR_X1 port map( D => n8124, CK => CLK, RN => 
                           n12638, Q => n_2214, QN => n10031);
   REGISTERS_reg_56_14_inst : DFFR_X1 port map( D => n8125, CK => CLK, RN => 
                           n12466, Q => n_2215, QN => n10063);
   REGISTERS_reg_56_13_inst : DFFR_X1 port map( D => n8126, CK => CLK, RN => 
                           n12473, Q => n_2216, QN => n10095);
   REGISTERS_reg_56_12_inst : DFFR_X1 port map( D => n8127, CK => CLK, RN => 
                           n12480, Q => n_2217, QN => n10127);
   REGISTERS_reg_56_11_inst : DFFR_X1 port map( D => n8128, CK => CLK, RN => 
                           n12572, Q => n_2218, QN => n10159);
   REGISTERS_reg_56_10_inst : DFFR_X1 port map( D => n8129, CK => CLK, RN => 
                           n12550, Q => n_2219, QN => n10191);
   REGISTERS_reg_56_9_inst : DFFR_X1 port map( D => n8130, CK => CLK, RN => 
                           n12557, Q => n_2220, QN => n10225);
   REGISTERS_reg_56_8_inst : DFFR_X1 port map( D => n8131, CK => CLK, RN => 
                           n12535, Q => n_2221, QN => n10257);
   REGISTERS_reg_56_7_inst : DFFR_X1 port map( D => n8132, CK => CLK, RN => 
                           n12645, Q => n_2222, QN => n10289);
   REGISTERS_reg_56_6_inst : DFFR_X1 port map( D => n8133, CK => CLK, RN => 
                           n12601, Q => n_2223, QN => n10324);
   REGISTERS_reg_56_5_inst : DFFR_X1 port map( D => n8134, CK => CLK, RN => 
                           n12488, Q => n_2224, QN => n10356);
   REGISTERS_reg_56_4_inst : DFFR_X1 port map( D => n8135, CK => CLK, RN => 
                           n12495, Q => n_2225, QN => n10388);
   REGISTERS_reg_56_3_inst : DFFR_X1 port map( D => n8136, CK => CLK, RN => 
                           n12579, Q => n_2226, QN => n10423);
   REGISTERS_reg_56_2_inst : DFFR_X1 port map( D => n8137, CK => CLK, RN => 
                           n12510, Q => n_2227, QN => n10455);
   REGISTERS_reg_56_1_inst : DFFR_X1 port map( D => n8138, CK => CLK, RN => 
                           n12437, Q => n_2228, QN => n10487);
   REGISTERS_reg_56_0_inst : DFFR_X1 port map( D => n8139, CK => CLK, RN => 
                           n12652, Q => n_2229, QN => n10519);
   REGISTERS_reg_57_31_inst : DFFR_X1 port map( D => n8140, CK => CLK, RN => 
                           n12660, Q => n_2230, QN => n5718);
   REGISTERS_reg_57_30_inst : DFFR_X1 port map( D => n8141, CK => CLK, RN => 
                           n12623, Q => n_2231, QN => n5750);
   REGISTERS_reg_57_29_inst : DFFR_X1 port map( D => n8142, CK => CLK, RN => 
                           n12608, Q => n_2232, QN => n5782);
   REGISTERS_reg_57_28_inst : DFFR_X1 port map( D => n8143, CK => CLK, RN => 
                           n12616, Q => n_2233, QN => n5814);
   REGISTERS_reg_57_27_inst : DFFR_X1 port map( D => n8144, CK => CLK, RN => 
                           n12586, Q => n_2234, QN => n5846);
   REGISTERS_reg_57_26_inst : DFFR_X1 port map( D => n8145, CK => CLK, RN => 
                           n12564, Q => n_2235, QN => n5878);
   REGISTERS_reg_57_25_inst : DFFR_X1 port map( D => n8146, CK => CLK, RN => 
                           n12542, Q => n_2236, QN => n5910);
   REGISTERS_reg_57_24_inst : DFFR_X1 port map( D => n8147, CK => CLK, RN => 
                           n12478, Q => n_2237, QN => n5942);
   REGISTERS_reg_57_23_inst : DFFR_X1 port map( D => n8148, CK => CLK, RN => 
                           n12630, Q => n_2238, QN => n6006);
   REGISTERS_reg_57_22_inst : DFFR_X1 port map( D => n8149, CK => CLK, RN => 
                           n12520, Q => n_2239, QN => n9141);
   REGISTERS_reg_57_21_inst : DFFR_X1 port map( D => n8150, CK => CLK, RN => 
                           n12528, Q => n_2240, QN => n9173);
   REGISTERS_reg_57_20_inst : DFFR_X1 port map( D => n8151, CK => CLK, RN => 
                           n12502, Q => n_2241, QN => n9205);
   REGISTERS_reg_57_19_inst : DFFR_X1 port map( D => n8152, CK => CLK, RN => 
                           n12594, Q => n_2242, QN => n9571);
   REGISTERS_reg_57_18_inst : DFFR_X1 port map( D => n8153, CK => CLK, RN => 
                           n12445, Q => n_2243, QN => n9603);
   REGISTERS_reg_57_17_inst : DFFR_X1 port map( D => n8154, CK => CLK, RN => 
                           n12452, Q => n_2244, QN => n9635);
   REGISTERS_reg_57_16_inst : DFFR_X1 port map( D => n8155, CK => CLK, RN => 
                           n12458, Q => n_2245, QN => n9699);
   REGISTERS_reg_57_15_inst : DFFR_X1 port map( D => n8156, CK => CLK, RN => 
                           n12638, Q => n_2246, QN => n10029);
   REGISTERS_reg_57_14_inst : DFFR_X1 port map( D => n8157, CK => CLK, RN => 
                           n12466, Q => n_2247, QN => n10061);
   REGISTERS_reg_57_13_inst : DFFR_X1 port map( D => n8158, CK => CLK, RN => 
                           n12473, Q => n_2248, QN => n10093);
   REGISTERS_reg_57_12_inst : DFFR_X1 port map( D => n8159, CK => CLK, RN => 
                           n12480, Q => n_2249, QN => n10125);
   REGISTERS_reg_57_11_inst : DFFR_X1 port map( D => n8160, CK => CLK, RN => 
                           n12572, Q => n_2250, QN => n10157);
   REGISTERS_reg_57_10_inst : DFFR_X1 port map( D => n8161, CK => CLK, RN => 
                           n12550, Q => n_2251, QN => n10189);
   REGISTERS_reg_57_9_inst : DFFR_X1 port map( D => n8162, CK => CLK, RN => 
                           n12557, Q => n_2252, QN => n10223);
   REGISTERS_reg_57_8_inst : DFFR_X1 port map( D => n8163, CK => CLK, RN => 
                           n12535, Q => n_2253, QN => n10255);
   REGISTERS_reg_57_7_inst : DFFR_X1 port map( D => n8164, CK => CLK, RN => 
                           n12645, Q => n_2254, QN => n10287);
   REGISTERS_reg_57_6_inst : DFFR_X1 port map( D => n8165, CK => CLK, RN => 
                           n12601, Q => n_2255, QN => n10322);
   REGISTERS_reg_57_5_inst : DFFR_X1 port map( D => n8166, CK => CLK, RN => 
                           n12488, Q => n_2256, QN => n10354);
   REGISTERS_reg_57_4_inst : DFFR_X1 port map( D => n8167, CK => CLK, RN => 
                           n12495, Q => n_2257, QN => n10386);
   REGISTERS_reg_57_3_inst : DFFR_X1 port map( D => n8168, CK => CLK, RN => 
                           n12579, Q => n_2258, QN => n10421);
   REGISTERS_reg_57_2_inst : DFFR_X1 port map( D => n8169, CK => CLK, RN => 
                           n12510, Q => n_2259, QN => n10453);
   REGISTERS_reg_57_1_inst : DFFR_X1 port map( D => n8170, CK => CLK, RN => 
                           n12437, Q => n_2260, QN => n10485);
   REGISTERS_reg_57_0_inst : DFFR_X1 port map( D => n8171, CK => CLK, RN => 
                           n12652, Q => n_2261, QN => n10517);
   REGISTERS_reg_58_31_inst : DFFR_X1 port map( D => n8172, CK => CLK, RN => 
                           n12660, Q => n_2262, QN => n5719);
   REGISTERS_reg_58_30_inst : DFFR_X1 port map( D => n8173, CK => CLK, RN => 
                           n12623, Q => n_2263, QN => n5751);
   REGISTERS_reg_58_29_inst : DFFR_X1 port map( D => n8174, CK => CLK, RN => 
                           n12608, Q => n_2264, QN => n5783);
   REGISTERS_reg_58_28_inst : DFFR_X1 port map( D => n8175, CK => CLK, RN => 
                           n12616, Q => n_2265, QN => n5815);
   REGISTERS_reg_58_27_inst : DFFR_X1 port map( D => n8176, CK => CLK, RN => 
                           n12586, Q => n_2266, QN => n5847);
   REGISTERS_reg_58_26_inst : DFFR_X1 port map( D => n8177, CK => CLK, RN => 
                           n12564, Q => n_2267, QN => n5879);
   REGISTERS_reg_58_25_inst : DFFR_X1 port map( D => n8178, CK => CLK, RN => 
                           n12542, Q => n_2268, QN => n5911);
   REGISTERS_reg_58_24_inst : DFFR_X1 port map( D => n8179, CK => CLK, RN => 
                           n12477, Q => n_2269, QN => n5943);
   REGISTERS_reg_58_23_inst : DFFR_X1 port map( D => n8180, CK => CLK, RN => 
                           n12630, Q => n_2270, QN => n6007);
   REGISTERS_reg_58_22_inst : DFFR_X1 port map( D => n8181, CK => CLK, RN => 
                           n12520, Q => n_2271, QN => n9142);
   REGISTERS_reg_58_21_inst : DFFR_X1 port map( D => n8182, CK => CLK, RN => 
                           n12528, Q => n_2272, QN => n9174);
   REGISTERS_reg_58_20_inst : DFFR_X1 port map( D => n8183, CK => CLK, RN => 
                           n12502, Q => n_2273, QN => n9206);
   REGISTERS_reg_58_19_inst : DFFR_X1 port map( D => n8184, CK => CLK, RN => 
                           n12594, Q => n_2274, QN => n9572);
   REGISTERS_reg_58_18_inst : DFFR_X1 port map( D => n8185, CK => CLK, RN => 
                           n12445, Q => n_2275, QN => n9604);
   REGISTERS_reg_58_17_inst : DFFR_X1 port map( D => n8186, CK => CLK, RN => 
                           n12452, Q => n_2276, QN => n9636);
   REGISTERS_reg_58_16_inst : DFFR_X1 port map( D => n8187, CK => CLK, RN => 
                           n12458, Q => n_2277, QN => n9700);
   REGISTERS_reg_58_15_inst : DFFR_X1 port map( D => n8188, CK => CLK, RN => 
                           n12638, Q => n_2278, QN => n10030);
   REGISTERS_reg_58_14_inst : DFFR_X1 port map( D => n8189, CK => CLK, RN => 
                           n12466, Q => n_2279, QN => n10062);
   REGISTERS_reg_58_13_inst : DFFR_X1 port map( D => n8190, CK => CLK, RN => 
                           n12473, Q => n_2280, QN => n10094);
   REGISTERS_reg_58_12_inst : DFFR_X1 port map( D => n8191, CK => CLK, RN => 
                           n12480, Q => n_2281, QN => n10126);
   REGISTERS_reg_58_11_inst : DFFR_X1 port map( D => n8192, CK => CLK, RN => 
                           n12572, Q => n_2282, QN => n10158);
   REGISTERS_reg_58_10_inst : DFFR_X1 port map( D => n8193, CK => CLK, RN => 
                           n12550, Q => n_2283, QN => n10190);
   REGISTERS_reg_58_9_inst : DFFR_X1 port map( D => n8194, CK => CLK, RN => 
                           n12557, Q => n_2284, QN => n10224);
   REGISTERS_reg_58_8_inst : DFFR_X1 port map( D => n8195, CK => CLK, RN => 
                           n12535, Q => n_2285, QN => n10256);
   REGISTERS_reg_58_7_inst : DFFR_X1 port map( D => n8196, CK => CLK, RN => 
                           n12645, Q => n_2286, QN => n10288);
   REGISTERS_reg_58_6_inst : DFFR_X1 port map( D => n8197, CK => CLK, RN => 
                           n12601, Q => n_2287, QN => n10323);
   REGISTERS_reg_58_5_inst : DFFR_X1 port map( D => n8198, CK => CLK, RN => 
                           n12488, Q => n_2288, QN => n10355);
   REGISTERS_reg_58_4_inst : DFFR_X1 port map( D => n8199, CK => CLK, RN => 
                           n12495, Q => n_2289, QN => n10387);
   REGISTERS_reg_58_3_inst : DFFR_X1 port map( D => n8200, CK => CLK, RN => 
                           n12579, Q => n_2290, QN => n10422);
   REGISTERS_reg_58_2_inst : DFFR_X1 port map( D => n8201, CK => CLK, RN => 
                           n12510, Q => n_2291, QN => n10454);
   REGISTERS_reg_58_1_inst : DFFR_X1 port map( D => n8202, CK => CLK, RN => 
                           n12437, Q => n_2292, QN => n10486);
   REGISTERS_reg_58_0_inst : DFFR_X1 port map( D => n8203, CK => CLK, RN => 
                           n12652, Q => n_2293, QN => n10518);
   REGISTERS_reg_59_31_inst : DFFR_X1 port map( D => n8204, CK => CLK, RN => 
                           n12660, Q => n_2294, QN => n5717);
   REGISTERS_reg_59_30_inst : DFFR_X1 port map( D => n8205, CK => CLK, RN => 
                           n12623, Q => n_2295, QN => n5749);
   REGISTERS_reg_59_29_inst : DFFR_X1 port map( D => n8206, CK => CLK, RN => 
                           n12608, Q => n_2296, QN => n5781);
   REGISTERS_reg_59_28_inst : DFFR_X1 port map( D => n8207, CK => CLK, RN => 
                           n12616, Q => n_2297, QN => n5813);
   REGISTERS_reg_59_27_inst : DFFR_X1 port map( D => n8208, CK => CLK, RN => 
                           n12586, Q => n_2298, QN => n5845);
   REGISTERS_reg_59_26_inst : DFFR_X1 port map( D => n8209, CK => CLK, RN => 
                           n12564, Q => n_2299, QN => n5877);
   REGISTERS_reg_59_25_inst : DFFR_X1 port map( D => n8210, CK => CLK, RN => 
                           n12542, Q => n_2300, QN => n5909);
   REGISTERS_reg_59_24_inst : DFFR_X1 port map( D => n8211, CK => CLK, RN => 
                           n12476, Q => n_2301, QN => n5941);
   REGISTERS_reg_59_23_inst : DFFR_X1 port map( D => n8212, CK => CLK, RN => 
                           n12630, Q => n_2302, QN => n6005);
   REGISTERS_reg_59_22_inst : DFFR_X1 port map( D => n8213, CK => CLK, RN => 
                           n12520, Q => n_2303, QN => n9140);
   REGISTERS_reg_59_21_inst : DFFR_X1 port map( D => n8214, CK => CLK, RN => 
                           n12528, Q => n_2304, QN => n9172);
   REGISTERS_reg_59_20_inst : DFFR_X1 port map( D => n8215, CK => CLK, RN => 
                           n12502, Q => n_2305, QN => n9204);
   REGISTERS_reg_59_19_inst : DFFR_X1 port map( D => n8216, CK => CLK, RN => 
                           n12594, Q => n_2306, QN => n9570);
   REGISTERS_reg_59_18_inst : DFFR_X1 port map( D => n8217, CK => CLK, RN => 
                           n12445, Q => n_2307, QN => n9602);
   REGISTERS_reg_59_17_inst : DFFR_X1 port map( D => n8218, CK => CLK, RN => 
                           n12452, Q => n_2308, QN => n9634);
   REGISTERS_reg_59_16_inst : DFFR_X1 port map( D => n8219, CK => CLK, RN => 
                           n12458, Q => n_2309, QN => n9698);
   REGISTERS_reg_59_15_inst : DFFR_X1 port map( D => n8220, CK => CLK, RN => 
                           n12638, Q => n_2310, QN => n10028);
   REGISTERS_reg_59_14_inst : DFFR_X1 port map( D => n8221, CK => CLK, RN => 
                           n12466, Q => n_2311, QN => n10060);
   REGISTERS_reg_59_13_inst : DFFR_X1 port map( D => n8222, CK => CLK, RN => 
                           n12473, Q => n_2312, QN => n10092);
   REGISTERS_reg_59_12_inst : DFFR_X1 port map( D => n8223, CK => CLK, RN => 
                           n12480, Q => n_2313, QN => n10124);
   REGISTERS_reg_59_11_inst : DFFR_X1 port map( D => n8224, CK => CLK, RN => 
                           n12572, Q => n_2314, QN => n10156);
   REGISTERS_reg_59_10_inst : DFFR_X1 port map( D => n8225, CK => CLK, RN => 
                           n12550, Q => n_2315, QN => n10188);
   REGISTERS_reg_59_9_inst : DFFR_X1 port map( D => n8226, CK => CLK, RN => 
                           n12557, Q => n_2316, QN => n10222);
   REGISTERS_reg_59_8_inst : DFFR_X1 port map( D => n8227, CK => CLK, RN => 
                           n12535, Q => n_2317, QN => n10254);
   REGISTERS_reg_59_7_inst : DFFR_X1 port map( D => n8228, CK => CLK, RN => 
                           n12645, Q => n_2318, QN => n10286);
   REGISTERS_reg_59_6_inst : DFFR_X1 port map( D => n8229, CK => CLK, RN => 
                           n12601, Q => n_2319, QN => n10321);
   REGISTERS_reg_59_5_inst : DFFR_X1 port map( D => n8230, CK => CLK, RN => 
                           n12488, Q => n_2320, QN => n10353);
   REGISTERS_reg_59_4_inst : DFFR_X1 port map( D => n8231, CK => CLK, RN => 
                           n12495, Q => n_2321, QN => n10385);
   REGISTERS_reg_59_3_inst : DFFR_X1 port map( D => n8232, CK => CLK, RN => 
                           n12579, Q => n_2322, QN => n10420);
   REGISTERS_reg_59_2_inst : DFFR_X1 port map( D => n8233, CK => CLK, RN => 
                           n12510, Q => n_2323, QN => n10452);
   REGISTERS_reg_59_1_inst : DFFR_X1 port map( D => n8234, CK => CLK, RN => 
                           n12437, Q => n_2324, QN => n10484);
   REGISTERS_reg_59_0_inst : DFFR_X1 port map( D => n8235, CK => CLK, RN => 
                           n12652, Q => n_2325, QN => n10516);
   REGISTERS_reg_60_31_inst : DFFR_X1 port map( D => n8236, CK => CLK, RN => 
                           n12660, Q => n_2326, QN => n5715);
   REGISTERS_reg_60_30_inst : DFFR_X1 port map( D => n8237, CK => CLK, RN => 
                           n12623, Q => n_2327, QN => n5747);
   REGISTERS_reg_60_29_inst : DFFR_X1 port map( D => n8238, CK => CLK, RN => 
                           n12609, Q => n_2328, QN => n5779);
   REGISTERS_reg_60_28_inst : DFFR_X1 port map( D => n8239, CK => CLK, RN => 
                           n12616, Q => n_2329, QN => n5811);
   REGISTERS_reg_60_27_inst : DFFR_X1 port map( D => n8240, CK => CLK, RN => 
                           n12587, Q => n_2330, QN => n5843);
   REGISTERS_reg_60_26_inst : DFFR_X1 port map( D => n8241, CK => CLK, RN => 
                           n12565, Q => n_2331, QN => n5875);
   REGISTERS_reg_60_25_inst : DFFR_X1 port map( D => n8242, CK => CLK, RN => 
                           n12543, Q => n_2332, QN => n5907);
   REGISTERS_reg_60_24_inst : DFFR_X1 port map( D => n8243, CK => CLK, RN => 
                           n12475, Q => n_2333, QN => n5939);
   REGISTERS_reg_60_23_inst : DFFR_X1 port map( D => n8244, CK => CLK, RN => 
                           n12631, Q => n_2334, QN => n6003);
   REGISTERS_reg_60_22_inst : DFFR_X1 port map( D => n8245, CK => CLK, RN => 
                           n12521, Q => n_2335, QN => n9138);
   REGISTERS_reg_60_21_inst : DFFR_X1 port map( D => n8246, CK => CLK, RN => 
                           n12528, Q => n_2336, QN => n9170);
   REGISTERS_reg_60_20_inst : DFFR_X1 port map( D => n8247, CK => CLK, RN => 
                           n12503, Q => n_2337, QN => n9202);
   REGISTERS_reg_60_19_inst : DFFR_X1 port map( D => n8248, CK => CLK, RN => 
                           n12594, Q => n_2338, QN => n9568);
   REGISTERS_reg_60_18_inst : DFFR_X1 port map( D => n8249, CK => CLK, RN => 
                           n12445, Q => n_2339, QN => n9600);
   REGISTERS_reg_60_17_inst : DFFR_X1 port map( D => n8250, CK => CLK, RN => 
                           n12452, Q => n_2340, QN => n9632);
   REGISTERS_reg_60_16_inst : DFFR_X1 port map( D => n8251, CK => CLK, RN => 
                           n12459, Q => n_2341, QN => n9696);
   REGISTERS_reg_60_15_inst : DFFR_X1 port map( D => n8252, CK => CLK, RN => 
                           n12638, Q => n_2342, QN => n10026);
   REGISTERS_reg_60_14_inst : DFFR_X1 port map( D => n8253, CK => CLK, RN => 
                           n12466, Q => n_2343, QN => n10058);
   REGISTERS_reg_60_13_inst : DFFR_X1 port map( D => n8254, CK => CLK, RN => 
                           n12473, Q => n_2344, QN => n10090);
   REGISTERS_reg_60_12_inst : DFFR_X1 port map( D => n8255, CK => CLK, RN => 
                           n12481, Q => n_2345, QN => n10122);
   REGISTERS_reg_60_11_inst : DFFR_X1 port map( D => n8256, CK => CLK, RN => 
                           n12572, Q => n_2346, QN => n10154);
   REGISTERS_reg_60_10_inst : DFFR_X1 port map( D => n8257, CK => CLK, RN => 
                           n12550, Q => n_2347, QN => n10186);
   REGISTERS_reg_60_9_inst : DFFR_X1 port map( D => n8258, CK => CLK, RN => 
                           n12557, Q => n_2348, QN => n10220);
   REGISTERS_reg_60_8_inst : DFFR_X1 port map( D => n8259, CK => CLK, RN => 
                           n12535, Q => n_2349, QN => n10252);
   REGISTERS_reg_60_7_inst : DFFR_X1 port map( D => n8260, CK => CLK, RN => 
                           n12645, Q => n_2350, QN => n10284);
   REGISTERS_reg_60_6_inst : DFFR_X1 port map( D => n8261, CK => CLK, RN => 
                           n12601, Q => n_2351, QN => n10319);
   REGISTERS_reg_60_5_inst : DFFR_X1 port map( D => n8262, CK => CLK, RN => 
                           n12488, Q => n_2352, QN => n10351);
   REGISTERS_reg_60_4_inst : DFFR_X1 port map( D => n8263, CK => CLK, RN => 
                           n12495, Q => n_2353, QN => n10383);
   REGISTERS_reg_60_3_inst : DFFR_X1 port map( D => n8264, CK => CLK, RN => 
                           n12579, Q => n_2354, QN => n10418);
   REGISTERS_reg_60_2_inst : DFFR_X1 port map( D => n8265, CK => CLK, RN => 
                           n12510, Q => n_2355, QN => n10450);
   REGISTERS_reg_60_1_inst : DFFR_X1 port map( D => n8266, CK => CLK, RN => 
                           n12438, Q => n_2356, QN => n10482);
   REGISTERS_reg_60_0_inst : DFFR_X1 port map( D => n8267, CK => CLK, RN => 
                           n12653, Q => n_2357, QN => n10514);
   REGISTERS_reg_61_31_inst : DFFR_X1 port map( D => n8268, CK => CLK, RN => 
                           n12660, Q => n_2358, QN => n13844);
   REGISTERS_reg_61_30_inst : DFFR_X1 port map( D => n8269, CK => CLK, RN => 
                           n12623, Q => n_2359, QN => n13845);
   REGISTERS_reg_61_29_inst : DFFR_X1 port map( D => n8270, CK => CLK, RN => 
                           n12609, Q => n_2360, QN => n13846);
   REGISTERS_reg_61_28_inst : DFFR_X1 port map( D => n8271, CK => CLK, RN => 
                           n12616, Q => n_2361, QN => n13847);
   REGISTERS_reg_61_27_inst : DFFR_X1 port map( D => n8272, CK => CLK, RN => 
                           n12587, Q => n_2362, QN => n13848);
   REGISTERS_reg_61_26_inst : DFFR_X1 port map( D => n8273, CK => CLK, RN => 
                           n12565, Q => n_2363, QN => n13849);
   REGISTERS_reg_61_25_inst : DFFR_X1 port map( D => n8274, CK => CLK, RN => 
                           n12543, Q => n_2364, QN => n13850);
   REGISTERS_reg_61_24_inst : DFFR_X1 port map( D => n8275, CK => CLK, RN => 
                           n12488, Q => n_2365, QN => n13851);
   REGISTERS_reg_61_23_inst : DFFR_X1 port map( D => n8276, CK => CLK, RN => 
                           n12631, Q => n_2366, QN => n13852);
   REGISTERS_reg_61_22_inst : DFFR_X1 port map( D => n8277, CK => CLK, RN => 
                           n12521, Q => n_2367, QN => n13853);
   REGISTERS_reg_61_21_inst : DFFR_X1 port map( D => n8278, CK => CLK, RN => 
                           n12528, Q => n_2368, QN => n13854);
   REGISTERS_reg_61_20_inst : DFFR_X1 port map( D => n8279, CK => CLK, RN => 
                           n12503, Q => n_2369, QN => n13855);
   REGISTERS_reg_61_19_inst : DFFR_X1 port map( D => n8280, CK => CLK, RN => 
                           n12594, Q => n_2370, QN => n13856);
   REGISTERS_reg_61_18_inst : DFFR_X1 port map( D => n8281, CK => CLK, RN => 
                           n12445, Q => n_2371, QN => n13857);
   REGISTERS_reg_61_17_inst : DFFR_X1 port map( D => n8282, CK => CLK, RN => 
                           n12452, Q => n_2372, QN => n13858);
   REGISTERS_reg_61_16_inst : DFFR_X1 port map( D => n8283, CK => CLK, RN => 
                           n12459, Q => n_2373, QN => n13859);
   REGISTERS_reg_61_15_inst : DFFR_X1 port map( D => n8284, CK => CLK, RN => 
                           n12638, Q => n_2374, QN => n13860);
   REGISTERS_reg_61_14_inst : DFFR_X1 port map( D => n8285, CK => CLK, RN => 
                           n12466, Q => n_2375, QN => n13861);
   REGISTERS_reg_61_13_inst : DFFR_X1 port map( D => n8286, CK => CLK, RN => 
                           n12473, Q => n_2376, QN => n13862);
   REGISTERS_reg_61_12_inst : DFFR_X1 port map( D => n8287, CK => CLK, RN => 
                           n12481, Q => n_2377, QN => n13863);
   REGISTERS_reg_61_11_inst : DFFR_X1 port map( D => n8288, CK => CLK, RN => 
                           n12572, Q => n_2378, QN => n13864);
   REGISTERS_reg_61_10_inst : DFFR_X1 port map( D => n8289, CK => CLK, RN => 
                           n12550, Q => n_2379, QN => n13865);
   REGISTERS_reg_61_9_inst : DFFR_X1 port map( D => n8290, CK => CLK, RN => 
                           n12557, Q => n_2380, QN => n13866);
   REGISTERS_reg_61_8_inst : DFFR_X1 port map( D => n8291, CK => CLK, RN => 
                           n12535, Q => n_2381, QN => n13867);
   REGISTERS_reg_61_7_inst : DFFR_X1 port map( D => n8292, CK => CLK, RN => 
                           n12645, Q => n_2382, QN => n13868);
   REGISTERS_reg_61_6_inst : DFFR_X1 port map( D => n8293, CK => CLK, RN => 
                           n12601, Q => n_2383, QN => n13869);
   REGISTERS_reg_61_5_inst : DFFR_X1 port map( D => n8294, CK => CLK, RN => 
                           n12488, Q => n_2384, QN => n13870);
   REGISTERS_reg_61_4_inst : DFFR_X1 port map( D => n8295, CK => CLK, RN => 
                           n12495, Q => n_2385, QN => n13871);
   REGISTERS_reg_61_3_inst : DFFR_X1 port map( D => n8296, CK => CLK, RN => 
                           n12579, Q => n_2386, QN => n13872);
   REGISTERS_reg_61_2_inst : DFFR_X1 port map( D => n8297, CK => CLK, RN => 
                           n12510, Q => n_2387, QN => n13873);
   REGISTERS_reg_61_1_inst : DFFR_X1 port map( D => n8298, CK => CLK, RN => 
                           n12438, Q => n_2388, QN => n13874);
   REGISTERS_reg_61_0_inst : DFFR_X1 port map( D => n8299, CK => CLK, RN => 
                           n12653, Q => n_2389, QN => n13875);
   REGISTERS_reg_62_31_inst : DFFR_X1 port map( D => n8300, CK => CLK, RN => 
                           n12660, Q => n_2390, QN => n5716);
   REGISTERS_reg_62_30_inst : DFFR_X1 port map( D => n8301, CK => CLK, RN => 
                           n12623, Q => n_2391, QN => n5748);
   REGISTERS_reg_62_29_inst : DFFR_X1 port map( D => n8302, CK => CLK, RN => 
                           n12609, Q => n_2392, QN => n5780);
   REGISTERS_reg_62_28_inst : DFFR_X1 port map( D => n8303, CK => CLK, RN => 
                           n12616, Q => n_2393, QN => n5812);
   REGISTERS_reg_62_27_inst : DFFR_X1 port map( D => n8304, CK => CLK, RN => 
                           n12587, Q => n_2394, QN => n5844);
   REGISTERS_reg_62_26_inst : DFFR_X1 port map( D => n8305, CK => CLK, RN => 
                           n12565, Q => n_2395, QN => n5876);
   REGISTERS_reg_62_25_inst : DFFR_X1 port map( D => n8306, CK => CLK, RN => 
                           n12543, Q => n_2396, QN => n5908);
   REGISTERS_reg_62_24_inst : DFFR_X1 port map( D => n8307, CK => CLK, RN => 
                           n12487, Q => n_2397, QN => n5940);
   REGISTERS_reg_62_23_inst : DFFR_X1 port map( D => n8308, CK => CLK, RN => 
                           n12631, Q => n_2398, QN => n6004);
   REGISTERS_reg_62_22_inst : DFFR_X1 port map( D => n8309, CK => CLK, RN => 
                           n12521, Q => n_2399, QN => n9139);
   REGISTERS_reg_62_21_inst : DFFR_X1 port map( D => n8310, CK => CLK, RN => 
                           n12528, Q => n_2400, QN => n9171);
   REGISTERS_reg_62_20_inst : DFFR_X1 port map( D => n8311, CK => CLK, RN => 
                           n12503, Q => n_2401, QN => n9203);
   REGISTERS_reg_62_19_inst : DFFR_X1 port map( D => n8312, CK => CLK, RN => 
                           n12594, Q => n_2402, QN => n9569);
   REGISTERS_reg_62_18_inst : DFFR_X1 port map( D => n8313, CK => CLK, RN => 
                           n12445, Q => n_2403, QN => n9601);
   REGISTERS_reg_62_17_inst : DFFR_X1 port map( D => n8314, CK => CLK, RN => 
                           n12452, Q => n_2404, QN => n9633);
   REGISTERS_reg_62_16_inst : DFFR_X1 port map( D => n8315, CK => CLK, RN => 
                           n12459, Q => n_2405, QN => n9697);
   REGISTERS_reg_62_15_inst : DFFR_X1 port map( D => n8316, CK => CLK, RN => 
                           n12638, Q => n_2406, QN => n10027);
   REGISTERS_reg_62_14_inst : DFFR_X1 port map( D => n8317, CK => CLK, RN => 
                           n12466, Q => n_2407, QN => n10059);
   REGISTERS_reg_62_13_inst : DFFR_X1 port map( D => n8318, CK => CLK, RN => 
                           n12473, Q => n_2408, QN => n10091);
   REGISTERS_reg_62_12_inst : DFFR_X1 port map( D => n8319, CK => CLK, RN => 
                           n12481, Q => n_2409, QN => n10123);
   REGISTERS_reg_62_11_inst : DFFR_X1 port map( D => n8320, CK => CLK, RN => 
                           n12572, Q => n_2410, QN => n10155);
   REGISTERS_reg_62_10_inst : DFFR_X1 port map( D => n8321, CK => CLK, RN => 
                           n12550, Q => n_2411, QN => n10187);
   REGISTERS_reg_62_9_inst : DFFR_X1 port map( D => n8322, CK => CLK, RN => 
                           n12557, Q => n_2412, QN => n10221);
   REGISTERS_reg_62_8_inst : DFFR_X1 port map( D => n8323, CK => CLK, RN => 
                           n12535, Q => n_2413, QN => n10253);
   REGISTERS_reg_62_7_inst : DFFR_X1 port map( D => n8324, CK => CLK, RN => 
                           n12645, Q => n_2414, QN => n10285);
   REGISTERS_reg_62_6_inst : DFFR_X1 port map( D => n8325, CK => CLK, RN => 
                           n12601, Q => n_2415, QN => n10320);
   REGISTERS_reg_62_5_inst : DFFR_X1 port map( D => n8326, CK => CLK, RN => 
                           n12488, Q => n_2416, QN => n10352);
   REGISTERS_reg_62_4_inst : DFFR_X1 port map( D => n8327, CK => CLK, RN => 
                           n12495, Q => n_2417, QN => n10384);
   REGISTERS_reg_62_3_inst : DFFR_X1 port map( D => n8328, CK => CLK, RN => 
                           n12579, Q => n_2418, QN => n10419);
   REGISTERS_reg_62_2_inst : DFFR_X1 port map( D => n8329, CK => CLK, RN => 
                           n12510, Q => n_2419, QN => n10451);
   REGISTERS_reg_62_1_inst : DFFR_X1 port map( D => n8330, CK => CLK, RN => 
                           n12438, Q => n_2420, QN => n10483);
   REGISTERS_reg_62_0_inst : DFFR_X1 port map( D => n8331, CK => CLK, RN => 
                           n12653, Q => n_2421, QN => n10515);
   REGISTERS_reg_63_31_inst : DFFR_X1 port map( D => n8332, CK => CLK, RN => 
                           n12660, Q => n_2422, QN => n13876);
   REGISTERS_reg_63_30_inst : DFFR_X1 port map( D => n8333, CK => CLK, RN => 
                           n12623, Q => n_2423, QN => n13877);
   REGISTERS_reg_63_29_inst : DFFR_X1 port map( D => n8334, CK => CLK, RN => 
                           n12609, Q => n_2424, QN => n13878);
   REGISTERS_reg_63_28_inst : DFFR_X1 port map( D => n8335, CK => CLK, RN => 
                           n12616, Q => n_2425, QN => n13879);
   REGISTERS_reg_63_27_inst : DFFR_X1 port map( D => n8336, CK => CLK, RN => 
                           n12587, Q => n_2426, QN => n13880);
   REGISTERS_reg_63_26_inst : DFFR_X1 port map( D => n8337, CK => CLK, RN => 
                           n12565, Q => n_2427, QN => n13881);
   REGISTERS_reg_63_25_inst : DFFR_X1 port map( D => n8338, CK => CLK, RN => 
                           n12543, Q => n_2428, QN => n13882);
   REGISTERS_reg_63_24_inst : DFFR_X1 port map( D => n8339, CK => CLK, RN => 
                           n12464, Q => n_2429, QN => n13883);
   REGISTERS_reg_63_23_inst : DFFR_X1 port map( D => n8340, CK => CLK, RN => 
                           n12631, Q => n_2430, QN => n13884);
   REGISTERS_reg_63_22_inst : DFFR_X1 port map( D => n8341, CK => CLK, RN => 
                           n12521, Q => n_2431, QN => n13885);
   REGISTERS_reg_63_21_inst : DFFR_X1 port map( D => n8342, CK => CLK, RN => 
                           n12528, Q => n_2432, QN => n13886);
   REGISTERS_reg_63_20_inst : DFFR_X1 port map( D => n8343, CK => CLK, RN => 
                           n12503, Q => n_2433, QN => n13887);
   REGISTERS_reg_63_19_inst : DFFR_X1 port map( D => n8344, CK => CLK, RN => 
                           n12594, Q => n_2434, QN => n13888);
   REGISTERS_reg_63_18_inst : DFFR_X1 port map( D => n8345, CK => CLK, RN => 
                           n12445, Q => n_2435, QN => n13889);
   REGISTERS_reg_63_17_inst : DFFR_X1 port map( D => n8346, CK => CLK, RN => 
                           n12452, Q => n_2436, QN => n13890);
   REGISTERS_reg_63_16_inst : DFFR_X1 port map( D => n8347, CK => CLK, RN => 
                           n12459, Q => n_2437, QN => n13891);
   REGISTERS_reg_63_15_inst : DFFR_X1 port map( D => n8348, CK => CLK, RN => 
                           n12638, Q => n_2438, QN => n13892);
   REGISTERS_reg_63_14_inst : DFFR_X1 port map( D => n8349, CK => CLK, RN => 
                           n12466, Q => n_2439, QN => n13893);
   REGISTERS_reg_63_13_inst : DFFR_X1 port map( D => n8350, CK => CLK, RN => 
                           n12473, Q => n_2440, QN => n13894);
   REGISTERS_reg_63_12_inst : DFFR_X1 port map( D => n8351, CK => CLK, RN => 
                           n12481, Q => n_2441, QN => n13895);
   REGISTERS_reg_63_11_inst : DFFR_X1 port map( D => n8352, CK => CLK, RN => 
                           n12572, Q => n_2442, QN => n13896);
   REGISTERS_reg_63_10_inst : DFFR_X1 port map( D => n8353, CK => CLK, RN => 
                           n12550, Q => n_2443, QN => n13897);
   REGISTERS_reg_63_9_inst : DFFR_X1 port map( D => n8354, CK => CLK, RN => 
                           n12557, Q => n_2444, QN => n13898);
   REGISTERS_reg_63_8_inst : DFFR_X1 port map( D => n8355, CK => CLK, RN => 
                           n12535, Q => n_2445, QN => n13899);
   REGISTERS_reg_63_7_inst : DFFR_X1 port map( D => n8356, CK => CLK, RN => 
                           n12645, Q => n_2446, QN => n13900);
   REGISTERS_reg_63_6_inst : DFFR_X1 port map( D => n8357, CK => CLK, RN => 
                           n12601, Q => n_2447, QN => n13901);
   REGISTERS_reg_63_5_inst : DFFR_X1 port map( D => n8358, CK => CLK, RN => 
                           n12488, Q => n_2448, QN => n13902);
   REGISTERS_reg_63_4_inst : DFFR_X1 port map( D => n8359, CK => CLK, RN => 
                           n12495, Q => n_2449, QN => n13903);
   REGISTERS_reg_63_3_inst : DFFR_X1 port map( D => n8360, CK => CLK, RN => 
                           n12579, Q => n_2450, QN => n13904);
   REGISTERS_reg_63_2_inst : DFFR_X1 port map( D => n8361, CK => CLK, RN => 
                           n12510, Q => n_2451, QN => n13905);
   REGISTERS_reg_63_1_inst : DFFR_X1 port map( D => n8362, CK => CLK, RN => 
                           n12438, Q => n_2452, QN => n13906);
   REGISTERS_reg_63_0_inst : DFFR_X1 port map( D => n8363, CK => CLK, RN => 
                           n12653, Q => n_2453, QN => n13907);
   REGISTERS_reg_64_31_inst : DFFR_X1 port map( D => n8364, CK => CLK, RN => 
                           n12660, Q => n_2454, QN => n5722);
   REGISTERS_reg_64_30_inst : DFFR_X1 port map( D => n8365, CK => CLK, RN => 
                           n12624, Q => n_2455, QN => n5754);
   REGISTERS_reg_64_29_inst : DFFR_X1 port map( D => n8366, CK => CLK, RN => 
                           n12609, Q => n_2456, QN => n5786);
   REGISTERS_reg_64_28_inst : DFFR_X1 port map( D => n8367, CK => CLK, RN => 
                           n12616, Q => n_2457, QN => n5818);
   REGISTERS_reg_64_27_inst : DFFR_X1 port map( D => n8368, CK => CLK, RN => 
                           n12587, Q => n_2458, QN => n5850);
   REGISTERS_reg_64_26_inst : DFFR_X1 port map( D => n8369, CK => CLK, RN => 
                           n12565, Q => n_2459, QN => n5882);
   REGISTERS_reg_64_25_inst : DFFR_X1 port map( D => n8370, CK => CLK, RN => 
                           n12543, Q => n_2460, QN => n5914);
   REGISTERS_reg_64_24_inst : DFFR_X1 port map( D => n8371, CK => CLK, RN => 
                           n12449, Q => n_2461, QN => n5946);
   REGISTERS_reg_64_23_inst : DFFR_X1 port map( D => n8372, CK => CLK, RN => 
                           n12631, Q => n_2462, QN => n6010);
   REGISTERS_reg_64_22_inst : DFFR_X1 port map( D => n8373, CK => CLK, RN => 
                           n12521, Q => n_2463, QN => n9145);
   REGISTERS_reg_64_21_inst : DFFR_X1 port map( D => n8374, CK => CLK, RN => 
                           n12528, Q => n_2464, QN => n9177);
   REGISTERS_reg_64_20_inst : DFFR_X1 port map( D => n8375, CK => CLK, RN => 
                           n12503, Q => n_2465, QN => n9209);
   REGISTERS_reg_64_19_inst : DFFR_X1 port map( D => n8376, CK => CLK, RN => 
                           n12594, Q => n_2466, QN => n9575);
   REGISTERS_reg_64_18_inst : DFFR_X1 port map( D => n8377, CK => CLK, RN => 
                           n12445, Q => n_2467, QN => n9607);
   REGISTERS_reg_64_17_inst : DFFR_X1 port map( D => n8378, CK => CLK, RN => 
                           n12453, Q => n_2468, QN => n9639);
   REGISTERS_reg_64_16_inst : DFFR_X1 port map( D => n8379, CK => CLK, RN => 
                           n12459, Q => n_2469, QN => n10001);
   REGISTERS_reg_64_15_inst : DFFR_X1 port map( D => n8380, CK => CLK, RN => 
                           n12638, Q => n_2470, QN => n10033);
   REGISTERS_reg_64_14_inst : DFFR_X1 port map( D => n8381, CK => CLK, RN => 
                           n12466, Q => n_2471, QN => n10065);
   REGISTERS_reg_64_13_inst : DFFR_X1 port map( D => n8382, CK => CLK, RN => 
                           n12474, Q => n_2472, QN => n10097);
   REGISTERS_reg_64_12_inst : DFFR_X1 port map( D => n8383, CK => CLK, RN => 
                           n12481, Q => n_2473, QN => n10129);
   REGISTERS_reg_64_11_inst : DFFR_X1 port map( D => n8384, CK => CLK, RN => 
                           n12572, Q => n_2474, QN => n10161);
   REGISTERS_reg_64_10_inst : DFFR_X1 port map( D => n8385, CK => CLK, RN => 
                           n12550, Q => n_2475, QN => n10193);
   REGISTERS_reg_64_9_inst : DFFR_X1 port map( D => n8386, CK => CLK, RN => 
                           n12558, Q => n_2476, QN => n10227);
   REGISTERS_reg_64_8_inst : DFFR_X1 port map( D => n8387, CK => CLK, RN => 
                           n12536, Q => n_2477, QN => n10259);
   REGISTERS_reg_64_7_inst : DFFR_X1 port map( D => n8388, CK => CLK, RN => 
                           n12646, Q => n_2478, QN => n10291);
   REGISTERS_reg_64_6_inst : DFFR_X1 port map( D => n8389, CK => CLK, RN => 
                           n12602, Q => n_2479, QN => n10326);
   REGISTERS_reg_64_5_inst : DFFR_X1 port map( D => n8390, CK => CLK, RN => 
                           n12488, Q => n_2480, QN => n10358);
   REGISTERS_reg_64_4_inst : DFFR_X1 port map( D => n8391, CK => CLK, RN => 
                           n12496, Q => n_2481, QN => n10390);
   REGISTERS_reg_64_3_inst : DFFR_X1 port map( D => n8392, CK => CLK, RN => 
                           n12580, Q => n_2482, QN => n10425);
   REGISTERS_reg_64_2_inst : DFFR_X1 port map( D => n8393, CK => CLK, RN => 
                           n12510, Q => n_2483, QN => n10457);
   REGISTERS_reg_64_1_inst : DFFR_X1 port map( D => n8394, CK => CLK, RN => 
                           n12438, Q => n_2484, QN => n10489);
   REGISTERS_reg_64_0_inst : DFFR_X1 port map( D => n8395, CK => CLK, RN => 
                           n12653, Q => n_2485, QN => n10521);
   REGISTERS_reg_65_31_inst : DFFR_X1 port map( D => n8396, CK => CLK, RN => 
                           n12660, Q => n_2486, QN => n13908);
   REGISTERS_reg_65_30_inst : DFFR_X1 port map( D => n8397, CK => CLK, RN => 
                           n12624, Q => n_2487, QN => n13909);
   REGISTERS_reg_65_29_inst : DFFR_X1 port map( D => n8398, CK => CLK, RN => 
                           n12609, Q => n_2488, QN => n13910);
   REGISTERS_reg_65_28_inst : DFFR_X1 port map( D => n8399, CK => CLK, RN => 
                           n12616, Q => n_2489, QN => n13911);
   REGISTERS_reg_65_27_inst : DFFR_X1 port map( D => n8400, CK => CLK, RN => 
                           n12587, Q => n_2490, QN => n13912);
   REGISTERS_reg_65_26_inst : DFFR_X1 port map( D => n8401, CK => CLK, RN => 
                           n12565, Q => n_2491, QN => n13913);
   REGISTERS_reg_65_25_inst : DFFR_X1 port map( D => n8402, CK => CLK, RN => 
                           n12543, Q => n_2492, QN => n13914);
   REGISTERS_reg_65_24_inst : DFFR_X1 port map( D => n8403, CK => CLK, RN => 
                           n12461, Q => n_2493, QN => n13915);
   REGISTERS_reg_65_23_inst : DFFR_X1 port map( D => n8404, CK => CLK, RN => 
                           n12631, Q => n_2494, QN => n13916);
   REGISTERS_reg_65_22_inst : DFFR_X1 port map( D => n8405, CK => CLK, RN => 
                           n12521, Q => n_2495, QN => n13917);
   REGISTERS_reg_65_21_inst : DFFR_X1 port map( D => n8406, CK => CLK, RN => 
                           n12528, Q => n_2496, QN => n13918);
   REGISTERS_reg_65_20_inst : DFFR_X1 port map( D => n8407, CK => CLK, RN => 
                           n12503, Q => n_2497, QN => n13919);
   REGISTERS_reg_65_19_inst : DFFR_X1 port map( D => n8408, CK => CLK, RN => 
                           n12594, Q => n_2498, QN => n13920);
   REGISTERS_reg_65_18_inst : DFFR_X1 port map( D => n8409, CK => CLK, RN => 
                           n12445, Q => n_2499, QN => n13921);
   REGISTERS_reg_65_17_inst : DFFR_X1 port map( D => n8410, CK => CLK, RN => 
                           n12453, Q => n_2500, QN => n13922);
   REGISTERS_reg_65_16_inst : DFFR_X1 port map( D => n8411, CK => CLK, RN => 
                           n12459, Q => n_2501, QN => n13923);
   REGISTERS_reg_65_15_inst : DFFR_X1 port map( D => n8412, CK => CLK, RN => 
                           n12638, Q => n_2502, QN => n13924);
   REGISTERS_reg_65_14_inst : DFFR_X1 port map( D => n8413, CK => CLK, RN => 
                           n12466, Q => n_2503, QN => n13925);
   REGISTERS_reg_65_13_inst : DFFR_X1 port map( D => n8414, CK => CLK, RN => 
                           n12474, Q => n_2504, QN => n13926);
   REGISTERS_reg_65_12_inst : DFFR_X1 port map( D => n8415, CK => CLK, RN => 
                           n12481, Q => n_2505, QN => n13927);
   REGISTERS_reg_65_11_inst : DFFR_X1 port map( D => n8416, CK => CLK, RN => 
                           n12572, Q => n_2506, QN => n13928);
   REGISTERS_reg_65_10_inst : DFFR_X1 port map( D => n8417, CK => CLK, RN => 
                           n12550, Q => n_2507, QN => n13929);
   REGISTERS_reg_65_9_inst : DFFR_X1 port map( D => n8418, CK => CLK, RN => 
                           n12558, Q => n_2508, QN => n13930);
   REGISTERS_reg_65_8_inst : DFFR_X1 port map( D => n8419, CK => CLK, RN => 
                           n12536, Q => n_2509, QN => n13931);
   REGISTERS_reg_65_7_inst : DFFR_X1 port map( D => n8420, CK => CLK, RN => 
                           n12646, Q => n_2510, QN => n13932);
   REGISTERS_reg_65_6_inst : DFFR_X1 port map( D => n8421, CK => CLK, RN => 
                           n12602, Q => n_2511, QN => n13933);
   REGISTERS_reg_65_5_inst : DFFR_X1 port map( D => n8422, CK => CLK, RN => 
                           n12488, Q => n_2512, QN => n13934);
   REGISTERS_reg_65_4_inst : DFFR_X1 port map( D => n8423, CK => CLK, RN => 
                           n12496, Q => n_2513, QN => n13935);
   REGISTERS_reg_65_3_inst : DFFR_X1 port map( D => n8424, CK => CLK, RN => 
                           n12580, Q => n_2514, QN => n13936);
   REGISTERS_reg_65_2_inst : DFFR_X1 port map( D => n8425, CK => CLK, RN => 
                           n12510, Q => n_2515, QN => n13937);
   REGISTERS_reg_65_1_inst : DFFR_X1 port map( D => n8426, CK => CLK, RN => 
                           n12438, Q => n_2516, QN => n13938);
   REGISTERS_reg_65_0_inst : DFFR_X1 port map( D => n8427, CK => CLK, RN => 
                           n12653, Q => n_2517, QN => n13939);
   REGISTERS_reg_66_31_inst : DFFR_X1 port map( D => n8428, CK => CLK, RN => 
                           n12660, Q => n_2518, QN => n13940);
   REGISTERS_reg_66_30_inst : DFFR_X1 port map( D => n8429, CK => CLK, RN => 
                           n12624, Q => n_2519, QN => n13941);
   REGISTERS_reg_66_29_inst : DFFR_X1 port map( D => n8430, CK => CLK, RN => 
                           n12609, Q => n_2520, QN => n13942);
   REGISTERS_reg_66_28_inst : DFFR_X1 port map( D => n8431, CK => CLK, RN => 
                           n12616, Q => n_2521, QN => n13943);
   REGISTERS_reg_66_27_inst : DFFR_X1 port map( D => n8432, CK => CLK, RN => 
                           n12587, Q => n_2522, QN => n13944);
   REGISTERS_reg_66_26_inst : DFFR_X1 port map( D => n8433, CK => CLK, RN => 
                           n12565, Q => n_2523, QN => n13945);
   REGISTERS_reg_66_25_inst : DFFR_X1 port map( D => n8434_port, CK => CLK, RN 
                           => n12543, Q => n_2524, QN => n13946);
   REGISTERS_reg_66_24_inst : DFFR_X1 port map( D => n8435_port, CK => CLK, RN 
                           => n12460, Q => n_2525, QN => n13947);
   REGISTERS_reg_66_23_inst : DFFR_X1 port map( D => n8436_port, CK => CLK, RN 
                           => n12631, Q => n_2526, QN => n13948);
   REGISTERS_reg_66_22_inst : DFFR_X1 port map( D => n8437_port, CK => CLK, RN 
                           => n12521, Q => n_2527, QN => n13949);
   REGISTERS_reg_66_21_inst : DFFR_X1 port map( D => n8438, CK => CLK, RN => 
                           n12528, Q => n_2528, QN => n13950);
   REGISTERS_reg_66_20_inst : DFFR_X1 port map( D => n8439, CK => CLK, RN => 
                           n12503, Q => n_2529, QN => n13951);
   REGISTERS_reg_66_19_inst : DFFR_X1 port map( D => n8440, CK => CLK, RN => 
                           n12594, Q => n_2530, QN => n13952);
   REGISTERS_reg_66_18_inst : DFFR_X1 port map( D => n8441, CK => CLK, RN => 
                           n12445, Q => n_2531, QN => n13953);
   REGISTERS_reg_66_17_inst : DFFR_X1 port map( D => n8442, CK => CLK, RN => 
                           n12453, Q => n_2532, QN => n13954);
   REGISTERS_reg_66_16_inst : DFFR_X1 port map( D => n8443, CK => CLK, RN => 
                           n12459, Q => n_2533, QN => n13955);
   REGISTERS_reg_66_15_inst : DFFR_X1 port map( D => n8444, CK => CLK, RN => 
                           n12638, Q => n_2534, QN => n13956);
   REGISTERS_reg_66_14_inst : DFFR_X1 port map( D => n8445, CK => CLK, RN => 
                           n12466, Q => n_2535, QN => n13957);
   REGISTERS_reg_66_13_inst : DFFR_X1 port map( D => n8446, CK => CLK, RN => 
                           n12474, Q => n_2536, QN => n13958);
   REGISTERS_reg_66_12_inst : DFFR_X1 port map( D => n8447, CK => CLK, RN => 
                           n12481, Q => n_2537, QN => n13959);
   REGISTERS_reg_66_11_inst : DFFR_X1 port map( D => n8448, CK => CLK, RN => 
                           n12572, Q => n_2538, QN => n13960);
   REGISTERS_reg_66_10_inst : DFFR_X1 port map( D => n8449, CK => CLK, RN => 
                           n12550, Q => n_2539, QN => n13961);
   REGISTERS_reg_66_9_inst : DFFR_X1 port map( D => n8450, CK => CLK, RN => 
                           n12558, Q => n_2540, QN => n13962);
   REGISTERS_reg_66_8_inst : DFFR_X1 port map( D => n8451, CK => CLK, RN => 
                           n12536, Q => n_2541, QN => n13963);
   REGISTERS_reg_66_7_inst : DFFR_X1 port map( D => n8452, CK => CLK, RN => 
                           n12646, Q => n_2542, QN => n13964);
   REGISTERS_reg_66_6_inst : DFFR_X1 port map( D => n8453, CK => CLK, RN => 
                           n12602, Q => n_2543, QN => n13965);
   REGISTERS_reg_66_5_inst : DFFR_X1 port map( D => n8454, CK => CLK, RN => 
                           n12488, Q => n_2544, QN => n13966);
   REGISTERS_reg_66_4_inst : DFFR_X1 port map( D => n8455, CK => CLK, RN => 
                           n12496, Q => n_2545, QN => n13967);
   REGISTERS_reg_66_3_inst : DFFR_X1 port map( D => n8456, CK => CLK, RN => 
                           n12580, Q => n_2546, QN => n13968);
   REGISTERS_reg_66_2_inst : DFFR_X1 port map( D => n8457, CK => CLK, RN => 
                           n12510, Q => n_2547, QN => n13969);
   REGISTERS_reg_66_1_inst : DFFR_X1 port map( D => n8458, CK => CLK, RN => 
                           n12438, Q => n_2548, QN => n13970);
   REGISTERS_reg_66_0_inst : DFFR_X1 port map( D => n8459, CK => CLK, RN => 
                           n12653, Q => n_2549, QN => n13971);
   REGISTERS_reg_67_31_inst : DFFR_X1 port map( D => n8460, CK => CLK, RN => 
                           n12660, Q => n_2550, QN => n13972);
   REGISTERS_reg_67_30_inst : DFFR_X1 port map( D => n8461, CK => CLK, RN => 
                           n12624, Q => n_2551, QN => n13973);
   REGISTERS_reg_67_29_inst : DFFR_X1 port map( D => n8462, CK => CLK, RN => 
                           n12609, Q => n_2552, QN => n13974);
   REGISTERS_reg_67_28_inst : DFFR_X1 port map( D => n8463, CK => CLK, RN => 
                           n12616, Q => n_2553, QN => n13975);
   REGISTERS_reg_67_27_inst : DFFR_X1 port map( D => n8464, CK => CLK, RN => 
                           n12587, Q => n_2554, QN => n13976);
   REGISTERS_reg_67_26_inst : DFFR_X1 port map( D => n8465, CK => CLK, RN => 
                           n12565, Q => n_2555, QN => n13977);
   REGISTERS_reg_67_25_inst : DFFR_X1 port map( D => n8466, CK => CLK, RN => 
                           n12543, Q => n_2556, QN => n13978);
   REGISTERS_reg_67_24_inst : DFFR_X1 port map( D => n8467, CK => CLK, RN => 
                           n12459, Q => n_2557, QN => n13979);
   REGISTERS_reg_67_23_inst : DFFR_X1 port map( D => n8468, CK => CLK, RN => 
                           n12631, Q => n_2558, QN => n13980);
   REGISTERS_reg_67_22_inst : DFFR_X1 port map( D => n8469, CK => CLK, RN => 
                           n12521, Q => n_2559, QN => n13981);
   REGISTERS_reg_67_21_inst : DFFR_X1 port map( D => n8470, CK => CLK, RN => 
                           n12528, Q => n_2560, QN => n13982);
   REGISTERS_reg_67_20_inst : DFFR_X1 port map( D => n8471, CK => CLK, RN => 
                           n12503, Q => n_2561, QN => n13983);
   REGISTERS_reg_67_19_inst : DFFR_X1 port map( D => n8472, CK => CLK, RN => 
                           n12594, Q => n_2562, QN => n13984);
   REGISTERS_reg_67_18_inst : DFFR_X1 port map( D => n8473, CK => CLK, RN => 
                           n12445, Q => n_2563, QN => n13985);
   REGISTERS_reg_67_17_inst : DFFR_X1 port map( D => n8474, CK => CLK, RN => 
                           n12453, Q => n_2564, QN => n13986);
   REGISTERS_reg_67_16_inst : DFFR_X1 port map( D => n8475, CK => CLK, RN => 
                           n12459, Q => n_2565, QN => n13987);
   REGISTERS_reg_67_15_inst : DFFR_X1 port map( D => n8476, CK => CLK, RN => 
                           n12638, Q => n_2566, QN => n13988);
   REGISTERS_reg_67_14_inst : DFFR_X1 port map( D => n8477, CK => CLK, RN => 
                           n12466, Q => n_2567, QN => n13989);
   REGISTERS_reg_67_13_inst : DFFR_X1 port map( D => n8478, CK => CLK, RN => 
                           n12474, Q => n_2568, QN => n13990);
   REGISTERS_reg_67_12_inst : DFFR_X1 port map( D => n8479, CK => CLK, RN => 
                           n12481, Q => n_2569, QN => n13991);
   REGISTERS_reg_67_11_inst : DFFR_X1 port map( D => n8480, CK => CLK, RN => 
                           n12572, Q => n_2570, QN => n13992);
   REGISTERS_reg_67_10_inst : DFFR_X1 port map( D => n8481, CK => CLK, RN => 
                           n12550, Q => n_2571, QN => n13993);
   REGISTERS_reg_67_9_inst : DFFR_X1 port map( D => n8482, CK => CLK, RN => 
                           n12558, Q => n_2572, QN => n13994);
   REGISTERS_reg_67_8_inst : DFFR_X1 port map( D => n8483, CK => CLK, RN => 
                           n12536, Q => n_2573, QN => n13995);
   REGISTERS_reg_67_7_inst : DFFR_X1 port map( D => n8484, CK => CLK, RN => 
                           n12646, Q => n_2574, QN => n13996);
   REGISTERS_reg_67_6_inst : DFFR_X1 port map( D => n8485, CK => CLK, RN => 
                           n12602, Q => n_2575, QN => n13997);
   REGISTERS_reg_67_5_inst : DFFR_X1 port map( D => n8486, CK => CLK, RN => 
                           n12488, Q => n_2576, QN => n13998);
   REGISTERS_reg_67_4_inst : DFFR_X1 port map( D => n8487, CK => CLK, RN => 
                           n12496, Q => n_2577, QN => n13999);
   REGISTERS_reg_67_3_inst : DFFR_X1 port map( D => n8488, CK => CLK, RN => 
                           n12580, Q => n_2578, QN => n14000);
   REGISTERS_reg_67_2_inst : DFFR_X1 port map( D => n8489, CK => CLK, RN => 
                           n12510, Q => n_2579, QN => n14001);
   REGISTERS_reg_67_1_inst : DFFR_X1 port map( D => n8490, CK => CLK, RN => 
                           n12438, Q => n_2580, QN => n14002);
   REGISTERS_reg_67_0_inst : DFFR_X1 port map( D => n8491, CK => CLK, RN => 
                           n12653, Q => n_2581, QN => n14003);
   REGISTERS_reg_68_31_inst : DFFR_X1 port map( D => n8492, CK => CLK, RN => 
                           n12661, Q => n_2582, QN => n998);
   REGISTERS_reg_68_30_inst : DFFR_X1 port map( D => n8493, CK => CLK, RN => 
                           n12624, Q => n_2583, QN => n14004);
   REGISTERS_reg_68_29_inst : DFFR_X1 port map( D => n8494, CK => CLK, RN => 
                           n12609, Q => n_2584, QN => n14005);
   REGISTERS_reg_68_28_inst : DFFR_X1 port map( D => n8495, CK => CLK, RN => 
                           n12617, Q => n_2585, QN => n14006);
   REGISTERS_reg_68_27_inst : DFFR_X1 port map( D => n8496, CK => CLK, RN => 
                           n12587, Q => n_2586, QN => n14007);
   REGISTERS_reg_68_26_inst : DFFR_X1 port map( D => n8497, CK => CLK, RN => 
                           n12565, Q => n_2587, QN => n14008);
   REGISTERS_reg_68_25_inst : DFFR_X1 port map( D => n8498, CK => CLK, RN => 
                           n12543, Q => n_2588, QN => n14009);
   REGISTERS_reg_68_24_inst : DFFR_X1 port map( D => n8499, CK => CLK, RN => 
                           n12458, Q => n_2589, QN => n14010);
   REGISTERS_reg_68_23_inst : DFFR_X1 port map( D => n8500, CK => CLK, RN => 
                           n12631, Q => n_2590, QN => n14011);
   REGISTERS_reg_68_22_inst : DFFR_X1 port map( D => n8501, CK => CLK, RN => 
                           n12521, Q => n_2591, QN => n14012);
   REGISTERS_reg_68_21_inst : DFFR_X1 port map( D => n8502, CK => CLK, RN => 
                           n12529, Q => n_2592, QN => n14013);
   REGISTERS_reg_68_20_inst : DFFR_X1 port map( D => n8503, CK => CLK, RN => 
                           n12503, Q => n_2593, QN => n14014);
   REGISTERS_reg_68_19_inst : DFFR_X1 port map( D => n8504, CK => CLK, RN => 
                           n12595, Q => n_2594, QN => n14015);
   REGISTERS_reg_68_18_inst : DFFR_X1 port map( D => n8505, CK => CLK, RN => 
                           n12446, Q => n_2595, QN => n14016);
   REGISTERS_reg_68_17_inst : DFFR_X1 port map( D => n8506, CK => CLK, RN => 
                           n12453, Q => n_2596, QN => n14017);
   REGISTERS_reg_68_16_inst : DFFR_X1 port map( D => n8507, CK => CLK, RN => 
                           n12459, Q => n_2597, QN => n14018);
   REGISTERS_reg_68_15_inst : DFFR_X1 port map( D => n8508, CK => CLK, RN => 
                           n12639, Q => n_2598, QN => n14019);
   REGISTERS_reg_68_14_inst : DFFR_X1 port map( D => n8509, CK => CLK, RN => 
                           n12467, Q => n_2599, QN => n14020);
   REGISTERS_reg_68_13_inst : DFFR_X1 port map( D => n8510, CK => CLK, RN => 
                           n12474, Q => n_2600, QN => n14021);
   REGISTERS_reg_68_12_inst : DFFR_X1 port map( D => n8511, CK => CLK, RN => 
                           n12481, Q => n_2601, QN => n14022);
   REGISTERS_reg_68_11_inst : DFFR_X1 port map( D => n8512, CK => CLK, RN => 
                           n12573, Q => n_2602, QN => n14023);
   REGISTERS_reg_68_10_inst : DFFR_X1 port map( D => n8513, CK => CLK, RN => 
                           n12551, Q => n_2603, QN => n14024);
   REGISTERS_reg_68_9_inst : DFFR_X1 port map( D => n8514, CK => CLK, RN => 
                           n12558, Q => n_2604, QN => n14025);
   REGISTERS_reg_68_8_inst : DFFR_X1 port map( D => n8515, CK => CLK, RN => 
                           n12536, Q => n_2605, QN => n14026);
   REGISTERS_reg_68_7_inst : DFFR_X1 port map( D => n8516, CK => CLK, RN => 
                           n12646, Q => n_2606, QN => n14027);
   REGISTERS_reg_68_6_inst : DFFR_X1 port map( D => n8517, CK => CLK, RN => 
                           n12602, Q => n_2607, QN => n14028);
   REGISTERS_reg_68_5_inst : DFFR_X1 port map( D => n8518, CK => CLK, RN => 
                           n12489, Q => n_2608, QN => n14029);
   REGISTERS_reg_68_4_inst : DFFR_X1 port map( D => n8519, CK => CLK, RN => 
                           n12496, Q => n_2609, QN => n14030);
   REGISTERS_reg_68_3_inst : DFFR_X1 port map( D => n8520, CK => CLK, RN => 
                           n12580, Q => n_2610, QN => n14031);
   REGISTERS_reg_68_2_inst : DFFR_X1 port map( D => n8521, CK => CLK, RN => 
                           n12511, Q => n_2611, QN => n14032);
   REGISTERS_reg_68_1_inst : DFFR_X1 port map( D => n8522, CK => CLK, RN => 
                           n12438, Q => n_2612, QN => n14033);
   REGISTERS_reg_68_0_inst : DFFR_X1 port map( D => n8523, CK => CLK, RN => 
                           n12653, Q => n_2613, QN => n14034);
   REGISTERS_reg_69_31_inst : DFFR_X1 port map( D => n8524, CK => CLK, RN => 
                           n12661, Q => n_2614, QN => n14035);
   REGISTERS_reg_69_30_inst : DFFR_X1 port map( D => n8525, CK => CLK, RN => 
                           n12624, Q => n_2615, QN => n14036);
   REGISTERS_reg_69_29_inst : DFFR_X1 port map( D => n8526, CK => CLK, RN => 
                           n12609, Q => n_2616, QN => n14037);
   REGISTERS_reg_69_28_inst : DFFR_X1 port map( D => n8527, CK => CLK, RN => 
                           n12617, Q => n_2617, QN => n14038);
   REGISTERS_reg_69_27_inst : DFFR_X1 port map( D => n8528, CK => CLK, RN => 
                           n12587, Q => n_2618, QN => n14039);
   REGISTERS_reg_69_26_inst : DFFR_X1 port map( D => n8529, CK => CLK, RN => 
                           n12565, Q => n_2619, QN => n14040);
   REGISTERS_reg_69_25_inst : DFFR_X1 port map( D => n8530, CK => CLK, RN => 
                           n12543, Q => n_2620, QN => n14041);
   REGISTERS_reg_69_24_inst : DFFR_X1 port map( D => n8531, CK => CLK, RN => 
                           n12467, Q => n_2621, QN => n14042);
   REGISTERS_reg_69_23_inst : DFFR_X1 port map( D => n8532, CK => CLK, RN => 
                           n12631, Q => n_2622, QN => n14043);
   REGISTERS_reg_69_22_inst : DFFR_X1 port map( D => n8533, CK => CLK, RN => 
                           n12521, Q => n_2623, QN => n14044);
   REGISTERS_reg_69_21_inst : DFFR_X1 port map( D => n8534, CK => CLK, RN => 
                           n12529, Q => n_2624, QN => n14045);
   REGISTERS_reg_69_20_inst : DFFR_X1 port map( D => n8535, CK => CLK, RN => 
                           n12503, Q => n_2625, QN => n14046);
   REGISTERS_reg_69_19_inst : DFFR_X1 port map( D => n8536, CK => CLK, RN => 
                           n12595, Q => n_2626, QN => n14047);
   REGISTERS_reg_69_18_inst : DFFR_X1 port map( D => n8537, CK => CLK, RN => 
                           n12446, Q => n_2627, QN => n14048);
   REGISTERS_reg_69_17_inst : DFFR_X1 port map( D => n8538, CK => CLK, RN => 
                           n12453, Q => n_2628, QN => n14049);
   REGISTERS_reg_69_16_inst : DFFR_X1 port map( D => n8539, CK => CLK, RN => 
                           n12459, Q => n_2629, QN => n14050);
   REGISTERS_reg_69_15_inst : DFFR_X1 port map( D => n8540, CK => CLK, RN => 
                           n12639, Q => n_2630, QN => n14051);
   REGISTERS_reg_69_14_inst : DFFR_X1 port map( D => n8541, CK => CLK, RN => 
                           n12467, Q => n_2631, QN => n14052);
   REGISTERS_reg_69_13_inst : DFFR_X1 port map( D => n8542, CK => CLK, RN => 
                           n12474, Q => n_2632, QN => n14053);
   REGISTERS_reg_69_12_inst : DFFR_X1 port map( D => n8543, CK => CLK, RN => 
                           n12481, Q => n_2633, QN => n14054);
   REGISTERS_reg_69_11_inst : DFFR_X1 port map( D => n8544, CK => CLK, RN => 
                           n12573, Q => n_2634, QN => n14055);
   REGISTERS_reg_69_10_inst : DFFR_X1 port map( D => n8545, CK => CLK, RN => 
                           n12551, Q => n_2635, QN => n14056);
   REGISTERS_reg_69_9_inst : DFFR_X1 port map( D => n8546, CK => CLK, RN => 
                           n12558, Q => n_2636, QN => n14057);
   REGISTERS_reg_69_8_inst : DFFR_X1 port map( D => n8547, CK => CLK, RN => 
                           n12536, Q => n_2637, QN => n14058);
   REGISTERS_reg_69_7_inst : DFFR_X1 port map( D => n8548, CK => CLK, RN => 
                           n12646, Q => n_2638, QN => n14059);
   REGISTERS_reg_69_6_inst : DFFR_X1 port map( D => n8549, CK => CLK, RN => 
                           n12602, Q => n_2639, QN => n14060);
   REGISTERS_reg_69_5_inst : DFFR_X1 port map( D => n8550, CK => CLK, RN => 
                           n12489, Q => n_2640, QN => n14061);
   REGISTERS_reg_69_4_inst : DFFR_X1 port map( D => n8551, CK => CLK, RN => 
                           n12496, Q => n_2641, QN => n14062);
   REGISTERS_reg_69_3_inst : DFFR_X1 port map( D => n8552, CK => CLK, RN => 
                           n12580, Q => n_2642, QN => n14063);
   REGISTERS_reg_69_2_inst : DFFR_X1 port map( D => n8553, CK => CLK, RN => 
                           n12511, Q => n_2643, QN => n14064);
   REGISTERS_reg_69_1_inst : DFFR_X1 port map( D => n8554, CK => CLK, RN => 
                           n12438, Q => n_2644, QN => n14065);
   REGISTERS_reg_69_0_inst : DFFR_X1 port map( D => n8555, CK => CLK, RN => 
                           n12653, Q => n_2645, QN => n14066);
   REGISTERS_reg_70_31_inst : DFFR_X1 port map( D => n8556, CK => CLK, RN => 
                           n12661, Q => n_2646, QN => n14067);
   REGISTERS_reg_70_30_inst : DFFR_X1 port map( D => n8557, CK => CLK, RN => 
                           n12624, Q => n_2647, QN => n14068);
   REGISTERS_reg_70_29_inst : DFFR_X1 port map( D => n8558, CK => CLK, RN => 
                           n12609, Q => n_2648, QN => n14069);
   REGISTERS_reg_70_28_inst : DFFR_X1 port map( D => n8559, CK => CLK, RN => 
                           n12617, Q => n_2649, QN => n14070);
   REGISTERS_reg_70_27_inst : DFFR_X1 port map( D => n8560, CK => CLK, RN => 
                           n12587, Q => n_2650, QN => n14071);
   REGISTERS_reg_70_26_inst : DFFR_X1 port map( D => n8561, CK => CLK, RN => 
                           n12565, Q => n_2651, QN => n14072);
   REGISTERS_reg_70_25_inst : DFFR_X1 port map( D => n8562, CK => CLK, RN => 
                           n12543, Q => n_2652, QN => n14073);
   REGISTERS_reg_70_24_inst : DFFR_X1 port map( D => n8563, CK => CLK, RN => 
                           n12457, Q => n_2653, QN => n14074);
   REGISTERS_reg_70_23_inst : DFFR_X1 port map( D => n8564, CK => CLK, RN => 
                           n12631, Q => n_2654, QN => n14075);
   REGISTERS_reg_70_22_inst : DFFR_X1 port map( D => n8565, CK => CLK, RN => 
                           n12521, Q => n_2655, QN => n14076);
   REGISTERS_reg_70_21_inst : DFFR_X1 port map( D => n8566, CK => CLK, RN => 
                           n12529, Q => n_2656, QN => n14077);
   REGISTERS_reg_70_20_inst : DFFR_X1 port map( D => n8567, CK => CLK, RN => 
                           n12503, Q => n_2657, QN => n14078);
   REGISTERS_reg_70_19_inst : DFFR_X1 port map( D => n8568, CK => CLK, RN => 
                           n12595, Q => n_2658, QN => n14079);
   REGISTERS_reg_70_18_inst : DFFR_X1 port map( D => n8569, CK => CLK, RN => 
                           n12446, Q => n_2659, QN => n14080);
   REGISTERS_reg_70_17_inst : DFFR_X1 port map( D => n8570, CK => CLK, RN => 
                           n12453, Q => n_2660, QN => n14081);
   REGISTERS_reg_70_16_inst : DFFR_X1 port map( D => n8571, CK => CLK, RN => 
                           n12459, Q => n_2661, QN => n14082);
   REGISTERS_reg_70_15_inst : DFFR_X1 port map( D => n8572, CK => CLK, RN => 
                           n12639, Q => n_2662, QN => n14083);
   REGISTERS_reg_70_14_inst : DFFR_X1 port map( D => n8573, CK => CLK, RN => 
                           n12467, Q => n_2663, QN => n14084);
   REGISTERS_reg_70_13_inst : DFFR_X1 port map( D => n8574, CK => CLK, RN => 
                           n12474, Q => n_2664, QN => n14085);
   REGISTERS_reg_70_12_inst : DFFR_X1 port map( D => n8575, CK => CLK, RN => 
                           n12481, Q => n_2665, QN => n14086);
   REGISTERS_reg_70_11_inst : DFFR_X1 port map( D => n8576, CK => CLK, RN => 
                           n12573, Q => n_2666, QN => n14087);
   REGISTERS_reg_70_10_inst : DFFR_X1 port map( D => n8577, CK => CLK, RN => 
                           n12551, Q => n_2667, QN => n14088);
   REGISTERS_reg_70_9_inst : DFFR_X1 port map( D => n8578_port, CK => CLK, RN 
                           => n12558, Q => n_2668, QN => n14089);
   REGISTERS_reg_70_8_inst : DFFR_X1 port map( D => n8579_port, CK => CLK, RN 
                           => n12536, Q => n_2669, QN => n14090);
   REGISTERS_reg_70_7_inst : DFFR_X1 port map( D => n8580_port, CK => CLK, RN 
                           => n12646, Q => n_2670, QN => n14091);
   REGISTERS_reg_70_6_inst : DFFR_X1 port map( D => n8581_port, CK => CLK, RN 
                           => n12602, Q => n_2671, QN => n14092);
   REGISTERS_reg_70_5_inst : DFFR_X1 port map( D => n8582, CK => CLK, RN => 
                           n12489, Q => n_2672, QN => n14093);
   REGISTERS_reg_70_4_inst : DFFR_X1 port map( D => n8583, CK => CLK, RN => 
                           n12496, Q => n_2673, QN => n14094);
   REGISTERS_reg_70_3_inst : DFFR_X1 port map( D => n8584, CK => CLK, RN => 
                           n12580, Q => n_2674, QN => n14095);
   REGISTERS_reg_70_2_inst : DFFR_X1 port map( D => n8585, CK => CLK, RN => 
                           n12511, Q => n_2675, QN => n14096);
   REGISTERS_reg_70_1_inst : DFFR_X1 port map( D => n8586, CK => CLK, RN => 
                           n12438, Q => n_2676, QN => n14097);
   REGISTERS_reg_70_0_inst : DFFR_X1 port map( D => n8587, CK => CLK, RN => 
                           n12653, Q => n_2677, QN => n14098);
   REGISTERS_reg_71_31_inst : DFFR_X1 port map( D => n8588, CK => CLK, RN => 
                           n12661, Q => n_2678, QN => n997);
   REGISTERS_reg_71_30_inst : DFFR_X1 port map( D => n8589, CK => CLK, RN => 
                           n12624, Q => n_2679, QN => n14099);
   REGISTERS_reg_71_29_inst : DFFR_X1 port map( D => n8590, CK => CLK, RN => 
                           n12609, Q => n_2680, QN => n14100);
   REGISTERS_reg_71_28_inst : DFFR_X1 port map( D => n8591, CK => CLK, RN => 
                           n12617, Q => n_2681, QN => n14101);
   REGISTERS_reg_71_27_inst : DFFR_X1 port map( D => n8592, CK => CLK, RN => 
                           n12587, Q => n_2682, QN => n14102);
   REGISTERS_reg_71_26_inst : DFFR_X1 port map( D => n8593, CK => CLK, RN => 
                           n12565, Q => n_2683, QN => n14103);
   REGISTERS_reg_71_25_inst : DFFR_X1 port map( D => n8594, CK => CLK, RN => 
                           n12543, Q => n_2684, QN => n14104);
   REGISTERS_reg_71_24_inst : DFFR_X1 port map( D => n8595, CK => CLK, RN => 
                           n12456, Q => n_2685, QN => n14105);
   REGISTERS_reg_71_23_inst : DFFR_X1 port map( D => n8596, CK => CLK, RN => 
                           n12631, Q => n_2686, QN => n14106);
   REGISTERS_reg_71_22_inst : DFFR_X1 port map( D => n8597, CK => CLK, RN => 
                           n12521, Q => n_2687, QN => n14107);
   REGISTERS_reg_71_21_inst : DFFR_X1 port map( D => n8598, CK => CLK, RN => 
                           n12529, Q => n_2688, QN => n14108);
   REGISTERS_reg_71_20_inst : DFFR_X1 port map( D => n8599, CK => CLK, RN => 
                           n12503, Q => n_2689, QN => n14109);
   REGISTERS_reg_71_19_inst : DFFR_X1 port map( D => n8600, CK => CLK, RN => 
                           n12595, Q => n_2690, QN => n14110);
   REGISTERS_reg_71_18_inst : DFFR_X1 port map( D => n8601, CK => CLK, RN => 
                           n12446, Q => n_2691, QN => n14111);
   REGISTERS_reg_71_17_inst : DFFR_X1 port map( D => n8602, CK => CLK, RN => 
                           n12453, Q => n_2692, QN => n14112);
   REGISTERS_reg_71_16_inst : DFFR_X1 port map( D => n8603, CK => CLK, RN => 
                           n12459, Q => n_2693, QN => n14113);
   REGISTERS_reg_71_15_inst : DFFR_X1 port map( D => n8604, CK => CLK, RN => 
                           n12639, Q => n_2694, QN => n14114);
   REGISTERS_reg_71_14_inst : DFFR_X1 port map( D => n8605, CK => CLK, RN => 
                           n12467, Q => n_2695, QN => n14115);
   REGISTERS_reg_71_13_inst : DFFR_X1 port map( D => n8606, CK => CLK, RN => 
                           n12474, Q => n_2696, QN => n14116);
   REGISTERS_reg_71_12_inst : DFFR_X1 port map( D => n8607, CK => CLK, RN => 
                           n12481, Q => n_2697, QN => n14117);
   REGISTERS_reg_71_11_inst : DFFR_X1 port map( D => n8608, CK => CLK, RN => 
                           n12573, Q => n_2698, QN => n14118);
   REGISTERS_reg_71_10_inst : DFFR_X1 port map( D => n8609, CK => CLK, RN => 
                           n12551, Q => n_2699, QN => n14119);
   REGISTERS_reg_71_9_inst : DFFR_X1 port map( D => n8610, CK => CLK, RN => 
                           n12558, Q => n_2700, QN => n14120);
   REGISTERS_reg_71_8_inst : DFFR_X1 port map( D => n8611, CK => CLK, RN => 
                           n12536, Q => n_2701, QN => n14121);
   REGISTERS_reg_71_7_inst : DFFR_X1 port map( D => n8612, CK => CLK, RN => 
                           n12646, Q => n_2702, QN => n14122);
   REGISTERS_reg_71_6_inst : DFFR_X1 port map( D => n8613, CK => CLK, RN => 
                           n12602, Q => n_2703, QN => n14123);
   REGISTERS_reg_71_5_inst : DFFR_X1 port map( D => n8614, CK => CLK, RN => 
                           n12489, Q => n_2704, QN => n14124);
   REGISTERS_reg_71_4_inst : DFFR_X1 port map( D => n8615, CK => CLK, RN => 
                           n12496, Q => n_2705, QN => n14125);
   REGISTERS_reg_71_3_inst : DFFR_X1 port map( D => n8616, CK => CLK, RN => 
                           n12580, Q => n_2706, QN => n14126);
   REGISTERS_reg_71_2_inst : DFFR_X1 port map( D => n8617, CK => CLK, RN => 
                           n12511, Q => n_2707, QN => n14127);
   REGISTERS_reg_71_1_inst : DFFR_X1 port map( D => n8618, CK => CLK, RN => 
                           n12438, Q => n_2708, QN => n14128);
   REGISTERS_reg_71_0_inst : DFFR_X1 port map( D => n8619, CK => CLK, RN => 
                           n12653, Q => n_2709, QN => n14129);
   REGISTERS_reg_72_31_inst : DFFR_X1 port map( D => n8620, CK => CLK, RN => 
                           n12661, Q => n_2710, QN => n14130);
   REGISTERS_reg_72_30_inst : DFFR_X1 port map( D => n8621, CK => CLK, RN => 
                           n12624, Q => n_2711, QN => n14131);
   REGISTERS_reg_72_29_inst : DFFR_X1 port map( D => n8622, CK => CLK, RN => 
                           n12610, Q => n_2712, QN => n14132);
   REGISTERS_reg_72_28_inst : DFFR_X1 port map( D => n8623, CK => CLK, RN => 
                           n12617, Q => n_2713, QN => n14133);
   REGISTERS_reg_72_27_inst : DFFR_X1 port map( D => n8624, CK => CLK, RN => 
                           n12588, Q => n_2714, QN => n14134);
   REGISTERS_reg_72_26_inst : DFFR_X1 port map( D => n8625, CK => CLK, RN => 
                           n12566, Q => n_2715, QN => n14135);
   REGISTERS_reg_72_25_inst : DFFR_X1 port map( D => n8626, CK => CLK, RN => 
                           n12544, Q => n_2716, QN => n14136);
   REGISTERS_reg_72_24_inst : DFFR_X1 port map( D => n8627, CK => CLK, RN => 
                           n12466, Q => n_2717, QN => n14137);
   REGISTERS_reg_72_23_inst : DFFR_X1 port map( D => n8628, CK => CLK, RN => 
                           n12632, Q => n_2718, QN => n14138);
   REGISTERS_reg_72_22_inst : DFFR_X1 port map( D => n8629, CK => CLK, RN => 
                           n12522, Q => n_2719, QN => n14139);
   REGISTERS_reg_72_21_inst : DFFR_X1 port map( D => n8630, CK => CLK, RN => 
                           n12529, Q => n_2720, QN => n14140);
   REGISTERS_reg_72_20_inst : DFFR_X1 port map( D => n8631, CK => CLK, RN => 
                           n12504, Q => n_2721, QN => n14141);
   REGISTERS_reg_72_19_inst : DFFR_X1 port map( D => n8632, CK => CLK, RN => 
                           n12595, Q => n_2722, QN => n14142);
   REGISTERS_reg_72_18_inst : DFFR_X1 port map( D => n8633, CK => CLK, RN => 
                           n12446, Q => n_2723, QN => n14143);
   REGISTERS_reg_72_17_inst : DFFR_X1 port map( D => n8634, CK => CLK, RN => 
                           n12453, Q => n_2724, QN => n14144);
   REGISTERS_reg_72_16_inst : DFFR_X1 port map( D => n8635, CK => CLK, RN => 
                           n12460, Q => n_2725, QN => n14145);
   REGISTERS_reg_72_15_inst : DFFR_X1 port map( D => n8636, CK => CLK, RN => 
                           n12639, Q => n_2726, QN => n14146);
   REGISTERS_reg_72_14_inst : DFFR_X1 port map( D => n8637, CK => CLK, RN => 
                           n12467, Q => n_2727, QN => n14147);
   REGISTERS_reg_72_13_inst : DFFR_X1 port map( D => n8638, CK => CLK, RN => 
                           n12474, Q => n_2728, QN => n14148);
   REGISTERS_reg_72_12_inst : DFFR_X1 port map( D => n8639, CK => CLK, RN => 
                           n12482, Q => n_2729, QN => n14149);
   REGISTERS_reg_72_11_inst : DFFR_X1 port map( D => n8640, CK => CLK, RN => 
                           n12573, Q => n_2730, QN => n14150);
   REGISTERS_reg_72_10_inst : DFFR_X1 port map( D => n8641, CK => CLK, RN => 
                           n12551, Q => n_2731, QN => n14151);
   REGISTERS_reg_72_9_inst : DFFR_X1 port map( D => n8642, CK => CLK, RN => 
                           n12558, Q => n_2732, QN => n14152);
   REGISTERS_reg_72_8_inst : DFFR_X1 port map( D => n8643, CK => CLK, RN => 
                           n12536, Q => n_2733, QN => n14153);
   REGISTERS_reg_72_7_inst : DFFR_X1 port map( D => n8644, CK => CLK, RN => 
                           n12646, Q => n_2734, QN => n14154);
   REGISTERS_reg_72_6_inst : DFFR_X1 port map( D => n8645, CK => CLK, RN => 
                           n12602, Q => n_2735, QN => n14155);
   REGISTERS_reg_72_5_inst : DFFR_X1 port map( D => n8646, CK => CLK, RN => 
                           n12489, Q => n_2736, QN => n14156);
   REGISTERS_reg_72_4_inst : DFFR_X1 port map( D => n8647, CK => CLK, RN => 
                           n12496, Q => n_2737, QN => n14157);
   REGISTERS_reg_72_3_inst : DFFR_X1 port map( D => n8648, CK => CLK, RN => 
                           n12580, Q => n_2738, QN => n14158);
   REGISTERS_reg_72_2_inst : DFFR_X1 port map( D => n8649, CK => CLK, RN => 
                           n12511, Q => n_2739, QN => n14159);
   REGISTERS_reg_72_1_inst : DFFR_X1 port map( D => n8650, CK => CLK, RN => 
                           n12439, Q => n_2740, QN => n14160);
   REGISTERS_reg_72_0_inst : DFFR_X1 port map( D => n8651, CK => CLK, RN => 
                           n12654, Q => n_2741, QN => n14161);
   REGISTERS_reg_73_31_inst : DFFR_X1 port map( D => n8652, CK => CLK, RN => 
                           n12661, Q => n_2742, QN => n14162);
   REGISTERS_reg_73_30_inst : DFFR_X1 port map( D => n8653, CK => CLK, RN => 
                           n12624, Q => n_2743, QN => n14163);
   REGISTERS_reg_73_29_inst : DFFR_X1 port map( D => n8654, CK => CLK, RN => 
                           n12610, Q => n_2744, QN => n14164);
   REGISTERS_reg_73_28_inst : DFFR_X1 port map( D => n8655, CK => CLK, RN => 
                           n12617, Q => n_2745, QN => n14165);
   REGISTERS_reg_73_27_inst : DFFR_X1 port map( D => n8656, CK => CLK, RN => 
                           n12588, Q => n_2746, QN => n14166);
   REGISTERS_reg_73_26_inst : DFFR_X1 port map( D => n8657, CK => CLK, RN => 
                           n12566, Q => n_2747, QN => n14167);
   REGISTERS_reg_73_25_inst : DFFR_X1 port map( D => n8658, CK => CLK, RN => 
                           n12544, Q => n_2748, QN => n14168);
   REGISTERS_reg_73_24_inst : DFFR_X1 port map( D => n8659, CK => CLK, RN => 
                           n12455, Q => n_2749, QN => n14169);
   REGISTERS_reg_73_23_inst : DFFR_X1 port map( D => n8660, CK => CLK, RN => 
                           n12632, Q => n_2750, QN => n14170);
   REGISTERS_reg_73_22_inst : DFFR_X1 port map( D => n8661, CK => CLK, RN => 
                           n12522, Q => n_2751, QN => n14171);
   REGISTERS_reg_73_21_inst : DFFR_X1 port map( D => n8662, CK => CLK, RN => 
                           n12529, Q => n_2752, QN => n14172);
   REGISTERS_reg_73_20_inst : DFFR_X1 port map( D => n8663, CK => CLK, RN => 
                           n12504, Q => n_2753, QN => n14173);
   REGISTERS_reg_73_19_inst : DFFR_X1 port map( D => n8664, CK => CLK, RN => 
                           n12595, Q => n_2754, QN => n14174);
   REGISTERS_reg_73_18_inst : DFFR_X1 port map( D => n8665, CK => CLK, RN => 
                           n12446, Q => n_2755, QN => n14175);
   REGISTERS_reg_73_17_inst : DFFR_X1 port map( D => n8666, CK => CLK, RN => 
                           n12453, Q => n_2756, QN => n14176);
   REGISTERS_reg_73_16_inst : DFFR_X1 port map( D => n8667, CK => CLK, RN => 
                           n12460, Q => n_2757, QN => n14177);
   REGISTERS_reg_73_15_inst : DFFR_X1 port map( D => n8668, CK => CLK, RN => 
                           n12639, Q => n_2758, QN => n14178);
   REGISTERS_reg_73_14_inst : DFFR_X1 port map( D => n8669, CK => CLK, RN => 
                           n12467, Q => n_2759, QN => n14179);
   REGISTERS_reg_73_13_inst : DFFR_X1 port map( D => n8670, CK => CLK, RN => 
                           n12474, Q => n_2760, QN => n14180);
   REGISTERS_reg_73_12_inst : DFFR_X1 port map( D => n8671, CK => CLK, RN => 
                           n12482, Q => n_2761, QN => n14181);
   REGISTERS_reg_73_11_inst : DFFR_X1 port map( D => n8672, CK => CLK, RN => 
                           n12573, Q => n_2762, QN => n14182);
   REGISTERS_reg_73_10_inst : DFFR_X1 port map( D => n8673, CK => CLK, RN => 
                           n12551, Q => n_2763, QN => n14183);
   REGISTERS_reg_73_9_inst : DFFR_X1 port map( D => n8674, CK => CLK, RN => 
                           n12558, Q => n_2764, QN => n14184);
   REGISTERS_reg_73_8_inst : DFFR_X1 port map( D => n8675, CK => CLK, RN => 
                           n12536, Q => n_2765, QN => n14185);
   REGISTERS_reg_73_7_inst : DFFR_X1 port map( D => n8676, CK => CLK, RN => 
                           n12646, Q => n_2766, QN => n14186);
   REGISTERS_reg_73_6_inst : DFFR_X1 port map( D => n8677, CK => CLK, RN => 
                           n12602, Q => n_2767, QN => n14187);
   REGISTERS_reg_73_5_inst : DFFR_X1 port map( D => n8678, CK => CLK, RN => 
                           n12489, Q => n_2768, QN => n14188);
   REGISTERS_reg_73_4_inst : DFFR_X1 port map( D => n8679, CK => CLK, RN => 
                           n12496, Q => n_2769, QN => n14189);
   REGISTERS_reg_73_3_inst : DFFR_X1 port map( D => n8680, CK => CLK, RN => 
                           n12580, Q => n_2770, QN => n14190);
   REGISTERS_reg_73_2_inst : DFFR_X1 port map( D => n8681, CK => CLK, RN => 
                           n12511, Q => n_2771, QN => n14191);
   REGISTERS_reg_73_1_inst : DFFR_X1 port map( D => n8682, CK => CLK, RN => 
                           n12439, Q => n_2772, QN => n14192);
   REGISTERS_reg_73_0_inst : DFFR_X1 port map( D => n8683, CK => CLK, RN => 
                           n12654, Q => n_2773, QN => n14193);
   REGISTERS_reg_74_31_inst : DFFR_X1 port map( D => n8684, CK => CLK, RN => 
                           n12661, Q => n_2774, QN => n996);
   REGISTERS_reg_74_30_inst : DFFR_X1 port map( D => n8685, CK => CLK, RN => 
                           n12624, Q => n_2775, QN => n14194);
   REGISTERS_reg_74_29_inst : DFFR_X1 port map( D => n8686, CK => CLK, RN => 
                           n12610, Q => n_2776, QN => n14195);
   REGISTERS_reg_74_28_inst : DFFR_X1 port map( D => n8687, CK => CLK, RN => 
                           n12617, Q => n_2777, QN => n14196);
   REGISTERS_reg_74_27_inst : DFFR_X1 port map( D => n8688, CK => CLK, RN => 
                           n12588, Q => n_2778, QN => n14197);
   REGISTERS_reg_74_26_inst : DFFR_X1 port map( D => n8689, CK => CLK, RN => 
                           n12566, Q => n_2779, QN => n14198);
   REGISTERS_reg_74_25_inst : DFFR_X1 port map( D => n8690, CK => CLK, RN => 
                           n12544, Q => n_2780, QN => n14199);
   REGISTERS_reg_74_24_inst : DFFR_X1 port map( D => n8691, CK => CLK, RN => 
                           n12468, Q => n_2781, QN => n14200);
   REGISTERS_reg_74_23_inst : DFFR_X1 port map( D => n8692, CK => CLK, RN => 
                           n12632, Q => n_2782, QN => n14201);
   REGISTERS_reg_74_22_inst : DFFR_X1 port map( D => n8693, CK => CLK, RN => 
                           n12522, Q => n_2783, QN => n14202);
   REGISTERS_reg_74_21_inst : DFFR_X1 port map( D => n8694, CK => CLK, RN => 
                           n12529, Q => n_2784, QN => n14203);
   REGISTERS_reg_74_20_inst : DFFR_X1 port map( D => n8695, CK => CLK, RN => 
                           n12504, Q => n_2785, QN => n14204);
   REGISTERS_reg_74_19_inst : DFFR_X1 port map( D => n8696, CK => CLK, RN => 
                           n12595, Q => n_2786, QN => n14205);
   REGISTERS_reg_74_18_inst : DFFR_X1 port map( D => n8697, CK => CLK, RN => 
                           n12446, Q => n_2787, QN => n14206);
   REGISTERS_reg_74_17_inst : DFFR_X1 port map( D => n8698, CK => CLK, RN => 
                           n12453, Q => n_2788, QN => n14207);
   REGISTERS_reg_74_16_inst : DFFR_X1 port map( D => n8699, CK => CLK, RN => 
                           n12460, Q => n_2789, QN => n14208);
   REGISTERS_reg_74_15_inst : DFFR_X1 port map( D => n8700, CK => CLK, RN => 
                           n12639, Q => n_2790, QN => n14209);
   REGISTERS_reg_74_14_inst : DFFR_X1 port map( D => n8701, CK => CLK, RN => 
                           n12467, Q => n_2791, QN => n14210);
   REGISTERS_reg_74_13_inst : DFFR_X1 port map( D => n8702_port, CK => CLK, RN 
                           => n12474, Q => n_2792, QN => n14211);
   REGISTERS_reg_74_12_inst : DFFR_X1 port map( D => n8703_port, CK => CLK, RN 
                           => n12482, Q => n_2793, QN => n14212);
   REGISTERS_reg_74_11_inst : DFFR_X1 port map( D => n8704_port, CK => CLK, RN 
                           => n12573, Q => n_2794, QN => n14213);
   REGISTERS_reg_74_10_inst : DFFR_X1 port map( D => n8705_port, CK => CLK, RN 
                           => n12551, Q => n_2795, QN => n14214);
   REGISTERS_reg_74_9_inst : DFFR_X1 port map( D => n8706_port, CK => CLK, RN 
                           => n12558, Q => n_2796, QN => n14215);
   REGISTERS_reg_74_8_inst : DFFR_X1 port map( D => n8707_port, CK => CLK, RN 
                           => n12536, Q => n_2797, QN => n14216);
   REGISTERS_reg_74_7_inst : DFFR_X1 port map( D => n8708_port, CK => CLK, RN 
                           => n12646, Q => n_2798, QN => n14217);
   REGISTERS_reg_74_6_inst : DFFR_X1 port map( D => n8709_port, CK => CLK, RN 
                           => n12602, Q => n_2799, QN => n14218);
   REGISTERS_reg_74_5_inst : DFFR_X1 port map( D => n8710_port, CK => CLK, RN 
                           => n12489, Q => n_2800, QN => n14219);
   REGISTERS_reg_74_4_inst : DFFR_X1 port map( D => n8711_port, CK => CLK, RN 
                           => n12496, Q => n_2801, QN => n14220);
   REGISTERS_reg_74_3_inst : DFFR_X1 port map( D => n8712_port, CK => CLK, RN 
                           => n12580, Q => n_2802, QN => n14221);
   REGISTERS_reg_74_2_inst : DFFR_X1 port map( D => n8713_port, CK => CLK, RN 
                           => n12511, Q => n_2803, QN => n14222);
   REGISTERS_reg_74_1_inst : DFFR_X1 port map( D => n8714_port, CK => CLK, RN 
                           => n12439, Q => n_2804, QN => n14223);
   REGISTERS_reg_74_0_inst : DFFR_X1 port map( D => n8715_port, CK => CLK, RN 
                           => n12654, Q => n_2805, QN => n14224);
   REGISTERS_reg_75_31_inst : DFFR_X1 port map( D => n8716_port, CK => CLK, RN 
                           => n12661, Q => n_2806, QN => n868);
   REGISTERS_reg_75_30_inst : DFFR_X1 port map( D => n8717_port, CK => CLK, RN 
                           => n12624, Q => n_2807, QN => n872);
   REGISTERS_reg_75_29_inst : DFFR_X1 port map( D => n8718_port, CK => CLK, RN 
                           => n12610, Q => n_2808, QN => n876);
   REGISTERS_reg_75_28_inst : DFFR_X1 port map( D => n8719_port, CK => CLK, RN 
                           => n12617, Q => n_2809, QN => n880);
   REGISTERS_reg_75_27_inst : DFFR_X1 port map( D => n8720_port, CK => CLK, RN 
                           => n12588, Q => n_2810, QN => n884);
   REGISTERS_reg_75_26_inst : DFFR_X1 port map( D => n8721_port, CK => CLK, RN 
                           => n12566, Q => n_2811, QN => n888);
   REGISTERS_reg_75_25_inst : DFFR_X1 port map( D => n8722_port, CK => CLK, RN 
                           => n12544, Q => n_2812, QN => n892);
   REGISTERS_reg_75_24_inst : DFFR_X1 port map( D => n8723_port, CK => CLK, RN 
                           => n12465, Q => n_2813, QN => n896);
   REGISTERS_reg_75_23_inst : DFFR_X1 port map( D => n8724_port, CK => CLK, RN 
                           => n12632, Q => n_2814, QN => n900);
   REGISTERS_reg_75_22_inst : DFFR_X1 port map( D => n8725_port, CK => CLK, RN 
                           => n12522, Q => n_2815, QN => n904);
   REGISTERS_reg_75_21_inst : DFFR_X1 port map( D => n8726_port, CK => CLK, RN 
                           => n12529, Q => n_2816, QN => n908);
   REGISTERS_reg_75_20_inst : DFFR_X1 port map( D => n8727_port, CK => CLK, RN 
                           => n12504, Q => n_2817, QN => n912);
   REGISTERS_reg_75_19_inst : DFFR_X1 port map( D => n8728_port, CK => CLK, RN 
                           => n12595, Q => n_2818, QN => n916);
   REGISTERS_reg_75_18_inst : DFFR_X1 port map( D => n8729_port, CK => CLK, RN 
                           => n12446, Q => n_2819, QN => n920);
   REGISTERS_reg_75_17_inst : DFFR_X1 port map( D => n8730_port, CK => CLK, RN 
                           => n12453, Q => n_2820, QN => n924);
   REGISTERS_reg_75_16_inst : DFFR_X1 port map( D => n8731_port, CK => CLK, RN 
                           => n12460, Q => n_2821, QN => n928);
   REGISTERS_reg_75_15_inst : DFFR_X1 port map( D => n8732_port, CK => CLK, RN 
                           => n12639, Q => n_2822, QN => n932);
   REGISTERS_reg_75_14_inst : DFFR_X1 port map( D => n8733_port, CK => CLK, RN 
                           => n12467, Q => n_2823, QN => n936);
   REGISTERS_reg_75_13_inst : DFFR_X1 port map( D => n8734_port, CK => CLK, RN 
                           => n12474, Q => n_2824, QN => n940);
   REGISTERS_reg_75_12_inst : DFFR_X1 port map( D => n8735_port, CK => CLK, RN 
                           => n12482, Q => n_2825, QN => n944);
   REGISTERS_reg_75_11_inst : DFFR_X1 port map( D => n8736_port, CK => CLK, RN 
                           => n12573, Q => n_2826, QN => n948);
   REGISTERS_reg_75_10_inst : DFFR_X1 port map( D => n8737_port, CK => CLK, RN 
                           => n12551, Q => n_2827, QN => n952);
   REGISTERS_reg_75_9_inst : DFFR_X1 port map( D => n8738_port, CK => CLK, RN 
                           => n12558, Q => n_2828, QN => n956);
   REGISTERS_reg_75_8_inst : DFFR_X1 port map( D => n8739_port, CK => CLK, RN 
                           => n12536, Q => n_2829, QN => n960);
   REGISTERS_reg_75_7_inst : DFFR_X1 port map( D => n8740_port, CK => CLK, RN 
                           => n12646, Q => n_2830, QN => n964);
   REGISTERS_reg_75_6_inst : DFFR_X1 port map( D => n8741_port, CK => CLK, RN 
                           => n12602, Q => n_2831, QN => n968);
   REGISTERS_reg_75_5_inst : DFFR_X1 port map( D => n8742_port, CK => CLK, RN 
                           => n12489, Q => n_2832, QN => n972);
   REGISTERS_reg_75_4_inst : DFFR_X1 port map( D => n8743_port, CK => CLK, RN 
                           => n12496, Q => n_2833, QN => n976);
   REGISTERS_reg_75_3_inst : DFFR_X1 port map( D => n8744_port, CK => CLK, RN 
                           => n12580, Q => n_2834, QN => n980);
   REGISTERS_reg_75_2_inst : DFFR_X1 port map( D => n8745_port, CK => CLK, RN 
                           => n12511, Q => n_2835, QN => n984);
   REGISTERS_reg_75_1_inst : DFFR_X1 port map( D => n8746_port, CK => CLK, RN 
                           => n12439, Q => n_2836, QN => n988);
   REGISTERS_reg_75_0_inst : DFFR_X1 port map( D => n8747_port, CK => CLK, RN 
                           => n12654, Q => n_2837, QN => n992);
   REGISTERS_reg_76_31_inst : DFFR_X1 port map( D => n8748_port, CK => CLK, RN 
                           => n12661, Q => n_2838, QN => n14225);
   REGISTERS_reg_76_30_inst : DFFR_X1 port map( D => n8749_port, CK => CLK, RN 
                           => n12625, Q => n_2839, QN => n14226);
   REGISTERS_reg_76_29_inst : DFFR_X1 port map( D => n8750_port, CK => CLK, RN 
                           => n12610, Q => n_2840, QN => n14227);
   REGISTERS_reg_76_28_inst : DFFR_X1 port map( D => n8751_port, CK => CLK, RN 
                           => n12617, Q => n_2841, QN => n14228);
   REGISTERS_reg_76_27_inst : DFFR_X1 port map( D => n8752_port, CK => CLK, RN 
                           => n12588, Q => n_2842, QN => n14229);
   REGISTERS_reg_76_26_inst : DFFR_X1 port map( D => n8753_port, CK => CLK, RN 
                           => n12566, Q => n_2843, QN => n14230);
   REGISTERS_reg_76_25_inst : DFFR_X1 port map( D => n8754_port, CK => CLK, RN 
                           => n12544, Q => n_2844, QN => n14231);
   REGISTERS_reg_76_24_inst : DFFR_X1 port map( D => n8755_port, CK => CLK, RN 
                           => n12508, Q => n_2845, QN => n14232);
   REGISTERS_reg_76_23_inst : DFFR_X1 port map( D => n8756_port, CK => CLK, RN 
                           => n12632, Q => n_2846, QN => n14233);
   REGISTERS_reg_76_22_inst : DFFR_X1 port map( D => n8757_port, CK => CLK, RN 
                           => n12522, Q => n_2847, QN => n14234);
   REGISTERS_reg_76_21_inst : DFFR_X1 port map( D => n8758_port, CK => CLK, RN 
                           => n12529, Q => n_2848, QN => n14235);
   REGISTERS_reg_76_20_inst : DFFR_X1 port map( D => n8759_port, CK => CLK, RN 
                           => n12504, Q => n_2849, QN => n14236);
   REGISTERS_reg_76_19_inst : DFFR_X1 port map( D => n8760_port, CK => CLK, RN 
                           => n12595, Q => n_2850, QN => n14237);
   REGISTERS_reg_76_18_inst : DFFR_X1 port map( D => n8761_port, CK => CLK, RN 
                           => n12446, Q => n_2851, QN => n14238);
   REGISTERS_reg_76_17_inst : DFFR_X1 port map( D => n8762_port, CK => CLK, RN 
                           => n12454, Q => n_2852, QN => n14239);
   REGISTERS_reg_76_16_inst : DFFR_X1 port map( D => n8763_port, CK => CLK, RN 
                           => n12460, Q => n_2853, QN => n14240);
   REGISTERS_reg_76_15_inst : DFFR_X1 port map( D => n8764_port, CK => CLK, RN 
                           => n12639, Q => n_2854, QN => n14241);
   REGISTERS_reg_76_14_inst : DFFR_X1 port map( D => n8765_port, CK => CLK, RN 
                           => n12467, Q => n_2855, QN => n14242);
   REGISTERS_reg_76_13_inst : DFFR_X1 port map( D => n8766_port, CK => CLK, RN 
                           => n12475, Q => n_2856, QN => n14243);
   REGISTERS_reg_76_12_inst : DFFR_X1 port map( D => n8767_port, CK => CLK, RN 
                           => n12482, Q => n_2857, QN => n14244);
   REGISTERS_reg_76_11_inst : DFFR_X1 port map( D => n8768, CK => CLK, RN => 
                           n12573, Q => n_2858, QN => n14245);
   REGISTERS_reg_76_10_inst : DFFR_X1 port map( D => n8769, CK => CLK, RN => 
                           n12551, Q => n_2859, QN => n14246);
   REGISTERS_reg_76_9_inst : DFFR_X1 port map( D => n8770, CK => CLK, RN => 
                           n12559, Q => n_2860, QN => n14247);
   REGISTERS_reg_76_8_inst : DFFR_X1 port map( D => n8771, CK => CLK, RN => 
                           n12537, Q => n_2861, QN => n14248);
   REGISTERS_reg_76_7_inst : DFFR_X1 port map( D => n8772, CK => CLK, RN => 
                           n12647, Q => n_2862, QN => n14249);
   REGISTERS_reg_76_6_inst : DFFR_X1 port map( D => n8773, CK => CLK, RN => 
                           n12603, Q => n_2863, QN => n14250);
   REGISTERS_reg_76_5_inst : DFFR_X1 port map( D => n8774, CK => CLK, RN => 
                           n12489, Q => n_2864, QN => n14251);
   REGISTERS_reg_76_4_inst : DFFR_X1 port map( D => n8775, CK => CLK, RN => 
                           n12497, Q => n_2865, QN => n14252);
   REGISTERS_reg_76_3_inst : DFFR_X1 port map( D => n8776, CK => CLK, RN => 
                           n12581, Q => n_2866, QN => n14253);
   REGISTERS_reg_76_2_inst : DFFR_X1 port map( D => n8777, CK => CLK, RN => 
                           n12511, Q => n_2867, QN => n14254);
   REGISTERS_reg_76_1_inst : DFFR_X1 port map( D => n8778, CK => CLK, RN => 
                           n12439, Q => n_2868, QN => n14255);
   REGISTERS_reg_76_0_inst : DFFR_X1 port map( D => n8779, CK => CLK, RN => 
                           n12654, Q => n_2869, QN => n14256);
   REGISTERS_reg_78_31_inst : DFFR_X1 port map( D => n8812, CK => CLK, RN => 
                           n12661, Q => n_2870, QN => n5712);
   REGISTERS_reg_78_30_inst : DFFR_X1 port map( D => n8813, CK => CLK, RN => 
                           n12625, Q => n_2871, QN => n5744);
   REGISTERS_reg_78_29_inst : DFFR_X1 port map( D => n8814, CK => CLK, RN => 
                           n12610, Q => n_2872, QN => n5776);
   REGISTERS_reg_78_28_inst : DFFR_X1 port map( D => n8815, CK => CLK, RN => 
                           n12617, Q => n_2873, QN => n5808);
   REGISTERS_reg_78_27_inst : DFFR_X1 port map( D => n8816, CK => CLK, RN => 
                           n12588, Q => n_2874, QN => n5840);
   REGISTERS_reg_78_26_inst : DFFR_X1 port map( D => n8817, CK => CLK, RN => 
                           n12566, Q => n_2875, QN => n5872);
   REGISTERS_reg_78_25_inst : DFFR_X1 port map( D => n8818, CK => CLK, RN => 
                           n12544, Q => n_2876, QN => n5904);
   REGISTERS_reg_78_24_inst : DFFR_X1 port map( D => n8819, CK => CLK, RN => 
                           n12507, Q => n_2877, QN => n5936);
   REGISTERS_reg_78_23_inst : DFFR_X1 port map( D => n8820, CK => CLK, RN => 
                           n12632, Q => n_2878, QN => n6000);
   REGISTERS_reg_78_22_inst : DFFR_X1 port map( D => n8821, CK => CLK, RN => 
                           n12522, Q => n_2879, QN => n9135);
   REGISTERS_reg_78_21_inst : DFFR_X1 port map( D => n8822, CK => CLK, RN => 
                           n12529, Q => n_2880, QN => n9167);
   REGISTERS_reg_78_20_inst : DFFR_X1 port map( D => n8823, CK => CLK, RN => 
                           n12504, Q => n_2881, QN => n9199);
   REGISTERS_reg_78_19_inst : DFFR_X1 port map( D => n8824, CK => CLK, RN => 
                           n12595, Q => n_2882, QN => n9263);
   REGISTERS_reg_78_18_inst : DFFR_X1 port map( D => n8825, CK => CLK, RN => 
                           n12446, Q => n_2883, QN => n9597);
   REGISTERS_reg_78_17_inst : DFFR_X1 port map( D => n8826, CK => CLK, RN => 
                           n12454, Q => n_2884, QN => n9629);
   REGISTERS_reg_78_16_inst : DFFR_X1 port map( D => n8827, CK => CLK, RN => 
                           n12460, Q => n_2885, QN => n9661);
   REGISTERS_reg_78_15_inst : DFFR_X1 port map( D => n8828, CK => CLK, RN => 
                           n12639, Q => n_2886, QN => n10023);
   REGISTERS_reg_78_14_inst : DFFR_X1 port map( D => n8829, CK => CLK, RN => 
                           n12467, Q => n_2887, QN => n10055);
   REGISTERS_reg_78_13_inst : DFFR_X1 port map( D => n8830, CK => CLK, RN => 
                           n12475, Q => n_2888, QN => n10087);
   REGISTERS_reg_78_12_inst : DFFR_X1 port map( D => n8831, CK => CLK, RN => 
                           n12482, Q => n_2889, QN => n10119);
   REGISTERS_reg_78_11_inst : DFFR_X1 port map( D => n8832, CK => CLK, RN => 
                           n12573, Q => n_2890, QN => n10151);
   REGISTERS_reg_78_10_inst : DFFR_X1 port map( D => n8833, CK => CLK, RN => 
                           n12551, Q => n_2891, QN => n10183);
   REGISTERS_reg_78_9_inst : DFFR_X1 port map( D => n8834, CK => CLK, RN => 
                           n12559, Q => n_2892, QN => n10217);
   REGISTERS_reg_78_8_inst : DFFR_X1 port map( D => n8835, CK => CLK, RN => 
                           n12537, Q => n_2893, QN => n10249);
   REGISTERS_reg_78_7_inst : DFFR_X1 port map( D => n8836, CK => CLK, RN => 
                           n12647, Q => n_2894, QN => n10281);
   REGISTERS_reg_78_6_inst : DFFR_X1 port map( D => n8837, CK => CLK, RN => 
                           n12603, Q => n_2895, QN => n10316);
   REGISTERS_reg_78_5_inst : DFFR_X1 port map( D => n8838, CK => CLK, RN => 
                           n12489, Q => n_2896, QN => n10348);
   REGISTERS_reg_78_4_inst : DFFR_X1 port map( D => n8839, CK => CLK, RN => 
                           n12497, Q => n_2897, QN => n10380);
   REGISTERS_reg_78_3_inst : DFFR_X1 port map( D => n8840, CK => CLK, RN => 
                           n12581, Q => n_2898, QN => n10415);
   REGISTERS_reg_78_2_inst : DFFR_X1 port map( D => n8841, CK => CLK, RN => 
                           n12511, Q => n_2899, QN => n10447);
   REGISTERS_reg_78_1_inst : DFFR_X1 port map( D => n8842, CK => CLK, RN => 
                           n12439, Q => n_2900, QN => n10479);
   REGISTERS_reg_78_0_inst : DFFR_X1 port map( D => n8843, CK => CLK, RN => 
                           n12654, Q => n_2901, QN => n10511);
   REGISTERS_reg_79_31_inst : DFFR_X1 port map( D => n8844, CK => CLK, RN => 
                           n12661, Q => n_2902, QN => n5710);
   REGISTERS_reg_79_30_inst : DFFR_X1 port map( D => n8845, CK => CLK, RN => 
                           n12625, Q => n_2903, QN => n5742);
   REGISTERS_reg_79_29_inst : DFFR_X1 port map( D => n8846, CK => CLK, RN => 
                           n12610, Q => n_2904, QN => n5774);
   REGISTERS_reg_79_28_inst : DFFR_X1 port map( D => n8847, CK => CLK, RN => 
                           n12617, Q => n_2905, QN => n5806);
   REGISTERS_reg_79_27_inst : DFFR_X1 port map( D => n8848, CK => CLK, RN => 
                           n12588, Q => n_2906, QN => n5838);
   REGISTERS_reg_79_26_inst : DFFR_X1 port map( D => n8849, CK => CLK, RN => 
                           n12566, Q => n_2907, QN => n5870);
   REGISTERS_reg_79_25_inst : DFFR_X1 port map( D => n8850, CK => CLK, RN => 
                           n12544, Q => n_2908, QN => n5902);
   REGISTERS_reg_79_24_inst : DFFR_X1 port map( D => n8851, CK => CLK, RN => 
                           n12506, Q => n_2909, QN => n5934);
   REGISTERS_reg_79_23_inst : DFFR_X1 port map( D => n8852, CK => CLK, RN => 
                           n12632, Q => n_2910, QN => n5998);
   REGISTERS_reg_79_22_inst : DFFR_X1 port map( D => n8853, CK => CLK, RN => 
                           n12522, Q => n_2911, QN => n6315);
   REGISTERS_reg_79_21_inst : DFFR_X1 port map( D => n8854, CK => CLK, RN => 
                           n12529, Q => n_2912, QN => n9165);
   REGISTERS_reg_79_20_inst : DFFR_X1 port map( D => n8855, CK => CLK, RN => 
                           n12504, Q => n_2913, QN => n9197);
   REGISTERS_reg_79_19_inst : DFFR_X1 port map( D => n8856, CK => CLK, RN => 
                           n12595, Q => n_2914, QN => n9261);
   REGISTERS_reg_79_18_inst : DFFR_X1 port map( D => n8857, CK => CLK, RN => 
                           n12446, Q => n_2915, QN => n9595);
   REGISTERS_reg_79_17_inst : DFFR_X1 port map( D => n8858, CK => CLK, RN => 
                           n12454, Q => n_2916, QN => n9627);
   REGISTERS_reg_79_16_inst : DFFR_X1 port map( D => n8859, CK => CLK, RN => 
                           n12460, Q => n_2917, QN => n9659);
   REGISTERS_reg_79_15_inst : DFFR_X1 port map( D => n8860, CK => CLK, RN => 
                           n12639, Q => n_2918, QN => n10021);
   REGISTERS_reg_79_14_inst : DFFR_X1 port map( D => n8861, CK => CLK, RN => 
                           n12467, Q => n_2919, QN => n10053);
   REGISTERS_reg_79_13_inst : DFFR_X1 port map( D => n8862, CK => CLK, RN => 
                           n12475, Q => n_2920, QN => n10085);
   REGISTERS_reg_79_12_inst : DFFR_X1 port map( D => n8863, CK => CLK, RN => 
                           n12482, Q => n_2921, QN => n10117);
   REGISTERS_reg_79_11_inst : DFFR_X1 port map( D => n8864, CK => CLK, RN => 
                           n12573, Q => n_2922, QN => n10149);
   REGISTERS_reg_79_10_inst : DFFR_X1 port map( D => n8865, CK => CLK, RN => 
                           n12551, Q => n_2923, QN => n10181);
   REGISTERS_reg_79_9_inst : DFFR_X1 port map( D => n8866, CK => CLK, RN => 
                           n12559, Q => n_2924, QN => n10215);
   REGISTERS_reg_79_8_inst : DFFR_X1 port map( D => n8867, CK => CLK, RN => 
                           n12537, Q => n_2925, QN => n10247);
   REGISTERS_reg_79_7_inst : DFFR_X1 port map( D => n8868, CK => CLK, RN => 
                           n12647, Q => n_2926, QN => n10279);
   REGISTERS_reg_79_6_inst : DFFR_X1 port map( D => n8869, CK => CLK, RN => 
                           n12603, Q => n_2927, QN => n10314);
   REGISTERS_reg_79_5_inst : DFFR_X1 port map( D => n8870, CK => CLK, RN => 
                           n12489, Q => n_2928, QN => n10346);
   REGISTERS_reg_79_4_inst : DFFR_X1 port map( D => n8871, CK => CLK, RN => 
                           n12497, Q => n_2929, QN => n10378);
   REGISTERS_reg_79_3_inst : DFFR_X1 port map( D => n8872, CK => CLK, RN => 
                           n12581, Q => n_2930, QN => n10413);
   REGISTERS_reg_79_2_inst : DFFR_X1 port map( D => n8873, CK => CLK, RN => 
                           n12511, Q => n_2931, QN => n10445);
   REGISTERS_reg_79_1_inst : DFFR_X1 port map( D => n8874, CK => CLK, RN => 
                           n12439, Q => n_2932, QN => n10477);
   REGISTERS_reg_79_0_inst : DFFR_X1 port map( D => n8875, CK => CLK, RN => 
                           n12654, Q => n_2933, QN => n10509);
   REGISTERS_reg_80_6_inst : DFFR_X1 port map( D => n8901, CK => CLK, RN => 
                           n12603, Q => n_2934, QN => n10315);
   REGISTERS_reg_80_5_inst : DFFR_X1 port map( D => n8902, CK => CLK, RN => 
                           n12490, Q => n_2935, QN => n10347);
   REGISTERS_reg_80_4_inst : DFFR_X1 port map( D => n8903, CK => CLK, RN => 
                           n12497, Q => n_2936, QN => n10379);
   REGISTERS_reg_80_3_inst : DFFR_X1 port map( D => n8904, CK => CLK, RN => 
                           n12581, Q => n_2937, QN => n10414);
   REGISTERS_reg_80_2_inst : DFFR_X1 port map( D => n8905, CK => CLK, RN => 
                           n12512, Q => n_2938, QN => n10446);
   REGISTERS_reg_80_1_inst : DFFR_X1 port map( D => n8906, CK => CLK, RN => 
                           n12439, Q => n_2939, QN => n10478);
   REGISTERS_reg_80_0_inst : DFFR_X1 port map( D => n8907, CK => CLK, RN => 
                           n12654, Q => n_2940, QN => n10510);
   OUT2_reg_31_inst : DLH_X1 port map( G => n12426, D => N8767, Q => OUT2(31));
   OUT1_reg_31_inst : DLH_X1 port map( G => n12429, D => N8734, Q => OUT1(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => n12428, D => N8766, Q => OUT2(30));
   OUT1_reg_30_inst : DLH_X1 port map( G => n12429, D => N8733, Q => OUT1(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => n12428, D => N8765, Q => OUT2(29));
   OUT1_reg_29_inst : DLH_X1 port map( G => n12429, D => N8732, Q => OUT1(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => n12426, D => N8764, Q => OUT2(28));
   OUT1_reg_28_inst : DLH_X1 port map( G => n12429, D => N8731, Q => OUT1(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => n12428, D => N8763, Q => OUT2(27));
   OUT1_reg_27_inst : DLH_X1 port map( G => n12429, D => N8730, Q => OUT1(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => n12428, D => N8762, Q => OUT2(26));
   OUT1_reg_26_inst : DLH_X1 port map( G => n12430, D => N8729, Q => OUT1(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => n12428, D => N8761, Q => OUT2(25));
   OUT1_reg_25_inst : DLH_X1 port map( G => n12430, D => N8728, Q => OUT1(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => n12428, D => N8760, Q => OUT2(24));
   OUT1_reg_24_inst : DLH_X1 port map( G => n12430, D => N8727, Q => OUT1(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => n12426, D => N8759, Q => OUT2(23));
   OUT1_reg_23_inst : DLH_X1 port map( G => n12429, D => N8726, Q => OUT1(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => n12428, D => N8758, Q => OUT2(22));
   OUT1_reg_22_inst : DLH_X1 port map( G => n12430, D => N8725, Q => OUT1(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => n12426, D => N8757, Q => OUT2(21));
   OUT1_reg_21_inst : DLH_X1 port map( G => n12430, D => N8724, Q => OUT1(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => n12427, D => N8756, Q => OUT2(20));
   OUT1_reg_20_inst : DLH_X1 port map( G => n12431, D => N8723, Q => OUT1(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => n12426, D => N8755, Q => OUT2(19));
   OUT1_reg_19_inst : DLH_X1 port map( G => n12429, D => N8722, Q => OUT1(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => n12427, D => N8754, Q => OUT2(18));
   OUT1_reg_18_inst : DLH_X1 port map( G => n12431, D => N8721, Q => OUT1(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => n12427, D => N8753, Q => OUT2(17));
   OUT1_reg_17_inst : DLH_X1 port map( G => n12431, D => N8720, Q => OUT1(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => n12427, D => N8752, Q => OUT2(16));
   OUT1_reg_16_inst : DLH_X1 port map( G => n12431, D => N8719, Q => OUT1(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => n12426, D => N8751, Q => OUT2(15));
   OUT1_reg_15_inst : DLH_X1 port map( G => n12429, D => N8718, Q => OUT1(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => n12427, D => N8750, Q => OUT2(14));
   OUT1_reg_14_inst : DLH_X1 port map( G => n12431, D => N8717, Q => OUT1(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => n12427, D => N8749, Q => OUT2(13));
   OUT1_reg_13_inst : DLH_X1 port map( G => n12431, D => N8716, Q => OUT1(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => n12427, D => N8748, Q => OUT2(12));
   OUT1_reg_12_inst : DLH_X1 port map( G => n12431, D => N8715, Q => OUT1(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => n12428, D => N8747, Q => OUT2(11));
   OUT1_reg_11_inst : DLH_X1 port map( G => n12430, D => N8714, Q => OUT1(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => n12428, D => N8746, Q => OUT2(10));
   OUT1_reg_10_inst : DLH_X1 port map( G => n12430, D => N8713, Q => OUT1(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => n12426, D => N8745, Q => OUT2(9));
   OUT1_reg_9_inst : DLH_X1 port map( G => n12430, D => N8712, Q => OUT1(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => n12428, D => N8744, Q => OUT2(8));
   OUT1_reg_8_inst : DLH_X1 port map( G => n12430, D => N8711, Q => OUT1(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => n12426, D => N8743, Q => OUT2(7));
   OUT1_reg_7_inst : DLH_X1 port map( G => n12429, D => N8710, Q => OUT1(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => n12426, D => N8742, Q => OUT2(6));
   OUT1_reg_6_inst : DLH_X1 port map( G => n12429, D => N8709, Q => OUT1(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => n12427, D => N8741, Q => OUT2(5));
   OUT1_reg_5_inst : DLH_X1 port map( G => n12431, D => N8708, Q => OUT1(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => n12427, D => N8740, Q => OUT2(4));
   OUT1_reg_4_inst : DLH_X1 port map( G => n12431, D => N8707, Q => OUT1(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => n12426, D => N8739, Q => OUT2(3));
   OUT1_reg_3_inst : DLH_X1 port map( G => n12430, D => N8706, Q => OUT1(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => n12427, D => N8738, Q => OUT2(2));
   OUT1_reg_2_inst : DLH_X1 port map( G => n12430, D => N8705, Q => OUT1(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => n12427, D => N8737, Q => OUT2(1));
   OUT1_reg_1_inst : DLH_X1 port map( G => n12431, D => N8704, Q => OUT1(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => n12426, D => N8736, Q => OUT2(0));
   OUT1_reg_0_inst : DLH_X1 port map( G => n12429, D => N8703, Q => OUT1(0));
   FILL <= '0';
   SPILL <= '0';
   BUSout(31) <= '0';
   BUSout(30) <= '0';
   BUSout(29) <= '0';
   BUSout(28) <= '0';
   BUSout(27) <= '0';
   BUSout(26) <= '0';
   BUSout(25) <= '0';
   BUSout(24) <= '0';
   BUSout(23) <= '0';
   BUSout(22) <= '0';
   BUSout(21) <= '0';
   BUSout(20) <= '0';
   BUSout(19) <= '0';
   BUSout(18) <= '0';
   BUSout(17) <= '0';
   BUSout(16) <= '0';
   BUSout(15) <= '0';
   BUSout(14) <= '0';
   BUSout(13) <= '0';
   BUSout(12) <= '0';
   BUSout(11) <= '0';
   BUSout(10) <= '0';
   BUSout(9) <= '0';
   BUSout(8) <= '0';
   BUSout(7) <= '0';
   BUSout(6) <= '0';
   BUSout(5) <= '0';
   BUSout(4) <= '0';
   BUSout(3) <= '0';
   BUSout(2) <= '0';
   BUSout(1) <= '0';
   BUSout(0) <= '0';
   U4359 : NOR3_X2 port map( A1 => N8580, A2 => N8581, A3 => N8579, ZN => n4219
                           );
   U5825 : NOR3_X2 port map( A1 => N8436, A2 => N8437, A3 => N8435, ZN => n5652
                           );
   U7835 : NAND3_X1 port map( A1 => n14517, A2 => n2483, A3 => RETRN, ZN => 
                           n2480);
   U7836 : NAND3_X1 port map( A1 => n2489, A2 => n14518, A3 => n14517, ZN => 
                           n2481);
   U7837 : NAND3_X1 port map( A1 => n2936, A2 => n2935, A3 => n2937, ZN => 
                           n2483);
   U7838 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => wr_signal, ZN => 
                           n2597);
   r486_U4 : XOR2_X1 port map( A => U3_U99_Z_5, B => r486_carry_5_port, Z => 
                           N8580);
   r486_U1_4 : FA_X1 port map( A => U3_U99_Z_4, B => ADD_RD2(4), CI => 
                           r486_carry_4_port, CO => r486_carry_5_port, S => 
                           N8579);
   r480_U4 : XOR2_X1 port map( A => U3_U98_Z_5, B => r480_carry_5_port, Z => 
                           N8436);
   r480_U1_4 : FA_X1 port map( A => U3_U98_Z_4, B => ADD_RD1(4), CI => 
                           r480_carry_4_port, CO => r480_carry_5_port, S => 
                           N8435);
   r472_U3 : XOR2_X1 port map( A => U3_U97_Z_5, B => r472_carry_5_port, Z => 
                           N2172);
   r472_U1_4 : FA_X1 port map( A => ADD_WR(4), B => U3_U97_Z_4, CI => 
                           r472_carry_4_port, CO => r472_carry_5_port, S => 
                           N2171);
   REGISTERS_reg_87_31_inst : DFFR_X1 port map( D => n9100, CK => CLK, RN => 
                           RESET, Q => n14481, QN => n2882);
   REGISTERS_reg_87_30_inst : DFFR_X1 port map( D => n9101, CK => CLK, RN => 
                           n12625, Q => n14482, QN => n2883);
   REGISTERS_reg_87_29_inst : DFFR_X1 port map( D => n9102, CK => CLK, RN => 
                           n12611, Q => n14483, QN => n2884);
   REGISTERS_reg_87_28_inst : DFFR_X1 port map( D => n9103, CK => CLK, RN => 
                           n12618, Q => n14484, QN => n2885);
   REGISTERS_reg_87_27_inst : DFFR_X1 port map( D => n9104, CK => CLK, RN => 
                           n12589, Q => n14485, QN => n2886);
   REGISTERS_reg_87_26_inst : DFFR_X1 port map( D => n9105, CK => CLK, RN => 
                           n12567, Q => n14486, QN => n2887);
   REGISTERS_reg_87_25_inst : DFFR_X1 port map( D => n9106, CK => CLK, RN => 
                           n12545, Q => n14487, QN => n2888);
   REGISTERS_reg_87_24_inst : DFFR_X1 port map( D => n9107, CK => CLK, RN => 
                           n12505, Q => n14488, QN => n2889);
   REGISTERS_reg_87_23_inst : DFFR_X1 port map( D => n9108, CK => CLK, RN => 
                           n12633, Q => n14489, QN => n2890);
   REGISTERS_reg_87_22_inst : DFFR_X1 port map( D => n9109, CK => CLK, RN => 
                           n12523, Q => n14490, QN => n2891);
   REGISTERS_reg_87_21_inst : DFFR_X1 port map( D => n9110, CK => CLK, RN => 
                           n12530, Q => n14491, QN => n2892);
   REGISTERS_reg_87_20_inst : DFFR_X1 port map( D => n9111, CK => CLK, RN => 
                           n12505, Q => n14492, QN => n2893);
   REGISTERS_reg_87_19_inst : DFFR_X1 port map( D => n9112, CK => CLK, RN => 
                           n12596, Q => n14493, QN => n2894);
   REGISTERS_reg_87_18_inst : DFFR_X1 port map( D => n9113, CK => CLK, RN => 
                           n12447, Q => n14494, QN => n2895);
   REGISTERS_reg_87_17_inst : DFFR_X1 port map( D => n9114, CK => CLK, RN => 
                           n12454, Q => n14495, QN => n2896);
   REGISTERS_reg_87_16_inst : DFFR_X1 port map( D => n9115, CK => CLK, RN => 
                           n12461, Q => n14496, QN => n2897);
   REGISTERS_reg_87_15_inst : DFFR_X1 port map( D => n9116, CK => CLK, RN => 
                           n12640, Q => n14497, QN => n2898);
   REGISTERS_reg_87_14_inst : DFFR_X1 port map( D => n9117, CK => CLK, RN => 
                           n12468, Q => n14498, QN => n2899);
   REGISTERS_reg_87_13_inst : DFFR_X1 port map( D => n9118, CK => CLK, RN => 
                           n12475, Q => n14499, QN => n2900);
   REGISTERS_reg_87_12_inst : DFFR_X1 port map( D => n9119, CK => CLK, RN => 
                           n12483, Q => n14500, QN => n2901);
   REGISTERS_reg_87_11_inst : DFFR_X1 port map( D => n9120, CK => CLK, RN => 
                           n12574, Q => n14501, QN => n2902);
   REGISTERS_reg_87_10_inst : DFFR_X1 port map( D => n9121, CK => CLK, RN => 
                           n12552, Q => n14502, QN => n2903);
   REGISTERS_reg_87_9_inst : DFFR_X1 port map( D => n9122, CK => CLK, RN => 
                           n12559, Q => n14503, QN => n2904);
   REGISTERS_reg_87_8_inst : DFFR_X1 port map( D => n9123, CK => CLK, RN => 
                           n12537, Q => n14504, QN => n2905);
   REGISTERS_reg_87_7_inst : DFFR_X1 port map( D => n9124, CK => CLK, RN => 
                           n12647, Q => n14505, QN => n2906);
   REGISTERS_reg_87_6_inst : DFFR_X1 port map( D => n9125, CK => CLK, RN => 
                           n12603, Q => n14506, QN => n2907);
   REGISTERS_reg_87_5_inst : DFFR_X1 port map( D => n9126, CK => CLK, RN => 
                           n12490, Q => n14507, QN => n2908);
   REGISTERS_reg_87_4_inst : DFFR_X1 port map( D => n9127, CK => CLK, RN => 
                           n12497, Q => n14508, QN => n2909);
   REGISTERS_reg_87_3_inst : DFFR_X1 port map( D => n9128, CK => CLK, RN => 
                           n12581, Q => n14509, QN => n2910);
   REGISTERS_reg_87_2_inst : DFFR_X1 port map( D => n9129, CK => CLK, RN => 
                           n12512, Q => n14510, QN => n2911);
   REGISTERS_reg_87_1_inst : DFFR_X1 port map( D => n9130, CK => CLK, RN => 
                           n12440, Q => n14511, QN => n2912);
   REGISTERS_reg_87_0_inst : DFFR_X1 port map( D => n9131, CK => CLK, RN => 
                           n12655, Q => n14512, QN => n2913);
   REGISTERS_reg_86_31_inst : DFFR_X1 port map( D => n9068, CK => CLK, RN => 
                           n12662, Q => n14449, QN => n5714);
   REGISTERS_reg_86_30_inst : DFFR_X1 port map( D => n9069, CK => CLK, RN => 
                           n12625, Q => n14450, QN => n5746);
   REGISTERS_reg_86_29_inst : DFFR_X1 port map( D => n9070, CK => CLK, RN => 
                           n12611, Q => n14451, QN => n5778);
   REGISTERS_reg_86_28_inst : DFFR_X1 port map( D => n9071, CK => CLK, RN => 
                           n12618, Q => n14452, QN => n5810);
   REGISTERS_reg_86_27_inst : DFFR_X1 port map( D => n9072, CK => CLK, RN => 
                           n12589, Q => n14453, QN => n5842);
   REGISTERS_reg_86_26_inst : DFFR_X1 port map( D => n9073, CK => CLK, RN => 
                           n12567, Q => n14454, QN => n5874);
   REGISTERS_reg_86_25_inst : DFFR_X1 port map( D => n9074, CK => CLK, RN => 
                           n12545, Q => n14455, QN => n5906);
   REGISTERS_reg_86_24_inst : DFFR_X1 port map( D => n9075, CK => CLK, RN => 
                           n12504, Q => n14456, QN => n5938);
   REGISTERS_reg_86_23_inst : DFFR_X1 port map( D => n9076, CK => CLK, RN => 
                           n12633, Q => n14457, QN => n6002);
   REGISTERS_reg_86_22_inst : DFFR_X1 port map( D => n9077, CK => CLK, RN => 
                           n12523, Q => n14458, QN => n9137);
   REGISTERS_reg_86_21_inst : DFFR_X1 port map( D => n9078, CK => CLK, RN => 
                           n12530, Q => n14459, QN => n9169);
   REGISTERS_reg_86_20_inst : DFFR_X1 port map( D => n9079, CK => CLK, RN => 
                           n12505, Q => n14460, QN => n9201);
   REGISTERS_reg_86_19_inst : DFFR_X1 port map( D => n9080, CK => CLK, RN => 
                           n12596, Q => n14461, QN => n9311);
   REGISTERS_reg_86_18_inst : DFFR_X1 port map( D => n9081, CK => CLK, RN => 
                           n12447, Q => n14462, QN => n9599);
   REGISTERS_reg_86_17_inst : DFFR_X1 port map( D => n9082, CK => CLK, RN => 
                           n12454, Q => n14463, QN => n9631);
   REGISTERS_reg_86_16_inst : DFFR_X1 port map( D => n9083, CK => CLK, RN => 
                           n12461, Q => n14464, QN => n9663);
   REGISTERS_reg_86_15_inst : DFFR_X1 port map( D => n9084, CK => CLK, RN => 
                           n12640, Q => n14465, QN => n10025);
   REGISTERS_reg_86_14_inst : DFFR_X1 port map( D => n9085, CK => CLK, RN => 
                           n12468, Q => n14466, QN => n10057);
   REGISTERS_reg_86_13_inst : DFFR_X1 port map( D => n9086, CK => CLK, RN => 
                           n12475, Q => n14467, QN => n10089);
   REGISTERS_reg_86_12_inst : DFFR_X1 port map( D => n9087, CK => CLK, RN => 
                           n12483, Q => n14468, QN => n10121);
   REGISTERS_reg_86_11_inst : DFFR_X1 port map( D => n9088, CK => CLK, RN => 
                           n12574, Q => n14469, QN => n10153);
   REGISTERS_reg_86_10_inst : DFFR_X1 port map( D => n9089, CK => CLK, RN => 
                           n12552, Q => n14470, QN => n10185);
   REGISTERS_reg_86_9_inst : DFFR_X1 port map( D => n9090, CK => CLK, RN => 
                           n12559, Q => n14471, QN => n10219);
   REGISTERS_reg_86_8_inst : DFFR_X1 port map( D => n9091, CK => CLK, RN => 
                           n12537, Q => n14472, QN => n10251);
   REGISTERS_reg_86_7_inst : DFFR_X1 port map( D => n9092, CK => CLK, RN => 
                           n12647, Q => n14473, QN => n10283);
   REGISTERS_reg_86_6_inst : DFFR_X1 port map( D => n9093, CK => CLK, RN => 
                           n12603, Q => n14474, QN => n10318);
   REGISTERS_reg_86_5_inst : DFFR_X1 port map( D => n9094, CK => CLK, RN => 
                           n12490, Q => n14475, QN => n10350);
   REGISTERS_reg_86_4_inst : DFFR_X1 port map( D => n9095, CK => CLK, RN => 
                           n12497, Q => n14476, QN => n10382);
   REGISTERS_reg_86_3_inst : DFFR_X1 port map( D => n9096, CK => CLK, RN => 
                           n12581, Q => n14477, QN => n10417);
   REGISTERS_reg_86_2_inst : DFFR_X1 port map( D => n9097, CK => CLK, RN => 
                           n12512, Q => n14478, QN => n10449);
   REGISTERS_reg_86_1_inst : DFFR_X1 port map( D => n9098, CK => CLK, RN => 
                           n12440, Q => n14479, QN => n10481);
   REGISTERS_reg_86_0_inst : DFFR_X1 port map( D => n9099, CK => CLK, RN => 
                           n12655, Q => n14480, QN => n10513);
   REGISTERS_reg_85_31_inst : DFFR_X1 port map( D => n9036, CK => CLK, RN => 
                           n12662, Q => n14417, QN => n2818);
   REGISTERS_reg_85_30_inst : DFFR_X1 port map( D => n9037, CK => CLK, RN => 
                           n12625, Q => n14418, QN => n2819);
   REGISTERS_reg_85_29_inst : DFFR_X1 port map( D => n9038, CK => CLK, RN => 
                           n12611, Q => n14419, QN => n2820);
   REGISTERS_reg_85_28_inst : DFFR_X1 port map( D => n9039, CK => CLK, RN => 
                           n12618, Q => n14420, QN => n2821);
   REGISTERS_reg_85_27_inst : DFFR_X1 port map( D => n9040, CK => CLK, RN => 
                           n12589, Q => n14421, QN => n2822);
   REGISTERS_reg_85_26_inst : DFFR_X1 port map( D => n9041, CK => CLK, RN => 
                           n12567, Q => n14422, QN => n2823);
   REGISTERS_reg_85_25_inst : DFFR_X1 port map( D => n9042, CK => CLK, RN => 
                           n12545, Q => n14423, QN => n2824);
   REGISTERS_reg_85_24_inst : DFFR_X1 port map( D => n9043, CK => CLK, RN => 
                           n12503, Q => n14424, QN => n2825);
   REGISTERS_reg_85_23_inst : DFFR_X1 port map( D => n9044, CK => CLK, RN => 
                           n12633, Q => n14425, QN => n2826);
   REGISTERS_reg_85_22_inst : DFFR_X1 port map( D => n9045, CK => CLK, RN => 
                           n12523, Q => n14426, QN => n2827);
   REGISTERS_reg_85_21_inst : DFFR_X1 port map( D => n9046, CK => CLK, RN => 
                           n12530, Q => n14427, QN => n2828);
   REGISTERS_reg_85_20_inst : DFFR_X1 port map( D => n9047, CK => CLK, RN => 
                           n12505, Q => n14428, QN => n2829);
   REGISTERS_reg_85_19_inst : DFFR_X1 port map( D => n9048, CK => CLK, RN => 
                           n12596, Q => n14429, QN => n2830);
   REGISTERS_reg_85_18_inst : DFFR_X1 port map( D => n9049, CK => CLK, RN => 
                           n12447, Q => n14430, QN => n2831);
   REGISTERS_reg_85_17_inst : DFFR_X1 port map( D => n9050, CK => CLK, RN => 
                           n12454, Q => n14431, QN => n2832);
   REGISTERS_reg_85_16_inst : DFFR_X1 port map( D => n9051, CK => CLK, RN => 
                           n12461, Q => n14432, QN => n2833);
   REGISTERS_reg_85_15_inst : DFFR_X1 port map( D => n9052, CK => CLK, RN => 
                           n12640, Q => n14433, QN => n2834);
   REGISTERS_reg_85_14_inst : DFFR_X1 port map( D => n9053, CK => CLK, RN => 
                           n12468, Q => n14434, QN => n2835);
   REGISTERS_reg_85_13_inst : DFFR_X1 port map( D => n9054, CK => CLK, RN => 
                           n12475, Q => n14435, QN => n2836);
   REGISTERS_reg_85_12_inst : DFFR_X1 port map( D => n9055, CK => CLK, RN => 
                           n12483, Q => n14436, QN => n2837);
   REGISTERS_reg_85_11_inst : DFFR_X1 port map( D => n9056, CK => CLK, RN => 
                           n12574, Q => n14437, QN => n2838);
   REGISTERS_reg_85_10_inst : DFFR_X1 port map( D => n9057, CK => CLK, RN => 
                           n12552, Q => n14438, QN => n2839);
   REGISTERS_reg_85_9_inst : DFFR_X1 port map( D => n9058, CK => CLK, RN => 
                           n12559, Q => n14439, QN => n2840);
   REGISTERS_reg_85_8_inst : DFFR_X1 port map( D => n9059, CK => CLK, RN => 
                           n12537, Q => n14440, QN => n2841);
   REGISTERS_reg_85_7_inst : DFFR_X1 port map( D => n9060, CK => CLK, RN => 
                           n12647, Q => n14441, QN => n2842);
   REGISTERS_reg_85_6_inst : DFFR_X1 port map( D => n9061, CK => CLK, RN => 
                           n12603, Q => n14442, QN => n2843);
   REGISTERS_reg_85_5_inst : DFFR_X1 port map( D => n9062, CK => CLK, RN => 
                           n12490, Q => n14443, QN => n2844);
   REGISTERS_reg_85_4_inst : DFFR_X1 port map( D => n9063, CK => CLK, RN => 
                           n12497, Q => n14444, QN => n2845);
   REGISTERS_reg_85_3_inst : DFFR_X1 port map( D => n9064, CK => CLK, RN => 
                           n12581, Q => n14445, QN => n2846);
   REGISTERS_reg_85_2_inst : DFFR_X1 port map( D => n9065, CK => CLK, RN => 
                           n12512, Q => n14446, QN => n2847);
   REGISTERS_reg_85_1_inst : DFFR_X1 port map( D => n9066, CK => CLK, RN => 
                           n12440, Q => n14447, QN => n2848);
   REGISTERS_reg_85_0_inst : DFFR_X1 port map( D => n9067, CK => CLK, RN => 
                           n12655, Q => n14448, QN => n2849);
   REGISTERS_reg_84_31_inst : DFFR_X1 port map( D => n9004, CK => CLK, RN => 
                           n12662, Q => n14385, QN => n5708);
   REGISTERS_reg_84_30_inst : DFFR_X1 port map( D => n9005, CK => CLK, RN => 
                           n12625, Q => n14386, QN => n5740);
   REGISTERS_reg_84_29_inst : DFFR_X1 port map( D => n9006, CK => CLK, RN => 
                           n12611, Q => n14387, QN => n5772);
   REGISTERS_reg_84_28_inst : DFFR_X1 port map( D => n9007, CK => CLK, RN => 
                           n12618, Q => n14388, QN => n5804);
   REGISTERS_reg_84_27_inst : DFFR_X1 port map( D => n9008, CK => CLK, RN => 
                           n12589, Q => n14389, QN => n5836);
   REGISTERS_reg_84_26_inst : DFFR_X1 port map( D => n9009, CK => CLK, RN => 
                           n12567, Q => n14390, QN => n5868);
   REGISTERS_reg_84_25_inst : DFFR_X1 port map( D => n9010, CK => CLK, RN => 
                           n12545, Q => n14391, QN => n5900);
   REGISTERS_reg_84_24_inst : DFFR_X1 port map( D => n9011, CK => CLK, RN => 
                           n12509, Q => n14392, QN => n5932);
   REGISTERS_reg_84_23_inst : DFFR_X1 port map( D => n9012, CK => CLK, RN => 
                           n12633, Q => n14393, QN => n5996);
   REGISTERS_reg_84_22_inst : DFFR_X1 port map( D => n9013, CK => CLK, RN => 
                           n12523, Q => n14394, QN => n6313);
   REGISTERS_reg_84_21_inst : DFFR_X1 port map( D => n9014, CK => CLK, RN => 
                           n12530, Q => n14395, QN => n9163);
   REGISTERS_reg_84_20_inst : DFFR_X1 port map( D => n9015, CK => CLK, RN => 
                           n12505, Q => n14396, QN => n9195);
   REGISTERS_reg_84_19_inst : DFFR_X1 port map( D => n9016, CK => CLK, RN => 
                           n12596, Q => n14397, QN => n9259);
   REGISTERS_reg_84_18_inst : DFFR_X1 port map( D => n9017, CK => CLK, RN => 
                           n12447, Q => n14398, QN => n9593);
   REGISTERS_reg_84_17_inst : DFFR_X1 port map( D => n9018, CK => CLK, RN => 
                           n12454, Q => n14399, QN => n9625);
   REGISTERS_reg_84_16_inst : DFFR_X1 port map( D => n9019, CK => CLK, RN => 
                           n12461, Q => n14400, QN => n9657);
   REGISTERS_reg_84_15_inst : DFFR_X1 port map( D => n9020, CK => CLK, RN => 
                           n12640, Q => n14401, QN => n10019);
   REGISTERS_reg_84_14_inst : DFFR_X1 port map( D => n9021, CK => CLK, RN => 
                           n12468, Q => n14402, QN => n10051);
   REGISTERS_reg_84_13_inst : DFFR_X1 port map( D => n9022, CK => CLK, RN => 
                           n12475, Q => n14403, QN => n10083);
   REGISTERS_reg_84_12_inst : DFFR_X1 port map( D => n9023, CK => CLK, RN => 
                           n12483, Q => n14404, QN => n10115);
   REGISTERS_reg_84_11_inst : DFFR_X1 port map( D => n9024, CK => CLK, RN => 
                           n12574, Q => n14405, QN => n10147);
   REGISTERS_reg_84_10_inst : DFFR_X1 port map( D => n9025, CK => CLK, RN => 
                           n12552, Q => n14406, QN => n10179);
   REGISTERS_reg_84_9_inst : DFFR_X1 port map( D => n9026, CK => CLK, RN => 
                           n12559, Q => n14407, QN => n10213);
   REGISTERS_reg_84_8_inst : DFFR_X1 port map( D => n9027, CK => CLK, RN => 
                           n12537, Q => n14408, QN => n10245);
   REGISTERS_reg_84_7_inst : DFFR_X1 port map( D => n9028, CK => CLK, RN => 
                           n12647, Q => n14409, QN => n10277);
   REGISTERS_reg_84_6_inst : DFFR_X1 port map( D => n9029, CK => CLK, RN => 
                           n12603, Q => n14410, QN => n10312);
   REGISTERS_reg_84_5_inst : DFFR_X1 port map( D => n9030, CK => CLK, RN => 
                           n12490, Q => n14411, QN => n10344);
   REGISTERS_reg_84_4_inst : DFFR_X1 port map( D => n9031, CK => CLK, RN => 
                           n12497, Q => n14412, QN => n10376);
   REGISTERS_reg_84_3_inst : DFFR_X1 port map( D => n9032, CK => CLK, RN => 
                           n12581, Q => n14413, QN => n10411);
   REGISTERS_reg_84_2_inst : DFFR_X1 port map( D => n9033, CK => CLK, RN => 
                           n12512, Q => n14414, QN => n10443);
   REGISTERS_reg_84_1_inst : DFFR_X1 port map( D => n9034, CK => CLK, RN => 
                           n12440, Q => n14415, QN => n10475);
   REGISTERS_reg_84_0_inst : DFFR_X1 port map( D => n9035, CK => CLK, RN => 
                           n12655, Q => n14416, QN => n10507);
   REGISTERS_reg_83_31_inst : DFFR_X1 port map( D => n8972, CK => CLK, RN => 
                           n12662, Q => n14353, QN => n2754);
   REGISTERS_reg_83_30_inst : DFFR_X1 port map( D => n8973, CK => CLK, RN => 
                           n12625, Q => n14354, QN => n2755);
   REGISTERS_reg_83_29_inst : DFFR_X1 port map( D => n8974, CK => CLK, RN => 
                           n12610, Q => n14355, QN => n2756);
   REGISTERS_reg_83_28_inst : DFFR_X1 port map( D => n8975, CK => CLK, RN => 
                           n12618, Q => n14356, QN => n2757);
   REGISTERS_reg_83_27_inst : DFFR_X1 port map( D => n8976, CK => CLK, RN => 
                           n12588, Q => n14357, QN => n2758);
   REGISTERS_reg_83_26_inst : DFFR_X1 port map( D => n8977, CK => CLK, RN => 
                           n12566, Q => n14358, QN => n2759);
   REGISTERS_reg_83_25_inst : DFFR_X1 port map( D => n8978, CK => CLK, RN => 
                           n12544, Q => n14359, QN => n2760);
   REGISTERS_reg_83_24_inst : DFFR_X1 port map( D => n8979, CK => CLK, RN => 
                           n12454, Q => n14360, QN => n2761);
   REGISTERS_reg_83_23_inst : DFFR_X1 port map( D => n8980, CK => CLK, RN => 
                           n12632, Q => n14361, QN => n2762);
   REGISTERS_reg_83_22_inst : DFFR_X1 port map( D => n8981, CK => CLK, RN => 
                           n12522, Q => n14362, QN => n2763);
   REGISTERS_reg_83_21_inst : DFFR_X1 port map( D => n8982, CK => CLK, RN => 
                           n12530, Q => n14363, QN => n2764);
   REGISTERS_reg_83_20_inst : DFFR_X1 port map( D => n8983, CK => CLK, RN => 
                           n12504, Q => n14364, QN => n2765);
   REGISTERS_reg_83_19_inst : DFFR_X1 port map( D => n8984, CK => CLK, RN => 
                           n12596, Q => n14365, QN => n2766);
   REGISTERS_reg_83_18_inst : DFFR_X1 port map( D => n8985, CK => CLK, RN => 
                           n12447, Q => n14366, QN => n2767);
   REGISTERS_reg_83_17_inst : DFFR_X1 port map( D => n8986, CK => CLK, RN => 
                           n12454, Q => n14367, QN => n2768);
   REGISTERS_reg_83_16_inst : DFFR_X1 port map( D => n8987, CK => CLK, RN => 
                           n12460, Q => n14368, QN => n2769);
   REGISTERS_reg_83_15_inst : DFFR_X1 port map( D => n8988, CK => CLK, RN => 
                           n12640, Q => n14369, QN => n2770);
   REGISTERS_reg_83_14_inst : DFFR_X1 port map( D => n8989, CK => CLK, RN => 
                           n12468, Q => n14370, QN => n2771);
   REGISTERS_reg_83_13_inst : DFFR_X1 port map( D => n8990, CK => CLK, RN => 
                           n12475, Q => n14371, QN => n2772);
   REGISTERS_reg_83_12_inst : DFFR_X1 port map( D => n8991, CK => CLK, RN => 
                           n12482, Q => n14372, QN => n2773);
   REGISTERS_reg_83_11_inst : DFFR_X1 port map( D => n8992, CK => CLK, RN => 
                           n12574, Q => n14373, QN => n2774);
   REGISTERS_reg_83_10_inst : DFFR_X1 port map( D => n8993, CK => CLK, RN => 
                           n12552, Q => n14374, QN => n2775);
   REGISTERS_reg_83_9_inst : DFFR_X1 port map( D => n8994, CK => CLK, RN => 
                           n12559, Q => n14375, QN => n2776);
   REGISTERS_reg_83_8_inst : DFFR_X1 port map( D => n8995, CK => CLK, RN => 
                           n12537, Q => n14376, QN => n2777);
   REGISTERS_reg_83_7_inst : DFFR_X1 port map( D => n8996, CK => CLK, RN => 
                           n12647, Q => n14377, QN => n2778);
   REGISTERS_reg_83_6_inst : DFFR_X1 port map( D => n8997, CK => CLK, RN => 
                           n12603, Q => n14378, QN => n2779);
   REGISTERS_reg_83_5_inst : DFFR_X1 port map( D => n8998, CK => CLK, RN => 
                           n12490, Q => n14379, QN => n2780);
   REGISTERS_reg_83_4_inst : DFFR_X1 port map( D => n8999, CK => CLK, RN => 
                           n12497, Q => n14380, QN => n2781);
   REGISTERS_reg_83_3_inst : DFFR_X1 port map( D => n9000, CK => CLK, RN => 
                           n12581, Q => n14381, QN => n2782);
   REGISTERS_reg_83_2_inst : DFFR_X1 port map( D => n9001, CK => CLK, RN => 
                           n12512, Q => n14382, QN => n2783);
   REGISTERS_reg_83_1_inst : DFFR_X1 port map( D => n9002, CK => CLK, RN => 
                           n12439, Q => n14383, QN => n2784);
   REGISTERS_reg_83_0_inst : DFFR_X1 port map( D => n9003, CK => CLK, RN => 
                           n12654, Q => n14384, QN => n2785);
   REGISTERS_reg_82_31_inst : DFFR_X1 port map( D => n8940, CK => CLK, RN => 
                           n12662, Q => n14321, QN => n5707);
   REGISTERS_reg_82_30_inst : DFFR_X1 port map( D => n8941, CK => CLK, RN => 
                           n12625, Q => n14322, QN => n5739);
   REGISTERS_reg_82_29_inst : DFFR_X1 port map( D => n8942, CK => CLK, RN => 
                           n12610, Q => n14323, QN => n5771);
   REGISTERS_reg_82_28_inst : DFFR_X1 port map( D => n8943, CK => CLK, RN => 
                           n12618, Q => n14324, QN => n5803);
   REGISTERS_reg_82_27_inst : DFFR_X1 port map( D => n8944, CK => CLK, RN => 
                           n12588, Q => n14325, QN => n5835);
   REGISTERS_reg_82_26_inst : DFFR_X1 port map( D => n8945, CK => CLK, RN => 
                           n12566, Q => n14326, QN => n5867);
   REGISTERS_reg_82_25_inst : DFFR_X1 port map( D => n8946, CK => CLK, RN => 
                           n12544, Q => n14327, QN => n5899);
   REGISTERS_reg_82_24_inst : DFFR_X1 port map( D => n8947, CK => CLK, RN => 
                           n12453, Q => n14328, QN => n5931);
   REGISTERS_reg_82_23_inst : DFFR_X1 port map( D => n8948, CK => CLK, RN => 
                           n12632, Q => n14329, QN => n5995);
   REGISTERS_reg_82_22_inst : DFFR_X1 port map( D => n8949, CK => CLK, RN => 
                           n12522, Q => n14330, QN => n6312);
   REGISTERS_reg_82_21_inst : DFFR_X1 port map( D => n8950, CK => CLK, RN => 
                           n12530, Q => n14331, QN => n9162);
   REGISTERS_reg_82_20_inst : DFFR_X1 port map( D => n8951, CK => CLK, RN => 
                           n12504, Q => n14332, QN => n9194);
   REGISTERS_reg_82_19_inst : DFFR_X1 port map( D => n8952, CK => CLK, RN => 
                           n12596, Q => n14333, QN => n9258);
   REGISTERS_reg_82_18_inst : DFFR_X1 port map( D => n8953, CK => CLK, RN => 
                           n12447, Q => n14334, QN => n9592);
   REGISTERS_reg_82_17_inst : DFFR_X1 port map( D => n8954, CK => CLK, RN => 
                           n12454, Q => n14335, QN => n9624);
   REGISTERS_reg_82_16_inst : DFFR_X1 port map( D => n8955, CK => CLK, RN => 
                           n12460, Q => n14336, QN => n9656);
   REGISTERS_reg_82_15_inst : DFFR_X1 port map( D => n8956, CK => CLK, RN => 
                           n12640, Q => n14337, QN => n10018);
   REGISTERS_reg_82_14_inst : DFFR_X1 port map( D => n8957, CK => CLK, RN => 
                           n12468, Q => n14338, QN => n10050);
   REGISTERS_reg_82_13_inst : DFFR_X1 port map( D => n8958, CK => CLK, RN => 
                           n12475, Q => n14339, QN => n10082);
   REGISTERS_reg_82_12_inst : DFFR_X1 port map( D => n8959, CK => CLK, RN => 
                           n12482, Q => n14340, QN => n10114);
   REGISTERS_reg_82_11_inst : DFFR_X1 port map( D => n8960, CK => CLK, RN => 
                           n12574, Q => n14341, QN => n10146);
   REGISTERS_reg_82_10_inst : DFFR_X1 port map( D => n8961, CK => CLK, RN => 
                           n12552, Q => n14342, QN => n10178);
   REGISTERS_reg_82_9_inst : DFFR_X1 port map( D => n8962, CK => CLK, RN => 
                           n12559, Q => n14343, QN => n10212);
   REGISTERS_reg_82_8_inst : DFFR_X1 port map( D => n8963, CK => CLK, RN => 
                           n12537, Q => n14344, QN => n10244);
   REGISTERS_reg_82_7_inst : DFFR_X1 port map( D => n8964, CK => CLK, RN => 
                           n12647, Q => n14345, QN => n10276);
   REGISTERS_reg_82_6_inst : DFFR_X1 port map( D => n8965, CK => CLK, RN => 
                           n12603, Q => n14346, QN => n10311);
   REGISTERS_reg_82_5_inst : DFFR_X1 port map( D => n8966, CK => CLK, RN => 
                           n12490, Q => n14347, QN => n10343);
   REGISTERS_reg_82_4_inst : DFFR_X1 port map( D => n8967, CK => CLK, RN => 
                           n12497, Q => n14348, QN => n10375);
   REGISTERS_reg_82_3_inst : DFFR_X1 port map( D => n8968, CK => CLK, RN => 
                           n12581, Q => n14349, QN => n10410);
   REGISTERS_reg_82_2_inst : DFFR_X1 port map( D => n8969, CK => CLK, RN => 
                           n12512, Q => n14350, QN => n10442);
   REGISTERS_reg_82_1_inst : DFFR_X1 port map( D => n8970, CK => CLK, RN => 
                           n12439, Q => n14351, QN => n10474);
   REGISTERS_reg_82_0_inst : DFFR_X1 port map( D => n8971, CK => CLK, RN => 
                           n12654, Q => n14352, QN => n10506);
   REGISTERS_reg_81_31_inst : DFFR_X1 port map( D => n8908, CK => CLK, RN => 
                           n12662, Q => n14289, QN => n5709);
   REGISTERS_reg_81_30_inst : DFFR_X1 port map( D => n8909, CK => CLK, RN => 
                           n12625, Q => n14290, QN => n5741);
   REGISTERS_reg_81_29_inst : DFFR_X1 port map( D => n8910, CK => CLK, RN => 
                           n12610, Q => n14291, QN => n5773);
   REGISTERS_reg_81_28_inst : DFFR_X1 port map( D => n8911, CK => CLK, RN => 
                           n12618, Q => n14292, QN => n5805);
   REGISTERS_reg_81_27_inst : DFFR_X1 port map( D => n8912, CK => CLK, RN => 
                           n12588, Q => n14293, QN => n5837);
   REGISTERS_reg_81_26_inst : DFFR_X1 port map( D => n8913, CK => CLK, RN => 
                           n12566, Q => n14294, QN => n5869);
   REGISTERS_reg_81_25_inst : DFFR_X1 port map( D => n8914, CK => CLK, RN => 
                           n12544, Q => n14295, QN => n5901);
   REGISTERS_reg_81_24_inst : DFFR_X1 port map( D => n8915, CK => CLK, RN => 
                           n12452, Q => n14296, QN => n5933);
   REGISTERS_reg_81_23_inst : DFFR_X1 port map( D => n8916, CK => CLK, RN => 
                           n12632, Q => n14297, QN => n5997);
   REGISTERS_reg_81_22_inst : DFFR_X1 port map( D => n8917, CK => CLK, RN => 
                           n12522, Q => n14298, QN => n6314);
   REGISTERS_reg_81_21_inst : DFFR_X1 port map( D => n8918, CK => CLK, RN => 
                           n12530, Q => n14299, QN => n9164);
   REGISTERS_reg_81_20_inst : DFFR_X1 port map( D => n8919, CK => CLK, RN => 
                           n12504, Q => n14300, QN => n9196);
   REGISTERS_reg_81_19_inst : DFFR_X1 port map( D => n8920, CK => CLK, RN => 
                           n12596, Q => n14301, QN => n9260);
   REGISTERS_reg_81_18_inst : DFFR_X1 port map( D => n8921, CK => CLK, RN => 
                           n12447, Q => n14302, QN => n9594);
   REGISTERS_reg_81_17_inst : DFFR_X1 port map( D => n8922, CK => CLK, RN => 
                           n12454, Q => n14303, QN => n9626);
   REGISTERS_reg_81_16_inst : DFFR_X1 port map( D => n8923, CK => CLK, RN => 
                           n12460, Q => n14304, QN => n9658);
   REGISTERS_reg_81_15_inst : DFFR_X1 port map( D => n8924, CK => CLK, RN => 
                           n12640, Q => n14305, QN => n10020);
   REGISTERS_reg_81_14_inst : DFFR_X1 port map( D => n8925, CK => CLK, RN => 
                           n12468, Q => n14306, QN => n10052);
   REGISTERS_reg_81_13_inst : DFFR_X1 port map( D => n8926, CK => CLK, RN => 
                           n12475, Q => n14307, QN => n10084);
   REGISTERS_reg_81_12_inst : DFFR_X1 port map( D => n8927, CK => CLK, RN => 
                           n12482, Q => n14308, QN => n10116);
   REGISTERS_reg_81_11_inst : DFFR_X1 port map( D => n8928, CK => CLK, RN => 
                           n12574, Q => n14309, QN => n10148);
   REGISTERS_reg_81_10_inst : DFFR_X1 port map( D => n8929, CK => CLK, RN => 
                           n12552, Q => n14310, QN => n10180);
   REGISTERS_reg_81_9_inst : DFFR_X1 port map( D => n8930, CK => CLK, RN => 
                           n12559, Q => n14311, QN => n10214);
   REGISTERS_reg_81_8_inst : DFFR_X1 port map( D => n8931, CK => CLK, RN => 
                           n12537, Q => n14312, QN => n10246);
   REGISTERS_reg_81_7_inst : DFFR_X1 port map( D => n8932, CK => CLK, RN => 
                           n12647, Q => n14313, QN => n10278);
   REGISTERS_reg_81_6_inst : DFFR_X1 port map( D => n8933, CK => CLK, RN => 
                           n12603, Q => n14314, QN => n10313);
   REGISTERS_reg_81_5_inst : DFFR_X1 port map( D => n8934, CK => CLK, RN => 
                           n12490, Q => n14315, QN => n10345);
   REGISTERS_reg_81_4_inst : DFFR_X1 port map( D => n8935, CK => CLK, RN => 
                           n12497, Q => n14316, QN => n10377);
   REGISTERS_reg_81_3_inst : DFFR_X1 port map( D => n8936, CK => CLK, RN => 
                           n12581, Q => n14317, QN => n10412);
   REGISTERS_reg_81_2_inst : DFFR_X1 port map( D => n8937, CK => CLK, RN => 
                           n12512, Q => n14318, QN => n10444);
   REGISTERS_reg_81_1_inst : DFFR_X1 port map( D => n8938, CK => CLK, RN => 
                           n12439, Q => n14319, QN => n10476);
   REGISTERS_reg_81_0_inst : DFFR_X1 port map( D => n8939, CK => CLK, RN => 
                           n12654, Q => n14320, QN => n10508);
   REGISTERS_reg_77_31_inst : DFFR_X1 port map( D => n8780, CK => CLK, RN => 
                           n12661, Q => n14257, QN => n5713);
   REGISTERS_reg_77_30_inst : DFFR_X1 port map( D => n8781, CK => CLK, RN => 
                           n12625, Q => n14258, QN => n5745);
   REGISTERS_reg_77_29_inst : DFFR_X1 port map( D => n8782, CK => CLK, RN => 
                           n12610, Q => n14259, QN => n5777);
   REGISTERS_reg_77_28_inst : DFFR_X1 port map( D => n8783, CK => CLK, RN => 
                           n12617, Q => n14260, QN => n5809);
   REGISTERS_reg_77_27_inst : DFFR_X1 port map( D => n8784, CK => CLK, RN => 
                           n12588, Q => n14261, QN => n5841);
   REGISTERS_reg_77_26_inst : DFFR_X1 port map( D => n8785, CK => CLK, RN => 
                           n12566, Q => n14262, QN => n5873);
   REGISTERS_reg_77_25_inst : DFFR_X1 port map( D => n8786, CK => CLK, RN => 
                           n12544, Q => n14263, QN => n5905);
   REGISTERS_reg_77_24_inst : DFFR_X1 port map( D => n8787, CK => CLK, RN => 
                           n12451, Q => n14264, QN => n5937);
   REGISTERS_reg_77_23_inst : DFFR_X1 port map( D => n8788, CK => CLK, RN => 
                           n12632, Q => n14265, QN => n6001);
   REGISTERS_reg_77_22_inst : DFFR_X1 port map( D => n8789, CK => CLK, RN => 
                           n12522, Q => n14266, QN => n9136);
   REGISTERS_reg_77_21_inst : DFFR_X1 port map( D => n8790, CK => CLK, RN => 
                           n12529, Q => n14267, QN => n9168);
   REGISTERS_reg_77_20_inst : DFFR_X1 port map( D => n8791, CK => CLK, RN => 
                           n12504, Q => n14268, QN => n9200);
   REGISTERS_reg_77_19_inst : DFFR_X1 port map( D => n8792, CK => CLK, RN => 
                           n12595, Q => n14269, QN => n9264);
   REGISTERS_reg_77_18_inst : DFFR_X1 port map( D => n8793, CK => CLK, RN => 
                           n12446, Q => n14270, QN => n9598);
   REGISTERS_reg_77_17_inst : DFFR_X1 port map( D => n8794, CK => CLK, RN => 
                           n12454, Q => n14271, QN => n9630);
   REGISTERS_reg_77_16_inst : DFFR_X1 port map( D => n8795, CK => CLK, RN => 
                           n12460, Q => n14272, QN => n9662);
   REGISTERS_reg_77_15_inst : DFFR_X1 port map( D => n8796, CK => CLK, RN => 
                           n12639, Q => n14273, QN => n10024);
   REGISTERS_reg_77_14_inst : DFFR_X1 port map( D => n8797, CK => CLK, RN => 
                           n12467, Q => n14274, QN => n10056);
   REGISTERS_reg_77_13_inst : DFFR_X1 port map( D => n8798, CK => CLK, RN => 
                           n12475, Q => n14275, QN => n10088);
   REGISTERS_reg_77_12_inst : DFFR_X1 port map( D => n8799, CK => CLK, RN => 
                           n12482, Q => n14276, QN => n10120);
   REGISTERS_reg_77_11_inst : DFFR_X1 port map( D => n8800, CK => CLK, RN => 
                           n12573, Q => n14277, QN => n10152);
   REGISTERS_reg_77_10_inst : DFFR_X1 port map( D => n8801, CK => CLK, RN => 
                           n12551, Q => n14278, QN => n10184);
   REGISTERS_reg_77_9_inst : DFFR_X1 port map( D => n8802, CK => CLK, RN => 
                           n12559, Q => n14279, QN => n10218);
   REGISTERS_reg_77_8_inst : DFFR_X1 port map( D => n8803, CK => CLK, RN => 
                           n12537, Q => n14280, QN => n10250);
   REGISTERS_reg_77_7_inst : DFFR_X1 port map( D => n8804, CK => CLK, RN => 
                           n12647, Q => n14281, QN => n10282);
   REGISTERS_reg_77_6_inst : DFFR_X1 port map( D => n8805, CK => CLK, RN => 
                           n12603, Q => n14282, QN => n10317);
   REGISTERS_reg_77_5_inst : DFFR_X1 port map( D => n8806, CK => CLK, RN => 
                           n12489, Q => n14283, QN => n10349);
   REGISTERS_reg_77_4_inst : DFFR_X1 port map( D => n8807, CK => CLK, RN => 
                           n12497, Q => n14284, QN => n10381);
   REGISTERS_reg_77_3_inst : DFFR_X1 port map( D => n8808, CK => CLK, RN => 
                           n12581, Q => n14285, QN => n10416);
   REGISTERS_reg_77_2_inst : DFFR_X1 port map( D => n8809, CK => CLK, RN => 
                           n12511, Q => n14286, QN => n10448);
   REGISTERS_reg_77_1_inst : DFFR_X1 port map( D => n8810, CK => CLK, RN => 
                           n12439, Q => n14287, QN => n10480);
   REGISTERS_reg_77_0_inst : DFFR_X1 port map( D => n8811, CK => CLK, RN => 
                           n12654, Q => n14288, QN => n10512);
   REGISTERS_reg_53_16_inst : DFFR_X1 port map( D => n8027, CK => CLK, RN => 
                           n12458, Q => n13795, QN => n929);
   REGISTERS_reg_53_15_inst : DFFR_X1 port map( D => n8028, CK => CLK, RN => 
                           n12637, Q => n13796, QN => n933);
   REGISTERS_reg_53_14_inst : DFFR_X1 port map( D => n8029, CK => CLK, RN => 
                           n12465, Q => n13797, QN => n937);
   REGISTERS_reg_53_13_inst : DFFR_X1 port map( D => n8030, CK => CLK, RN => 
                           n12473, Q => n13798, QN => n941);
   REGISTERS_reg_53_12_inst : DFFR_X1 port map( D => n8031, CK => CLK, RN => 
                           n12480, Q => n13799, QN => n945);
   REGISTERS_reg_53_11_inst : DFFR_X1 port map( D => n8032, CK => CLK, RN => 
                           n12571, Q => n13800, QN => n949);
   REGISTERS_reg_53_10_inst : DFFR_X1 port map( D => n8033, CK => CLK, RN => 
                           n12549, Q => n13801, QN => n953);
   REGISTERS_reg_53_9_inst : DFFR_X1 port map( D => n8034, CK => CLK, RN => 
                           n12557, Q => n13802, QN => n957);
   REGISTERS_reg_53_8_inst : DFFR_X1 port map( D => n8035, CK => CLK, RN => 
                           n12535, Q => n13803, QN => n961);
   REGISTERS_reg_53_7_inst : DFFR_X1 port map( D => n8036, CK => CLK, RN => 
                           n12645, Q => n13804, QN => n965);
   REGISTERS_reg_53_6_inst : DFFR_X1 port map( D => n8037, CK => CLK, RN => 
                           n12601, Q => n13805, QN => n969);
   REGISTERS_reg_53_5_inst : DFFR_X1 port map( D => n8038, CK => CLK, RN => 
                           n12487, Q => n13806, QN => n973);
   REGISTERS_reg_53_4_inst : DFFR_X1 port map( D => n8039, CK => CLK, RN => 
                           n12495, Q => n13807, QN => n977);
   REGISTERS_reg_53_3_inst : DFFR_X1 port map( D => n8040, CK => CLK, RN => 
                           n12579, Q => n13808, QN => n981);
   REGISTERS_reg_53_2_inst : DFFR_X1 port map( D => n8041, CK => CLK, RN => 
                           n12509, Q => n13809, QN => n985);
   REGISTERS_reg_53_1_inst : DFFR_X1 port map( D => n8042, CK => CLK, RN => 
                           n12437, Q => n13810, QN => n989);
   REGISTERS_reg_53_0_inst : DFFR_X1 port map( D => n8043, CK => CLK, RN => 
                           n12652, Q => n13811, QN => n993);
   REGISTERS_reg_52_31_inst : DFFR_X1 port map( D => n7980, CK => CLK, RN => 
                           n12659, Q => n13748, QN => n999);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n7334, CK => CLK, RN => 
                           n12485, Q => n13358, QN => n974);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n7335, CK => CLK, RN => 
                           n12493, Q => n13359, QN => n978);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n7336, CK => CLK, RN => 
                           n12577, Q => n13360, QN => n982);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n7337, CK => CLK, RN => 
                           n12507, Q => n13361, QN => n986);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n7338, CK => CLK, RN => 
                           n12435, Q => n13362, QN => n990);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n7339, CK => CLK, RN => 
                           n12650, Q => n13363, QN => n994);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n7020, CK => CLK, RN => 
                           n12657, Q => n13044, QN => n1868);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n7021, CK => CLK, RN => 
                           n12620, Q => n13045, QN => n1880);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n7022, CK => CLK, RN => 
                           n12605, Q => n13046, QN => n1892);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n7023, CK => CLK, RN => 
                           n12613, Q => n13047, QN => n1904);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n7024, CK => CLK, RN => 
                           n12583, Q => n13048, QN => n1916);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n7025, CK => CLK, RN => 
                           n12561, Q => n13049, QN => n1928);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n7026, CK => CLK, RN => 
                           n12539, Q => n13050, QN => n1940);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n7027, CK => CLK, RN => 
                           n12514, Q => n13051, QN => n1952);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n7028, CK => CLK, RN => 
                           n12627, Q => n13052, QN => n1964);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n7029, CK => CLK, RN => 
                           n12517, Q => n13053, QN => n1976);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n7030, CK => CLK, RN => 
                           n12525, Q => n13054, QN => n1988);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n7031, CK => CLK, RN => 
                           n12499, Q => n13055, QN => n2000);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n7032, CK => CLK, RN => 
                           n12591, Q => n13056, QN => n2012);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n7033, CK => CLK, RN => 
                           n12442, Q => n13057, QN => n2024);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n7034, CK => CLK, RN => 
                           n12449, Q => n13058, QN => n2036);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n7035, CK => CLK, RN => 
                           n12455, Q => n13059, QN => n2048);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n6988, CK => CLK, RN => 
                           n12657, Q => n13012, QN => n770);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n6989, CK => CLK, RN => 
                           n12620, Q => n13013, QN => n771);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n6990, CK => CLK, RN => 
                           n12605, Q => n13014, QN => n772);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n6991, CK => CLK, RN => 
                           n12613, Q => n13015, QN => n773);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n6992, CK => CLK, RN => 
                           n12583, Q => n13016, QN => n774);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n6993, CK => CLK, RN => 
                           n12561, Q => n13017, QN => n775);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n6994, CK => CLK, RN => 
                           n12539, Q => n13018, QN => n776);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n6995, CK => CLK, RN => 
                           n12514, Q => n13019, QN => n777);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n6996, CK => CLK, RN => 
                           n12627, Q => n13020, QN => n778);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n6997, CK => CLK, RN => 
                           n12517, Q => n13021, QN => n779);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n6998, CK => CLK, RN => 
                           n12525, Q => n13022, QN => n780);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n6999, CK => CLK, RN => 
                           n12499, Q => n13023, QN => n781);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n7000, CK => CLK, RN => 
                           n12591, Q => n13024, QN => n782);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n7001, CK => CLK, RN => 
                           n12442, Q => n13025, QN => n783);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n7002, CK => CLK, RN => 
                           n12449, Q => n13026, QN => n784);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n7003, CK => CLK, RN => 
                           n12455, Q => n13027, QN => n785);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n7004, CK => CLK, RN => 
                           n12635, Q => n13028, QN => n786);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n7005, CK => CLK, RN => 
                           n12463, Q => n13029, QN => n787);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n7006, CK => CLK, RN => 
                           n12470, Q => n13030, QN => n788);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n7007, CK => CLK, RN => 
                           n12477, Q => n13031, QN => n789);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n7008, CK => CLK, RN => 
                           n12569, Q => n13032, QN => n790);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n7009, CK => CLK, RN => 
                           n12547, Q => n13033, QN => n791);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n7010, CK => CLK, RN => 
                           n12554, Q => n13034, QN => n792);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n7011, CK => CLK, RN => 
                           n12532, Q => n13035, QN => n793);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n7012, CK => CLK, RN => 
                           n12642, Q => n13036, QN => n794);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n7013, CK => CLK, RN => 
                           n12598, Q => n13037, QN => n795);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n7014, CK => CLK, RN => 
                           n12485, Q => n13038, QN => n796);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n7015, CK => CLK, RN => 
                           n12492, Q => n13039, QN => n797);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n7016, CK => CLK, RN => 
                           n12576, Q => n13040, QN => n798);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n7017, CK => CLK, RN => 
                           n12507, Q => n13041, QN => n799);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n7018, CK => CLK, RN => 
                           n12434, Q => n13042, QN => n800);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n7019, CK => CLK, RN => 
                           n12649, Q => n13043, QN => n801);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n6956, CK => CLK, RN => 
                           n12657, Q => n12980, QN => n5738);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n6957, CK => CLK, RN => 
                           n12620, Q => n12981, QN => n5770);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n6958, CK => CLK, RN => 
                           n12605, Q => n12982, QN => n5802);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n6959, CK => CLK, RN => 
                           n12613, Q => n12983, QN => n5834);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n6960, CK => CLK, RN => 
                           n12583, Q => n12984, QN => n5866);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n6961, CK => CLK, RN => 
                           n12561, Q => n12985, QN => n5898);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n6962, CK => CLK, RN => 
                           n12539, Q => n12986, QN => n5930);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n6963, CK => CLK, RN => 
                           n12514, Q => n12987, QN => n5994);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n6964, CK => CLK, RN => 
                           n12627, Q => n12988, QN => n6311);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n6965, CK => CLK, RN => 
                           n12517, Q => n12989, QN => n9161);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n6966, CK => CLK, RN => 
                           n12525, Q => n12990, QN => n9193);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n6967, CK => CLK, RN => 
                           n12499, Q => n12991, QN => n9257);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n6968, CK => CLK, RN => 
                           n12591, Q => n12992, QN => n9591);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n6969, CK => CLK, RN => 
                           n12442, Q => n12993, QN => n9623);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n6970, CK => CLK, RN => 
                           n12449, Q => n12994, QN => n9655);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n6971, CK => CLK, RN => 
                           n12455, Q => n12995, QN => n10017);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n6972, CK => CLK, RN => 
                           n12635, Q => n12996, QN => n10049);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n6973, CK => CLK, RN => 
                           n12463, Q => n12997, QN => n10081);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n6974, CK => CLK, RN => 
                           n12470, Q => n12998, QN => n10113);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n6975, CK => CLK, RN => 
                           n12477, Q => n12999, QN => n10145);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n6976, CK => CLK, RN => 
                           n12569, Q => n13000, QN => n10177);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n6977, CK => CLK, RN => 
                           n12547, Q => n13001, QN => n10211);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n6978, CK => CLK, RN => 
                           n12554, Q => n13002, QN => n10243);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n6979, CK => CLK, RN => 
                           n12532, Q => n13003, QN => n10275);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n6980, CK => CLK, RN => 
                           n12642, Q => n13004, QN => n10310);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n6981, CK => CLK, RN => 
                           n12598, Q => n13005, QN => n10342);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n6982, CK => CLK, RN => 
                           n12485, Q => n13006, QN => n10374);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n6983, CK => CLK, RN => 
                           n12492, Q => n13007, QN => n10409);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n6984, CK => CLK, RN => 
                           n12576, Q => n13008, QN => n10441);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n6985, CK => CLK, RN => 
                           n12507, Q => n13009, QN => n10473);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n6986, CK => CLK, RN => 
                           n12434, Q => n13010, QN => n10505);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n6987, CK => CLK, RN => 
                           n12649, Q => n13011, QN => n10537);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n6924, CK => CLK, RN => 
                           n12656, Q => n12948, QN => n706);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n6925, CK => CLK, RN => 
                           n12620, Q => n12949, QN => n707);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n6926, CK => CLK, RN => 
                           n12605, Q => n12950, QN => n708);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n6927, CK => CLK, RN => 
                           n12612, Q => n12951, QN => n709);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n6928, CK => CLK, RN => 
                           n12583, Q => n12952, QN => n710);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n6929, CK => CLK, RN => 
                           n12561, Q => n12953, QN => n711);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n6930, CK => CLK, RN => 
                           n12539, Q => n12954, QN => n712);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n6931, CK => CLK, RN => 
                           n12514, Q => n12955, QN => n713);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n6932, CK => CLK, RN => 
                           n12627, Q => n12956, QN => n714);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n6933, CK => CLK, RN => 
                           n12517, Q => n12957, QN => n715);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n6934, CK => CLK, RN => 
                           n12524, Q => n12958, QN => n716);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n6935, CK => CLK, RN => 
                           n12499, Q => n12959, QN => n717);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n6936, CK => CLK, RN => 
                           n12590, Q => n12960, QN => n718);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n6937, CK => CLK, RN => 
                           n12441, Q => n12961, QN => n719);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n6938, CK => CLK, RN => 
                           n12449, Q => n12962, QN => n720);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n6939, CK => CLK, RN => 
                           n12455, Q => n12963, QN => n721);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n6940, CK => CLK, RN => 
                           n12634, Q => n12964, QN => n722);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n6941, CK => CLK, RN => 
                           n12462, Q => n12965, QN => n723);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n6942, CK => CLK, RN => 
                           n12470, Q => n12966, QN => n724);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n6943, CK => CLK, RN => 
                           n12477, Q => n12967, QN => n725);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n6944, CK => CLK, RN => 
                           n12568, Q => n12968, QN => n726);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n6945, CK => CLK, RN => 
                           n12546, Q => n12969, QN => n727);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n6946, CK => CLK, RN => 
                           n12554, Q => n12970, QN => n728);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n6947, CK => CLK, RN => 
                           n12532, Q => n12971, QN => n729);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n6948, CK => CLK, RN => 
                           n12642, Q => n12972, QN => n730);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n6949, CK => CLK, RN => 
                           n12598, Q => n12973, QN => n731);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n6950, CK => CLK, RN => 
                           n12484, Q => n12974, QN => n732);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n6951, CK => CLK, RN => 
                           n12492, Q => n12975, QN => n733);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n6952, CK => CLK, RN => 
                           n12576, Q => n12976, QN => n734);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n6953, CK => CLK, RN => 
                           n12506, Q => n12977, QN => n735);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n6954, CK => CLK, RN => 
                           n12434, Q => n12978, QN => n736);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n6955, CK => CLK, RN => 
                           n12649, Q => n12979, QN => n737);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n6892, CK => CLK, RN => 
                           n12656, Q => n12916, QN => n5732);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n6893, CK => CLK, RN => 
                           n12620, Q => n12917, QN => n5764);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n6894, CK => CLK, RN => 
                           n12605, Q => n12918, QN => n5796);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n6895, CK => CLK, RN => 
                           n12612, Q => n12919, QN => n5828);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n6896, CK => CLK, RN => 
                           n12583, Q => n12920, QN => n5860);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n6897, CK => CLK, RN => 
                           n12561, Q => n12921, QN => n5892);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n6898, CK => CLK, RN => 
                           n12539, Q => n12922, QN => n5924);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n6899, CK => CLK, RN => 
                           n12514, Q => n12923, QN => n5988);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n6900, CK => CLK, RN => 
                           n12627, Q => n12924, QN => n6305);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n6901, CK => CLK, RN => 
                           n12517, Q => n12925, QN => n9155);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n6902, CK => CLK, RN => 
                           n12524, Q => n12926, QN => n9187);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n6903, CK => CLK, RN => 
                           n12499, Q => n12927, QN => n9251);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n6904, CK => CLK, RN => 
                           n12590, Q => n12928, QN => n9585);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n6905, CK => CLK, RN => 
                           n12441, Q => n12929, QN => n9617);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n6906, CK => CLK, RN => 
                           n12449, Q => n12930, QN => n9649);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n6907, CK => CLK, RN => 
                           n12455, Q => n12931, QN => n10011);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n6908, CK => CLK, RN => 
                           n12634, Q => n12932, QN => n10043);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n6909, CK => CLK, RN => 
                           n12462, Q => n12933, QN => n10075);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n6910, CK => CLK, RN => 
                           n12470, Q => n12934, QN => n10107);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n6911, CK => CLK, RN => 
                           n12477, Q => n12935, QN => n10139);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n6912, CK => CLK, RN => 
                           n12568, Q => n12936, QN => n10171);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n6913, CK => CLK, RN => 
                           n12546, Q => n12937, QN => n10203);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n6914, CK => CLK, RN => 
                           n12554, Q => n12938, QN => n10237);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n6915, CK => CLK, RN => 
                           n12532, Q => n12939, QN => n10269);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n6916, CK => CLK, RN => 
                           n12642, Q => n12940, QN => n10304);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n6917, CK => CLK, RN => 
                           n12598, Q => n12941, QN => n10336);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n6918, CK => CLK, RN => 
                           n12484, Q => n12942, QN => n10368);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n6919, CK => CLK, RN => 
                           n12492, Q => n12943, QN => n10403);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n6920, CK => CLK, RN => 
                           n12576, Q => n12944, QN => n10435);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n6921, CK => CLK, RN => 
                           n12506, Q => n12945, QN => n10467);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n6922, CK => CLK, RN => 
                           n12434, Q => n12946, QN => n10499);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n6923, CK => CLK, RN => 
                           n12649, Q => n12947, QN => n10531);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n6860, CK => CLK, RN => 
                           n12656, Q => n12884, QN => n642);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n6861, CK => CLK, RN => 
                           n12620, Q => n12885, QN => n643);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n6862, CK => CLK, RN => 
                           n12605, Q => n12886, QN => n644);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n6863, CK => CLK, RN => 
                           n12612, Q => n12887, QN => n645);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n6864, CK => CLK, RN => 
                           n12583, Q => n12888, QN => n646);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n6865, CK => CLK, RN => 
                           n12561, Q => n12889, QN => n647);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n6866, CK => CLK, RN => 
                           n12539, Q => n12890, QN => n648);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n6867, CK => CLK, RN => 
                           n12514, Q => n12891, QN => n649);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n6868, CK => CLK, RN => 
                           n12627, Q => n12892, QN => n650);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n6869, CK => CLK, RN => 
                           n12517, Q => n12893, QN => n651);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n6870, CK => CLK, RN => 
                           n12524, Q => n12894, QN => n652);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n6871, CK => CLK, RN => 
                           n12499, Q => n12895, QN => n653);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n6872, CK => CLK, RN => 
                           n12590, Q => n12896, QN => n654);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n6873, CK => CLK, RN => 
                           n12441, Q => n12897, QN => n655);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n6874, CK => CLK, RN => 
                           n12449, Q => n12898, QN => n656);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n6875, CK => CLK, RN => 
                           n12455, Q => n12899, QN => n657);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n6876, CK => CLK, RN => 
                           n12634, Q => n12900, QN => n658);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n6877, CK => CLK, RN => 
                           n12462, Q => n12901, QN => n659);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n6878, CK => CLK, RN => 
                           n12470, Q => n12902, QN => n660);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n6879, CK => CLK, RN => 
                           n12477, Q => n12903, QN => n661);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n6880, CK => CLK, RN => 
                           n12568, Q => n12904, QN => n662);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n6881, CK => CLK, RN => 
                           n12546, Q => n12905, QN => n663);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n6882, CK => CLK, RN => 
                           n12554, Q => n12906, QN => n664);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n6883, CK => CLK, RN => 
                           n12532, Q => n12907, QN => n665);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n6884, CK => CLK, RN => 
                           n12642, Q => n12908, QN => n666);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n6885, CK => CLK, RN => 
                           n12598, Q => n12909, QN => n667);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n6886, CK => CLK, RN => 
                           n12484, Q => n12910, QN => n668);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n6887, CK => CLK, RN => 
                           n12492, Q => n12911, QN => n669);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n6888, CK => CLK, RN => 
                           n12576, Q => n12912, QN => n670);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n6889, CK => CLK, RN => 
                           n12506, Q => n12913, QN => n671);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n6890, CK => CLK, RN => 
                           n12434, Q => n12914, QN => n672);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n6891, CK => CLK, RN => 
                           n12649, Q => n12915, QN => n673);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n6828, CK => CLK, RN => 
                           n12656, Q => n12852, QN => n5731);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n6829, CK => CLK, RN => 
                           n12620, Q => n12853, QN => n5763);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n6830, CK => CLK, RN => 
                           n12605, Q => n12854, QN => n5795);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n6831, CK => CLK, RN => 
                           n12612, Q => n12855, QN => n5827);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n6832, CK => CLK, RN => 
                           n12583, Q => n12856, QN => n5859);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n6833, CK => CLK, RN => 
                           n12561, Q => n12857, QN => n5891);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n6834, CK => CLK, RN => 
                           n12539, Q => n12858, QN => n5923);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n6835, CK => CLK, RN => 
                           n12514, Q => n12859, QN => n5987);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n6836, CK => CLK, RN => 
                           n12627, Q => n12860, QN => n6304);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n6837, CK => CLK, RN => 
                           n12517, Q => n12861, QN => n9154);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n6838, CK => CLK, RN => 
                           n12524, Q => n12862, QN => n9186);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n6839, CK => CLK, RN => 
                           n12499, Q => n12863, QN => n9250);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n6840, CK => CLK, RN => 
                           n12590, Q => n12864, QN => n9584);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n6841, CK => CLK, RN => 
                           n12441, Q => n12865, QN => n9616);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n6842, CK => CLK, RN => 
                           n12449, Q => n12866, QN => n9648);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n6843, CK => CLK, RN => 
                           n12455, Q => n12867, QN => n10010);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n6844, CK => CLK, RN => 
                           n12634, Q => n12868, QN => n10042);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n6845, CK => CLK, RN => 
                           n12462, Q => n12869, QN => n10074);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n6846, CK => CLK, RN => 
                           n12470, Q => n12870, QN => n10106);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n6847, CK => CLK, RN => 
                           n12477, Q => n12871, QN => n10138);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n6848, CK => CLK, RN => 
                           n12568, Q => n12872, QN => n10170);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n6849, CK => CLK, RN => 
                           n12546, Q => n12873, QN => n10202);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n6850, CK => CLK, RN => 
                           n12554, Q => n12874, QN => n10236);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n6851, CK => CLK, RN => 
                           n12532, Q => n12875, QN => n10268);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n6852, CK => CLK, RN => 
                           n12642, Q => n12876, QN => n10300);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n6853, CK => CLK, RN => 
                           n12598, Q => n12877, QN => n10335);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n6854, CK => CLK, RN => 
                           n12484, Q => n12878, QN => n10367);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n6855, CK => CLK, RN => 
                           n12492, Q => n12879, QN => n10402);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n6856, CK => CLK, RN => 
                           n12576, Q => n12880, QN => n10434);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n6857, CK => CLK, RN => 
                           n12506, Q => n12881, QN => n10466);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n6858, CK => CLK, RN => 
                           n12434, Q => n12882, QN => n10498);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n6859, CK => CLK, RN => 
                           n12649, Q => n12883, QN => n10530);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n6796, CK => CLK, RN => 
                           n12656, Q => n12820, QN => n5733);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n6797, CK => CLK, RN => 
                           n12619, Q => n12821, QN => n5765);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n6798, CK => CLK, RN => 
                           n12605, Q => n12822, QN => n5797);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n6799, CK => CLK, RN => 
                           n12612, Q => n12823, QN => n5829);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n6800, CK => CLK, RN => 
                           n12583, Q => n12824, QN => n5861);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n6801, CK => CLK, RN => 
                           n12561, Q => n12825, QN => n5893);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n6802, CK => CLK, RN => 
                           n12539, Q => n12826, QN => n5925);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n6803, CK => CLK, RN => 
                           n12513, Q => n12827, QN => n5989);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n6804, CK => CLK, RN => 
                           n12627, Q => n12828, QN => n6306);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n6805, CK => CLK, RN => 
                           n12517, Q => n12829, QN => n9156);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n6806, CK => CLK, RN => 
                           n12524, Q => n12830, QN => n9188);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n6807, CK => CLK, RN => 
                           n12499, Q => n12831, QN => n9252);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n6808, CK => CLK, RN => 
                           n12590, Q => n12832, QN => n9586);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n6809, CK => CLK, RN => 
                           n12441, Q => n12833, QN => n9618);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n6810, CK => CLK, RN => 
                           n12448, Q => n12834, QN => n9650);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n6811, CK => CLK, RN => 
                           n12455, Q => n12835, QN => n10012);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n6812, CK => CLK, RN => 
                           n12634, Q => n12836, QN => n10044);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n6813, CK => CLK, RN => 
                           n12462, Q => n12837, QN => n10076);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n6814, CK => CLK, RN => 
                           n12469, Q => n12838, QN => n10108);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n6815, CK => CLK, RN => 
                           n12477, Q => n12839, QN => n10140);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n6816, CK => CLK, RN => 
                           n12568, Q => n12840, QN => n10172);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n6817, CK => CLK, RN => 
                           n12546, Q => n12841, QN => n10204);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n6818, CK => CLK, RN => 
                           n12553, Q => n12842, QN => n10238);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n6819, CK => CLK, RN => 
                           n12531, Q => n12843, QN => n10270);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n6820, CK => CLK, RN => 
                           n12641, Q => n12844, QN => n10305);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n6821, CK => CLK, RN => 
                           n12597, Q => n12845, QN => n10337);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n6822, CK => CLK, RN => 
                           n12484, Q => n12846, QN => n10369);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n6823, CK => CLK, RN => 
                           n12491, Q => n12847, QN => n10404);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n6824, CK => CLK, RN => 
                           n12575, Q => n12848, QN => n10436);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n6825, CK => CLK, RN => 
                           n12506, Q => n12849, QN => n10468);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n6826, CK => CLK, RN => 
                           n12434, Q => n12850, QN => n10500);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n6827, CK => CLK, RN => 
                           n12649, Q => n12851, QN => n10532);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n6668, CK => CLK, RN => 
                           n12656, Q => n12788, QN => n5737);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n6669, CK => CLK, RN => 
                           n12619, Q => n12789, QN => n5769);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n6670, CK => CLK, RN => 
                           n12604, Q => n12790, QN => n5801);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n6671, CK => CLK, RN => 
                           n12612, Q => n12791, QN => n5833);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n6672, CK => CLK, RN => 
                           n12582, Q => n12792, QN => n5865);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n6673, CK => CLK, RN => 
                           n12560, Q => n12793, QN => n5897);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n6674, CK => CLK, RN => 
                           n12538, Q => n12794, QN => n5929);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n6675, CK => CLK, RN => 
                           n12513, Q => n12795, QN => n5993);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n6676, CK => CLK, RN => 
                           n12626, Q => n12796, QN => n6310);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n6677, CK => CLK, RN => 
                           n12469, Q => n12797, QN => n9160);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n6678, CK => CLK, RN => 
                           n12524, Q => n12798, QN => n9192);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n6679, CK => CLK, RN => 
                           n12498, Q => n12799, QN => n9256);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n6680, CK => CLK, RN => 
                           n12590, Q => n12800, QN => n9590);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n6681, CK => CLK, RN => 
                           n12441, Q => n12801, QN => n9622);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n6682, CK => CLK, RN => 
                           n12448, Q => n12802, QN => n9654);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n6683, CK => CLK, RN => 
                           n12489, Q => n12803, QN => n10016);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n6684, CK => CLK, RN => 
                           n12634, Q => n12804, QN => n10048);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n6685, CK => CLK, RN => 
                           n12462, Q => n12805, QN => n10080);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n6686, CK => CLK, RN => 
                           n12469, Q => n12806, QN => n10112);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n6687, CK => CLK, RN => 
                           n12476, Q => n12807, QN => n10144);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n6688, CK => CLK, RN => 
                           n12568, Q => n12808, QN => n10176);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n6689, CK => CLK, RN => 
                           n12546, Q => n12809, QN => n10210);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n6690, CK => CLK, RN => 
                           n12553, Q => n12810, QN => n10242);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n6691, CK => CLK, RN => 
                           n12531, Q => n12811, QN => n10274);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n6692, CK => CLK, RN => 
                           n12641, Q => n12812, QN => n10309);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n6693, CK => CLK, RN => 
                           n12597, Q => n12813, QN => n10341);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n6694, CK => CLK, RN => 
                           n12484, Q => n12814, QN => n10373);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n6695, CK => CLK, RN => 
                           n12491, Q => n12815, QN => n10408);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n6696, CK => CLK, RN => 
                           n12575, Q => n12816, QN => n10440);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n6697, CK => CLK, RN => 
                           n12506, Q => n12817, QN => n10472);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n6698, CK => CLK, RN => 
                           n12433, Q => n12818, QN => n10504);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n6699, CK => CLK, RN => 
                           n12648, Q => n12819, QN => n10536);
   REGISTERS_reg_80_31_inst : DFFR_X1 port map( D => n8876, CK => CLK, RN => 
                           n12662, Q => n_2941, QN => n5711);
   REGISTERS_reg_80_30_inst : DFFR_X1 port map( D => n8877, CK => CLK, RN => 
                           n12625, Q => n_2942, QN => n5743);
   REGISTERS_reg_80_29_inst : DFFR_X1 port map( D => n8878, CK => CLK, RN => 
                           n12610, Q => n_2943, QN => n5775);
   REGISTERS_reg_80_28_inst : DFFR_X1 port map( D => n8879, CK => CLK, RN => 
                           n12618, Q => n_2944, QN => n5807);
   REGISTERS_reg_80_27_inst : DFFR_X1 port map( D => n8880, CK => CLK, RN => 
                           n12588, Q => n_2945, QN => n5839);
   REGISTERS_reg_80_26_inst : DFFR_X1 port map( D => n8881, CK => CLK, RN => 
                           n12566, Q => n_2946, QN => n5871);
   REGISTERS_reg_80_25_inst : DFFR_X1 port map( D => n8882, CK => CLK, RN => 
                           n12544, Q => n_2947, QN => n5903);
   REGISTERS_reg_80_24_inst : DFFR_X1 port map( D => n8883, CK => CLK, RN => 
                           n12450, Q => n_2948, QN => n5935);
   REGISTERS_reg_80_23_inst : DFFR_X1 port map( D => n8884, CK => CLK, RN => 
                           n12632, Q => n_2949, QN => n5999);
   REGISTERS_reg_80_22_inst : DFFR_X1 port map( D => n8885, CK => CLK, RN => 
                           n12522, Q => n_2950, QN => n9134);
   REGISTERS_reg_80_21_inst : DFFR_X1 port map( D => n8886, CK => CLK, RN => 
                           n12530, Q => n_2951, QN => n9166);
   REGISTERS_reg_80_20_inst : DFFR_X1 port map( D => n8887, CK => CLK, RN => 
                           n12504, Q => n_2952, QN => n9198);
   REGISTERS_reg_80_19_inst : DFFR_X1 port map( D => n8888, CK => CLK, RN => 
                           n12596, Q => n_2953, QN => n9262);
   REGISTERS_reg_80_18_inst : DFFR_X1 port map( D => n8889, CK => CLK, RN => 
                           n12447, Q => n_2954, QN => n9596);
   REGISTERS_reg_80_17_inst : DFFR_X1 port map( D => n8890, CK => CLK, RN => 
                           n12454, Q => n_2955, QN => n9628);
   REGISTERS_reg_80_16_inst : DFFR_X1 port map( D => n8891, CK => CLK, RN => 
                           n12460, Q => n_2956, QN => n9660);
   REGISTERS_reg_80_15_inst : DFFR_X1 port map( D => n8892, CK => CLK, RN => 
                           n12640, Q => n_2957, QN => n10022);
   REGISTERS_reg_80_14_inst : DFFR_X1 port map( D => n8893, CK => CLK, RN => 
                           n12468, Q => n_2958, QN => n10054);
   REGISTERS_reg_80_13_inst : DFFR_X1 port map( D => n8894, CK => CLK, RN => 
                           n12475, Q => n_2959, QN => n10086);
   REGISTERS_reg_80_12_inst : DFFR_X1 port map( D => n8895, CK => CLK, RN => 
                           n12482, Q => n_2960, QN => n10118);
   REGISTERS_reg_80_11_inst : DFFR_X1 port map( D => n8896, CK => CLK, RN => 
                           n12574, Q => n_2961, QN => n10150);
   REGISTERS_reg_80_10_inst : DFFR_X1 port map( D => n8897, CK => CLK, RN => 
                           n12552, Q => n_2962, QN => n10182);
   REGISTERS_reg_80_9_inst : DFFR_X1 port map( D => n8898, CK => CLK, RN => 
                           n12559, Q => n_2963, QN => n10216);
   REGISTERS_reg_80_8_inst : DFFR_X1 port map( D => n8899, CK => CLK, RN => 
                           n12537, Q => n_2964, QN => n10248);
   REGISTERS_reg_80_7_inst : DFFR_X1 port map( D => n8900, CK => CLK, RN => 
                           n12647, Q => n_2965, QN => n10280);
   U3 : XNOR2_X1 port map( A => U3_U98_Z_6, B => r480_n4, ZN => N8437);
   U4 : XNOR2_X1 port map( A => U3_U99_Z_6, B => r486_n4, ZN => N8581);
   U5 : AND2_X1 port map( A1 => n2574, A2 => n2491, ZN => n10538);
   U6 : AND2_X1 port map( A1 => n2574, A2 => n2494, ZN => n10539);
   U7 : AND2_X1 port map( A1 => n2574, A2 => n2496, ZN => n10540);
   U8 : AND2_X1 port map( A1 => n2574, A2 => n2498, ZN => n10541);
   U9 : AND2_X1 port map( A1 => n2574, A2 => n2500, ZN => n10542);
   U10 : AND2_X1 port map( A1 => n2574, A2 => n2566, ZN => n10543);
   U11 : AND2_X1 port map( A1 => n2574, A2 => n2568, ZN => n10544);
   U12 : AND2_X1 port map( A1 => n2574, A2 => n2570, ZN => n10545);
   U13 : AND2_X1 port map( A1 => n2599, A2 => n2573, ZN => n10546);
   U14 : AND2_X1 port map( A1 => n2599, A2 => n2578, ZN => n10547);
   U15 : AND2_X1 port map( A1 => n2599, A2 => n2570, ZN => n10548);
   U16 : AND2_X1 port map( A1 => n2617, A2 => n2573, ZN => n10549);
   U17 : AND2_X1 port map( A1 => n2617, A2 => n2576, ZN => n10550);
   U18 : AND2_X1 port map( A1 => n2617, A2 => n2582, ZN => n10551);
   U19 : AND2_X1 port map( A1 => n2617, A2 => n2586, ZN => n10552);
   U20 : AND2_X1 port map( A1 => n2617, A2 => n2491, ZN => n10553);
   U21 : AND2_X1 port map( A1 => n2698, A2 => n2584, ZN => n10554);
   U22 : AND2_X1 port map( A1 => n2698, A2 => n2586, ZN => n10555);
   U23 : AND2_X1 port map( A1 => n2698, A2 => n2588, ZN => n10556);
   U24 : AND2_X1 port map( A1 => n2599, A2 => n2582, ZN => n10557);
   U25 : AND2_X1 port map( A1 => n2599, A2 => n2588, ZN => n10558);
   U26 : AND2_X1 port map( A1 => n2617, A2 => n2496, ZN => n10559);
   U27 : AND2_X1 port map( A1 => n2617, A2 => n2566, ZN => n10560);
   U28 : AND2_X1 port map( A1 => n2715, A2 => n2580, ZN => n10561);
   U29 : AND2_X1 port map( A1 => n2715, A2 => n2588, ZN => n10562);
   U30 : AND2_X1 port map( A1 => n2715, A2 => n2496, ZN => n10563);
   U31 : AND2_X1 port map( A1 => n2715, A2 => n2566, ZN => n10564);
   U32 : AND2_X1 port map( A1 => n2599, A2 => n2580, ZN => n10565);
   U33 : AND2_X1 port map( A1 => n2599, A2 => n2586, ZN => n10566);
   U34 : AND2_X1 port map( A1 => n2617, A2 => n2494, ZN => n10567);
   U35 : AND2_X1 port map( A1 => n2617, A2 => n2500, ZN => n10568);
   U36 : AND2_X1 port map( A1 => n2715, A2 => n2578, ZN => n10569);
   U37 : AND2_X1 port map( A1 => n2715, A2 => n2584, ZN => n10570);
   U38 : AND2_X1 port map( A1 => n2715, A2 => n2491, ZN => n10571);
   U39 : AND2_X1 port map( A1 => n2715, A2 => n2498, ZN => n10572);
   U40 : AND2_X1 port map( A1 => n2599, A2 => n2576, ZN => n10573);
   U41 : AND2_X1 port map( A1 => n2599, A2 => n2584, ZN => n10574);
   U42 : AND2_X1 port map( A1 => n2617, A2 => n2588, ZN => n10575);
   U43 : AND2_X1 port map( A1 => n2617, A2 => n2498, ZN => n10576);
   U44 : AND2_X1 port map( A1 => n2715, A2 => n2576, ZN => n10577);
   U45 : AND2_X1 port map( A1 => n2715, A2 => n2586, ZN => n10578);
   U46 : AND2_X1 port map( A1 => n2715, A2 => n2494, ZN => n10579);
   U47 : AND2_X1 port map( A1 => n2715, A2 => n2500, ZN => n10580);
   U48 : AND2_X1 port map( A1 => n2599, A2 => n2491, ZN => n10581);
   U49 : AND2_X1 port map( A1 => n2617, A2 => n2568, ZN => n10582);
   U50 : AND2_X1 port map( A1 => n2715, A2 => n2568, ZN => n10583);
   U51 : AND2_X1 port map( A1 => n2617, A2 => n2584, ZN => n10584);
   U52 : AND2_X1 port map( A1 => n2715, A2 => n2570, ZN => n10585);
   U53 : AND2_X1 port map( A1 => n2599, A2 => n2496, ZN => n10586);
   U54 : AND2_X1 port map( A1 => n2698, A2 => n2496, ZN => n10587);
   U55 : AND2_X1 port map( A1 => n2698, A2 => n2498, ZN => n10588);
   U56 : AND2_X1 port map( A1 => n2698, A2 => n2500, ZN => n10589);
   U57 : AND2_X1 port map( A1 => n2698, A2 => n2566, ZN => n10590);
   U58 : AND2_X1 port map( A1 => n2698, A2 => n2568, ZN => n10591);
   U59 : AND2_X1 port map( A1 => n2698, A2 => n2570, ZN => n10592);
   U60 : AND2_X1 port map( A1 => n2715, A2 => n2573, ZN => n10593);
   U61 : AND2_X1 port map( A1 => n2715, A2 => n2582, ZN => n10594);
   U62 : AND2_X1 port map( A1 => n2599, A2 => n2494, ZN => n10595);
   U63 : AND2_X1 port map( A1 => n2599, A2 => n2498, ZN => n10596);
   U64 : AND2_X1 port map( A1 => n2599, A2 => n2500, ZN => n10597);
   U65 : AND2_X1 port map( A1 => n2599, A2 => n2566, ZN => n10598);
   U66 : AND2_X1 port map( A1 => n2599, A2 => n2568, ZN => n10599);
   U67 : AND2_X1 port map( A1 => n2617, A2 => n2578, ZN => n10600);
   U68 : AND2_X1 port map( A1 => n2617, A2 => n2580, ZN => n10601);
   U69 : AND2_X1 port map( A1 => n2617, A2 => n2570, ZN => n10602);
   U70 : AND2_X1 port map( A1 => n2698, A2 => n2573, ZN => n10603);
   U71 : AND2_X1 port map( A1 => n2698, A2 => n2576, ZN => n10604);
   U72 : AND2_X1 port map( A1 => n2698, A2 => n2578, ZN => n10605);
   U73 : AND2_X1 port map( A1 => n2698, A2 => n2580, ZN => n10606);
   U74 : AND2_X1 port map( A1 => n2698, A2 => n2582, ZN => n10607);
   U75 : AND2_X1 port map( A1 => n2698, A2 => n2491, ZN => n10608);
   U76 : AND2_X1 port map( A1 => n2698, A2 => n2494, ZN => n10609);
   U77 : AND2_X1 port map( A1 => n2580, A2 => n2574, ZN => n10610);
   U78 : AND2_X1 port map( A1 => n2584, A2 => n2574, ZN => n10611);
   U79 : AND2_X1 port map( A1 => n2586, A2 => n2574, ZN => n10612);
   U80 : AND2_X1 port map( A1 => n2588, A2 => n2574, ZN => n10613);
   U81 : AND2_X1 port map( A1 => n2576, A2 => n2574, ZN => n10614);
   U82 : AND2_X1 port map( A1 => n2573, A2 => n2574, ZN => n10615);
   U83 : AND2_X1 port map( A1 => n2582, A2 => n2574, ZN => n10616);
   U84 : AND2_X1 port map( A1 => n2578, A2 => n2574, ZN => n10617);
   U85 : AND2_X1 port map( A1 => n2570, A2 => n2492, ZN => n10618);
   U86 : AND2_X1 port map( A1 => n2494, A2 => n2492, ZN => n10619);
   U87 : AND2_X1 port map( A1 => n2496, A2 => n2492, ZN => n10620);
   U88 : AND2_X1 port map( A1 => n2498, A2 => n2492, ZN => n10621);
   U89 : AND2_X1 port map( A1 => n2500, A2 => n2492, ZN => n10622);
   U90 : AND2_X1 port map( A1 => n2566, A2 => n2492, ZN => n10623);
   U91 : AND2_X1 port map( A1 => n2568, A2 => n2492, ZN => n10624);
   U92 : NOR2_X1 port map( A1 => n12770, A2 => N8435, ZN => n5675);
   U93 : NOR2_X1 port map( A1 => n12774, A2 => N8579, ZN => n4242);
   U94 : AND3_X1 port map( A1 => n2615, A2 => N2171, A3 => N2172, ZN => n2599);
   U95 : AND3_X1 port map( A1 => N2171, A2 => n12732, A3 => n2615, ZN => n2698)
                           ;
   U96 : INV_X1 port map( A => n12290, ZN => n12280);
   U97 : INV_X1 port map( A => n12290, ZN => n12279);
   U98 : INV_X1 port map( A => n12242, ZN => n12232);
   U99 : INV_X1 port map( A => n12242, ZN => n12231);
   U100 : INV_X1 port map( A => n11906, ZN => n11896);
   U101 : INV_X1 port map( A => n11906, ZN => n11895);
   U102 : INV_X1 port map( A => n11858, ZN => n11848);
   U103 : INV_X1 port map( A => n11858, ZN => n11847);
   U104 : INV_X1 port map( A => n11522, ZN => n11512);
   U105 : INV_X1 port map( A => n11522, ZN => n11511);
   U106 : INV_X1 port map( A => n11474, ZN => n11464);
   U107 : INV_X1 port map( A => n11474, ZN => n11463);
   U108 : INV_X1 port map( A => n12415, ZN => n12406);
   U109 : INV_X1 port map( A => n12415, ZN => n12405);
   U110 : INV_X1 port map( A => n12404, ZN => n12395);
   U111 : INV_X1 port map( A => n12404, ZN => n12394);
   U112 : INV_X1 port map( A => n12393, ZN => n12384);
   U113 : INV_X1 port map( A => n12393, ZN => n12383);
   U114 : INV_X1 port map( A => n12382, ZN => n12373);
   U115 : INV_X1 port map( A => n12382, ZN => n12372);
   U116 : INV_X1 port map( A => n12371, ZN => n12362);
   U117 : INV_X1 port map( A => n12371, ZN => n12361);
   U118 : INV_X1 port map( A => n12360, ZN => n12351);
   U119 : INV_X1 port map( A => n12360, ZN => n12350);
   U120 : INV_X1 port map( A => n12349, ZN => n12340);
   U121 : INV_X1 port map( A => n12349, ZN => n12339);
   U122 : INV_X1 port map( A => n12338, ZN => n12328);
   U123 : INV_X1 port map( A => n12338, ZN => n12327);
   U124 : INV_X1 port map( A => n12326, ZN => n12316);
   U125 : INV_X1 port map( A => n12326, ZN => n12315);
   U126 : INV_X1 port map( A => n12314, ZN => n12304);
   U127 : INV_X1 port map( A => n12314, ZN => n12303);
   U128 : INV_X1 port map( A => n12302, ZN => n12292);
   U129 : INV_X1 port map( A => n12302, ZN => n12291);
   U130 : INV_X1 port map( A => n12278, ZN => n12268);
   U131 : INV_X1 port map( A => n12278, ZN => n12267);
   U132 : INV_X1 port map( A => n12266, ZN => n12256);
   U133 : INV_X1 port map( A => n12266, ZN => n12255);
   U134 : INV_X1 port map( A => n12254, ZN => n12244);
   U135 : INV_X1 port map( A => n12254, ZN => n12243);
   U136 : INV_X1 port map( A => n12230, ZN => n12220);
   U137 : INV_X1 port map( A => n12230, ZN => n12219);
   U138 : INV_X1 port map( A => n12218, ZN => n12208);
   U139 : INV_X1 port map( A => n12218, ZN => n12207);
   U140 : INV_X1 port map( A => n12206, ZN => n12196);
   U141 : INV_X1 port map( A => n12206, ZN => n12195);
   U142 : INV_X1 port map( A => n12194, ZN => n12184);
   U143 : INV_X1 port map( A => n12194, ZN => n12183);
   U144 : INV_X1 port map( A => n12182, ZN => n12172);
   U145 : INV_X1 port map( A => n12182, ZN => n12171);
   U146 : INV_X1 port map( A => n12170, ZN => n12160);
   U147 : INV_X1 port map( A => n12170, ZN => n12159);
   U148 : INV_X1 port map( A => n12158, ZN => n12148);
   U149 : INV_X1 port map( A => n12158, ZN => n12147);
   U150 : INV_X1 port map( A => n12146, ZN => n12136);
   U151 : INV_X1 port map( A => n12146, ZN => n12135);
   U152 : INV_X1 port map( A => n12134, ZN => n12124);
   U153 : INV_X1 port map( A => n12134, ZN => n12123);
   U154 : INV_X1 port map( A => n12122, ZN => n12112);
   U155 : INV_X1 port map( A => n12122, ZN => n12111);
   U156 : INV_X1 port map( A => n12110, ZN => n12100);
   U157 : INV_X1 port map( A => n12110, ZN => n12099);
   U158 : INV_X1 port map( A => n12098, ZN => n12088);
   U159 : INV_X1 port map( A => n12098, ZN => n12087);
   U160 : INV_X1 port map( A => n12086, ZN => n12076);
   U161 : INV_X1 port map( A => n12086, ZN => n12075);
   U162 : INV_X1 port map( A => n12074, ZN => n12064);
   U163 : INV_X1 port map( A => n12074, ZN => n12063);
   U164 : INV_X1 port map( A => n12062, ZN => n12052);
   U165 : INV_X1 port map( A => n12062, ZN => n12051);
   U166 : INV_X1 port map( A => n12050, ZN => n12040);
   U167 : INV_X1 port map( A => n12050, ZN => n12039);
   U168 : INV_X1 port map( A => n12038, ZN => n12028);
   U169 : INV_X1 port map( A => n12038, ZN => n12027);
   U170 : INV_X1 port map( A => n12026, ZN => n12016);
   U171 : INV_X1 port map( A => n12026, ZN => n12015);
   U172 : INV_X1 port map( A => n12014, ZN => n12004);
   U173 : INV_X1 port map( A => n12014, ZN => n12003);
   U174 : INV_X1 port map( A => n12002, ZN => n11992);
   U175 : INV_X1 port map( A => n12002, ZN => n11991);
   U176 : INV_X1 port map( A => n11990, ZN => n11980);
   U177 : INV_X1 port map( A => n11990, ZN => n11979);
   U178 : INV_X1 port map( A => n11978, ZN => n11968);
   U179 : INV_X1 port map( A => n11978, ZN => n11967);
   U180 : INV_X1 port map( A => n11966, ZN => n11956);
   U181 : INV_X1 port map( A => n11966, ZN => n11955);
   U182 : INV_X1 port map( A => n11954, ZN => n11944);
   U183 : INV_X1 port map( A => n11954, ZN => n11943);
   U184 : INV_X1 port map( A => n11942, ZN => n11932);
   U185 : INV_X1 port map( A => n11942, ZN => n11931);
   U186 : INV_X1 port map( A => n11930, ZN => n11920);
   U187 : INV_X1 port map( A => n11930, ZN => n11919);
   U188 : INV_X1 port map( A => n11918, ZN => n11908);
   U189 : INV_X1 port map( A => n11918, ZN => n11907);
   U191 : INV_X1 port map( A => n11894, ZN => n11884);
   U192 : INV_X1 port map( A => n11894, ZN => n11883);
   U193 : INV_X1 port map( A => n11882, ZN => n11872);
   U194 : INV_X1 port map( A => n11882, ZN => n11871);
   U195 : INV_X1 port map( A => n11870, ZN => n11860);
   U196 : INV_X1 port map( A => n11870, ZN => n11859);
   U197 : INV_X1 port map( A => n11846, ZN => n11836);
   U198 : INV_X1 port map( A => n11846, ZN => n11835);
   U199 : INV_X1 port map( A => n11834, ZN => n11824);
   U200 : INV_X1 port map( A => n11834, ZN => n11823);
   U201 : INV_X1 port map( A => n11822, ZN => n11812);
   U202 : INV_X1 port map( A => n11822, ZN => n11811);
   U203 : INV_X1 port map( A => n11810, ZN => n11800);
   U204 : INV_X1 port map( A => n11810, ZN => n11799);
   U205 : INV_X1 port map( A => n11798, ZN => n11788);
   U206 : INV_X1 port map( A => n11798, ZN => n11787);
   U207 : INV_X1 port map( A => n11786, ZN => n11776);
   U208 : INV_X1 port map( A => n11786, ZN => n11775);
   U209 : INV_X1 port map( A => n11774, ZN => n11764);
   U210 : INV_X1 port map( A => n11774, ZN => n11763);
   U211 : INV_X1 port map( A => n11762, ZN => n11752);
   U212 : INV_X1 port map( A => n11762, ZN => n11751);
   U213 : INV_X1 port map( A => n11750, ZN => n11740);
   U214 : INV_X1 port map( A => n11750, ZN => n11739);
   U215 : INV_X1 port map( A => n11738, ZN => n11728);
   U216 : INV_X1 port map( A => n11738, ZN => n11727);
   U217 : INV_X1 port map( A => n11726, ZN => n11716);
   U218 : INV_X1 port map( A => n11726, ZN => n11715);
   U219 : INV_X1 port map( A => n11714, ZN => n11704);
   U220 : INV_X1 port map( A => n11714, ZN => n11703);
   U221 : INV_X1 port map( A => n11702, ZN => n11692);
   U222 : INV_X1 port map( A => n11702, ZN => n11691);
   U223 : INV_X1 port map( A => n11690, ZN => n11680);
   U225 : INV_X1 port map( A => n11690, ZN => n11679);
   U226 : INV_X1 port map( A => n11678, ZN => n11668);
   U227 : INV_X1 port map( A => n11678, ZN => n11667);
   U228 : INV_X1 port map( A => n11666, ZN => n11656);
   U229 : INV_X1 port map( A => n11666, ZN => n11655);
   U230 : INV_X1 port map( A => n11654, ZN => n11644);
   U231 : INV_X1 port map( A => n11654, ZN => n11643);
   U232 : INV_X1 port map( A => n11642, ZN => n11632);
   U233 : INV_X1 port map( A => n11642, ZN => n11631);
   U234 : INV_X1 port map( A => n11630, ZN => n11620);
   U235 : INV_X1 port map( A => n11630, ZN => n11619);
   U236 : INV_X1 port map( A => n11618, ZN => n11608);
   U237 : INV_X1 port map( A => n11618, ZN => n11607);
   U238 : INV_X1 port map( A => n11606, ZN => n11596);
   U239 : INV_X1 port map( A => n11606, ZN => n11595);
   U240 : INV_X1 port map( A => n11594, ZN => n11584);
   U241 : INV_X1 port map( A => n11594, ZN => n11583);
   U242 : INV_X1 port map( A => n11582, ZN => n11572);
   U243 : INV_X1 port map( A => n11582, ZN => n11571);
   U244 : INV_X1 port map( A => n11570, ZN => n11560);
   U245 : INV_X1 port map( A => n11570, ZN => n11559);
   U246 : INV_X1 port map( A => n11558, ZN => n11548);
   U247 : INV_X1 port map( A => n11558, ZN => n11547);
   U248 : INV_X1 port map( A => n11546, ZN => n11536);
   U249 : INV_X1 port map( A => n11546, ZN => n11535);
   U250 : INV_X1 port map( A => n11534, ZN => n11524);
   U251 : INV_X1 port map( A => n11534, ZN => n11523);
   U252 : INV_X1 port map( A => n11510, ZN => n11500);
   U253 : INV_X1 port map( A => n11510, ZN => n11499);
   U254 : INV_X1 port map( A => n11498, ZN => n11488);
   U255 : INV_X1 port map( A => n11498, ZN => n11487);
   U256 : INV_X1 port map( A => n11486, ZN => n11476);
   U257 : INV_X1 port map( A => n11486, ZN => n11475);
   U258 : INV_X1 port map( A => n11462, ZN => n11452);
   U259 : INV_X1 port map( A => n11462, ZN => n11451);
   U260 : INV_X1 port map( A => n11450, ZN => n11440);
   U261 : INV_X1 port map( A => n11450, ZN => n11439);
   U262 : INV_X1 port map( A => n11438, ZN => n11428);
   U263 : INV_X1 port map( A => n11438, ZN => n11427);
   U264 : INV_X1 port map( A => n11426, ZN => n11416);
   U265 : INV_X1 port map( A => n11426, ZN => n11415);
   U266 : INV_X1 port map( A => n11414, ZN => n11404);
   U267 : INV_X1 port map( A => n11414, ZN => n11403);
   U268 : INV_X1 port map( A => n11402, ZN => n11392);
   U269 : INV_X1 port map( A => n11402, ZN => n11391);
   U270 : INV_X1 port map( A => n11390, ZN => n11380);
   U271 : INV_X1 port map( A => n11390, ZN => n11379);
   U272 : BUF_X1 port map( A => n10594, Z => n11514);
   U273 : BUF_X1 port map( A => n10594, Z => n11515);
   U274 : BUF_X1 port map( A => n10594, Z => n11516);
   U275 : BUF_X1 port map( A => n10594, Z => n11517);
   U276 : BUF_X1 port map( A => n11522, Z => n11518);
   U277 : BUF_X1 port map( A => n11520, Z => n11519);
   U278 : BUF_X1 port map( A => n10594, Z => n11520);
   U279 : BUF_X1 port map( A => n11522, Z => n11521);
   U280 : BUF_X1 port map( A => n10571, Z => n11466);
   U281 : BUF_X1 port map( A => n10571, Z => n11467);
   U282 : BUF_X1 port map( A => n10571, Z => n11468);
   U283 : BUF_X1 port map( A => n10571, Z => n11469);
   U284 : BUF_X1 port map( A => n11474, Z => n11470);
   U285 : BUF_X1 port map( A => n11472, Z => n11471);
   U286 : BUF_X1 port map( A => n10571, Z => n11472);
   U287 : BUF_X1 port map( A => n11474, Z => n11473);
   U288 : BUF_X1 port map( A => n10616, Z => n12282);
   U289 : BUF_X1 port map( A => n10616, Z => n12283);
   U290 : BUF_X1 port map( A => n10616, Z => n12284);
   U291 : BUF_X1 port map( A => n10616, Z => n12285);
   U292 : BUF_X1 port map( A => n12290, Z => n12286);
   U293 : BUF_X1 port map( A => n12288, Z => n12287);
   U294 : BUF_X1 port map( A => n10616, Z => n12288);
   U295 : BUF_X1 port map( A => n12290, Z => n12289);
   U296 : BUF_X1 port map( A => n10538, Z => n12234);
   U297 : BUF_X1 port map( A => n10538, Z => n12235);
   U298 : BUF_X1 port map( A => n10538, Z => n12236);
   U299 : BUF_X1 port map( A => n10538, Z => n12237);
   U300 : BUF_X1 port map( A => n10538, Z => n12238);
   U301 : BUF_X1 port map( A => n10538, Z => n12239);
   U302 : BUF_X1 port map( A => n12234, Z => n12240);
   U303 : BUF_X1 port map( A => n12236, Z => n12241);
   U304 : BUF_X1 port map( A => n10551, Z => n11898);
   U305 : BUF_X1 port map( A => n10551, Z => n11899);
   U338 : BUF_X1 port map( A => n10551, Z => n11900);
   U339 : BUF_X1 port map( A => n10551, Z => n11901);
   U340 : BUF_X1 port map( A => n11906, Z => n11902);
   U341 : BUF_X1 port map( A => n11904, Z => n11903);
   U342 : BUF_X1 port map( A => n10551, Z => n11904);
   U343 : BUF_X1 port map( A => n11906, Z => n11905);
   U344 : BUF_X1 port map( A => n10553, Z => n11850);
   U345 : BUF_X1 port map( A => n10553, Z => n11851);
   U346 : BUF_X1 port map( A => n10553, Z => n11852);
   U347 : BUF_X1 port map( A => n10553, Z => n11853);
   U348 : BUF_X1 port map( A => n11858, Z => n11854);
   U349 : BUF_X1 port map( A => n11856, Z => n11855);
   U350 : BUF_X1 port map( A => n10553, Z => n11856);
   U351 : BUF_X1 port map( A => n11858, Z => n11857);
   U352 : BUF_X1 port map( A => n12237, Z => n12242);
   U353 : BUF_X1 port map( A => n10551, Z => n11906);
   U354 : BUF_X1 port map( A => n10553, Z => n11858);
   U355 : BUF_X1 port map( A => n10594, Z => n11522);
   U356 : BUF_X1 port map( A => n10571, Z => n11474);
   U357 : BUF_X1 port map( A => n10616, Z => n12290);
   U358 : INV_X1 port map( A => n12425, ZN => n12417);
   U359 : INV_X1 port map( A => n12425, ZN => n12416);
   U360 : BUF_X1 port map( A => n12714, Z => n12708);
   U361 : BUF_X1 port map( A => n12713, Z => n12711);
   U362 : BUF_X1 port map( A => n12722, Z => n12685);
   U363 : BUF_X1 port map( A => n12719, Z => n12693);
   U364 : BUF_X1 port map( A => n12723, Z => n12680);
   U365 : BUF_X1 port map( A => n12716, Z => n12703);
   U366 : BUF_X1 port map( A => n12723, Z => n12682);
   U367 : BUF_X1 port map( A => n12722, Z => n12683);
   U368 : BUF_X1 port map( A => n12717, Z => n12700);
   U369 : BUF_X1 port map( A => n12719, Z => n12694);
   U370 : BUF_X1 port map( A => n12715, Z => n12706);
   U371 : BUF_X1 port map( A => n12714, Z => n12707);
   U372 : BUF_X1 port map( A => n12715, Z => n12704);
   U373 : BUF_X1 port map( A => n12722, Z => n12684);
   U374 : BUF_X1 port map( A => n12721, Z => n12686);
   U375 : BUF_X1 port map( A => n12721, Z => n12687);
   U376 : BUF_X1 port map( A => n12718, Z => n12695);
   U377 : BUF_X1 port map( A => n12721, Z => n12688);
   U378 : BUF_X1 port map( A => n12720, Z => n12689);
   U379 : BUF_X1 port map( A => n12720, Z => n12690);
   U380 : BUF_X1 port map( A => n12716, Z => n12701);
   U381 : BUF_X1 port map( A => n12723, Z => n12681);
   U382 : BUF_X1 port map( A => n12713, Z => n12710);
   U383 : BUF_X1 port map( A => n12718, Z => n12696);
   U384 : BUF_X1 port map( A => n12724, Z => n12679);
   U385 : BUF_X1 port map( A => n12714, Z => n12709);
   U386 : BUF_X1 port map( A => n12715, Z => n12705);
   U387 : BUF_X1 port map( A => n12716, Z => n12702);
   U388 : BUF_X1 port map( A => n12717, Z => n12698);
   U389 : BUF_X1 port map( A => n12717, Z => n12699);
   U390 : BUF_X1 port map( A => n12718, Z => n12697);
   U391 : BUF_X1 port map( A => n12719, Z => n12692);
   U392 : BUF_X1 port map( A => n12720, Z => n12691);
   U393 : BUF_X1 port map( A => n12726, Z => n12672);
   U394 : BUF_X1 port map( A => n12726, Z => n12673);
   U395 : BUF_X1 port map( A => n12728, Z => n12665);
   U396 : BUF_X1 port map( A => n12725, Z => n12674);
   U397 : BUF_X1 port map( A => n12728, Z => n12666);
   U398 : BUF_X1 port map( A => n12725, Z => n12675);
   U399 : BUF_X1 port map( A => n12728, Z => n12667);
   U400 : BUF_X1 port map( A => n12725, Z => n12676);
   U401 : BUF_X1 port map( A => n12727, Z => n12668);
   U402 : BUF_X1 port map( A => n12724, Z => n12677);
   U403 : BUF_X1 port map( A => n12727, Z => n12669);
   U404 : BUF_X1 port map( A => n12724, Z => n12678);
   U405 : BUF_X1 port map( A => n12727, Z => n12670);
   U406 : BUF_X1 port map( A => n12726, Z => n12671);
   U407 : BUF_X1 port map( A => n12729, Z => n12663);
   U408 : BUF_X1 port map( A => n12729, Z => n12664);
   U409 : BUF_X1 port map( A => n10545, Z => n12150);
   U410 : BUF_X1 port map( A => n10545, Z => n12151);
   U411 : BUF_X1 port map( A => n10545, Z => n12152);
   U412 : BUF_X1 port map( A => n10545, Z => n12153);
   U413 : BUF_X1 port map( A => n12158, Z => n12154);
   U414 : BUF_X1 port map( A => n12156, Z => n12155);
   U415 : BUF_X1 port map( A => n10545, Z => n12156);
   U416 : BUF_X1 port map( A => n12158, Z => n12157);
   U417 : BUF_X1 port map( A => n10573, Z => n12126);
   U418 : BUF_X1 port map( A => n10573, Z => n12127);
   U419 : BUF_X1 port map( A => n10573, Z => n12128);
   U420 : BUF_X1 port map( A => n10573, Z => n12129);
   U421 : BUF_X1 port map( A => n12134, Z => n12130);
   U422 : BUF_X1 port map( A => n12132, Z => n12131);
   U423 : BUF_X1 port map( A => n10573, Z => n12132);
   U424 : BUF_X1 port map( A => n12134, Z => n12133);
   U425 : BUF_X1 port map( A => n10565, Z => n12102);
   U426 : BUF_X1 port map( A => n10565, Z => n12103);
   U427 : BUF_X1 port map( A => n10565, Z => n12104);
   U428 : BUF_X1 port map( A => n10565, Z => n12105);
   U429 : BUF_X1 port map( A => n12110, Z => n12106);
   U430 : BUF_X1 port map( A => n12108, Z => n12107);
   U431 : BUF_X1 port map( A => n10565, Z => n12108);
   U432 : BUF_X1 port map( A => n12110, Z => n12109);
   U433 : BUF_X1 port map( A => n10557, Z => n12090);
   U434 : BUF_X1 port map( A => n10557, Z => n12091);
   U435 : BUF_X1 port map( A => n10557, Z => n12092);
   U436 : BUF_X1 port map( A => n10557, Z => n12093);
   U437 : BUF_X1 port map( A => n12098, Z => n12094);
   U438 : BUF_X1 port map( A => n12096, Z => n12095);
   U439 : BUF_X1 port map( A => n10557, Z => n12096);
   U440 : BUF_X1 port map( A => n12098, Z => n12097);
   U441 : BUF_X1 port map( A => n10574, Z => n12078);
   U442 : BUF_X1 port map( A => n10574, Z => n12079);
   U443 : BUF_X1 port map( A => n10574, Z => n12080);
   U444 : BUF_X1 port map( A => n10574, Z => n12081);
   U445 : BUF_X1 port map( A => n12086, Z => n12082);
   U446 : BUF_X1 port map( A => n12084, Z => n12083);
   U447 : BUF_X1 port map( A => n10574, Z => n12084);
   U448 : BUF_X1 port map( A => n12086, Z => n12085);
   U449 : BUF_X1 port map( A => n10566, Z => n12066);
   U450 : BUF_X1 port map( A => n10566, Z => n12067);
   U451 : BUF_X1 port map( A => n10566, Z => n12068);
   U452 : BUF_X1 port map( A => n10566, Z => n12069);
   U453 : BUF_X1 port map( A => n12074, Z => n12070);
   U454 : BUF_X1 port map( A => n12072, Z => n12071);
   U455 : BUF_X1 port map( A => n10566, Z => n12072);
   U456 : BUF_X1 port map( A => n12074, Z => n12073);
   U457 : BUF_X1 port map( A => n10558, Z => n12054);
   U458 : BUF_X1 port map( A => n10558, Z => n12055);
   U459 : BUF_X1 port map( A => n10558, Z => n12056);
   U460 : BUF_X1 port map( A => n10558, Z => n12057);
   U461 : BUF_X1 port map( A => n12062, Z => n12058);
   U462 : BUF_X1 port map( A => n12060, Z => n12059);
   U463 : BUF_X1 port map( A => n10558, Z => n12060);
   U464 : BUF_X1 port map( A => n12062, Z => n12061);
   U465 : BUF_X1 port map( A => n10581, Z => n12042);
   U466 : BUF_X1 port map( A => n10581, Z => n12043);
   U467 : BUF_X1 port map( A => n10581, Z => n12044);
   U468 : BUF_X1 port map( A => n10581, Z => n12045);
   U469 : BUF_X1 port map( A => n12050, Z => n12046);
   U470 : BUF_X1 port map( A => n12048, Z => n12047);
   U471 : BUF_X1 port map( A => n10581, Z => n12048);
   U472 : BUF_X1 port map( A => n12050, Z => n12049);
   U473 : BUF_X1 port map( A => n10586, Z => n12018);
   U474 : BUF_X1 port map( A => n10586, Z => n12019);
   U475 : BUF_X1 port map( A => n10586, Z => n12020);
   U476 : BUF_X1 port map( A => n10586, Z => n12021);
   U477 : BUF_X1 port map( A => n10584, Z => n11886);
   U478 : BUF_X1 port map( A => n10584, Z => n11887);
   U479 : BUF_X1 port map( A => n10584, Z => n11888);
   U480 : BUF_X1 port map( A => n10584, Z => n11889);
   U481 : BUF_X1 port map( A => n11894, Z => n11890);
   U482 : BUF_X1 port map( A => n11892, Z => n11891);
   U483 : BUF_X1 port map( A => n10584, Z => n11892);
   U484 : BUF_X1 port map( A => n11894, Z => n11893);
   U485 : BUF_X1 port map( A => n10575, Z => n11862);
   U486 : BUF_X1 port map( A => n10575, Z => n11863);
   U487 : BUF_X1 port map( A => n10575, Z => n11864);
   U488 : BUF_X1 port map( A => n10575, Z => n11865);
   U489 : BUF_X1 port map( A => n11870, Z => n11866);
   U490 : BUF_X1 port map( A => n11868, Z => n11867);
   U491 : BUF_X1 port map( A => n10575, Z => n11868);
   U492 : BUF_X1 port map( A => n11870, Z => n11869);
   U493 : BUF_X1 port map( A => n10567, Z => n11838);
   U494 : BUF_X1 port map( A => n10567, Z => n11839);
   U495 : BUF_X1 port map( A => n10567, Z => n11840);
   U496 : BUF_X1 port map( A => n10567, Z => n11841);
   U497 : BUF_X1 port map( A => n11846, Z => n11842);
   U498 : BUF_X1 port map( A => n11844, Z => n11843);
   U499 : BUF_X1 port map( A => n10567, Z => n11844);
   U500 : BUF_X1 port map( A => n11846, Z => n11845);
   U501 : BUF_X1 port map( A => n10559, Z => n11826);
   U502 : BUF_X1 port map( A => n10559, Z => n11827);
   U503 : BUF_X1 port map( A => n10559, Z => n11828);
   U504 : BUF_X1 port map( A => n10559, Z => n11829);
   U505 : BUF_X1 port map( A => n11834, Z => n11830);
   U506 : BUF_X1 port map( A => n11832, Z => n11831);
   U507 : BUF_X1 port map( A => n10559, Z => n11832);
   U508 : BUF_X1 port map( A => n11834, Z => n11833);
   U509 : BUF_X1 port map( A => n10576, Z => n11814);
   U510 : BUF_X1 port map( A => n10576, Z => n11815);
   U511 : BUF_X1 port map( A => n10576, Z => n11816);
   U512 : BUF_X1 port map( A => n10576, Z => n11817);
   U513 : BUF_X1 port map( A => n11822, Z => n11818);
   U514 : BUF_X1 port map( A => n11820, Z => n11819);
   U515 : BUF_X1 port map( A => n10576, Z => n11820);
   U516 : BUF_X1 port map( A => n11822, Z => n11821);
   U517 : BUF_X1 port map( A => n10568, Z => n11802);
   U518 : BUF_X1 port map( A => n10568, Z => n11803);
   U519 : BUF_X1 port map( A => n10568, Z => n11804);
   U520 : BUF_X1 port map( A => n10568, Z => n11805);
   U521 : BUF_X1 port map( A => n11810, Z => n11806);
   U522 : BUF_X1 port map( A => n11808, Z => n11807);
   U523 : BUF_X1 port map( A => n10568, Z => n11808);
   U524 : BUF_X1 port map( A => n11810, Z => n11809);
   U525 : BUF_X1 port map( A => n10560, Z => n11790);
   U526 : BUF_X1 port map( A => n10560, Z => n11791);
   U527 : BUF_X1 port map( A => n10560, Z => n11792);
   U528 : BUF_X1 port map( A => n10560, Z => n11793);
   U529 : BUF_X1 port map( A => n11798, Z => n11794);
   U530 : BUF_X1 port map( A => n11796, Z => n11795);
   U531 : BUF_X1 port map( A => n10560, Z => n11796);
   U532 : BUF_X1 port map( A => n11798, Z => n11797);
   U533 : BUF_X1 port map( A => n10582, Z => n11778);
   U534 : BUF_X1 port map( A => n10582, Z => n11779);
   U535 : BUF_X1 port map( A => n10582, Z => n11780);
   U536 : BUF_X1 port map( A => n10582, Z => n11781);
   U537 : BUF_X1 port map( A => n11786, Z => n11782);
   U538 : BUF_X1 port map( A => n11784, Z => n11783);
   U539 : BUF_X1 port map( A => n10582, Z => n11784);
   U540 : BUF_X1 port map( A => n11786, Z => n11785);
   U541 : BUF_X1 port map( A => n10603, Z => n11754);
   U542 : BUF_X1 port map( A => n10609, Z => n11646);
   U543 : BUF_X1 port map( A => n11654, Z => n11647);
   U544 : BUF_X1 port map( A => n11649, Z => n11648);
   U545 : BUF_X1 port map( A => n10609, Z => n11649);
   U546 : BUF_X1 port map( A => n10587, Z => n11634);
   U547 : BUF_X1 port map( A => n10587, Z => n11635);
   U548 : BUF_X1 port map( A => n10587, Z => n11636);
   U549 : BUF_X1 port map( A => n10587, Z => n11637);
   U550 : BUF_X1 port map( A => n11642, Z => n11638);
   U551 : BUF_X1 port map( A => n11640, Z => n11639);
   U552 : BUF_X1 port map( A => n10587, Z => n11640);
   U553 : BUF_X1 port map( A => n11642, Z => n11641);
   U554 : BUF_X1 port map( A => n10588, Z => n11622);
   U555 : BUF_X1 port map( A => n10588, Z => n11623);
   U556 : BUF_X1 port map( A => n10588, Z => n11624);
   U557 : BUF_X1 port map( A => n10588, Z => n11625);
   U558 : BUF_X1 port map( A => n11630, Z => n11626);
   U559 : BUF_X1 port map( A => n11628, Z => n11627);
   U560 : BUF_X1 port map( A => n10588, Z => n11628);
   U561 : BUF_X1 port map( A => n11630, Z => n11629);
   U562 : BUF_X1 port map( A => n10589, Z => n11610);
   U563 : BUF_X1 port map( A => n10589, Z => n11611);
   U564 : BUF_X1 port map( A => n10589, Z => n11612);
   U565 : BUF_X1 port map( A => n10589, Z => n11613);
   U566 : BUF_X1 port map( A => n11618, Z => n11614);
   U567 : BUF_X1 port map( A => n11616, Z => n11615);
   U568 : BUF_X1 port map( A => n10589, Z => n11616);
   U569 : BUF_X1 port map( A => n11618, Z => n11617);
   U570 : BUF_X1 port map( A => n10590, Z => n11598);
   U571 : BUF_X1 port map( A => n10590, Z => n11599);
   U572 : BUF_X1 port map( A => n10590, Z => n11600);
   U573 : BUF_X1 port map( A => n10590, Z => n11601);
   U574 : BUF_X1 port map( A => n11606, Z => n11602);
   U575 : BUF_X1 port map( A => n11604, Z => n11603);
   U576 : BUF_X1 port map( A => n10590, Z => n11604);
   U577 : BUF_X1 port map( A => n11606, Z => n11605);
   U578 : BUF_X1 port map( A => n10591, Z => n11586);
   U579 : BUF_X1 port map( A => n10591, Z => n11587);
   U580 : BUF_X1 port map( A => n10591, Z => n11588);
   U581 : BUF_X1 port map( A => n10591, Z => n11589);
   U582 : BUF_X1 port map( A => n11594, Z => n11590);
   U583 : BUF_X1 port map( A => n11592, Z => n11591);
   U584 : BUF_X1 port map( A => n10591, Z => n11592);
   U585 : BUF_X1 port map( A => n11594, Z => n11593);
   U586 : BUF_X1 port map( A => n10592, Z => n11574);
   U587 : BUF_X1 port map( A => n10592, Z => n11575);
   U588 : BUF_X1 port map( A => n10592, Z => n11576);
   U589 : BUF_X1 port map( A => n10592, Z => n11577);
   U590 : BUF_X1 port map( A => n11582, Z => n11578);
   U591 : BUF_X1 port map( A => n11580, Z => n11579);
   U592 : BUF_X1 port map( A => n10592, Z => n11580);
   U593 : BUF_X1 port map( A => n11582, Z => n11581);
   U594 : BUF_X1 port map( A => n10593, Z => n11562);
   U595 : BUF_X1 port map( A => n10593, Z => n11563);
   U596 : BUF_X1 port map( A => n10593, Z => n11564);
   U597 : BUF_X1 port map( A => n10593, Z => n11565);
   U598 : BUF_X1 port map( A => n11570, Z => n11566);
   U599 : BUF_X1 port map( A => n11568, Z => n11567);
   U600 : BUF_X1 port map( A => n10593, Z => n11568);
   U601 : BUF_X1 port map( A => n11570, Z => n11569);
   U602 : BUF_X1 port map( A => n10577, Z => n11550);
   U603 : BUF_X1 port map( A => n10577, Z => n11551);
   U604 : BUF_X1 port map( A => n10577, Z => n11552);
   U605 : BUF_X1 port map( A => n10577, Z => n11553);
   U606 : BUF_X1 port map( A => n11558, Z => n11554);
   U607 : BUF_X1 port map( A => n11556, Z => n11555);
   U608 : BUF_X1 port map( A => n10577, Z => n11556);
   U609 : BUF_X1 port map( A => n11558, Z => n11557);
   U610 : BUF_X1 port map( A => n10569, Z => n11538);
   U611 : BUF_X1 port map( A => n10569, Z => n11539);
   U612 : BUF_X1 port map( A => n10569, Z => n11540);
   U613 : BUF_X1 port map( A => n10569, Z => n11541);
   U614 : BUF_X1 port map( A => n11546, Z => n11542);
   U615 : BUF_X1 port map( A => n11544, Z => n11543);
   U616 : BUF_X1 port map( A => n10569, Z => n11544);
   U617 : BUF_X1 port map( A => n11546, Z => n11545);
   U618 : BUF_X1 port map( A => n10561, Z => n11526);
   U619 : BUF_X1 port map( A => n10561, Z => n11527);
   U620 : BUF_X1 port map( A => n10561, Z => n11528);
   U621 : BUF_X1 port map( A => n10561, Z => n11529);
   U622 : BUF_X1 port map( A => n11534, Z => n11530);
   U623 : BUF_X1 port map( A => n11532, Z => n11531);
   U624 : BUF_X1 port map( A => n10561, Z => n11532);
   U625 : BUF_X1 port map( A => n11534, Z => n11533);
   U626 : BUF_X1 port map( A => n10570, Z => n11502);
   U627 : BUF_X1 port map( A => n10570, Z => n11503);
   U628 : BUF_X1 port map( A => n10570, Z => n11504);
   U629 : BUF_X1 port map( A => n10570, Z => n11505);
   U630 : BUF_X1 port map( A => n11510, Z => n11506);
   U631 : BUF_X1 port map( A => n11508, Z => n11507);
   U632 : BUF_X1 port map( A => n10570, Z => n11508);
   U633 : BUF_X1 port map( A => n11510, Z => n11509);
   U634 : BUF_X1 port map( A => n10578, Z => n11490);
   U635 : BUF_X1 port map( A => n10578, Z => n11491);
   U636 : BUF_X1 port map( A => n10578, Z => n11492);
   U637 : BUF_X1 port map( A => n10578, Z => n11493);
   U638 : BUF_X1 port map( A => n11498, Z => n11494);
   U639 : BUF_X1 port map( A => n11496, Z => n11495);
   U640 : BUF_X1 port map( A => n10578, Z => n11496);
   U641 : BUF_X1 port map( A => n11498, Z => n11497);
   U642 : BUF_X1 port map( A => n10562, Z => n11478);
   U643 : BUF_X1 port map( A => n10562, Z => n11479);
   U644 : BUF_X1 port map( A => n10562, Z => n11480);
   U645 : BUF_X1 port map( A => n10562, Z => n11481);
   U646 : BUF_X1 port map( A => n11486, Z => n11482);
   U647 : BUF_X1 port map( A => n11484, Z => n11483);
   U648 : BUF_X1 port map( A => n10562, Z => n11484);
   U649 : BUF_X1 port map( A => n10579, Z => n11454);
   U650 : BUF_X1 port map( A => n10579, Z => n11455);
   U651 : BUF_X1 port map( A => n10579, Z => n11456);
   U652 : BUF_X1 port map( A => n10579, Z => n11457);
   U653 : BUF_X1 port map( A => n11462, Z => n11458);
   U654 : BUF_X1 port map( A => n11460, Z => n11459);
   U655 : BUF_X1 port map( A => n10579, Z => n11460);
   U656 : BUF_X1 port map( A => n11462, Z => n11461);
   U657 : BUF_X1 port map( A => n10563, Z => n11442);
   U658 : BUF_X1 port map( A => n10563, Z => n11443);
   U659 : BUF_X1 port map( A => n10563, Z => n11444);
   U660 : BUF_X1 port map( A => n10563, Z => n11445);
   U661 : BUF_X1 port map( A => n11450, Z => n11446);
   U662 : BUF_X1 port map( A => n11448, Z => n11447);
   U663 : BUF_X1 port map( A => n10563, Z => n11448);
   U664 : BUF_X1 port map( A => n10572, Z => n11430);
   U665 : BUF_X1 port map( A => n10572, Z => n11431);
   U666 : BUF_X1 port map( A => n10572, Z => n11432);
   U667 : BUF_X1 port map( A => n10572, Z => n11433);
   U668 : BUF_X1 port map( A => n11438, Z => n11434);
   U669 : BUF_X1 port map( A => n11436, Z => n11435);
   U670 : BUF_X1 port map( A => n10572, Z => n11436);
   U671 : BUF_X1 port map( A => n11438, Z => n11437);
   U672 : BUF_X1 port map( A => n10580, Z => n11418);
   U673 : BUF_X1 port map( A => n10580, Z => n11419);
   U674 : BUF_X1 port map( A => n10580, Z => n11420);
   U675 : BUF_X1 port map( A => n10580, Z => n11421);
   U676 : BUF_X1 port map( A => n11426, Z => n11422);
   U677 : BUF_X1 port map( A => n11424, Z => n11423);
   U678 : BUF_X1 port map( A => n10580, Z => n11424);
   U679 : BUF_X1 port map( A => n11426, Z => n11425);
   U680 : BUF_X1 port map( A => n10564, Z => n11406);
   U681 : BUF_X1 port map( A => n10564, Z => n11407);
   U682 : BUF_X1 port map( A => n10564, Z => n11408);
   U683 : BUF_X1 port map( A => n10564, Z => n11409);
   U684 : BUF_X1 port map( A => n11414, Z => n11410);
   U685 : BUF_X1 port map( A => n11412, Z => n11411);
   U686 : BUF_X1 port map( A => n10564, Z => n11412);
   U687 : BUF_X1 port map( A => n10583, Z => n11394);
   U688 : BUF_X1 port map( A => n10583, Z => n11395);
   U689 : BUF_X1 port map( A => n10583, Z => n11396);
   U690 : BUF_X1 port map( A => n10583, Z => n11397);
   U691 : BUF_X1 port map( A => n11402, Z => n11398);
   U692 : BUF_X1 port map( A => n11400, Z => n11399);
   U693 : BUF_X1 port map( A => n10583, Z => n11400);
   U694 : BUF_X1 port map( A => n11402, Z => n11401);
   U695 : BUF_X1 port map( A => n10585, Z => n11382);
   U696 : BUF_X1 port map( A => n10585, Z => n11383);
   U697 : BUF_X1 port map( A => n10585, Z => n11384);
   U698 : BUF_X1 port map( A => n10585, Z => n11385);
   U699 : BUF_X1 port map( A => n11390, Z => n11386);
   U700 : BUF_X1 port map( A => n11388, Z => n11387);
   U701 : BUF_X1 port map( A => n10585, Z => n11388);
   U702 : BUF_X1 port map( A => n11390, Z => n11389);
   U703 : BUF_X1 port map( A => n10619, Z => n12407);
   U704 : BUF_X1 port map( A => n10619, Z => n12408);
   U705 : BUF_X1 port map( A => n10619, Z => n12409);
   U706 : BUF_X1 port map( A => n10619, Z => n12410);
   U707 : BUF_X1 port map( A => n12415, Z => n12411);
   U708 : BUF_X1 port map( A => n12413, Z => n12412);
   U709 : BUF_X1 port map( A => n10619, Z => n12413);
   U710 : BUF_X1 port map( A => n12415, Z => n12414);
   U711 : BUF_X1 port map( A => n10620, Z => n12396);
   U712 : BUF_X1 port map( A => n10620, Z => n12397);
   U713 : BUF_X1 port map( A => n10620, Z => n12398);
   U714 : BUF_X1 port map( A => n10620, Z => n12399);
   U715 : BUF_X1 port map( A => n12404, Z => n12400);
   U716 : BUF_X1 port map( A => n12402, Z => n12401);
   U717 : BUF_X1 port map( A => n10620, Z => n12402);
   U718 : BUF_X1 port map( A => n12404, Z => n12403);
   U719 : BUF_X1 port map( A => n10621, Z => n12385);
   U720 : BUF_X1 port map( A => n10621, Z => n12386);
   U721 : BUF_X1 port map( A => n10621, Z => n12387);
   U722 : BUF_X1 port map( A => n10621, Z => n12388);
   U723 : BUF_X1 port map( A => n12393, Z => n12389);
   U724 : BUF_X1 port map( A => n12391, Z => n12390);
   U725 : BUF_X1 port map( A => n10621, Z => n12391);
   U726 : BUF_X1 port map( A => n12393, Z => n12392);
   U727 : BUF_X1 port map( A => n10622, Z => n12374);
   U728 : BUF_X1 port map( A => n10622, Z => n12375);
   U729 : BUF_X1 port map( A => n10622, Z => n12376);
   U730 : BUF_X1 port map( A => n10622, Z => n12377);
   U731 : BUF_X1 port map( A => n12382, Z => n12378);
   U732 : BUF_X1 port map( A => n12380, Z => n12379);
   U733 : BUF_X1 port map( A => n10622, Z => n12380);
   U734 : BUF_X1 port map( A => n12382, Z => n12381);
   U735 : BUF_X1 port map( A => n10623, Z => n12363);
   U736 : BUF_X1 port map( A => n10623, Z => n12364);
   U737 : BUF_X1 port map( A => n10623, Z => n12365);
   U738 : BUF_X1 port map( A => n10623, Z => n12366);
   U739 : BUF_X1 port map( A => n12371, Z => n12367);
   U740 : BUF_X1 port map( A => n12369, Z => n12368);
   U741 : BUF_X1 port map( A => n10623, Z => n12369);
   U742 : BUF_X1 port map( A => n12371, Z => n12370);
   U743 : BUF_X1 port map( A => n10624, Z => n12352);
   U744 : BUF_X1 port map( A => n10624, Z => n12353);
   U745 : BUF_X1 port map( A => n10624, Z => n12354);
   U746 : BUF_X1 port map( A => n10624, Z => n12355);
   U747 : BUF_X1 port map( A => n12360, Z => n12356);
   U748 : BUF_X1 port map( A => n12358, Z => n12357);
   U749 : BUF_X1 port map( A => n10624, Z => n12358);
   U750 : BUF_X1 port map( A => n12360, Z => n12359);
   U751 : BUF_X1 port map( A => n10618, Z => n12341);
   U752 : BUF_X1 port map( A => n10618, Z => n12342);
   U753 : BUF_X1 port map( A => n10618, Z => n12343);
   U754 : BUF_X1 port map( A => n10618, Z => n12344);
   U755 : BUF_X1 port map( A => n12349, Z => n12345);
   U756 : BUF_X1 port map( A => n12347, Z => n12346);
   U757 : BUF_X1 port map( A => n10618, Z => n12347);
   U758 : BUF_X1 port map( A => n12349, Z => n12348);
   U759 : BUF_X1 port map( A => n10615, Z => n12330);
   U760 : BUF_X1 port map( A => n10615, Z => n12331);
   U761 : BUF_X1 port map( A => n10615, Z => n12332);
   U762 : BUF_X1 port map( A => n10615, Z => n12333);
   U763 : BUF_X1 port map( A => n12338, Z => n12334);
   U764 : BUF_X1 port map( A => n12336, Z => n12335);
   U765 : BUF_X1 port map( A => n10615, Z => n12336);
   U766 : BUF_X1 port map( A => n12338, Z => n12337);
   U767 : BUF_X1 port map( A => n10614, Z => n12318);
   U768 : BUF_X1 port map( A => n10614, Z => n12319);
   U769 : BUF_X1 port map( A => n10614, Z => n12320);
   U770 : BUF_X1 port map( A => n10614, Z => n12321);
   U771 : BUF_X1 port map( A => n12326, Z => n12322);
   U772 : BUF_X1 port map( A => n12324, Z => n12323);
   U773 : BUF_X1 port map( A => n10614, Z => n12324);
   U774 : BUF_X1 port map( A => n12326, Z => n12325);
   U775 : BUF_X1 port map( A => n10617, Z => n12306);
   U776 : BUF_X1 port map( A => n10617, Z => n12307);
   U777 : BUF_X1 port map( A => n10617, Z => n12308);
   U778 : BUF_X1 port map( A => n10617, Z => n12309);
   U779 : BUF_X1 port map( A => n12314, Z => n12310);
   U780 : BUF_X1 port map( A => n12312, Z => n12311);
   U781 : BUF_X1 port map( A => n10617, Z => n12312);
   U782 : BUF_X1 port map( A => n12314, Z => n12313);
   U783 : BUF_X1 port map( A => n10603, Z => n11755);
   U784 : BUF_X1 port map( A => n11486, Z => n11485);
   U785 : BUF_X1 port map( A => n10541, Z => n12198);
   U786 : BUF_X1 port map( A => n12026, Z => n12022);
   U787 : BUF_X1 port map( A => n10596, Z => n12006);
   U788 : BUF_X1 port map( A => n11450, Z => n11449);
   U789 : BUF_X1 port map( A => n11414, Z => n11413);
   U790 : BUF_X1 port map( A => n10611, Z => n12270);
   U791 : BUF_X1 port map( A => n10539, Z => n12222);
   U792 : BUF_X1 port map( A => n10539, Z => n12223);
   U793 : BUF_X1 port map( A => n10539, Z => n12224);
   U794 : BUF_X1 port map( A => n10539, Z => n12225);
   U795 : BUF_X1 port map( A => n12230, Z => n12226);
   U796 : BUF_X1 port map( A => n12228, Z => n12227);
   U797 : BUF_X1 port map( A => n10539, Z => n12228);
   U798 : BUF_X1 port map( A => n12230, Z => n12229);
   U799 : BUF_X1 port map( A => n10540, Z => n12210);
   U800 : BUF_X1 port map( A => n10540, Z => n12211);
   U801 : BUF_X1 port map( A => n10540, Z => n12212);
   U802 : BUF_X1 port map( A => n10540, Z => n12213);
   U803 : BUF_X1 port map( A => n12218, Z => n12214);
   U804 : BUF_X1 port map( A => n12216, Z => n12215);
   U805 : BUF_X1 port map( A => n10540, Z => n12216);
   U806 : BUF_X1 port map( A => n12218, Z => n12217);
   U807 : BUF_X1 port map( A => n10541, Z => n12199);
   U808 : BUF_X1 port map( A => n10541, Z => n12200);
   U809 : BUF_X1 port map( A => n10541, Z => n12201);
   U810 : BUF_X1 port map( A => n10541, Z => n12202);
   U811 : BUF_X1 port map( A => n10541, Z => n12203);
   U812 : BUF_X1 port map( A => n12198, Z => n12204);
   U813 : BUF_X1 port map( A => n12200, Z => n12205);
   U814 : BUF_X1 port map( A => n10542, Z => n12186);
   U815 : BUF_X1 port map( A => n10542, Z => n12187);
   U816 : BUF_X1 port map( A => n10542, Z => n12188);
   U817 : BUF_X1 port map( A => n10542, Z => n12189);
   U818 : BUF_X1 port map( A => n12194, Z => n12190);
   U819 : BUF_X1 port map( A => n12192, Z => n12191);
   U820 : BUF_X1 port map( A => n10542, Z => n12192);
   U821 : BUF_X1 port map( A => n12194, Z => n12193);
   U822 : BUF_X1 port map( A => n10543, Z => n12174);
   U823 : BUF_X1 port map( A => n10543, Z => n12175);
   U824 : BUF_X1 port map( A => n10543, Z => n12176);
   U825 : BUF_X1 port map( A => n10543, Z => n12177);
   U826 : BUF_X1 port map( A => n12182, Z => n12178);
   U827 : BUF_X1 port map( A => n12180, Z => n12179);
   U828 : BUF_X1 port map( A => n10543, Z => n12180);
   U829 : BUF_X1 port map( A => n12182, Z => n12181);
   U830 : BUF_X1 port map( A => n10544, Z => n12162);
   U831 : BUF_X1 port map( A => n10544, Z => n12163);
   U832 : BUF_X1 port map( A => n10544, Z => n12164);
   U833 : BUF_X1 port map( A => n10544, Z => n12165);
   U834 : BUF_X1 port map( A => n12170, Z => n12166);
   U835 : BUF_X1 port map( A => n12168, Z => n12167);
   U836 : BUF_X1 port map( A => n10544, Z => n12168);
   U837 : BUF_X1 port map( A => n12170, Z => n12169);
   U838 : BUF_X1 port map( A => n10546, Z => n12138);
   U839 : BUF_X1 port map( A => n10546, Z => n12139);
   U840 : BUF_X1 port map( A => n10546, Z => n12140);
   U841 : BUF_X1 port map( A => n10546, Z => n12141);
   U842 : BUF_X1 port map( A => n12146, Z => n12142);
   U843 : BUF_X1 port map( A => n12144, Z => n12143);
   U844 : BUF_X1 port map( A => n10546, Z => n12144);
   U845 : BUF_X1 port map( A => n12146, Z => n12145);
   U846 : BUF_X1 port map( A => n10547, Z => n12114);
   U847 : BUF_X1 port map( A => n10547, Z => n12115);
   U848 : BUF_X1 port map( A => n10547, Z => n12116);
   U849 : BUF_X1 port map( A => n10547, Z => n12117);
   U850 : BUF_X1 port map( A => n12122, Z => n12118);
   U851 : BUF_X1 port map( A => n12120, Z => n12119);
   U852 : BUF_X1 port map( A => n10547, Z => n12120);
   U853 : BUF_X1 port map( A => n12122, Z => n12121);
   U854 : BUF_X1 port map( A => n10595, Z => n12030);
   U855 : BUF_X1 port map( A => n10595, Z => n12031);
   U856 : BUF_X1 port map( A => n10595, Z => n12032);
   U857 : BUF_X1 port map( A => n10595, Z => n12033);
   U858 : BUF_X1 port map( A => n12038, Z => n12034);
   U859 : BUF_X1 port map( A => n12036, Z => n12035);
   U860 : BUF_X1 port map( A => n10595, Z => n12036);
   U861 : BUF_X1 port map( A => n12038, Z => n12037);
   U862 : BUF_X1 port map( A => n12018, Z => n12023);
   U863 : BUF_X1 port map( A => n10586, Z => n12024);
   U864 : BUF_X1 port map( A => n12026, Z => n12025);
   U865 : BUF_X1 port map( A => n12014, Z => n12007);
   U866 : BUF_X1 port map( A => n12012, Z => n12008);
   U867 : BUF_X1 port map( A => n10596, Z => n12009);
   U868 : BUF_X1 port map( A => n10596, Z => n12010);
   U869 : BUF_X1 port map( A => n10596, Z => n12011);
   U870 : BUF_X1 port map( A => n10596, Z => n12012);
   U871 : BUF_X1 port map( A => n12014, Z => n12013);
   U872 : BUF_X1 port map( A => n10597, Z => n11994);
   U873 : BUF_X1 port map( A => n10597, Z => n11995);
   U874 : BUF_X1 port map( A => n10597, Z => n11996);
   U875 : BUF_X1 port map( A => n10597, Z => n11997);
   U876 : BUF_X1 port map( A => n12002, Z => n11998);
   U877 : BUF_X1 port map( A => n12000, Z => n11999);
   U878 : BUF_X1 port map( A => n10597, Z => n12000);
   U879 : BUF_X1 port map( A => n12002, Z => n12001);
   U880 : BUF_X1 port map( A => n10598, Z => n11982);
   U881 : BUF_X1 port map( A => n10598, Z => n11983);
   U882 : BUF_X1 port map( A => n10598, Z => n11984);
   U883 : BUF_X1 port map( A => n10598, Z => n11985);
   U884 : BUF_X1 port map( A => n11990, Z => n11986);
   U885 : BUF_X1 port map( A => n11988, Z => n11987);
   U886 : BUF_X1 port map( A => n10598, Z => n11988);
   U887 : BUF_X1 port map( A => n11990, Z => n11989);
   U888 : BUF_X1 port map( A => n10599, Z => n11970);
   U889 : BUF_X1 port map( A => n10599, Z => n11971);
   U890 : BUF_X1 port map( A => n10599, Z => n11972);
   U891 : BUF_X1 port map( A => n10599, Z => n11973);
   U892 : BUF_X1 port map( A => n11978, Z => n11974);
   U893 : BUF_X1 port map( A => n11976, Z => n11975);
   U894 : BUF_X1 port map( A => n10599, Z => n11976);
   U895 : BUF_X1 port map( A => n11978, Z => n11977);
   U896 : BUF_X1 port map( A => n10548, Z => n11958);
   U897 : BUF_X1 port map( A => n10548, Z => n11959);
   U898 : BUF_X1 port map( A => n10548, Z => n11960);
   U899 : BUF_X1 port map( A => n10548, Z => n11961);
   U900 : BUF_X1 port map( A => n11966, Z => n11962);
   U901 : BUF_X1 port map( A => n11964, Z => n11963);
   U902 : BUF_X1 port map( A => n10548, Z => n11964);
   U903 : BUF_X1 port map( A => n11966, Z => n11965);
   U904 : BUF_X1 port map( A => n10549, Z => n11946);
   U905 : BUF_X1 port map( A => n10549, Z => n11947);
   U906 : BUF_X1 port map( A => n10549, Z => n11948);
   U907 : BUF_X1 port map( A => n10549, Z => n11949);
   U908 : BUF_X1 port map( A => n11954, Z => n11950);
   U909 : BUF_X1 port map( A => n11952, Z => n11951);
   U910 : BUF_X1 port map( A => n10549, Z => n11952);
   U911 : BUF_X1 port map( A => n11954, Z => n11953);
   U912 : BUF_X1 port map( A => n10550, Z => n11934);
   U913 : BUF_X1 port map( A => n10550, Z => n11935);
   U914 : BUF_X1 port map( A => n10550, Z => n11936);
   U915 : BUF_X1 port map( A => n10550, Z => n11937);
   U916 : BUF_X1 port map( A => n11942, Z => n11938);
   U917 : BUF_X1 port map( A => n11940, Z => n11939);
   U918 : BUF_X1 port map( A => n10550, Z => n11940);
   U919 : BUF_X1 port map( A => n11942, Z => n11941);
   U920 : BUF_X1 port map( A => n10600, Z => n11922);
   U921 : BUF_X1 port map( A => n10600, Z => n11923);
   U922 : BUF_X1 port map( A => n10600, Z => n11924);
   U923 : BUF_X1 port map( A => n10600, Z => n11925);
   U924 : BUF_X1 port map( A => n11930, Z => n11926);
   U925 : BUF_X1 port map( A => n11928, Z => n11927);
   U926 : BUF_X1 port map( A => n10600, Z => n11928);
   U927 : BUF_X1 port map( A => n11930, Z => n11929);
   U928 : BUF_X1 port map( A => n10601, Z => n11910);
   U929 : BUF_X1 port map( A => n10601, Z => n11911);
   U930 : BUF_X1 port map( A => n10601, Z => n11912);
   U931 : BUF_X1 port map( A => n10601, Z => n11913);
   U932 : BUF_X1 port map( A => n11918, Z => n11914);
   U933 : BUF_X1 port map( A => n11916, Z => n11915);
   U934 : BUF_X1 port map( A => n10601, Z => n11916);
   U935 : BUF_X1 port map( A => n11918, Z => n11917);
   U936 : BUF_X1 port map( A => n10552, Z => n11874);
   U937 : BUF_X1 port map( A => n10552, Z => n11875);
   U938 : BUF_X1 port map( A => n10552, Z => n11876);
   U939 : BUF_X1 port map( A => n10552, Z => n11877);
   U940 : BUF_X1 port map( A => n11882, Z => n11878);
   U941 : BUF_X1 port map( A => n11880, Z => n11879);
   U942 : BUF_X1 port map( A => n10552, Z => n11880);
   U943 : BUF_X1 port map( A => n11882, Z => n11881);
   U944 : BUF_X1 port map( A => n10602, Z => n11766);
   U945 : BUF_X1 port map( A => n10602, Z => n11767);
   U946 : BUF_X1 port map( A => n10602, Z => n11768);
   U947 : BUF_X1 port map( A => n10602, Z => n11769);
   U948 : BUF_X1 port map( A => n11774, Z => n11770);
   U949 : BUF_X1 port map( A => n11772, Z => n11771);
   U950 : BUF_X1 port map( A => n10602, Z => n11772);
   U951 : BUF_X1 port map( A => n11774, Z => n11773);
   U952 : BUF_X1 port map( A => n10603, Z => n11756);
   U953 : BUF_X1 port map( A => n10603, Z => n11757);
   U954 : BUF_X1 port map( A => n11762, Z => n11758);
   U955 : BUF_X1 port map( A => n11754, Z => n11759);
   U956 : BUF_X1 port map( A => n10603, Z => n11760);
   U957 : BUF_X1 port map( A => n11762, Z => n11761);
   U958 : BUF_X1 port map( A => n10604, Z => n11742);
   U959 : BUF_X1 port map( A => n10604, Z => n11743);
   U960 : BUF_X1 port map( A => n10604, Z => n11744);
   U961 : BUF_X1 port map( A => n10604, Z => n11745);
   U962 : BUF_X1 port map( A => n11750, Z => n11746);
   U963 : BUF_X1 port map( A => n11748, Z => n11747);
   U964 : BUF_X1 port map( A => n10604, Z => n11748);
   U965 : BUF_X1 port map( A => n11750, Z => n11749);
   U966 : BUF_X1 port map( A => n10605, Z => n11730);
   U967 : BUF_X1 port map( A => n10605, Z => n11731);
   U968 : BUF_X1 port map( A => n10605, Z => n11732);
   U969 : BUF_X1 port map( A => n10605, Z => n11733);
   U970 : BUF_X1 port map( A => n11738, Z => n11734);
   U971 : BUF_X1 port map( A => n11736, Z => n11735);
   U972 : BUF_X1 port map( A => n10605, Z => n11736);
   U973 : BUF_X1 port map( A => n11738, Z => n11737);
   U974 : BUF_X1 port map( A => n10606, Z => n11718);
   U975 : BUF_X1 port map( A => n10606, Z => n11719);
   U976 : BUF_X1 port map( A => n10606, Z => n11720);
   U977 : BUF_X1 port map( A => n10606, Z => n11721);
   U978 : BUF_X1 port map( A => n11726, Z => n11722);
   U979 : BUF_X1 port map( A => n11724, Z => n11723);
   U980 : BUF_X1 port map( A => n10606, Z => n11724);
   U981 : BUF_X1 port map( A => n11726, Z => n11725);
   U982 : BUF_X1 port map( A => n10607, Z => n11706);
   U983 : BUF_X1 port map( A => n10607, Z => n11707);
   U984 : BUF_X1 port map( A => n10607, Z => n11708);
   U985 : BUF_X1 port map( A => n10607, Z => n11709);
   U986 : BUF_X1 port map( A => n11714, Z => n11710);
   U987 : BUF_X1 port map( A => n11712, Z => n11711);
   U988 : BUF_X1 port map( A => n10607, Z => n11712);
   U989 : BUF_X1 port map( A => n11714, Z => n11713);
   U990 : BUF_X1 port map( A => n10554, Z => n11694);
   U991 : BUF_X1 port map( A => n10554, Z => n11695);
   U992 : BUF_X1 port map( A => n10554, Z => n11696);
   U993 : BUF_X1 port map( A => n10554, Z => n11697);
   U994 : BUF_X1 port map( A => n11702, Z => n11698);
   U995 : BUF_X1 port map( A => n11700, Z => n11699);
   U996 : BUF_X1 port map( A => n10554, Z => n11700);
   U997 : BUF_X1 port map( A => n11702, Z => n11701);
   U998 : BUF_X1 port map( A => n10555, Z => n11682);
   U999 : BUF_X1 port map( A => n10555, Z => n11683);
   U1000 : BUF_X1 port map( A => n10555, Z => n11684);
   U1001 : BUF_X1 port map( A => n10555, Z => n11685);
   U1002 : BUF_X1 port map( A => n11690, Z => n11686);
   U1003 : BUF_X1 port map( A => n11688, Z => n11687);
   U1004 : BUF_X1 port map( A => n10555, Z => n11688);
   U1005 : BUF_X1 port map( A => n11690, Z => n11689);
   U1006 : BUF_X1 port map( A => n10556, Z => n11670);
   U1007 : BUF_X1 port map( A => n10556, Z => n11671);
   U1008 : BUF_X1 port map( A => n10556, Z => n11672);
   U1009 : BUF_X1 port map( A => n10556, Z => n11673);
   U1010 : BUF_X1 port map( A => n11678, Z => n11674);
   U1011 : BUF_X1 port map( A => n11676, Z => n11675);
   U1012 : BUF_X1 port map( A => n10556, Z => n11676);
   U1013 : BUF_X1 port map( A => n11678, Z => n11677);
   U1014 : BUF_X1 port map( A => n10608, Z => n11658);
   U1015 : BUF_X1 port map( A => n10608, Z => n11659);
   U1016 : BUF_X1 port map( A => n10608, Z => n11660);
   U1017 : BUF_X1 port map( A => n10608, Z => n11661);
   U1018 : BUF_X1 port map( A => n11666, Z => n11662);
   U1019 : BUF_X1 port map( A => n11664, Z => n11663);
   U1020 : BUF_X1 port map( A => n10608, Z => n11664);
   U1021 : BUF_X1 port map( A => n11666, Z => n11665);
   U1022 : BUF_X1 port map( A => n10609, Z => n11653);
   U1023 : BUF_X1 port map( A => n10609, Z => n11652);
   U1024 : BUF_X1 port map( A => n11654, Z => n11651);
   U1025 : BUF_X1 port map( A => n10609, Z => n11650);
   U1026 : BUF_X1 port map( A => n10610, Z => n12294);
   U1027 : BUF_X1 port map( A => n10610, Z => n12295);
   U1028 : BUF_X1 port map( A => n10610, Z => n12296);
   U1029 : BUF_X1 port map( A => n10610, Z => n12297);
   U1030 : BUF_X1 port map( A => n12302, Z => n12298);
   U1031 : BUF_X1 port map( A => n12300, Z => n12299);
   U1032 : BUF_X1 port map( A => n10610, Z => n12300);
   U1033 : BUF_X1 port map( A => n12302, Z => n12301);
   U1034 : BUF_X1 port map( A => n10611, Z => n12271);
   U1035 : BUF_X1 port map( A => n10611, Z => n12272);
   U1036 : BUF_X1 port map( A => n10611, Z => n12273);
   U1037 : BUF_X1 port map( A => n10611, Z => n12274);
   U1038 : BUF_X1 port map( A => n10611, Z => n12275);
   U1039 : BUF_X1 port map( A => n12270, Z => n12276);
   U1040 : BUF_X1 port map( A => n12272, Z => n12277);
   U1041 : BUF_X1 port map( A => n10612, Z => n12258);
   U1042 : BUF_X1 port map( A => n10612, Z => n12259);
   U1043 : BUF_X1 port map( A => n10612, Z => n12260);
   U1044 : BUF_X1 port map( A => n10612, Z => n12261);
   U1045 : BUF_X1 port map( A => n12266, Z => n12262);
   U1046 : BUF_X1 port map( A => n12264, Z => n12263);
   U1047 : BUF_X1 port map( A => n10612, Z => n12264);
   U1048 : BUF_X1 port map( A => n12266, Z => n12265);
   U1049 : BUF_X1 port map( A => n10613, Z => n12246);
   U1050 : BUF_X1 port map( A => n10613, Z => n12247);
   U1051 : BUF_X1 port map( A => n10613, Z => n12248);
   U1052 : BUF_X1 port map( A => n10613, Z => n12249);
   U1053 : BUF_X1 port map( A => n12254, Z => n12250);
   U1054 : BUF_X1 port map( A => n12252, Z => n12251);
   U1055 : BUF_X1 port map( A => n10613, Z => n12252);
   U1056 : BUF_X1 port map( A => n12254, Z => n12253);
   U1057 : BUF_X1 port map( A => n12713, Z => n12712);
   U1058 : BUF_X1 port map( A => n10539, Z => n12230);
   U1059 : BUF_X1 port map( A => n10540, Z => n12218);
   U1060 : BUF_X1 port map( A => n12201, Z => n12206);
   U1061 : BUF_X1 port map( A => n10542, Z => n12194);
   U1062 : BUF_X1 port map( A => n10543, Z => n12182);
   U1063 : BUF_X1 port map( A => n10544, Z => n12170);
   U1064 : BUF_X1 port map( A => n10545, Z => n12158);
   U1065 : BUF_X1 port map( A => n10546, Z => n12146);
   U1066 : BUF_X1 port map( A => n10573, Z => n12134);
   U1067 : BUF_X1 port map( A => n10547, Z => n12122);
   U1068 : BUF_X1 port map( A => n10565, Z => n12110);
   U1069 : BUF_X1 port map( A => n10557, Z => n12098);
   U1070 : BUF_X1 port map( A => n10574, Z => n12086);
   U1071 : BUF_X1 port map( A => n10566, Z => n12074);
   U1072 : BUF_X1 port map( A => n10558, Z => n12062);
   U1073 : BUF_X1 port map( A => n10581, Z => n12050);
   U1074 : BUF_X1 port map( A => n10595, Z => n12038);
   U1075 : BUF_X1 port map( A => n10586, Z => n12026);
   U1076 : BUF_X1 port map( A => n10596, Z => n12014);
   U1077 : BUF_X1 port map( A => n10597, Z => n12002);
   U1078 : BUF_X1 port map( A => n10598, Z => n11990);
   U1079 : BUF_X1 port map( A => n10599, Z => n11978);
   U1080 : BUF_X1 port map( A => n10548, Z => n11966);
   U1081 : BUF_X1 port map( A => n10549, Z => n11954);
   U1082 : BUF_X1 port map( A => n10550, Z => n11942);
   U1083 : BUF_X1 port map( A => n10600, Z => n11930);
   U1084 : BUF_X1 port map( A => n10601, Z => n11918);
   U1085 : BUF_X1 port map( A => n10584, Z => n11894);
   U1086 : BUF_X1 port map( A => n10552, Z => n11882);
   U1087 : BUF_X1 port map( A => n10575, Z => n11870);
   U1088 : BUF_X1 port map( A => n10567, Z => n11846);
   U1089 : BUF_X1 port map( A => n10559, Z => n11834);
   U1090 : BUF_X1 port map( A => n10576, Z => n11822);
   U1091 : BUF_X1 port map( A => n10568, Z => n11810);
   U1092 : BUF_X1 port map( A => n10560, Z => n11798);
   U1093 : BUF_X1 port map( A => n10582, Z => n11786);
   U1094 : BUF_X1 port map( A => n10602, Z => n11774);
   U1095 : BUF_X1 port map( A => n10603, Z => n11762);
   U1096 : BUF_X1 port map( A => n10604, Z => n11750);
   U1097 : BUF_X1 port map( A => n10605, Z => n11738);
   U1098 : BUF_X1 port map( A => n10606, Z => n11726);
   U1099 : BUF_X1 port map( A => n10607, Z => n11714);
   U1100 : BUF_X1 port map( A => n10554, Z => n11702);
   U1101 : BUF_X1 port map( A => n10555, Z => n11690);
   U1102 : BUF_X1 port map( A => n10556, Z => n11678);
   U1103 : BUF_X1 port map( A => n10608, Z => n11666);
   U1104 : BUF_X1 port map( A => n10609, Z => n11654);
   U1105 : BUF_X1 port map( A => n10587, Z => n11642);
   U1106 : BUF_X1 port map( A => n10588, Z => n11630);
   U1107 : BUF_X1 port map( A => n10589, Z => n11618);
   U1108 : BUF_X1 port map( A => n10590, Z => n11606);
   U1109 : BUF_X1 port map( A => n10591, Z => n11594);
   U1110 : BUF_X1 port map( A => n10592, Z => n11582);
   U1111 : BUF_X1 port map( A => n10593, Z => n11570);
   U1112 : BUF_X1 port map( A => n10577, Z => n11558);
   U1113 : BUF_X1 port map( A => n10569, Z => n11546);
   U1114 : BUF_X1 port map( A => n10561, Z => n11534);
   U1115 : BUF_X1 port map( A => n10570, Z => n11510);
   U1116 : BUF_X1 port map( A => n10578, Z => n11498);
   U1117 : BUF_X1 port map( A => n10562, Z => n11486);
   U1118 : BUF_X1 port map( A => n10579, Z => n11462);
   U1119 : BUF_X1 port map( A => n10563, Z => n11450);
   U1120 : BUF_X1 port map( A => n10572, Z => n11438);
   U1121 : BUF_X1 port map( A => n10580, Z => n11426);
   U1122 : BUF_X1 port map( A => n10564, Z => n11414);
   U1123 : BUF_X1 port map( A => n10583, Z => n11402);
   U1124 : BUF_X1 port map( A => n10585, Z => n11390);
   U1125 : BUF_X1 port map( A => n10619, Z => n12415);
   U1126 : BUF_X1 port map( A => n10620, Z => n12404);
   U1127 : BUF_X1 port map( A => n10621, Z => n12393);
   U1128 : BUF_X1 port map( A => n10622, Z => n12382);
   U1129 : BUF_X1 port map( A => n10623, Z => n12371);
   U1130 : BUF_X1 port map( A => n10624, Z => n12360);
   U1131 : BUF_X1 port map( A => n10618, Z => n12349);
   U1132 : BUF_X1 port map( A => n10615, Z => n12338);
   U1133 : BUF_X1 port map( A => n10614, Z => n12326);
   U1134 : BUF_X1 port map( A => n10617, Z => n12314);
   U1135 : BUF_X1 port map( A => n10610, Z => n12302);
   U1136 : BUF_X1 port map( A => n12273, Z => n12278);
   U1137 : BUF_X1 port map( A => n10612, Z => n12266);
   U1138 : BUF_X1 port map( A => n10613, Z => n12254);
   U1139 : BUF_X1 port map( A => n4339, Z => n10986);
   U1140 : BUF_X1 port map( A => n2871, Z => n11250);
   U1141 : BUF_X1 port map( A => n4339, Z => n10987);
   U1142 : BUF_X1 port map( A => n2871, Z => n11251);
   U1143 : BUF_X1 port map( A => n4337, Z => n10992);
   U1144 : BUF_X1 port map( A => n4340, Z => n10983);
   U1145 : BUF_X1 port map( A => n2869, Z => n11256);
   U1146 : BUF_X1 port map( A => n2872, Z => n11247);
   U1147 : BUF_X1 port map( A => n4337, Z => n10993);
   U1148 : BUF_X1 port map( A => n4340, Z => n10984);
   U1149 : BUF_X1 port map( A => n2869, Z => n11257);
   U1150 : BUF_X1 port map( A => n2872, Z => n11248);
   U1151 : BUF_X1 port map( A => n4318, Z => n11046);
   U1152 : BUF_X1 port map( A => n2850, Z => n11310);
   U1153 : BUF_X1 port map( A => n4318, Z => n11047);
   U1154 : BUF_X1 port map( A => n2850, Z => n11311);
   U1155 : BUF_X1 port map( A => n4298, Z => n11079);
   U1156 : BUF_X1 port map( A => n2798, Z => n11343);
   U1157 : BUF_X1 port map( A => n4298, Z => n11080);
   U1158 : BUF_X1 port map( A => n2798, Z => n11344);
   U1159 : BUF_X1 port map( A => n4360, Z => n10947);
   U1160 : BUF_X1 port map( A => n2924, Z => n11211);
   U1161 : BUF_X1 port map( A => n4360, Z => n10948);
   U1162 : BUF_X1 port map( A => n2924, Z => n11212);
   U1163 : BUF_X1 port map( A => n4307, Z => n11055);
   U1164 : BUF_X1 port map( A => n2807, Z => n11319);
   U1165 : BUF_X1 port map( A => n4307, Z => n11056);
   U1166 : BUF_X1 port map( A => n2807, Z => n11320);
   U1167 : BUF_X1 port map( A => n4335, Z => n10998);
   U1168 : BUF_X1 port map( A => n4338, Z => n10989);
   U1169 : BUF_X1 port map( A => n2867, Z => n11262);
   U1170 : BUF_X1 port map( A => n2870, Z => n11253);
   U1171 : BUF_X1 port map( A => n4335, Z => n10999);
   U1172 : BUF_X1 port map( A => n4338, Z => n10990);
   U1173 : BUF_X1 port map( A => n2867, Z => n11263);
   U1174 : BUF_X1 port map( A => n2870, Z => n11254);
   U1175 : BUF_X1 port map( A => n4361, Z => n10944);
   U1176 : BUF_X1 port map( A => n2925, Z => n11208);
   U1177 : BUF_X1 port map( A => n4361, Z => n10945);
   U1178 : BUF_X1 port map( A => n2925, Z => n11209);
   U1179 : BUF_X1 port map( A => n4297, Z => n11082);
   U1180 : BUF_X1 port map( A => n4303, Z => n11067);
   U1181 : BUF_X1 port map( A => n2797, Z => n11346);
   U1182 : BUF_X1 port map( A => n2803, Z => n11331);
   U1183 : BUF_X1 port map( A => n4297, Z => n11083);
   U1184 : BUF_X1 port map( A => n4303, Z => n11068);
   U1185 : BUF_X1 port map( A => n2797, Z => n11347);
   U1186 : BUF_X1 port map( A => n2803, Z => n11332);
   U1187 : BUF_X1 port map( A => n4334, Z => n11001);
   U1188 : BUF_X1 port map( A => n2866, Z => n11265);
   U1189 : BUF_X1 port map( A => n4334, Z => n11002);
   U1190 : BUF_X1 port map( A => n2866, Z => n11266);
   U1191 : BUF_X1 port map( A => n4328, Z => n11016);
   U1192 : BUF_X1 port map( A => n4353, Z => n10968);
   U1193 : BUF_X1 port map( A => n4356, Z => n10959);
   U1194 : BUF_X1 port map( A => n4359, Z => n10950);
   U1195 : BUF_X1 port map( A => n4365, Z => n10935);
   U1196 : BUF_X1 port map( A => n2860, Z => n11280);
   U1197 : BUF_X1 port map( A => n2917, Z => n11232);
   U1198 : BUF_X1 port map( A => n2920, Z => n11223);
   U1199 : BUF_X1 port map( A => n2923, Z => n11214);
   U1200 : BUF_X1 port map( A => n2929, Z => n11199);
   U1201 : BUF_X1 port map( A => n4328, Z => n11017);
   U1202 : BUF_X1 port map( A => n4353, Z => n10969);
   U1203 : BUF_X1 port map( A => n4356, Z => n10960);
   U1204 : BUF_X1 port map( A => n4359, Z => n10951);
   U1205 : BUF_X1 port map( A => n4365, Z => n10936);
   U1206 : BUF_X1 port map( A => n2860, Z => n11281);
   U1207 : BUF_X1 port map( A => n2917, Z => n11233);
   U1208 : BUF_X1 port map( A => n2920, Z => n11224);
   U1209 : BUF_X1 port map( A => n2923, Z => n11215);
   U1210 : BUF_X1 port map( A => n2929, Z => n11200);
   U1211 : BUF_X1 port map( A => n4295, Z => n11088);
   U1212 : BUF_X1 port map( A => n4301, Z => n11073);
   U1213 : BUF_X1 port map( A => n2795, Z => n11352);
   U1214 : BUF_X1 port map( A => n2801, Z => n11337);
   U1215 : BUF_X1 port map( A => n4295, Z => n11089);
   U1216 : BUF_X1 port map( A => n4301, Z => n11074);
   U1217 : BUF_X1 port map( A => n2795, Z => n11353);
   U1218 : BUF_X1 port map( A => n2801, Z => n11338);
   U1219 : BUF_X1 port map( A => n4296, Z => n11085);
   U1220 : BUF_X1 port map( A => n4302, Z => n11070);
   U1221 : BUF_X1 port map( A => n2796, Z => n11349);
   U1222 : BUF_X1 port map( A => n2802, Z => n11334);
   U1223 : BUF_X1 port map( A => n4296, Z => n11086);
   U1224 : BUF_X1 port map( A => n4302, Z => n11071);
   U1225 : BUF_X1 port map( A => n2796, Z => n11350);
   U1226 : BUF_X1 port map( A => n2802, Z => n11335);
   U1227 : BUF_X1 port map( A => n4332, Z => n11007);
   U1228 : BUF_X1 port map( A => n2864, Z => n11271);
   U1229 : BUF_X1 port map( A => n4332, Z => n11008);
   U1230 : BUF_X1 port map( A => n2864, Z => n11272);
   U1231 : BUF_X1 port map( A => n4323, Z => n11031);
   U1232 : BUF_X1 port map( A => n4326, Z => n11022);
   U1233 : BUF_X1 port map( A => n4351, Z => n10974);
   U1234 : BUF_X1 port map( A => n4354, Z => n10965);
   U1235 : BUF_X1 port map( A => n4363, Z => n10941);
   U1236 : BUF_X1 port map( A => n2855, Z => n11295);
   U1237 : BUF_X1 port map( A => n2858, Z => n11286);
   U1238 : BUF_X1 port map( A => n2915, Z => n11238);
   U1239 : BUF_X1 port map( A => n2918, Z => n11229);
   U1240 : BUF_X1 port map( A => n2927, Z => n11205);
   U1241 : BUF_X1 port map( A => n4323, Z => n11032);
   U1242 : BUF_X1 port map( A => n4326, Z => n11023);
   U1243 : BUF_X1 port map( A => n4351, Z => n10975);
   U1244 : BUF_X1 port map( A => n4354, Z => n10966);
   U1245 : BUF_X1 port map( A => n4363, Z => n10942);
   U1246 : BUF_X1 port map( A => n2855, Z => n11296);
   U1247 : BUF_X1 port map( A => n2858, Z => n11287);
   U1248 : BUF_X1 port map( A => n2915, Z => n11239);
   U1249 : BUF_X1 port map( A => n2918, Z => n11230);
   U1250 : BUF_X1 port map( A => n2927, Z => n11206);
   U1251 : BUF_X1 port map( A => n4333, Z => n11004);
   U1252 : BUF_X1 port map( A => n2865, Z => n11268);
   U1253 : BUF_X1 port map( A => n4333, Z => n11005);
   U1254 : BUF_X1 port map( A => n2865, Z => n11269);
   U1255 : BUF_X1 port map( A => n4352, Z => n10971);
   U1256 : BUF_X1 port map( A => n4355, Z => n10962);
   U1257 : BUF_X1 port map( A => n4358, Z => n10953);
   U1258 : BUF_X1 port map( A => n2916, Z => n11235);
   U1259 : BUF_X1 port map( A => n2919, Z => n11226);
   U1260 : BUF_X1 port map( A => n2922, Z => n11217);
   U1261 : BUF_X1 port map( A => n4352, Z => n10972);
   U1262 : BUF_X1 port map( A => n4355, Z => n10963);
   U1263 : BUF_X1 port map( A => n4358, Z => n10954);
   U1264 : BUF_X1 port map( A => n2916, Z => n11236);
   U1265 : BUF_X1 port map( A => n2919, Z => n11227);
   U1266 : BUF_X1 port map( A => n2922, Z => n11218);
   U1267 : BUF_X1 port map( A => n4318, Z => n11048);
   U1268 : BUF_X1 port map( A => n2850, Z => n11312);
   U1269 : BUF_X1 port map( A => n4298, Z => n11081);
   U1270 : BUF_X1 port map( A => n2798, Z => n11345);
   U1271 : BUF_X1 port map( A => n4360, Z => n10949);
   U1272 : BUF_X1 port map( A => n2924, Z => n11213);
   U1273 : BUF_X1 port map( A => n4307, Z => n11057);
   U1274 : BUF_X1 port map( A => n2807, Z => n11321);
   U1275 : BUF_X1 port map( A => n4335, Z => n11000);
   U1276 : BUF_X1 port map( A => n4338, Z => n10991);
   U1277 : BUF_X1 port map( A => n2867, Z => n11264);
   U1278 : BUF_X1 port map( A => n2870, Z => n11255);
   U1279 : BUF_X1 port map( A => n4361, Z => n10946);
   U1280 : BUF_X1 port map( A => n2925, Z => n11210);
   U1281 : BUF_X1 port map( A => n4297, Z => n11084);
   U1282 : BUF_X1 port map( A => n4303, Z => n11069);
   U1283 : BUF_X1 port map( A => n2797, Z => n11348);
   U1284 : BUF_X1 port map( A => n2803, Z => n11333);
   U1285 : BUF_X1 port map( A => n4334, Z => n11003);
   U1286 : BUF_X1 port map( A => n2866, Z => n11267);
   U1287 : BUF_X1 port map( A => n4328, Z => n11018);
   U1288 : BUF_X1 port map( A => n4353, Z => n10970);
   U1289 : BUF_X1 port map( A => n4356, Z => n10961);
   U1290 : BUF_X1 port map( A => n4359, Z => n10952);
   U1291 : BUF_X1 port map( A => n4365, Z => n10937);
   U1292 : BUF_X1 port map( A => n2860, Z => n11282);
   U1293 : BUF_X1 port map( A => n2917, Z => n11234);
   U1294 : BUF_X1 port map( A => n2920, Z => n11225);
   U1295 : BUF_X1 port map( A => n2923, Z => n11216);
   U1296 : BUF_X1 port map( A => n2929, Z => n11201);
   U1297 : BUF_X1 port map( A => n4339, Z => n10988);
   U1298 : BUF_X1 port map( A => n2871, Z => n11252);
   U1299 : BUF_X1 port map( A => n4295, Z => n11090);
   U1300 : BUF_X1 port map( A => n4301, Z => n11075);
   U1301 : BUF_X1 port map( A => n2795, Z => n11354);
   U1302 : BUF_X1 port map( A => n2801, Z => n11339);
   U1303 : BUF_X1 port map( A => n4296, Z => n11087);
   U1304 : BUF_X1 port map( A => n4302, Z => n11072);
   U1305 : BUF_X1 port map( A => n2796, Z => n11351);
   U1306 : BUF_X1 port map( A => n2802, Z => n11336);
   U1307 : BUF_X1 port map( A => n4332, Z => n11009);
   U1308 : BUF_X1 port map( A => n2864, Z => n11273);
   U1309 : BUF_X1 port map( A => n4323, Z => n11033);
   U1310 : BUF_X1 port map( A => n4326, Z => n11024);
   U1311 : BUF_X1 port map( A => n4351, Z => n10976);
   U1312 : BUF_X1 port map( A => n4354, Z => n10967);
   U1313 : BUF_X1 port map( A => n4363, Z => n10943);
   U1314 : BUF_X1 port map( A => n2855, Z => n11297);
   U1315 : BUF_X1 port map( A => n2858, Z => n11288);
   U1316 : BUF_X1 port map( A => n2915, Z => n11240);
   U1317 : BUF_X1 port map( A => n2918, Z => n11231);
   U1318 : BUF_X1 port map( A => n2927, Z => n11207);
   U1319 : BUF_X1 port map( A => n4333, Z => n11006);
   U1320 : BUF_X1 port map( A => n2865, Z => n11270);
   U1321 : BUF_X1 port map( A => n4352, Z => n10973);
   U1322 : BUF_X1 port map( A => n4355, Z => n10964);
   U1323 : BUF_X1 port map( A => n4358, Z => n10955);
   U1324 : BUF_X1 port map( A => n2916, Z => n11237);
   U1325 : BUF_X1 port map( A => n2919, Z => n11228);
   U1326 : BUF_X1 port map( A => n2922, Z => n11219);
   U1327 : BUF_X1 port map( A => n4337, Z => n10994);
   U1328 : BUF_X1 port map( A => n4340, Z => n10985);
   U1329 : BUF_X1 port map( A => n2869, Z => n11258);
   U1330 : BUF_X1 port map( A => n2872, Z => n11249);
   U1331 : BUF_X1 port map( A => n2490, Z => n12419);
   U1332 : BUF_X1 port map( A => n2490, Z => n12420);
   U1333 : BUF_X1 port map( A => n2490, Z => n12421);
   U1334 : BUF_X1 port map( A => n2490, Z => n12422);
   U1335 : BUF_X1 port map( A => n2490, Z => n12423);
   U1336 : BUF_X1 port map( A => n2490, Z => n12424);
   U1337 : BUF_X1 port map( A => n2490, Z => n12425);
   U1338 : BUF_X1 port map( A => n12726, Z => n12728);
   U1339 : BUF_X1 port map( A => n12730, Z => n12725);
   U1340 : BUF_X1 port map( A => n12724, Z => n12727);
   U1341 : BUF_X1 port map( A => n12722, Z => n12726);
   U1342 : BUF_X1 port map( A => n12730, Z => n12722);
   U1343 : BUF_X1 port map( A => n12730, Z => n12721);
   U1344 : BUF_X1 port map( A => n12730, Z => n12723);
   U1345 : BUF_X1 port map( A => n12721, Z => n12724);
   U1346 : BUF_X1 port map( A => n12728, Z => n12715);
   U1347 : BUF_X1 port map( A => n12727, Z => n12716);
   U1348 : BUF_X1 port map( A => n12729, Z => n12717);
   U1349 : BUF_X1 port map( A => n12714, Z => n12718);
   U1350 : BUF_X1 port map( A => n12715, Z => n12719);
   U1351 : BUF_X1 port map( A => n12716, Z => n12720);
   U1352 : BUF_X1 port map( A => n12729, Z => n12713);
   U1353 : BUF_X1 port map( A => n12725, Z => n12714);
   U1354 : BUF_X1 port map( A => n12723, Z => n12729);
   U1355 : NOR2_X1 port map( A1 => n12771, A2 => N8436, ZN => n5678);
   U1356 : NOR2_X1 port map( A1 => n12775, A2 => N8580, ZN => n4245);
   U1357 : NOR2_X1 port map( A1 => n12770, A2 => n12771, ZN => n5689);
   U1358 : NOR2_X1 port map( A1 => n12774, A2 => n12775, ZN => n4256);
   U1359 : AND2_X1 port map( A1 => n2571, A2 => n12733, ZN => n2574);
   U1360 : AND3_X1 port map( A1 => n2615, A2 => n12733, A3 => N2172, ZN => 
                           n2617);
   U1361 : AND3_X1 port map( A1 => n12733, A2 => n12732, A3 => n2615, ZN => 
                           n2715);
   U1362 : BUF_X1 port map( A => n4305, Z => n11061);
   U1363 : BUF_X1 port map( A => n4308, Z => n11052);
   U1364 : BUF_X1 port map( A => n4336, Z => n10995);
   U1365 : BUF_X1 port map( A => n4367, Z => n10929);
   U1366 : BUF_X1 port map( A => n4370, Z => n10920);
   U1367 : BUF_X1 port map( A => n4398, Z => n10863);
   U1368 : BUF_X1 port map( A => n4401, Z => n10854);
   U1369 : BUF_X1 port map( A => n2805, Z => n11325);
   U1370 : BUF_X1 port map( A => n2808, Z => n11316);
   U1371 : BUF_X1 port map( A => n2868, Z => n11259);
   U1372 : BUF_X1 port map( A => n2931, Z => n11193);
   U1373 : BUF_X1 port map( A => n2934, Z => n11184);
   U1374 : BUF_X1 port map( A => n2965, Z => n11127);
   U1375 : BUF_X1 port map( A => n2968, Z => n11118);
   U1376 : BUF_X1 port map( A => n4305, Z => n11062);
   U1377 : BUF_X1 port map( A => n4308, Z => n11053);
   U1378 : BUF_X1 port map( A => n4336, Z => n10996);
   U1379 : BUF_X1 port map( A => n4367, Z => n10930);
   U1380 : BUF_X1 port map( A => n4370, Z => n10921);
   U1381 : BUF_X1 port map( A => n4398, Z => n10864);
   U1382 : BUF_X1 port map( A => n4401, Z => n10855);
   U1383 : BUF_X1 port map( A => n2805, Z => n11326);
   U1384 : BUF_X1 port map( A => n2808, Z => n11317);
   U1385 : BUF_X1 port map( A => n2868, Z => n11260);
   U1386 : BUF_X1 port map( A => n2931, Z => n11194);
   U1387 : BUF_X1 port map( A => n2934, Z => n11185);
   U1388 : BUF_X1 port map( A => n2965, Z => n11128);
   U1389 : BUF_X1 port map( A => n2968, Z => n11119);
   U1390 : BUF_X1 port map( A => n4306, Z => n11058);
   U1391 : BUF_X1 port map( A => n4309, Z => n11049);
   U1392 : BUF_X1 port map( A => n4368, Z => n10926);
   U1393 : BUF_X1 port map( A => n4371, Z => n10917);
   U1394 : BUF_X1 port map( A => n4399, Z => n10860);
   U1395 : BUF_X1 port map( A => n4402, Z => n10851);
   U1396 : BUF_X1 port map( A => n2806, Z => n11322);
   U1397 : BUF_X1 port map( A => n2809, Z => n11313);
   U1398 : BUF_X1 port map( A => n2932, Z => n11190);
   U1399 : BUF_X1 port map( A => n2938, Z => n11181);
   U1400 : BUF_X1 port map( A => n2966, Z => n11124);
   U1401 : BUF_X1 port map( A => n2969, Z => n11115);
   U1402 : BUF_X1 port map( A => n4306, Z => n11059);
   U1403 : BUF_X1 port map( A => n4309, Z => n11050);
   U1404 : BUF_X1 port map( A => n4368, Z => n10927);
   U1405 : BUF_X1 port map( A => n4371, Z => n10918);
   U1406 : BUF_X1 port map( A => n4399, Z => n10861);
   U1407 : BUF_X1 port map( A => n4402, Z => n10852);
   U1408 : BUF_X1 port map( A => n2806, Z => n11323);
   U1409 : BUF_X1 port map( A => n2809, Z => n11314);
   U1410 : BUF_X1 port map( A => n2932, Z => n11191);
   U1411 : BUF_X1 port map( A => n2938, Z => n11182);
   U1412 : BUF_X1 port map( A => n2966, Z => n11125);
   U1413 : BUF_X1 port map( A => n2969, Z => n11116);
   U1414 : NAND2_X1 port map( A1 => n5652, A2 => n5655, ZN => n4297);
   U1415 : NAND2_X1 port map( A1 => n5652, A2 => n5657, ZN => n4295);
   U1416 : NAND2_X1 port map( A1 => n5652, A2 => n5656, ZN => n4296);
   U1417 : NAND2_X1 port map( A1 => n5652, A2 => n5659, ZN => n4303);
   U1418 : NAND2_X1 port map( A1 => n5652, A2 => n5661, ZN => n4301);
   U1419 : NAND2_X1 port map( A1 => n5652, A2 => n5660, ZN => n4302);
   U1420 : NAND2_X1 port map( A1 => n4219, A2 => n4222, ZN => n2797);
   U1421 : NAND2_X1 port map( A1 => n4219, A2 => n4224, ZN => n2795);
   U1422 : NAND2_X1 port map( A1 => n4219, A2 => n4223, ZN => n2796);
   U1423 : NAND2_X1 port map( A1 => n4219, A2 => n4226, ZN => n2803);
   U1424 : NAND2_X1 port map( A1 => n4219, A2 => n4228, ZN => n2801);
   U1425 : NAND2_X1 port map( A1 => n4219, A2 => n4227, ZN => n2802);
   U1426 : BUF_X1 port map( A => n4287, Z => n11112);
   U1427 : BUF_X1 port map( A => n4349, Z => n10980);
   U1428 : BUF_X1 port map( A => n4380, Z => n10914);
   U1429 : BUF_X1 port map( A => n2787, Z => n11376);
   U1430 : BUF_X1 port map( A => n2881, Z => n11244);
   U1431 : BUF_X1 port map( A => n2947, Z => n11178);
   U1432 : BUF_X1 port map( A => n4287, Z => n11113);
   U1433 : BUF_X1 port map( A => n4349, Z => n10981);
   U1434 : BUF_X1 port map( A => n4380, Z => n10915);
   U1435 : BUF_X1 port map( A => n2787, Z => n11377);
   U1436 : BUF_X1 port map( A => n2881, Z => n11245);
   U1437 : BUF_X1 port map( A => n2947, Z => n11179);
   U1438 : BUF_X1 port map( A => n4288, Z => n11109);
   U1439 : BUF_X1 port map( A => n4319, Z => n11043);
   U1440 : BUF_X1 port map( A => n4381, Z => n10911);
   U1441 : BUF_X1 port map( A => n2788, Z => n11373);
   U1442 : BUF_X1 port map( A => n2851, Z => n11307);
   U1443 : BUF_X1 port map( A => n2948, Z => n11175);
   U1444 : BUF_X1 port map( A => n4288, Z => n11110);
   U1445 : BUF_X1 port map( A => n4319, Z => n11044);
   U1446 : BUF_X1 port map( A => n4381, Z => n10912);
   U1447 : BUF_X1 port map( A => n2788, Z => n11374);
   U1448 : BUF_X1 port map( A => n2851, Z => n11308);
   U1449 : BUF_X1 port map( A => n2948, Z => n11176);
   U1450 : BUF_X1 port map( A => n4350, Z => n10977);
   U1451 : BUF_X1 port map( A => n2914, Z => n11241);
   U1452 : BUF_X1 port map( A => n4350, Z => n10978);
   U1453 : BUF_X1 port map( A => n2914, Z => n11242);
   U1454 : AND2_X1 port map( A1 => n2730, A2 => n2717, ZN => n2491);
   U1455 : BUF_X1 port map( A => n4329, Z => n11013);
   U1456 : BUF_X1 port map( A => n4391, Z => n10881);
   U1457 : BUF_X1 port map( A => n2861, Z => n11277);
   U1458 : BUF_X1 port map( A => n2958, Z => n11145);
   U1459 : BUF_X1 port map( A => n4329, Z => n11014);
   U1460 : BUF_X1 port map( A => n4391, Z => n10882);
   U1461 : BUF_X1 port map( A => n2861, Z => n11278);
   U1462 : BUF_X1 port map( A => n2958, Z => n11146);
   U1463 : BUF_X1 port map( A => n4304, Z => n11064);
   U1464 : BUF_X1 port map( A => n4366, Z => n10932);
   U1465 : BUF_X1 port map( A => n4369, Z => n10923);
   U1466 : BUF_X1 port map( A => n4397, Z => n10866);
   U1467 : BUF_X1 port map( A => n4400, Z => n10857);
   U1468 : BUF_X1 port map( A => n2804, Z => n11328);
   U1469 : BUF_X1 port map( A => n2930, Z => n11196);
   U1470 : BUF_X1 port map( A => n2933, Z => n11187);
   U1471 : BUF_X1 port map( A => n2964, Z => n11130);
   U1472 : BUF_X1 port map( A => n2967, Z => n11121);
   U1473 : BUF_X1 port map( A => n4304, Z => n11065);
   U1474 : BUF_X1 port map( A => n4366, Z => n10933);
   U1475 : BUF_X1 port map( A => n4369, Z => n10924);
   U1476 : BUF_X1 port map( A => n4397, Z => n10867);
   U1477 : BUF_X1 port map( A => n4400, Z => n10858);
   U1478 : BUF_X1 port map( A => n2804, Z => n11329);
   U1479 : BUF_X1 port map( A => n2930, Z => n11197);
   U1480 : BUF_X1 port map( A => n2933, Z => n11188);
   U1481 : BUF_X1 port map( A => n2964, Z => n11131);
   U1482 : BUF_X1 port map( A => n2967, Z => n11122);
   U1483 : BUF_X1 port map( A => n4299, Z => n11076);
   U1484 : BUF_X1 port map( A => n4330, Z => n11010);
   U1485 : BUF_X1 port map( A => n4392, Z => n10878);
   U1486 : BUF_X1 port map( A => n2799, Z => n11340);
   U1487 : BUF_X1 port map( A => n2862, Z => n11274);
   U1488 : BUF_X1 port map( A => n2959, Z => n11142);
   U1489 : BUF_X1 port map( A => n4299, Z => n11077);
   U1490 : BUF_X1 port map( A => n4330, Z => n11011);
   U1491 : BUF_X1 port map( A => n4392, Z => n10879);
   U1492 : BUF_X1 port map( A => n2799, Z => n11341);
   U1493 : BUF_X1 port map( A => n2862, Z => n11275);
   U1494 : BUF_X1 port map( A => n2959, Z => n11143);
   U1495 : BUF_X1 port map( A => n4390, Z => n10884);
   U1496 : BUF_X1 port map( A => n4396, Z => n10869);
   U1497 : BUF_X1 port map( A => n2957, Z => n11148);
   U1498 : BUF_X1 port map( A => n2963, Z => n11133);
   U1499 : BUF_X1 port map( A => n4390, Z => n10885);
   U1500 : BUF_X1 port map( A => n4396, Z => n10870);
   U1501 : BUF_X1 port map( A => n2957, Z => n11149);
   U1502 : BUF_X1 port map( A => n2963, Z => n11134);
   U1503 : BUF_X1 port map( A => n4291, Z => n11100);
   U1504 : BUF_X1 port map( A => n4322, Z => n11034);
   U1505 : BUF_X1 port map( A => n2791, Z => n11364);
   U1506 : BUF_X1 port map( A => n2854, Z => n11298);
   U1507 : BUF_X1 port map( A => n4291, Z => n11101);
   U1508 : BUF_X1 port map( A => n4322, Z => n11035);
   U1509 : BUF_X1 port map( A => n2791, Z => n11365);
   U1510 : BUF_X1 port map( A => n2854, Z => n11299);
   U1511 : BUF_X1 port map( A => n4294, Z => n11091);
   U1512 : BUF_X1 port map( A => n4325, Z => n11025);
   U1513 : BUF_X1 port map( A => n4384, Z => n10902);
   U1514 : BUF_X1 port map( A => n4387, Z => n10893);
   U1515 : BUF_X1 port map( A => n2794, Z => n11355);
   U1516 : BUF_X1 port map( A => n2857, Z => n11289);
   U1517 : BUF_X1 port map( A => n2951, Z => n11166);
   U1518 : BUF_X1 port map( A => n2954, Z => n11157);
   U1519 : BUF_X1 port map( A => n4294, Z => n11092);
   U1520 : BUF_X1 port map( A => n4325, Z => n11026);
   U1521 : BUF_X1 port map( A => n4384, Z => n10903);
   U1522 : BUF_X1 port map( A => n4387, Z => n10894);
   U1523 : BUF_X1 port map( A => n2794, Z => n11356);
   U1524 : BUF_X1 port map( A => n2857, Z => n11290);
   U1525 : BUF_X1 port map( A => n2951, Z => n11167);
   U1526 : BUF_X1 port map( A => n2954, Z => n11158);
   U1527 : BUF_X1 port map( A => n4385, Z => n10899);
   U1528 : BUF_X1 port map( A => n4388, Z => n10890);
   U1529 : BUF_X1 port map( A => n2952, Z => n11163);
   U1530 : BUF_X1 port map( A => n2955, Z => n11154);
   U1531 : BUF_X1 port map( A => n4385, Z => n10900);
   U1532 : BUF_X1 port map( A => n4388, Z => n10891);
   U1533 : BUF_X1 port map( A => n2952, Z => n11164);
   U1534 : BUF_X1 port map( A => n2955, Z => n11155);
   U1535 : BUF_X1 port map( A => n4386, Z => n10896);
   U1536 : BUF_X1 port map( A => n4395, Z => n10872);
   U1537 : BUF_X1 port map( A => n2953, Z => n11160);
   U1538 : BUF_X1 port map( A => n2962, Z => n11136);
   U1539 : BUF_X1 port map( A => n4386, Z => n10897);
   U1540 : BUF_X1 port map( A => n4395, Z => n10873);
   U1541 : BUF_X1 port map( A => n2953, Z => n11161);
   U1542 : BUF_X1 port map( A => n2962, Z => n11137);
   U1543 : BUF_X1 port map( A => n4389, Z => n10887);
   U1544 : BUF_X1 port map( A => n2956, Z => n11151);
   U1545 : BUF_X1 port map( A => n4389, Z => n10888);
   U1546 : BUF_X1 port map( A => n2956, Z => n11152);
   U1547 : BUF_X1 port map( A => n4289, Z => n11106);
   U1548 : BUF_X1 port map( A => n4357, Z => n10956);
   U1549 : BUF_X1 port map( A => n4394, Z => n10875);
   U1550 : BUF_X1 port map( A => n2789, Z => n11370);
   U1551 : BUF_X1 port map( A => n2921, Z => n11220);
   U1552 : BUF_X1 port map( A => n2961, Z => n11139);
   U1553 : BUF_X1 port map( A => n4289, Z => n11107);
   U1554 : BUF_X1 port map( A => n4357, Z => n10957);
   U1555 : BUF_X1 port map( A => n4394, Z => n10876);
   U1556 : BUF_X1 port map( A => n2789, Z => n11371);
   U1557 : BUF_X1 port map( A => n2921, Z => n11221);
   U1558 : BUF_X1 port map( A => n2961, Z => n11140);
   U1559 : BUF_X1 port map( A => n4292, Z => n11097);
   U1560 : BUF_X1 port map( A => n4320, Z => n11040);
   U1561 : BUF_X1 port map( A => n4382, Z => n10908);
   U1562 : BUF_X1 port map( A => n2792, Z => n11361);
   U1563 : BUF_X1 port map( A => n2852, Z => n11304);
   U1564 : BUF_X1 port map( A => n2949, Z => n11172);
   U1565 : BUF_X1 port map( A => n4292, Z => n11098);
   U1566 : BUF_X1 port map( A => n4320, Z => n11041);
   U1567 : BUF_X1 port map( A => n4382, Z => n10909);
   U1568 : BUF_X1 port map( A => n2792, Z => n11362);
   U1569 : BUF_X1 port map( A => n2852, Z => n11305);
   U1570 : BUF_X1 port map( A => n2949, Z => n11173);
   U1571 : BUF_X1 port map( A => n4321, Z => n11037);
   U1572 : BUF_X1 port map( A => n4364, Z => n10938);
   U1573 : BUF_X1 port map( A => n2853, Z => n11301);
   U1574 : BUF_X1 port map( A => n2928, Z => n11202);
   U1575 : BUF_X1 port map( A => n4321, Z => n11038);
   U1576 : BUF_X1 port map( A => n4364, Z => n10939);
   U1577 : BUF_X1 port map( A => n2853, Z => n11302);
   U1578 : BUF_X1 port map( A => n2928, Z => n11203);
   U1579 : BUF_X1 port map( A => n4290, Z => n11103);
   U1580 : BUF_X1 port map( A => n4293, Z => n11094);
   U1581 : BUF_X1 port map( A => n4324, Z => n11028);
   U1582 : BUF_X1 port map( A => n4327, Z => n11019);
   U1583 : BUF_X1 port map( A => n4383, Z => n10905);
   U1584 : BUF_X1 port map( A => n2790, Z => n11367);
   U1585 : BUF_X1 port map( A => n2793, Z => n11358);
   U1586 : BUF_X1 port map( A => n2856, Z => n11292);
   U1587 : BUF_X1 port map( A => n2859, Z => n11283);
   U1588 : BUF_X1 port map( A => n2950, Z => n11169);
   U1589 : BUF_X1 port map( A => n4290, Z => n11104);
   U1590 : BUF_X1 port map( A => n4293, Z => n11095);
   U1591 : BUF_X1 port map( A => n4324, Z => n11029);
   U1592 : BUF_X1 port map( A => n4327, Z => n11020);
   U1593 : BUF_X1 port map( A => n4383, Z => n10906);
   U1594 : BUF_X1 port map( A => n2790, Z => n11368);
   U1595 : BUF_X1 port map( A => n2793, Z => n11359);
   U1596 : BUF_X1 port map( A => n2856, Z => n11293);
   U1597 : BUF_X1 port map( A => n2859, Z => n11284);
   U1598 : BUF_X1 port map( A => n2950, Z => n11170);
   U1599 : BUF_X1 port map( A => n4287, Z => n11114);
   U1600 : BUF_X1 port map( A => n4349, Z => n10982);
   U1601 : BUF_X1 port map( A => n2787, Z => n11378);
   U1602 : BUF_X1 port map( A => n2881, Z => n11246);
   U1603 : BUF_X1 port map( A => n4380, Z => n10916);
   U1604 : BUF_X1 port map( A => n2947, Z => n11180);
   U1605 : BUF_X1 port map( A => n4288, Z => n11111);
   U1606 : BUF_X1 port map( A => n4319, Z => n11045);
   U1607 : BUF_X1 port map( A => n2788, Z => n11375);
   U1608 : BUF_X1 port map( A => n2851, Z => n11309);
   U1609 : BUF_X1 port map( A => n4381, Z => n10913);
   U1610 : BUF_X1 port map( A => n2948, Z => n11177);
   U1611 : BUF_X1 port map( A => n4350, Z => n10979);
   U1612 : BUF_X1 port map( A => n2914, Z => n11243);
   U1613 : BUF_X1 port map( A => n4391, Z => n10883);
   U1614 : BUF_X1 port map( A => n2958, Z => n11147);
   U1615 : BUF_X1 port map( A => n4329, Z => n11015);
   U1616 : BUF_X1 port map( A => n2861, Z => n11279);
   U1617 : BUF_X1 port map( A => n4304, Z => n11066);
   U1618 : BUF_X1 port map( A => n4366, Z => n10934);
   U1619 : BUF_X1 port map( A => n4369, Z => n10925);
   U1620 : BUF_X1 port map( A => n4397, Z => n10868);
   U1621 : BUF_X1 port map( A => n4400, Z => n10859);
   U1622 : BUF_X1 port map( A => n2804, Z => n11330);
   U1623 : BUF_X1 port map( A => n2930, Z => n11198);
   U1624 : BUF_X1 port map( A => n2933, Z => n11189);
   U1625 : BUF_X1 port map( A => n2964, Z => n11132);
   U1626 : BUF_X1 port map( A => n2967, Z => n11123);
   U1627 : BUF_X1 port map( A => n4299, Z => n11078);
   U1628 : BUF_X1 port map( A => n4330, Z => n11012);
   U1629 : BUF_X1 port map( A => n4392, Z => n10880);
   U1630 : BUF_X1 port map( A => n2799, Z => n11342);
   U1631 : BUF_X1 port map( A => n2862, Z => n11276);
   U1632 : BUF_X1 port map( A => n2959, Z => n11144);
   U1633 : BUF_X1 port map( A => n4390, Z => n10886);
   U1634 : BUF_X1 port map( A => n4396, Z => n10871);
   U1635 : BUF_X1 port map( A => n2957, Z => n11150);
   U1636 : BUF_X1 port map( A => n2963, Z => n11135);
   U1637 : BUF_X1 port map( A => n4291, Z => n11102);
   U1638 : BUF_X1 port map( A => n4322, Z => n11036);
   U1639 : BUF_X1 port map( A => n2791, Z => n11366);
   U1640 : BUF_X1 port map( A => n2854, Z => n11300);
   U1641 : BUF_X1 port map( A => n4294, Z => n11093);
   U1642 : BUF_X1 port map( A => n4325, Z => n11027);
   U1643 : BUF_X1 port map( A => n4384, Z => n10904);
   U1644 : BUF_X1 port map( A => n4387, Z => n10895);
   U1645 : BUF_X1 port map( A => n2794, Z => n11357);
   U1646 : BUF_X1 port map( A => n2857, Z => n11291);
   U1647 : BUF_X1 port map( A => n2951, Z => n11168);
   U1648 : BUF_X1 port map( A => n2954, Z => n11159);
   U1649 : BUF_X1 port map( A => n4305, Z => n11063);
   U1650 : BUF_X1 port map( A => n4308, Z => n11054);
   U1651 : BUF_X1 port map( A => n4336, Z => n10997);
   U1652 : BUF_X1 port map( A => n4367, Z => n10931);
   U1653 : BUF_X1 port map( A => n4370, Z => n10922);
   U1654 : BUF_X1 port map( A => n4398, Z => n10865);
   U1655 : BUF_X1 port map( A => n4401, Z => n10856);
   U1656 : BUF_X1 port map( A => n2805, Z => n11327);
   U1657 : BUF_X1 port map( A => n2808, Z => n11318);
   U1658 : BUF_X1 port map( A => n2868, Z => n11261);
   U1659 : BUF_X1 port map( A => n2931, Z => n11195);
   U1660 : BUF_X1 port map( A => n2934, Z => n11186);
   U1661 : BUF_X1 port map( A => n2965, Z => n11129);
   U1662 : BUF_X1 port map( A => n2968, Z => n11120);
   U1663 : BUF_X1 port map( A => n4385, Z => n10901);
   U1664 : BUF_X1 port map( A => n4388, Z => n10892);
   U1665 : BUF_X1 port map( A => n2952, Z => n11165);
   U1666 : BUF_X1 port map( A => n2955, Z => n11156);
   U1667 : BUF_X1 port map( A => n4386, Z => n10898);
   U1668 : BUF_X1 port map( A => n4395, Z => n10874);
   U1669 : BUF_X1 port map( A => n2953, Z => n11162);
   U1670 : BUF_X1 port map( A => n2962, Z => n11138);
   U1671 : BUF_X1 port map( A => n4389, Z => n10889);
   U1672 : BUF_X1 port map( A => n2956, Z => n11153);
   U1673 : BUF_X1 port map( A => n4357, Z => n10958);
   U1674 : BUF_X1 port map( A => n4394, Z => n10877);
   U1675 : BUF_X1 port map( A => n2921, Z => n11222);
   U1676 : BUF_X1 port map( A => n2961, Z => n11141);
   U1677 : BUF_X1 port map( A => n4289, Z => n11108);
   U1678 : BUF_X1 port map( A => n2789, Z => n11372);
   U1679 : BUF_X1 port map( A => n4292, Z => n11099);
   U1680 : BUF_X1 port map( A => n4320, Z => n11042);
   U1681 : BUF_X1 port map( A => n4382, Z => n10910);
   U1682 : BUF_X1 port map( A => n2792, Z => n11363);
   U1683 : BUF_X1 port map( A => n2852, Z => n11306);
   U1684 : BUF_X1 port map( A => n2949, Z => n11174);
   U1685 : BUF_X1 port map( A => n4364, Z => n10940);
   U1686 : BUF_X1 port map( A => n2928, Z => n11204);
   U1687 : BUF_X1 port map( A => n4321, Z => n11039);
   U1688 : BUF_X1 port map( A => n2853, Z => n11303);
   U1689 : BUF_X1 port map( A => n4290, Z => n11105);
   U1690 : BUF_X1 port map( A => n4293, Z => n11096);
   U1691 : BUF_X1 port map( A => n4324, Z => n11030);
   U1692 : BUF_X1 port map( A => n4327, Z => n11021);
   U1693 : BUF_X1 port map( A => n4383, Z => n10907);
   U1694 : BUF_X1 port map( A => n2790, Z => n11369);
   U1695 : BUF_X1 port map( A => n2793, Z => n11360);
   U1696 : BUF_X1 port map( A => n2856, Z => n11294);
   U1697 : BUF_X1 port map( A => n2859, Z => n11285);
   U1698 : BUF_X1 port map( A => n2950, Z => n11171);
   U1699 : AND2_X1 port map( A1 => n2725, A2 => n2717, ZN => n2582);
   U1700 : BUF_X1 port map( A => n4306, Z => n11060);
   U1701 : BUF_X1 port map( A => n4309, Z => n11051);
   U1702 : BUF_X1 port map( A => n4368, Z => n10928);
   U1703 : BUF_X1 port map( A => n4371, Z => n10919);
   U1704 : BUF_X1 port map( A => n4399, Z => n10862);
   U1705 : BUF_X1 port map( A => n4402, Z => n10853);
   U1706 : BUF_X1 port map( A => n2806, Z => n11324);
   U1707 : BUF_X1 port map( A => n2809, Z => n11315);
   U1708 : BUF_X1 port map( A => n2932, Z => n11192);
   U1709 : BUF_X1 port map( A => n2938, Z => n11183);
   U1710 : BUF_X1 port map( A => n2966, Z => n11126);
   U1711 : BUF_X1 port map( A => n2969, Z => n11117);
   U1712 : NAND2_X1 port map( A1 => n5678, A2 => n5655, ZN => n4334);
   U1713 : NAND2_X1 port map( A1 => n5678, A2 => n5657, ZN => n4332);
   U1714 : NAND2_X1 port map( A1 => n5678, A2 => n5656, ZN => n4333);
   U1715 : NAND2_X1 port map( A1 => n4245, A2 => n4222, ZN => n2866);
   U1716 : NAND2_X1 port map( A1 => n4245, A2 => n4224, ZN => n2864);
   U1717 : NAND2_X1 port map( A1 => n4245, A2 => n4223, ZN => n2865);
   U1718 : NAND2_X1 port map( A1 => n2491, A2 => n2492, ZN => n2490);
   U1719 : AND2_X1 port map( A1 => n5652, A2 => n5653, ZN => n5646);
   U1720 : AND2_X1 port map( A1 => n4219, A2 => n4220, ZN => n4213);
   U1721 : INV_X1 port map( A => N8436, ZN => n12770);
   U1722 : INV_X1 port map( A => N8580, ZN => n12774);
   U1723 : INV_X1 port map( A => N2172, ZN => n12732);
   U1724 : AND2_X1 port map( A1 => n5653, A2 => n5701, ZN => n5690);
   U1725 : AND2_X1 port map( A1 => n4220, A2 => n4268, ZN => n4257);
   U1726 : AND2_X1 port map( A1 => n5675, A2 => n5653, ZN => n5674);
   U1727 : AND2_X1 port map( A1 => n4242, A2 => n4220, ZN => n4241);
   U1728 : NAND2_X1 port map( A1 => n5689, A2 => n5655, ZN => n4353);
   U1729 : NAND2_X1 port map( A1 => n5689, A2 => n5656, ZN => n4351);
   U1730 : NAND2_X1 port map( A1 => n5689, A2 => n5657, ZN => n4352);
   U1731 : NAND2_X1 port map( A1 => n5689, A2 => n5663, ZN => n4356);
   U1732 : NAND2_X1 port map( A1 => n5689, A2 => n5661, ZN => n4354);
   U1733 : NAND2_X1 port map( A1 => n5689, A2 => n5659, ZN => n4355);
   U1734 : NAND2_X1 port map( A1 => n5689, A2 => n5665, ZN => n4359);
   U1735 : NAND2_X1 port map( A1 => n5689, A2 => n5660, ZN => n4358);
   U1736 : NAND2_X1 port map( A1 => n4256, A2 => n4222, ZN => n2917);
   U1737 : NAND2_X1 port map( A1 => n4256, A2 => n4223, ZN => n2915);
   U1738 : NAND2_X1 port map( A1 => n4256, A2 => n4224, ZN => n2916);
   U1739 : NAND2_X1 port map( A1 => n4256, A2 => n4230, ZN => n2920);
   U1740 : NAND2_X1 port map( A1 => n4256, A2 => n4228, ZN => n2918);
   U1741 : NAND2_X1 port map( A1 => n4256, A2 => n4226, ZN => n2919);
   U1742 : NAND2_X1 port map( A1 => n4256, A2 => n4232, ZN => n2923);
   U1743 : NAND2_X1 port map( A1 => n4256, A2 => n4227, ZN => n2922);
   U1744 : NAND2_X1 port map( A1 => n5675, A2 => n5655, ZN => n4323);
   U1745 : NAND2_X1 port map( A1 => n5675, A2 => n5657, ZN => n4328);
   U1746 : NAND2_X1 port map( A1 => n5675, A2 => n5663, ZN => n4326);
   U1747 : NAND2_X1 port map( A1 => n5675, A2 => n5656, ZN => n4318);
   U1748 : NAND2_X1 port map( A1 => n5675, A2 => n5661, ZN => n4365);
   U1749 : NAND2_X1 port map( A1 => n5675, A2 => n5665, ZN => n4363);
   U1750 : NAND2_X1 port map( A1 => n4242, A2 => n4222, ZN => n2855);
   U1751 : NAND2_X1 port map( A1 => n4242, A2 => n4224, ZN => n2860);
   U1752 : NAND2_X1 port map( A1 => n4242, A2 => n4230, ZN => n2858);
   U1753 : NAND2_X1 port map( A1 => n4242, A2 => n4223, ZN => n2850);
   U1754 : NAND2_X1 port map( A1 => n4242, A2 => n4228, ZN => n2929);
   U1755 : NAND2_X1 port map( A1 => n4242, A2 => n4232, ZN => n2927);
   U1756 : AND2_X1 port map( A1 => n5652, A2 => n5665, ZN => n4307);
   U1757 : AND2_X1 port map( A1 => n5652, A2 => n5663, ZN => n4298);
   U1758 : AND2_X1 port map( A1 => n4219, A2 => n4232, ZN => n2807);
   U1759 : AND2_X1 port map( A1 => n4219, A2 => n4230, ZN => n2798);
   U1760 : AND3_X1 port map( A1 => n5653, A2 => n12769, A3 => n5678, ZN => 
                           n5664);
   U1761 : AND3_X1 port map( A1 => n4220, A2 => n12773, A3 => n4245, ZN => 
                           n4231);
   U1762 : AND2_X1 port map( A1 => n5678, A2 => n5661, ZN => n4335);
   U1763 : AND2_X1 port map( A1 => n5678, A2 => n5663, ZN => n4338);
   U1764 : AND2_X1 port map( A1 => n4245, A2 => n4228, ZN => n2867);
   U1765 : AND2_X1 port map( A1 => n4245, A2 => n4230, ZN => n2870);
   U1766 : AND2_X1 port map( A1 => n5689, A2 => n5653, ZN => n5687);
   U1767 : AND2_X1 port map( A1 => n4256, A2 => n4220, ZN => n4254);
   U1768 : AND2_X1 port map( A1 => n5675, A2 => n5660, ZN => n4360);
   U1769 : AND2_X1 port map( A1 => n5675, A2 => n5659, ZN => n4361);
   U1770 : AND2_X1 port map( A1 => n4242, A2 => n4227, ZN => n2924);
   U1771 : AND2_X1 port map( A1 => n4242, A2 => n4226, ZN => n2925);
   U1772 : AND2_X1 port map( A1 => n5678, A2 => n5665, ZN => n4337);
   U1773 : AND2_X1 port map( A1 => n5678, A2 => n5660, ZN => n4339);
   U1774 : AND2_X1 port map( A1 => n5678, A2 => n5659, ZN => n4340);
   U1775 : AND2_X1 port map( A1 => n4245, A2 => n4232, ZN => n2869);
   U1776 : AND2_X1 port map( A1 => n4245, A2 => n4227, ZN => n2871);
   U1777 : AND2_X1 port map( A1 => n4245, A2 => n4226, ZN => n2872);
   U1778 : INV_X1 port map( A => n12432, ZN => n12730);
   U1779 : OAI22_X1 port map( A1 => n10844, A2 => n12293, B1 => n12294, B2 => 
                           n14256, ZN => n8779);
   U1780 : OAI22_X1 port map( A1 => n10837, A2 => n12293, B1 => n12294, B2 => 
                           n14255, ZN => n8778);
   U1781 : OAI22_X1 port map( A1 => n10830, A2 => n12293, B1 => n12294, B2 => 
                           n14254, ZN => n8777);
   U1782 : OAI22_X1 port map( A1 => n10823, A2 => n12293, B1 => n12294, B2 => 
                           n14253, ZN => n8776);
   U1783 : OAI22_X1 port map( A1 => n10816, A2 => n12293, B1 => n12295, B2 => 
                           n14252, ZN => n8775);
   U1784 : OAI22_X1 port map( A1 => n10809, A2 => n12293, B1 => n12295, B2 => 
                           n14251, ZN => n8774);
   U1785 : OAI22_X1 port map( A1 => n10802, A2 => n12293, B1 => n12295, B2 => 
                           n14250, ZN => n8773);
   U1786 : OAI22_X1 port map( A1 => n10795, A2 => n12293, B1 => n12295, B2 => 
                           n14249, ZN => n8772);
   U1787 : OAI22_X1 port map( A1 => n10788, A2 => n12292, B1 => n12296, B2 => 
                           n14248, ZN => n8771);
   U1788 : OAI22_X1 port map( A1 => n10781, A2 => n12292, B1 => n12296, B2 => 
                           n14247, ZN => n8770);
   U1789 : OAI22_X1 port map( A1 => n10774, A2 => n12292, B1 => n12296, B2 => 
                           n14246, ZN => n8769);
   U1790 : OAI22_X1 port map( A1 => n10767, A2 => n12292, B1 => n12296, B2 => 
                           n14245, ZN => n8768);
   U1791 : OAI22_X1 port map( A1 => n10760, A2 => n12292, B1 => n12297, B2 => 
                           n14244, ZN => n8767_port);
   U1792 : OAI22_X1 port map( A1 => n10753, A2 => n12292, B1 => n12297, B2 => 
                           n14243, ZN => n8766_port);
   U1793 : OAI22_X1 port map( A1 => n10746, A2 => n12292, B1 => n12297, B2 => 
                           n14242, ZN => n8765_port);
   U1794 : OAI22_X1 port map( A1 => n10739, A2 => n12292, B1 => n12297, B2 => 
                           n14241, ZN => n8764_port);
   U1795 : OAI22_X1 port map( A1 => n10732, A2 => n12292, B1 => n12298, B2 => 
                           n14240, ZN => n8763_port);
   U1796 : OAI22_X1 port map( A1 => n10725, A2 => n12292, B1 => n12298, B2 => 
                           n14239, ZN => n8762_port);
   U1797 : OAI22_X1 port map( A1 => n10718, A2 => n12292, B1 => n12298, B2 => 
                           n14238, ZN => n8761_port);
   U1798 : OAI22_X1 port map( A1 => n10711, A2 => n12292, B1 => n12298, B2 => 
                           n14237, ZN => n8760_port);
   U1799 : OAI22_X1 port map( A1 => n10704, A2 => n12291, B1 => n12299, B2 => 
                           n14236, ZN => n8759_port);
   U1800 : OAI22_X1 port map( A1 => n10697, A2 => n12291, B1 => n12299, B2 => 
                           n14235, ZN => n8758_port);
   U1801 : OAI22_X1 port map( A1 => n10690, A2 => n12291, B1 => n12299, B2 => 
                           n14234, ZN => n8757_port);
   U1802 : OAI22_X1 port map( A1 => n10683, A2 => n12291, B1 => n12299, B2 => 
                           n14233, ZN => n8756_port);
   U1803 : OAI22_X1 port map( A1 => n10676, A2 => n12291, B1 => n12300, B2 => 
                           n14232, ZN => n8755_port);
   U1804 : OAI22_X1 port map( A1 => n10669, A2 => n12291, B1 => n12300, B2 => 
                           n14231, ZN => n8754_port);
   U1805 : OAI22_X1 port map( A1 => n10662, A2 => n12291, B1 => n12300, B2 => 
                           n14230, ZN => n8753_port);
   U1806 : OAI22_X1 port map( A1 => n10655, A2 => n12291, B1 => n12300, B2 => 
                           n14229, ZN => n8752_port);
   U1807 : OAI22_X1 port map( A1 => n10648, A2 => n12291, B1 => n12301, B2 => 
                           n14228, ZN => n8751_port);
   U1808 : OAI22_X1 port map( A1 => n10641, A2 => n12291, B1 => n12301, B2 => 
                           n14227, ZN => n8750_port);
   U1809 : OAI22_X1 port map( A1 => n10634, A2 => n12291, B1 => n12301, B2 => 
                           n14226, ZN => n8749_port);
   U1810 : OAI22_X1 port map( A1 => n10627, A2 => n12291, B1 => n12301, B2 => 
                           n14225, ZN => n8748_port);
   U1811 : OAI22_X1 port map( A1 => n10845, A2 => n12269, B1 => n12274, B2 => 
                           n14224, ZN => n8715_port);
   U1812 : OAI22_X1 port map( A1 => n10838, A2 => n12269, B1 => n12270, B2 => 
                           n14223, ZN => n8714_port);
   U1813 : OAI22_X1 port map( A1 => n10831, A2 => n12269, B1 => n12270, B2 => 
                           n14222, ZN => n8713_port);
   U1814 : OAI22_X1 port map( A1 => n10824, A2 => n12269, B1 => n12270, B2 => 
                           n14221, ZN => n8712_port);
   U1815 : OAI22_X1 port map( A1 => n10817, A2 => n12269, B1 => n12271, B2 => 
                           n14220, ZN => n8711_port);
   U1816 : OAI22_X1 port map( A1 => n10810, A2 => n12269, B1 => n12271, B2 => 
                           n14219, ZN => n8710_port);
   U1817 : OAI22_X1 port map( A1 => n10803, A2 => n12269, B1 => n12271, B2 => 
                           n14218, ZN => n8709_port);
   U1818 : OAI22_X1 port map( A1 => n10796, A2 => n12269, B1 => n12271, B2 => 
                           n14217, ZN => n8708_port);
   U1819 : OAI22_X1 port map( A1 => n10789, A2 => n12268, B1 => n12272, B2 => 
                           n14216, ZN => n8707_port);
   U1820 : OAI22_X1 port map( A1 => n10782, A2 => n12268, B1 => n12272, B2 => 
                           n14215, ZN => n8706_port);
   U1821 : OAI22_X1 port map( A1 => n10775, A2 => n12268, B1 => n12272, B2 => 
                           n14214, ZN => n8705_port);
   U1822 : OAI22_X1 port map( A1 => n10768, A2 => n12268, B1 => n12272, B2 => 
                           n14213, ZN => n8704_port);
   U1823 : OAI22_X1 port map( A1 => n10761, A2 => n12268, B1 => n12273, B2 => 
                           n14212, ZN => n8703_port);
   U1824 : OAI22_X1 port map( A1 => n10754, A2 => n12268, B1 => n12273, B2 => 
                           n14211, ZN => n8702_port);
   U1825 : OAI22_X1 port map( A1 => n10747, A2 => n12268, B1 => n12273, B2 => 
                           n14210, ZN => n8701);
   U1826 : OAI22_X1 port map( A1 => n10740, A2 => n12268, B1 => n12273, B2 => 
                           n14209, ZN => n8700);
   U1827 : OAI22_X1 port map( A1 => n10733, A2 => n12268, B1 => n12274, B2 => 
                           n14208, ZN => n8699);
   U1828 : OAI22_X1 port map( A1 => n10726, A2 => n12268, B1 => n12274, B2 => 
                           n14207, ZN => n8698);
   U1829 : OAI22_X1 port map( A1 => n10719, A2 => n12268, B1 => n12274, B2 => 
                           n14206, ZN => n8697);
   U1830 : OAI22_X1 port map( A1 => n10712, A2 => n12268, B1 => n12275, B2 => 
                           n14205, ZN => n8696);
   U1831 : OAI22_X1 port map( A1 => n10705, A2 => n12267, B1 => n12275, B2 => 
                           n14204, ZN => n8695);
   U1832 : OAI22_X1 port map( A1 => n10698, A2 => n12267, B1 => n12275, B2 => 
                           n14203, ZN => n8694);
   U1833 : OAI22_X1 port map( A1 => n10691, A2 => n12267, B1 => n12275, B2 => 
                           n14202, ZN => n8693);
   U1834 : OAI22_X1 port map( A1 => n10684, A2 => n12267, B1 => n12276, B2 => 
                           n14201, ZN => n8692);
   U1835 : OAI22_X1 port map( A1 => n10677, A2 => n12267, B1 => n12276, B2 => 
                           n14200, ZN => n8691);
   U1836 : OAI22_X1 port map( A1 => n10670, A2 => n12267, B1 => n12276, B2 => 
                           n14199, ZN => n8690);
   U1837 : OAI22_X1 port map( A1 => n10663, A2 => n12267, B1 => n12276, B2 => 
                           n14198, ZN => n8689);
   U1838 : OAI22_X1 port map( A1 => n10656, A2 => n12267, B1 => n12277, B2 => 
                           n14197, ZN => n8688);
   U1839 : OAI22_X1 port map( A1 => n10649, A2 => n12267, B1 => n12277, B2 => 
                           n14196, ZN => n8687);
   U1840 : OAI22_X1 port map( A1 => n10642, A2 => n12267, B1 => n12277, B2 => 
                           n14195, ZN => n8686);
   U1841 : OAI22_X1 port map( A1 => n10635, A2 => n12267, B1 => n12277, B2 => 
                           n14194, ZN => n8685);
   U1842 : OAI22_X1 port map( A1 => n10845, A2 => n12257, B1 => n12258, B2 => 
                           n14193, ZN => n8683);
   U1843 : OAI22_X1 port map( A1 => n10838, A2 => n12257, B1 => n12258, B2 => 
                           n14192, ZN => n8682);
   U1844 : OAI22_X1 port map( A1 => n10831, A2 => n12257, B1 => n12258, B2 => 
                           n14191, ZN => n8681);
   U1845 : OAI22_X1 port map( A1 => n10824, A2 => n12257, B1 => n12258, B2 => 
                           n14190, ZN => n8680);
   U1846 : OAI22_X1 port map( A1 => n10817, A2 => n12257, B1 => n12259, B2 => 
                           n14189, ZN => n8679);
   U1847 : OAI22_X1 port map( A1 => n10810, A2 => n12257, B1 => n12259, B2 => 
                           n14188, ZN => n8678);
   U1848 : OAI22_X1 port map( A1 => n10803, A2 => n12257, B1 => n12259, B2 => 
                           n14187, ZN => n8677);
   U1849 : OAI22_X1 port map( A1 => n10796, A2 => n12257, B1 => n12259, B2 => 
                           n14186, ZN => n8676);
   U1850 : OAI22_X1 port map( A1 => n10789, A2 => n12256, B1 => n12260, B2 => 
                           n14185, ZN => n8675);
   U1851 : OAI22_X1 port map( A1 => n10782, A2 => n12256, B1 => n12260, B2 => 
                           n14184, ZN => n8674);
   U1852 : OAI22_X1 port map( A1 => n10775, A2 => n12256, B1 => n12260, B2 => 
                           n14183, ZN => n8673);
   U1853 : OAI22_X1 port map( A1 => n10768, A2 => n12256, B1 => n12260, B2 => 
                           n14182, ZN => n8672);
   U1854 : OAI22_X1 port map( A1 => n10761, A2 => n12256, B1 => n12261, B2 => 
                           n14181, ZN => n8671);
   U1855 : OAI22_X1 port map( A1 => n10754, A2 => n12256, B1 => n12261, B2 => 
                           n14180, ZN => n8670);
   U1856 : OAI22_X1 port map( A1 => n10747, A2 => n12256, B1 => n12261, B2 => 
                           n14179, ZN => n8669);
   U1857 : OAI22_X1 port map( A1 => n10740, A2 => n12256, B1 => n12261, B2 => 
                           n14178, ZN => n8668);
   U1858 : OAI22_X1 port map( A1 => n10733, A2 => n12256, B1 => n12262, B2 => 
                           n14177, ZN => n8667);
   U1859 : OAI22_X1 port map( A1 => n10726, A2 => n12256, B1 => n12262, B2 => 
                           n14176, ZN => n8666);
   U1860 : OAI22_X1 port map( A1 => n10719, A2 => n12256, B1 => n12262, B2 => 
                           n14175, ZN => n8665);
   U1861 : OAI22_X1 port map( A1 => n10712, A2 => n12256, B1 => n12262, B2 => 
                           n14174, ZN => n8664);
   U1862 : OAI22_X1 port map( A1 => n10705, A2 => n12255, B1 => n12263, B2 => 
                           n14173, ZN => n8663);
   U1863 : OAI22_X1 port map( A1 => n10698, A2 => n12255, B1 => n12263, B2 => 
                           n14172, ZN => n8662);
   U1864 : OAI22_X1 port map( A1 => n10691, A2 => n12255, B1 => n12263, B2 => 
                           n14171, ZN => n8661);
   U1865 : OAI22_X1 port map( A1 => n10684, A2 => n12255, B1 => n12263, B2 => 
                           n14170, ZN => n8660);
   U1866 : OAI22_X1 port map( A1 => n10677, A2 => n12255, B1 => n12264, B2 => 
                           n14169, ZN => n8659);
   U1867 : OAI22_X1 port map( A1 => n10670, A2 => n12255, B1 => n12264, B2 => 
                           n14168, ZN => n8658);
   U1868 : OAI22_X1 port map( A1 => n10663, A2 => n12255, B1 => n12264, B2 => 
                           n14167, ZN => n8657);
   U1869 : OAI22_X1 port map( A1 => n10656, A2 => n12255, B1 => n12264, B2 => 
                           n14166, ZN => n8656);
   U1870 : OAI22_X1 port map( A1 => n10649, A2 => n12255, B1 => n12265, B2 => 
                           n14165, ZN => n8655);
   U1871 : OAI22_X1 port map( A1 => n10642, A2 => n12255, B1 => n12265, B2 => 
                           n14164, ZN => n8654);
   U1872 : OAI22_X1 port map( A1 => n10635, A2 => n12255, B1 => n12265, B2 => 
                           n14163, ZN => n8653);
   U1873 : OAI22_X1 port map( A1 => n10628, A2 => n12255, B1 => n12265, B2 => 
                           n14162, ZN => n8652);
   U1874 : OAI22_X1 port map( A1 => n10845, A2 => n12245, B1 => n12246, B2 => 
                           n14161, ZN => n8651);
   U1875 : OAI22_X1 port map( A1 => n10838, A2 => n12245, B1 => n12246, B2 => 
                           n14160, ZN => n8650);
   U1876 : OAI22_X1 port map( A1 => n10831, A2 => n12245, B1 => n12246, B2 => 
                           n14159, ZN => n8649);
   U1877 : OAI22_X1 port map( A1 => n10824, A2 => n12245, B1 => n12246, B2 => 
                           n14158, ZN => n8648);
   U1878 : OAI22_X1 port map( A1 => n10817, A2 => n12245, B1 => n12247, B2 => 
                           n14157, ZN => n8647);
   U1879 : OAI22_X1 port map( A1 => n10810, A2 => n12245, B1 => n12247, B2 => 
                           n14156, ZN => n8646);
   U1880 : OAI22_X1 port map( A1 => n10803, A2 => n12245, B1 => n12247, B2 => 
                           n14155, ZN => n8645);
   U1881 : OAI22_X1 port map( A1 => n10796, A2 => n12245, B1 => n12247, B2 => 
                           n14154, ZN => n8644);
   U1882 : OAI22_X1 port map( A1 => n10789, A2 => n12244, B1 => n12248, B2 => 
                           n14153, ZN => n8643);
   U1883 : OAI22_X1 port map( A1 => n10782, A2 => n12244, B1 => n12248, B2 => 
                           n14152, ZN => n8642);
   U1884 : OAI22_X1 port map( A1 => n10775, A2 => n12244, B1 => n12248, B2 => 
                           n14151, ZN => n8641);
   U1885 : OAI22_X1 port map( A1 => n10768, A2 => n12244, B1 => n12248, B2 => 
                           n14150, ZN => n8640);
   U1886 : OAI22_X1 port map( A1 => n10761, A2 => n12244, B1 => n12249, B2 => 
                           n14149, ZN => n8639);
   U1887 : OAI22_X1 port map( A1 => n10754, A2 => n12244, B1 => n12249, B2 => 
                           n14148, ZN => n8638);
   U1888 : OAI22_X1 port map( A1 => n10747, A2 => n12244, B1 => n12249, B2 => 
                           n14147, ZN => n8637);
   U1889 : OAI22_X1 port map( A1 => n10740, A2 => n12244, B1 => n12249, B2 => 
                           n14146, ZN => n8636);
   U1890 : OAI22_X1 port map( A1 => n10733, A2 => n12244, B1 => n12250, B2 => 
                           n14145, ZN => n8635);
   U1891 : OAI22_X1 port map( A1 => n10726, A2 => n12244, B1 => n12250, B2 => 
                           n14144, ZN => n8634);
   U1892 : OAI22_X1 port map( A1 => n10719, A2 => n12244, B1 => n12250, B2 => 
                           n14143, ZN => n8633);
   U1893 : OAI22_X1 port map( A1 => n10712, A2 => n12244, B1 => n12250, B2 => 
                           n14142, ZN => n8632);
   U1894 : OAI22_X1 port map( A1 => n10705, A2 => n12243, B1 => n12251, B2 => 
                           n14141, ZN => n8631);
   U1895 : OAI22_X1 port map( A1 => n10698, A2 => n12243, B1 => n12251, B2 => 
                           n14140, ZN => n8630);
   U1896 : OAI22_X1 port map( A1 => n10691, A2 => n12243, B1 => n12251, B2 => 
                           n14139, ZN => n8629);
   U1897 : OAI22_X1 port map( A1 => n10684, A2 => n12243, B1 => n12251, B2 => 
                           n14138, ZN => n8628);
   U1898 : OAI22_X1 port map( A1 => n10677, A2 => n12243, B1 => n12252, B2 => 
                           n14137, ZN => n8627);
   U1899 : OAI22_X1 port map( A1 => n10670, A2 => n12243, B1 => n12252, B2 => 
                           n14136, ZN => n8626);
   U1900 : OAI22_X1 port map( A1 => n10663, A2 => n12243, B1 => n12252, B2 => 
                           n14135, ZN => n8625);
   U1901 : OAI22_X1 port map( A1 => n10656, A2 => n12243, B1 => n12252, B2 => 
                           n14134, ZN => n8624);
   U1902 : OAI22_X1 port map( A1 => n10649, A2 => n12243, B1 => n12253, B2 => 
                           n14133, ZN => n8623);
   U1903 : OAI22_X1 port map( A1 => n10642, A2 => n12243, B1 => n12253, B2 => 
                           n14132, ZN => n8622);
   U1904 : OAI22_X1 port map( A1 => n10635, A2 => n12243, B1 => n12253, B2 => 
                           n14131, ZN => n8621);
   U1905 : OAI22_X1 port map( A1 => n10628, A2 => n12243, B1 => n12253, B2 => 
                           n14130, ZN => n8620);
   U1906 : OAI22_X1 port map( A1 => n10845, A2 => n12233, B1 => n12238, B2 => 
                           n14129, ZN => n8619);
   U1907 : OAI22_X1 port map( A1 => n10838, A2 => n12233, B1 => n12234, B2 => 
                           n14128, ZN => n8618);
   U1908 : OAI22_X1 port map( A1 => n10831, A2 => n12233, B1 => n12234, B2 => 
                           n14127, ZN => n8617);
   U1909 : OAI22_X1 port map( A1 => n10824, A2 => n12233, B1 => n12234, B2 => 
                           n14126, ZN => n8616);
   U1910 : OAI22_X1 port map( A1 => n10817, A2 => n12233, B1 => n12235, B2 => 
                           n14125, ZN => n8615);
   U1911 : OAI22_X1 port map( A1 => n10810, A2 => n12233, B1 => n12235, B2 => 
                           n14124, ZN => n8614);
   U1912 : OAI22_X1 port map( A1 => n10803, A2 => n12233, B1 => n12235, B2 => 
                           n14123, ZN => n8613);
   U1913 : OAI22_X1 port map( A1 => n10796, A2 => n12233, B1 => n12235, B2 => 
                           n14122, ZN => n8612);
   U1914 : OAI22_X1 port map( A1 => n10789, A2 => n12232, B1 => n12236, B2 => 
                           n14121, ZN => n8611);
   U1915 : OAI22_X1 port map( A1 => n10782, A2 => n12232, B1 => n12236, B2 => 
                           n14120, ZN => n8610);
   U1916 : OAI22_X1 port map( A1 => n10775, A2 => n12232, B1 => n12236, B2 => 
                           n14119, ZN => n8609);
   U1917 : OAI22_X1 port map( A1 => n10768, A2 => n12232, B1 => n12236, B2 => 
                           n14118, ZN => n8608);
   U1918 : OAI22_X1 port map( A1 => n10761, A2 => n12232, B1 => n12237, B2 => 
                           n14117, ZN => n8607);
   U1919 : OAI22_X1 port map( A1 => n10754, A2 => n12232, B1 => n12237, B2 => 
                           n14116, ZN => n8606);
   U1920 : OAI22_X1 port map( A1 => n10747, A2 => n12232, B1 => n12237, B2 => 
                           n14115, ZN => n8605);
   U1921 : OAI22_X1 port map( A1 => n10740, A2 => n12232, B1 => n12237, B2 => 
                           n14114, ZN => n8604);
   U1922 : OAI22_X1 port map( A1 => n10733, A2 => n12232, B1 => n12238, B2 => 
                           n14113, ZN => n8603);
   U1923 : OAI22_X1 port map( A1 => n10726, A2 => n12232, B1 => n12238, B2 => 
                           n14112, ZN => n8602);
   U1924 : OAI22_X1 port map( A1 => n10719, A2 => n12232, B1 => n12238, B2 => 
                           n14111, ZN => n8601);
   U1925 : OAI22_X1 port map( A1 => n10712, A2 => n12232, B1 => n12239, B2 => 
                           n14110, ZN => n8600);
   U1926 : OAI22_X1 port map( A1 => n10705, A2 => n12231, B1 => n12239, B2 => 
                           n14109, ZN => n8599);
   U1927 : OAI22_X1 port map( A1 => n10698, A2 => n12231, B1 => n12239, B2 => 
                           n14108, ZN => n8598);
   U1928 : OAI22_X1 port map( A1 => n10691, A2 => n12231, B1 => n12239, B2 => 
                           n14107, ZN => n8597);
   U1929 : OAI22_X1 port map( A1 => n10684, A2 => n12231, B1 => n12240, B2 => 
                           n14106, ZN => n8596);
   U1930 : OAI22_X1 port map( A1 => n10677, A2 => n12231, B1 => n12240, B2 => 
                           n14105, ZN => n8595);
   U1931 : OAI22_X1 port map( A1 => n10670, A2 => n12231, B1 => n12240, B2 => 
                           n14104, ZN => n8594);
   U1932 : OAI22_X1 port map( A1 => n10663, A2 => n12231, B1 => n12240, B2 => 
                           n14103, ZN => n8593);
   U1933 : OAI22_X1 port map( A1 => n10656, A2 => n12231, B1 => n12241, B2 => 
                           n14102, ZN => n8592);
   U1934 : OAI22_X1 port map( A1 => n10649, A2 => n12231, B1 => n12241, B2 => 
                           n14101, ZN => n8591);
   U1935 : OAI22_X1 port map( A1 => n10642, A2 => n12231, B1 => n12241, B2 => 
                           n14100, ZN => n8590);
   U1936 : OAI22_X1 port map( A1 => n10635, A2 => n12231, B1 => n12241, B2 => 
                           n14099, ZN => n8589);
   U1937 : OAI22_X1 port map( A1 => n10845, A2 => n12221, B1 => n12222, B2 => 
                           n14098, ZN => n8587);
   U1938 : OAI22_X1 port map( A1 => n10838, A2 => n12221, B1 => n12222, B2 => 
                           n14097, ZN => n8586);
   U1939 : OAI22_X1 port map( A1 => n10831, A2 => n12221, B1 => n12222, B2 => 
                           n14096, ZN => n8585);
   U1940 : OAI22_X1 port map( A1 => n10824, A2 => n12221, B1 => n12222, B2 => 
                           n14095, ZN => n8584);
   U1941 : OAI22_X1 port map( A1 => n10817, A2 => n12221, B1 => n12223, B2 => 
                           n14094, ZN => n8583);
   U1942 : OAI22_X1 port map( A1 => n10810, A2 => n12221, B1 => n12223, B2 => 
                           n14093, ZN => n8582);
   U1943 : OAI22_X1 port map( A1 => n10803, A2 => n12221, B1 => n12223, B2 => 
                           n14092, ZN => n8581_port);
   U1944 : OAI22_X1 port map( A1 => n10796, A2 => n12221, B1 => n12223, B2 => 
                           n14091, ZN => n8580_port);
   U1945 : OAI22_X1 port map( A1 => n10789, A2 => n12220, B1 => n12224, B2 => 
                           n14090, ZN => n8579_port);
   U1946 : OAI22_X1 port map( A1 => n10782, A2 => n12220, B1 => n12224, B2 => 
                           n14089, ZN => n8578_port);
   U1947 : OAI22_X1 port map( A1 => n10775, A2 => n12220, B1 => n12224, B2 => 
                           n14088, ZN => n8577);
   U1948 : OAI22_X1 port map( A1 => n10768, A2 => n12220, B1 => n12224, B2 => 
                           n14087, ZN => n8576);
   U1949 : OAI22_X1 port map( A1 => n10761, A2 => n12220, B1 => n12225, B2 => 
                           n14086, ZN => n8575);
   U1950 : OAI22_X1 port map( A1 => n10754, A2 => n12220, B1 => n12225, B2 => 
                           n14085, ZN => n8574);
   U1951 : OAI22_X1 port map( A1 => n10747, A2 => n12220, B1 => n12225, B2 => 
                           n14084, ZN => n8573);
   U1952 : OAI22_X1 port map( A1 => n10740, A2 => n12220, B1 => n12225, B2 => 
                           n14083, ZN => n8572);
   U1953 : OAI22_X1 port map( A1 => n10733, A2 => n12220, B1 => n12226, B2 => 
                           n14082, ZN => n8571);
   U1954 : OAI22_X1 port map( A1 => n10726, A2 => n12220, B1 => n12226, B2 => 
                           n14081, ZN => n8570);
   U1955 : OAI22_X1 port map( A1 => n10719, A2 => n12220, B1 => n12226, B2 => 
                           n14080, ZN => n8569);
   U1956 : OAI22_X1 port map( A1 => n10712, A2 => n12220, B1 => n12226, B2 => 
                           n14079, ZN => n8568);
   U1957 : OAI22_X1 port map( A1 => n10705, A2 => n12219, B1 => n12227, B2 => 
                           n14078, ZN => n8567);
   U1958 : OAI22_X1 port map( A1 => n10698, A2 => n12219, B1 => n12227, B2 => 
                           n14077, ZN => n8566);
   U1959 : OAI22_X1 port map( A1 => n10691, A2 => n12219, B1 => n12227, B2 => 
                           n14076, ZN => n8565);
   U1960 : OAI22_X1 port map( A1 => n10684, A2 => n12219, B1 => n12227, B2 => 
                           n14075, ZN => n8564);
   U1961 : OAI22_X1 port map( A1 => n10677, A2 => n12219, B1 => n12228, B2 => 
                           n14074, ZN => n8563);
   U1962 : OAI22_X1 port map( A1 => n10670, A2 => n12219, B1 => n12228, B2 => 
                           n14073, ZN => n8562);
   U1963 : OAI22_X1 port map( A1 => n10663, A2 => n12219, B1 => n12228, B2 => 
                           n14072, ZN => n8561);
   U1964 : OAI22_X1 port map( A1 => n10656, A2 => n12219, B1 => n12228, B2 => 
                           n14071, ZN => n8560);
   U1965 : OAI22_X1 port map( A1 => n10649, A2 => n12219, B1 => n12229, B2 => 
                           n14070, ZN => n8559);
   U1966 : OAI22_X1 port map( A1 => n10642, A2 => n12219, B1 => n12229, B2 => 
                           n14069, ZN => n8558);
   U1967 : OAI22_X1 port map( A1 => n10635, A2 => n12219, B1 => n12229, B2 => 
                           n14068, ZN => n8557);
   U1968 : OAI22_X1 port map( A1 => n10628, A2 => n12219, B1 => n12229, B2 => 
                           n14067, ZN => n8556);
   U1969 : OAI22_X1 port map( A1 => n10845, A2 => n12209, B1 => n12210, B2 => 
                           n14066, ZN => n8555);
   U1970 : OAI22_X1 port map( A1 => n10838, A2 => n12209, B1 => n12210, B2 => 
                           n14065, ZN => n8554);
   U1971 : OAI22_X1 port map( A1 => n10831, A2 => n12209, B1 => n12210, B2 => 
                           n14064, ZN => n8553);
   U1972 : OAI22_X1 port map( A1 => n10824, A2 => n12209, B1 => n12210, B2 => 
                           n14063, ZN => n8552);
   U1973 : OAI22_X1 port map( A1 => n10817, A2 => n12209, B1 => n12211, B2 => 
                           n14062, ZN => n8551);
   U1974 : OAI22_X1 port map( A1 => n10810, A2 => n12209, B1 => n12211, B2 => 
                           n14061, ZN => n8550);
   U1975 : OAI22_X1 port map( A1 => n10803, A2 => n12209, B1 => n12211, B2 => 
                           n14060, ZN => n8549);
   U1976 : OAI22_X1 port map( A1 => n10796, A2 => n12209, B1 => n12211, B2 => 
                           n14059, ZN => n8548);
   U1977 : OAI22_X1 port map( A1 => n10789, A2 => n12208, B1 => n12212, B2 => 
                           n14058, ZN => n8547);
   U1978 : OAI22_X1 port map( A1 => n10782, A2 => n12208, B1 => n12212, B2 => 
                           n14057, ZN => n8546);
   U1979 : OAI22_X1 port map( A1 => n10775, A2 => n12208, B1 => n12212, B2 => 
                           n14056, ZN => n8545);
   U1980 : OAI22_X1 port map( A1 => n10768, A2 => n12208, B1 => n12212, B2 => 
                           n14055, ZN => n8544);
   U1981 : OAI22_X1 port map( A1 => n10761, A2 => n12208, B1 => n12213, B2 => 
                           n14054, ZN => n8543);
   U1982 : OAI22_X1 port map( A1 => n10754, A2 => n12208, B1 => n12213, B2 => 
                           n14053, ZN => n8542);
   U1983 : OAI22_X1 port map( A1 => n10747, A2 => n12208, B1 => n12213, B2 => 
                           n14052, ZN => n8541);
   U1984 : OAI22_X1 port map( A1 => n10740, A2 => n12208, B1 => n12213, B2 => 
                           n14051, ZN => n8540);
   U1985 : OAI22_X1 port map( A1 => n10733, A2 => n12208, B1 => n12214, B2 => 
                           n14050, ZN => n8539);
   U1986 : OAI22_X1 port map( A1 => n10726, A2 => n12208, B1 => n12214, B2 => 
                           n14049, ZN => n8538);
   U1987 : OAI22_X1 port map( A1 => n10719, A2 => n12208, B1 => n12214, B2 => 
                           n14048, ZN => n8537);
   U1988 : OAI22_X1 port map( A1 => n10712, A2 => n12208, B1 => n12214, B2 => 
                           n14047, ZN => n8536);
   U1989 : OAI22_X1 port map( A1 => n10705, A2 => n12207, B1 => n12215, B2 => 
                           n14046, ZN => n8535);
   U1990 : OAI22_X1 port map( A1 => n10698, A2 => n12207, B1 => n12215, B2 => 
                           n14045, ZN => n8534);
   U1991 : OAI22_X1 port map( A1 => n10691, A2 => n12207, B1 => n12215, B2 => 
                           n14044, ZN => n8533);
   U1992 : OAI22_X1 port map( A1 => n10684, A2 => n12207, B1 => n12215, B2 => 
                           n14043, ZN => n8532);
   U1993 : OAI22_X1 port map( A1 => n10677, A2 => n12207, B1 => n12216, B2 => 
                           n14042, ZN => n8531);
   U1994 : OAI22_X1 port map( A1 => n10670, A2 => n12207, B1 => n12216, B2 => 
                           n14041, ZN => n8530);
   U1995 : OAI22_X1 port map( A1 => n10663, A2 => n12207, B1 => n12216, B2 => 
                           n14040, ZN => n8529);
   U1996 : OAI22_X1 port map( A1 => n10656, A2 => n12207, B1 => n12216, B2 => 
                           n14039, ZN => n8528);
   U1997 : OAI22_X1 port map( A1 => n10649, A2 => n12207, B1 => n12217, B2 => 
                           n14038, ZN => n8527);
   U1998 : OAI22_X1 port map( A1 => n10642, A2 => n12207, B1 => n12217, B2 => 
                           n14037, ZN => n8526);
   U1999 : OAI22_X1 port map( A1 => n10635, A2 => n12207, B1 => n12217, B2 => 
                           n14036, ZN => n8525);
   U2000 : OAI22_X1 port map( A1 => n10628, A2 => n12207, B1 => n12217, B2 => 
                           n14035, ZN => n8524);
   U2001 : OAI22_X1 port map( A1 => n10845, A2 => n12197, B1 => n12202, B2 => 
                           n14034, ZN => n8523);
   U2002 : OAI22_X1 port map( A1 => n10838, A2 => n12197, B1 => n12198, B2 => 
                           n14033, ZN => n8522);
   U2003 : OAI22_X1 port map( A1 => n10831, A2 => n12197, B1 => n12198, B2 => 
                           n14032, ZN => n8521);
   U2004 : OAI22_X1 port map( A1 => n10824, A2 => n12197, B1 => n12198, B2 => 
                           n14031, ZN => n8520);
   U2005 : OAI22_X1 port map( A1 => n10817, A2 => n12197, B1 => n12199, B2 => 
                           n14030, ZN => n8519);
   U2006 : OAI22_X1 port map( A1 => n10810, A2 => n12197, B1 => n12199, B2 => 
                           n14029, ZN => n8518);
   U2007 : OAI22_X1 port map( A1 => n10803, A2 => n12197, B1 => n12199, B2 => 
                           n14028, ZN => n8517);
   U2008 : OAI22_X1 port map( A1 => n10796, A2 => n12197, B1 => n12199, B2 => 
                           n14027, ZN => n8516);
   U2009 : OAI22_X1 port map( A1 => n10789, A2 => n12196, B1 => n12200, B2 => 
                           n14026, ZN => n8515);
   U2010 : OAI22_X1 port map( A1 => n10782, A2 => n12196, B1 => n12200, B2 => 
                           n14025, ZN => n8514);
   U2011 : OAI22_X1 port map( A1 => n10775, A2 => n12196, B1 => n12200, B2 => 
                           n14024, ZN => n8513);
   U2012 : OAI22_X1 port map( A1 => n10768, A2 => n12196, B1 => n12200, B2 => 
                           n14023, ZN => n8512);
   U2013 : OAI22_X1 port map( A1 => n10761, A2 => n12196, B1 => n12201, B2 => 
                           n14022, ZN => n8511);
   U2014 : OAI22_X1 port map( A1 => n10754, A2 => n12196, B1 => n12201, B2 => 
                           n14021, ZN => n8510);
   U2015 : OAI22_X1 port map( A1 => n10747, A2 => n12196, B1 => n12201, B2 => 
                           n14020, ZN => n8509);
   U2016 : OAI22_X1 port map( A1 => n10740, A2 => n12196, B1 => n12201, B2 => 
                           n14019, ZN => n8508);
   U2017 : OAI22_X1 port map( A1 => n10733, A2 => n12196, B1 => n12202, B2 => 
                           n14018, ZN => n8507);
   U2018 : OAI22_X1 port map( A1 => n10726, A2 => n12196, B1 => n12202, B2 => 
                           n14017, ZN => n8506);
   U2019 : OAI22_X1 port map( A1 => n10719, A2 => n12196, B1 => n12202, B2 => 
                           n14016, ZN => n8505);
   U2020 : OAI22_X1 port map( A1 => n10712, A2 => n12196, B1 => n12203, B2 => 
                           n14015, ZN => n8504);
   U2021 : OAI22_X1 port map( A1 => n10705, A2 => n12195, B1 => n12203, B2 => 
                           n14014, ZN => n8503);
   U2022 : OAI22_X1 port map( A1 => n10698, A2 => n12195, B1 => n12203, B2 => 
                           n14013, ZN => n8502);
   U2023 : OAI22_X1 port map( A1 => n10691, A2 => n12195, B1 => n12203, B2 => 
                           n14012, ZN => n8501);
   U2024 : OAI22_X1 port map( A1 => n10684, A2 => n12195, B1 => n12204, B2 => 
                           n14011, ZN => n8500);
   U2025 : OAI22_X1 port map( A1 => n10677, A2 => n12195, B1 => n12204, B2 => 
                           n14010, ZN => n8499);
   U2026 : OAI22_X1 port map( A1 => n10670, A2 => n12195, B1 => n12204, B2 => 
                           n14009, ZN => n8498);
   U2027 : OAI22_X1 port map( A1 => n10663, A2 => n12195, B1 => n12204, B2 => 
                           n14008, ZN => n8497);
   U2028 : OAI22_X1 port map( A1 => n10656, A2 => n12195, B1 => n12205, B2 => 
                           n14007, ZN => n8496);
   U2029 : OAI22_X1 port map( A1 => n10649, A2 => n12195, B1 => n12205, B2 => 
                           n14006, ZN => n8495);
   U2030 : OAI22_X1 port map( A1 => n10642, A2 => n12195, B1 => n12205, B2 => 
                           n14005, ZN => n8494);
   U2031 : OAI22_X1 port map( A1 => n10635, A2 => n12195, B1 => n12205, B2 => 
                           n14004, ZN => n8493);
   U2032 : OAI22_X1 port map( A1 => n10845, A2 => n12185, B1 => n12186, B2 => 
                           n14003, ZN => n8491);
   U2033 : OAI22_X1 port map( A1 => n10838, A2 => n12185, B1 => n12186, B2 => 
                           n14002, ZN => n8490);
   U2034 : OAI22_X1 port map( A1 => n10831, A2 => n12185, B1 => n12186, B2 => 
                           n14001, ZN => n8489);
   U2035 : OAI22_X1 port map( A1 => n10824, A2 => n12185, B1 => n12186, B2 => 
                           n14000, ZN => n8488);
   U2036 : OAI22_X1 port map( A1 => n10817, A2 => n12185, B1 => n12187, B2 => 
                           n13999, ZN => n8487);
   U2037 : OAI22_X1 port map( A1 => n10810, A2 => n12185, B1 => n12187, B2 => 
                           n13998, ZN => n8486);
   U2038 : OAI22_X1 port map( A1 => n10803, A2 => n12185, B1 => n12187, B2 => 
                           n13997, ZN => n8485);
   U2039 : OAI22_X1 port map( A1 => n10796, A2 => n12185, B1 => n12187, B2 => 
                           n13996, ZN => n8484);
   U2040 : OAI22_X1 port map( A1 => n10789, A2 => n12184, B1 => n12188, B2 => 
                           n13995, ZN => n8483);
   U2041 : OAI22_X1 port map( A1 => n10782, A2 => n12184, B1 => n12188, B2 => 
                           n13994, ZN => n8482);
   U2042 : OAI22_X1 port map( A1 => n10775, A2 => n12184, B1 => n12188, B2 => 
                           n13993, ZN => n8481);
   U2043 : OAI22_X1 port map( A1 => n10768, A2 => n12184, B1 => n12188, B2 => 
                           n13992, ZN => n8480);
   U2044 : OAI22_X1 port map( A1 => n10761, A2 => n12184, B1 => n12189, B2 => 
                           n13991, ZN => n8479);
   U2045 : OAI22_X1 port map( A1 => n10754, A2 => n12184, B1 => n12189, B2 => 
                           n13990, ZN => n8478);
   U2046 : OAI22_X1 port map( A1 => n10747, A2 => n12184, B1 => n12189, B2 => 
                           n13989, ZN => n8477);
   U2047 : OAI22_X1 port map( A1 => n10740, A2 => n12184, B1 => n12189, B2 => 
                           n13988, ZN => n8476);
   U2048 : OAI22_X1 port map( A1 => n10733, A2 => n12184, B1 => n12190, B2 => 
                           n13987, ZN => n8475);
   U2049 : OAI22_X1 port map( A1 => n10726, A2 => n12184, B1 => n12190, B2 => 
                           n13986, ZN => n8474);
   U2050 : OAI22_X1 port map( A1 => n10719, A2 => n12184, B1 => n12190, B2 => 
                           n13985, ZN => n8473);
   U2051 : OAI22_X1 port map( A1 => n10712, A2 => n12184, B1 => n12190, B2 => 
                           n13984, ZN => n8472);
   U2052 : OAI22_X1 port map( A1 => n10705, A2 => n12183, B1 => n12191, B2 => 
                           n13983, ZN => n8471);
   U2053 : OAI22_X1 port map( A1 => n10698, A2 => n12183, B1 => n12191, B2 => 
                           n13982, ZN => n8470);
   U2054 : OAI22_X1 port map( A1 => n10691, A2 => n12183, B1 => n12191, B2 => 
                           n13981, ZN => n8469);
   U2055 : OAI22_X1 port map( A1 => n10684, A2 => n12183, B1 => n12191, B2 => 
                           n13980, ZN => n8468);
   U2056 : OAI22_X1 port map( A1 => n10677, A2 => n12183, B1 => n12192, B2 => 
                           n13979, ZN => n8467);
   U2057 : OAI22_X1 port map( A1 => n10670, A2 => n12183, B1 => n12192, B2 => 
                           n13978, ZN => n8466);
   U2058 : OAI22_X1 port map( A1 => n10663, A2 => n12183, B1 => n12192, B2 => 
                           n13977, ZN => n8465);
   U2059 : OAI22_X1 port map( A1 => n10656, A2 => n12183, B1 => n12192, B2 => 
                           n13976, ZN => n8464);
   U2060 : OAI22_X1 port map( A1 => n10649, A2 => n12183, B1 => n12193, B2 => 
                           n13975, ZN => n8463);
   U2061 : OAI22_X1 port map( A1 => n10642, A2 => n12183, B1 => n12193, B2 => 
                           n13974, ZN => n8462);
   U2062 : OAI22_X1 port map( A1 => n10635, A2 => n12183, B1 => n12193, B2 => 
                           n13973, ZN => n8461);
   U2063 : OAI22_X1 port map( A1 => n10628, A2 => n12183, B1 => n12193, B2 => 
                           n13972, ZN => n8460);
   U2064 : OAI22_X1 port map( A1 => n10845, A2 => n12173, B1 => n12174, B2 => 
                           n13971, ZN => n8459);
   U2065 : OAI22_X1 port map( A1 => n10838, A2 => n12173, B1 => n12174, B2 => 
                           n13970, ZN => n8458);
   U2066 : OAI22_X1 port map( A1 => n10831, A2 => n12173, B1 => n12174, B2 => 
                           n13969, ZN => n8457);
   U2067 : OAI22_X1 port map( A1 => n10824, A2 => n12173, B1 => n12174, B2 => 
                           n13968, ZN => n8456);
   U2068 : OAI22_X1 port map( A1 => n10817, A2 => n12173, B1 => n12175, B2 => 
                           n13967, ZN => n8455);
   U2069 : OAI22_X1 port map( A1 => n10810, A2 => n12173, B1 => n12175, B2 => 
                           n13966, ZN => n8454);
   U2070 : OAI22_X1 port map( A1 => n10803, A2 => n12173, B1 => n12175, B2 => 
                           n13965, ZN => n8453);
   U2071 : OAI22_X1 port map( A1 => n10796, A2 => n12173, B1 => n12175, B2 => 
                           n13964, ZN => n8452);
   U2072 : OAI22_X1 port map( A1 => n10789, A2 => n12172, B1 => n12176, B2 => 
                           n13963, ZN => n8451);
   U2073 : OAI22_X1 port map( A1 => n10782, A2 => n12172, B1 => n12176, B2 => 
                           n13962, ZN => n8450);
   U2074 : OAI22_X1 port map( A1 => n10775, A2 => n12172, B1 => n12176, B2 => 
                           n13961, ZN => n8449);
   U2075 : OAI22_X1 port map( A1 => n10768, A2 => n12172, B1 => n12176, B2 => 
                           n13960, ZN => n8448);
   U2076 : OAI22_X1 port map( A1 => n10761, A2 => n12172, B1 => n12177, B2 => 
                           n13959, ZN => n8447);
   U2077 : OAI22_X1 port map( A1 => n10754, A2 => n12172, B1 => n12177, B2 => 
                           n13958, ZN => n8446);
   U2078 : OAI22_X1 port map( A1 => n10747, A2 => n12172, B1 => n12177, B2 => 
                           n13957, ZN => n8445);
   U2079 : OAI22_X1 port map( A1 => n10740, A2 => n12172, B1 => n12177, B2 => 
                           n13956, ZN => n8444);
   U2080 : OAI22_X1 port map( A1 => n10733, A2 => n12172, B1 => n12178, B2 => 
                           n13955, ZN => n8443);
   U2081 : OAI22_X1 port map( A1 => n10726, A2 => n12172, B1 => n12178, B2 => 
                           n13954, ZN => n8442);
   U2082 : OAI22_X1 port map( A1 => n10719, A2 => n12172, B1 => n12178, B2 => 
                           n13953, ZN => n8441);
   U2083 : OAI22_X1 port map( A1 => n10712, A2 => n12172, B1 => n12178, B2 => 
                           n13952, ZN => n8440);
   U2084 : OAI22_X1 port map( A1 => n10705, A2 => n12171, B1 => n12179, B2 => 
                           n13951, ZN => n8439);
   U2085 : OAI22_X1 port map( A1 => n10698, A2 => n12171, B1 => n12179, B2 => 
                           n13950, ZN => n8438);
   U2086 : OAI22_X1 port map( A1 => n10691, A2 => n12171, B1 => n12179, B2 => 
                           n13949, ZN => n8437_port);
   U2087 : OAI22_X1 port map( A1 => n10684, A2 => n12171, B1 => n12179, B2 => 
                           n13948, ZN => n8436_port);
   U2088 : OAI22_X1 port map( A1 => n10677, A2 => n12171, B1 => n12180, B2 => 
                           n13947, ZN => n8435_port);
   U2089 : OAI22_X1 port map( A1 => n10670, A2 => n12171, B1 => n12180, B2 => 
                           n13946, ZN => n8434_port);
   U2090 : OAI22_X1 port map( A1 => n10663, A2 => n12171, B1 => n12180, B2 => 
                           n13945, ZN => n8433);
   U2091 : OAI22_X1 port map( A1 => n10656, A2 => n12171, B1 => n12180, B2 => 
                           n13944, ZN => n8432);
   U2092 : OAI22_X1 port map( A1 => n10649, A2 => n12171, B1 => n12181, B2 => 
                           n13943, ZN => n8431);
   U2093 : OAI22_X1 port map( A1 => n10642, A2 => n12171, B1 => n12181, B2 => 
                           n13942, ZN => n8430);
   U2094 : OAI22_X1 port map( A1 => n10635, A2 => n12171, B1 => n12181, B2 => 
                           n13941, ZN => n8429);
   U2095 : OAI22_X1 port map( A1 => n10628, A2 => n12171, B1 => n12181, B2 => 
                           n13940, ZN => n8428);
   U2096 : OAI22_X1 port map( A1 => n10845, A2 => n12161, B1 => n12162, B2 => 
                           n13939, ZN => n8427);
   U2097 : OAI22_X1 port map( A1 => n10838, A2 => n12161, B1 => n12162, B2 => 
                           n13938, ZN => n8426);
   U2098 : OAI22_X1 port map( A1 => n10831, A2 => n12161, B1 => n12162, B2 => 
                           n13937, ZN => n8425);
   U2099 : OAI22_X1 port map( A1 => n10824, A2 => n12161, B1 => n12162, B2 => 
                           n13936, ZN => n8424);
   U2100 : OAI22_X1 port map( A1 => n10817, A2 => n12161, B1 => n12163, B2 => 
                           n13935, ZN => n8423);
   U2101 : OAI22_X1 port map( A1 => n10810, A2 => n12161, B1 => n12163, B2 => 
                           n13934, ZN => n8422);
   U2102 : OAI22_X1 port map( A1 => n10803, A2 => n12161, B1 => n12163, B2 => 
                           n13933, ZN => n8421);
   U2103 : OAI22_X1 port map( A1 => n10796, A2 => n12161, B1 => n12163, B2 => 
                           n13932, ZN => n8420);
   U2104 : OAI22_X1 port map( A1 => n10789, A2 => n12160, B1 => n12164, B2 => 
                           n13931, ZN => n8419);
   U2105 : OAI22_X1 port map( A1 => n10782, A2 => n12160, B1 => n12164, B2 => 
                           n13930, ZN => n8418);
   U2106 : OAI22_X1 port map( A1 => n10775, A2 => n12160, B1 => n12164, B2 => 
                           n13929, ZN => n8417);
   U2107 : OAI22_X1 port map( A1 => n10768, A2 => n12160, B1 => n12164, B2 => 
                           n13928, ZN => n8416);
   U2108 : OAI22_X1 port map( A1 => n10761, A2 => n12160, B1 => n12165, B2 => 
                           n13927, ZN => n8415);
   U2109 : OAI22_X1 port map( A1 => n10754, A2 => n12160, B1 => n12165, B2 => 
                           n13926, ZN => n8414);
   U2110 : OAI22_X1 port map( A1 => n10747, A2 => n12160, B1 => n12165, B2 => 
                           n13925, ZN => n8413);
   U2111 : OAI22_X1 port map( A1 => n10740, A2 => n12160, B1 => n12165, B2 => 
                           n13924, ZN => n8412);
   U2112 : OAI22_X1 port map( A1 => n10733, A2 => n12160, B1 => n12166, B2 => 
                           n13923, ZN => n8411);
   U2113 : OAI22_X1 port map( A1 => n10726, A2 => n12160, B1 => n12166, B2 => 
                           n13922, ZN => n8410);
   U2114 : OAI22_X1 port map( A1 => n10719, A2 => n12160, B1 => n12166, B2 => 
                           n13921, ZN => n8409);
   U2115 : OAI22_X1 port map( A1 => n10712, A2 => n12160, B1 => n12166, B2 => 
                           n13920, ZN => n8408);
   U2116 : OAI22_X1 port map( A1 => n10705, A2 => n12159, B1 => n12167, B2 => 
                           n13919, ZN => n8407);
   U2117 : OAI22_X1 port map( A1 => n10698, A2 => n12159, B1 => n12167, B2 => 
                           n13918, ZN => n8406);
   U2118 : OAI22_X1 port map( A1 => n10691, A2 => n12159, B1 => n12167, B2 => 
                           n13917, ZN => n8405);
   U2119 : OAI22_X1 port map( A1 => n10684, A2 => n12159, B1 => n12167, B2 => 
                           n13916, ZN => n8404);
   U2120 : OAI22_X1 port map( A1 => n10677, A2 => n12159, B1 => n12168, B2 => 
                           n13915, ZN => n8403);
   U2121 : OAI22_X1 port map( A1 => n10670, A2 => n12159, B1 => n12168, B2 => 
                           n13914, ZN => n8402);
   U2122 : OAI22_X1 port map( A1 => n10663, A2 => n12159, B1 => n12168, B2 => 
                           n13913, ZN => n8401);
   U2123 : OAI22_X1 port map( A1 => n10656, A2 => n12159, B1 => n12168, B2 => 
                           n13912, ZN => n8400);
   U2124 : OAI22_X1 port map( A1 => n10649, A2 => n12159, B1 => n12169, B2 => 
                           n13911, ZN => n8399);
   U2125 : OAI22_X1 port map( A1 => n10642, A2 => n12159, B1 => n12169, B2 => 
                           n13910, ZN => n8398);
   U2126 : OAI22_X1 port map( A1 => n10635, A2 => n12159, B1 => n12169, B2 => 
                           n13909, ZN => n8397);
   U2127 : OAI22_X1 port map( A1 => n10628, A2 => n12159, B1 => n12169, B2 => 
                           n13908, ZN => n8396);
   U2128 : OAI22_X1 port map( A1 => n10845, A2 => n12137, B1 => n12138, B2 => 
                           n13907, ZN => n8363);
   U2129 : OAI22_X1 port map( A1 => n10838, A2 => n12137, B1 => n12138, B2 => 
                           n13906, ZN => n8362);
   U2130 : OAI22_X1 port map( A1 => n10831, A2 => n12137, B1 => n12138, B2 => 
                           n13905, ZN => n8361);
   U2131 : OAI22_X1 port map( A1 => n10824, A2 => n12137, B1 => n12138, B2 => 
                           n13904, ZN => n8360);
   U2132 : OAI22_X1 port map( A1 => n10817, A2 => n12137, B1 => n12139, B2 => 
                           n13903, ZN => n8359);
   U2133 : OAI22_X1 port map( A1 => n10810, A2 => n12137, B1 => n12139, B2 => 
                           n13902, ZN => n8358);
   U2134 : OAI22_X1 port map( A1 => n10803, A2 => n12137, B1 => n12139, B2 => 
                           n13901, ZN => n8357);
   U2135 : OAI22_X1 port map( A1 => n10796, A2 => n12137, B1 => n12139, B2 => 
                           n13900, ZN => n8356);
   U2136 : OAI22_X1 port map( A1 => n10789, A2 => n12136, B1 => n12140, B2 => 
                           n13899, ZN => n8355);
   U2137 : OAI22_X1 port map( A1 => n10782, A2 => n12136, B1 => n12140, B2 => 
                           n13898, ZN => n8354);
   U2138 : OAI22_X1 port map( A1 => n10775, A2 => n12136, B1 => n12140, B2 => 
                           n13897, ZN => n8353);
   U2139 : OAI22_X1 port map( A1 => n10768, A2 => n12136, B1 => n12140, B2 => 
                           n13896, ZN => n8352);
   U2140 : OAI22_X1 port map( A1 => n10761, A2 => n12136, B1 => n12141, B2 => 
                           n13895, ZN => n8351);
   U2141 : OAI22_X1 port map( A1 => n10754, A2 => n12136, B1 => n12141, B2 => 
                           n13894, ZN => n8350);
   U2142 : OAI22_X1 port map( A1 => n10747, A2 => n12136, B1 => n12141, B2 => 
                           n13893, ZN => n8349);
   U2143 : OAI22_X1 port map( A1 => n10740, A2 => n12136, B1 => n12141, B2 => 
                           n13892, ZN => n8348);
   U2144 : OAI22_X1 port map( A1 => n10733, A2 => n12136, B1 => n12142, B2 => 
                           n13891, ZN => n8347);
   U2145 : OAI22_X1 port map( A1 => n10726, A2 => n12136, B1 => n12142, B2 => 
                           n13890, ZN => n8346);
   U2146 : OAI22_X1 port map( A1 => n10719, A2 => n12136, B1 => n12142, B2 => 
                           n13889, ZN => n8345);
   U2147 : OAI22_X1 port map( A1 => n10712, A2 => n12136, B1 => n12142, B2 => 
                           n13888, ZN => n8344);
   U2148 : OAI22_X1 port map( A1 => n10705, A2 => n12135, B1 => n12143, B2 => 
                           n13887, ZN => n8343);
   U2149 : OAI22_X1 port map( A1 => n10698, A2 => n12135, B1 => n12143, B2 => 
                           n13886, ZN => n8342);
   U2150 : OAI22_X1 port map( A1 => n10691, A2 => n12135, B1 => n12143, B2 => 
                           n13885, ZN => n8341);
   U2151 : OAI22_X1 port map( A1 => n10684, A2 => n12135, B1 => n12143, B2 => 
                           n13884, ZN => n8340);
   U2152 : OAI22_X1 port map( A1 => n10677, A2 => n12135, B1 => n12144, B2 => 
                           n13883, ZN => n8339);
   U2153 : OAI22_X1 port map( A1 => n10670, A2 => n12135, B1 => n12144, B2 => 
                           n13882, ZN => n8338);
   U2154 : OAI22_X1 port map( A1 => n10663, A2 => n12135, B1 => n12144, B2 => 
                           n13881, ZN => n8337);
   U2155 : OAI22_X1 port map( A1 => n10656, A2 => n12135, B1 => n12144, B2 => 
                           n13880, ZN => n8336);
   U2156 : OAI22_X1 port map( A1 => n10649, A2 => n12135, B1 => n12145, B2 => 
                           n13879, ZN => n8335);
   U2157 : OAI22_X1 port map( A1 => n10642, A2 => n12135, B1 => n12145, B2 => 
                           n13878, ZN => n8334);
   U2158 : OAI22_X1 port map( A1 => n10635, A2 => n12135, B1 => n12145, B2 => 
                           n13877, ZN => n8333);
   U2159 : OAI22_X1 port map( A1 => n10628, A2 => n12135, B1 => n12145, B2 => 
                           n13876, ZN => n8332);
   U2160 : OAI22_X1 port map( A1 => n10846, A2 => n12113, B1 => n12114, B2 => 
                           n13875, ZN => n8299);
   U2161 : OAI22_X1 port map( A1 => n10839, A2 => n12113, B1 => n12114, B2 => 
                           n13874, ZN => n8298);
   U2162 : OAI22_X1 port map( A1 => n10832, A2 => n12113, B1 => n12114, B2 => 
                           n13873, ZN => n8297);
   U2163 : OAI22_X1 port map( A1 => n10825, A2 => n12113, B1 => n12114, B2 => 
                           n13872, ZN => n8296);
   U2164 : OAI22_X1 port map( A1 => n10818, A2 => n12113, B1 => n12115, B2 => 
                           n13871, ZN => n8295);
   U2165 : OAI22_X1 port map( A1 => n10811, A2 => n12113, B1 => n12115, B2 => 
                           n13870, ZN => n8294);
   U2166 : OAI22_X1 port map( A1 => n10804, A2 => n12113, B1 => n12115, B2 => 
                           n13869, ZN => n8293);
   U2167 : OAI22_X1 port map( A1 => n10797, A2 => n12113, B1 => n12115, B2 => 
                           n13868, ZN => n8292);
   U2168 : OAI22_X1 port map( A1 => n10790, A2 => n12112, B1 => n12116, B2 => 
                           n13867, ZN => n8291);
   U2169 : OAI22_X1 port map( A1 => n10783, A2 => n12112, B1 => n12116, B2 => 
                           n13866, ZN => n8290);
   U2170 : OAI22_X1 port map( A1 => n10776, A2 => n12112, B1 => n12116, B2 => 
                           n13865, ZN => n8289);
   U2171 : OAI22_X1 port map( A1 => n10769, A2 => n12112, B1 => n12116, B2 => 
                           n13864, ZN => n8288);
   U2172 : OAI22_X1 port map( A1 => n10762, A2 => n12112, B1 => n12117, B2 => 
                           n13863, ZN => n8287);
   U2173 : OAI22_X1 port map( A1 => n10755, A2 => n12112, B1 => n12117, B2 => 
                           n13862, ZN => n8286);
   U2174 : OAI22_X1 port map( A1 => n10748, A2 => n12112, B1 => n12117, B2 => 
                           n13861, ZN => n8285);
   U2175 : OAI22_X1 port map( A1 => n10741, A2 => n12112, B1 => n12117, B2 => 
                           n13860, ZN => n8284);
   U2176 : OAI22_X1 port map( A1 => n10734, A2 => n12112, B1 => n12118, B2 => 
                           n13859, ZN => n8283);
   U2177 : OAI22_X1 port map( A1 => n10727, A2 => n12112, B1 => n12118, B2 => 
                           n13858, ZN => n8282);
   U2178 : OAI22_X1 port map( A1 => n10720, A2 => n12112, B1 => n12118, B2 => 
                           n13857, ZN => n8281);
   U2179 : OAI22_X1 port map( A1 => n10713, A2 => n12112, B1 => n12118, B2 => 
                           n13856, ZN => n8280);
   U2180 : OAI22_X1 port map( A1 => n10706, A2 => n12111, B1 => n12119, B2 => 
                           n13855, ZN => n8279);
   U2181 : OAI22_X1 port map( A1 => n10699, A2 => n12111, B1 => n12119, B2 => 
                           n13854, ZN => n8278);
   U2182 : OAI22_X1 port map( A1 => n10692, A2 => n12111, B1 => n12119, B2 => 
                           n13853, ZN => n8277);
   U2183 : OAI22_X1 port map( A1 => n10685, A2 => n12111, B1 => n12119, B2 => 
                           n13852, ZN => n8276);
   U2184 : OAI22_X1 port map( A1 => n10678, A2 => n12111, B1 => n12120, B2 => 
                           n13851, ZN => n8275);
   U2185 : OAI22_X1 port map( A1 => n10671, A2 => n12111, B1 => n12120, B2 => 
                           n13850, ZN => n8274);
   U2186 : OAI22_X1 port map( A1 => n10664, A2 => n12111, B1 => n12120, B2 => 
                           n13849, ZN => n8273);
   U2187 : OAI22_X1 port map( A1 => n10657, A2 => n12111, B1 => n12120, B2 => 
                           n13848, ZN => n8272);
   U2188 : OAI22_X1 port map( A1 => n10650, A2 => n12111, B1 => n12121, B2 => 
                           n13847, ZN => n8271);
   U2189 : OAI22_X1 port map( A1 => n10643, A2 => n12111, B1 => n12121, B2 => 
                           n13846, ZN => n8270);
   U2190 : OAI22_X1 port map( A1 => n10636, A2 => n12111, B1 => n12121, B2 => 
                           n13845, ZN => n8269);
   U2191 : OAI22_X1 port map( A1 => n10629, A2 => n12111, B1 => n12121, B2 => 
                           n13844, ZN => n8268);
   U2192 : OAI22_X1 port map( A1 => n10847, A2 => n11957, B1 => n11958, B2 => 
                           n13651, ZN => n7883);
   U2193 : OAI22_X1 port map( A1 => n10840, A2 => n11957, B1 => n11958, B2 => 
                           n13650, ZN => n7882);
   U2194 : OAI22_X1 port map( A1 => n10833, A2 => n11957, B1 => n11958, B2 => 
                           n13649, ZN => n7881);
   U2195 : OAI22_X1 port map( A1 => n10826, A2 => n11957, B1 => n11958, B2 => 
                           n13648, ZN => n7880);
   U2196 : OAI22_X1 port map( A1 => n10819, A2 => n11957, B1 => n11959, B2 => 
                           n13647, ZN => n7879);
   U2197 : OAI22_X1 port map( A1 => n10812, A2 => n11957, B1 => n11959, B2 => 
                           n13646, ZN => n7878);
   U2198 : OAI22_X1 port map( A1 => n10805, A2 => n11957, B1 => n11959, B2 => 
                           n13645, ZN => n7877);
   U2199 : OAI22_X1 port map( A1 => n10798, A2 => n11957, B1 => n11959, B2 => 
                           n13644, ZN => n7876);
   U2200 : OAI22_X1 port map( A1 => n10791, A2 => n11956, B1 => n11960, B2 => 
                           n13643, ZN => n7875);
   U2201 : OAI22_X1 port map( A1 => n10784, A2 => n11956, B1 => n11960, B2 => 
                           n13642, ZN => n7874);
   U2202 : OAI22_X1 port map( A1 => n10777, A2 => n11956, B1 => n11960, B2 => 
                           n13641, ZN => n7873);
   U2203 : OAI22_X1 port map( A1 => n10770, A2 => n11956, B1 => n11960, B2 => 
                           n13640, ZN => n7872);
   U2204 : OAI22_X1 port map( A1 => n10763, A2 => n11956, B1 => n11961, B2 => 
                           n13639, ZN => n7871);
   U2205 : OAI22_X1 port map( A1 => n10756, A2 => n11956, B1 => n11961, B2 => 
                           n13638, ZN => n7870);
   U2206 : OAI22_X1 port map( A1 => n10749, A2 => n11956, B1 => n11961, B2 => 
                           n13637, ZN => n7869);
   U2207 : OAI22_X1 port map( A1 => n10742, A2 => n11956, B1 => n11961, B2 => 
                           n13636, ZN => n7868);
   U2208 : OAI22_X1 port map( A1 => n10735, A2 => n11956, B1 => n11962, B2 => 
                           n13635, ZN => n7867);
   U2209 : OAI22_X1 port map( A1 => n10728, A2 => n11956, B1 => n11962, B2 => 
                           n13634, ZN => n7866);
   U2210 : OAI22_X1 port map( A1 => n10721, A2 => n11956, B1 => n11962, B2 => 
                           n13633, ZN => n7865);
   U2211 : OAI22_X1 port map( A1 => n10714, A2 => n11956, B1 => n11962, B2 => 
                           n13632, ZN => n7864);
   U2212 : OAI22_X1 port map( A1 => n10707, A2 => n11955, B1 => n11963, B2 => 
                           n13631, ZN => n7863);
   U2213 : OAI22_X1 port map( A1 => n10700, A2 => n11955, B1 => n11963, B2 => 
                           n13630, ZN => n7862);
   U2214 : OAI22_X1 port map( A1 => n10693, A2 => n11955, B1 => n11963, B2 => 
                           n13629, ZN => n7861);
   U2215 : OAI22_X1 port map( A1 => n10686, A2 => n11955, B1 => n11963, B2 => 
                           n13628, ZN => n7860);
   U2216 : OAI22_X1 port map( A1 => n10679, A2 => n11955, B1 => n11964, B2 => 
                           n13627, ZN => n7859);
   U2217 : OAI22_X1 port map( A1 => n10672, A2 => n11955, B1 => n11964, B2 => 
                           n13626, ZN => n7858);
   U2218 : OAI22_X1 port map( A1 => n10665, A2 => n11955, B1 => n11964, B2 => 
                           n13625, ZN => n7857);
   U2219 : OAI22_X1 port map( A1 => n10658, A2 => n11955, B1 => n11964, B2 => 
                           n13624, ZN => n7856);
   U2220 : OAI22_X1 port map( A1 => n10651, A2 => n11955, B1 => n11965, B2 => 
                           n13623, ZN => n7855);
   U2221 : OAI22_X1 port map( A1 => n10644, A2 => n11955, B1 => n11965, B2 => 
                           n13622, ZN => n7854);
   U2222 : OAI22_X1 port map( A1 => n10637, A2 => n11955, B1 => n11965, B2 => 
                           n13621, ZN => n7853);
   U2223 : OAI22_X1 port map( A1 => n10630, A2 => n11955, B1 => n11965, B2 => 
                           n13620, ZN => n7852);
   U2224 : OAI22_X1 port map( A1 => n10847, A2 => n11945, B1 => n11946, B2 => 
                           n13619, ZN => n7851);
   U2225 : OAI22_X1 port map( A1 => n10840, A2 => n11945, B1 => n11946, B2 => 
                           n13618, ZN => n7850);
   U2226 : OAI22_X1 port map( A1 => n10833, A2 => n11945, B1 => n11946, B2 => 
                           n13617, ZN => n7849);
   U2227 : OAI22_X1 port map( A1 => n10826, A2 => n11945, B1 => n11946, B2 => 
                           n13616, ZN => n7848);
   U2228 : OAI22_X1 port map( A1 => n10819, A2 => n11945, B1 => n11947, B2 => 
                           n13615, ZN => n7847);
   U2229 : OAI22_X1 port map( A1 => n10812, A2 => n11945, B1 => n11947, B2 => 
                           n13614, ZN => n7846);
   U2230 : OAI22_X1 port map( A1 => n10805, A2 => n11945, B1 => n11947, B2 => 
                           n13613, ZN => n7845);
   U2231 : OAI22_X1 port map( A1 => n10798, A2 => n11945, B1 => n11947, B2 => 
                           n13612, ZN => n7844);
   U2232 : OAI22_X1 port map( A1 => n10791, A2 => n11944, B1 => n11948, B2 => 
                           n13611, ZN => n7843);
   U2233 : OAI22_X1 port map( A1 => n10784, A2 => n11944, B1 => n11948, B2 => 
                           n13610, ZN => n7842);
   U2234 : OAI22_X1 port map( A1 => n10777, A2 => n11944, B1 => n11948, B2 => 
                           n13609, ZN => n7841);
   U2235 : OAI22_X1 port map( A1 => n10770, A2 => n11944, B1 => n11948, B2 => 
                           n13608, ZN => n7840);
   U2236 : OAI22_X1 port map( A1 => n10763, A2 => n11944, B1 => n11949, B2 => 
                           n13607, ZN => n7839);
   U2237 : OAI22_X1 port map( A1 => n10756, A2 => n11944, B1 => n11949, B2 => 
                           n13606, ZN => n7838);
   U2238 : OAI22_X1 port map( A1 => n10749, A2 => n11944, B1 => n11949, B2 => 
                           n13605, ZN => n7837);
   U2239 : OAI22_X1 port map( A1 => n10742, A2 => n11944, B1 => n11949, B2 => 
                           n13604, ZN => n7836);
   U2240 : OAI22_X1 port map( A1 => n10735, A2 => n11944, B1 => n11950, B2 => 
                           n13603, ZN => n7835);
   U2241 : OAI22_X1 port map( A1 => n10728, A2 => n11944, B1 => n11950, B2 => 
                           n13602, ZN => n7834);
   U2242 : OAI22_X1 port map( A1 => n10721, A2 => n11944, B1 => n11950, B2 => 
                           n13601, ZN => n7833);
   U2243 : OAI22_X1 port map( A1 => n10714, A2 => n11944, B1 => n11950, B2 => 
                           n13600, ZN => n7832);
   U2244 : OAI22_X1 port map( A1 => n10707, A2 => n11943, B1 => n11951, B2 => 
                           n13599, ZN => n7831);
   U2245 : OAI22_X1 port map( A1 => n10700, A2 => n11943, B1 => n11951, B2 => 
                           n13598, ZN => n7830);
   U2246 : OAI22_X1 port map( A1 => n10693, A2 => n11943, B1 => n11951, B2 => 
                           n13597, ZN => n7829);
   U2247 : OAI22_X1 port map( A1 => n10686, A2 => n11943, B1 => n11951, B2 => 
                           n13596, ZN => n7828);
   U2248 : OAI22_X1 port map( A1 => n10679, A2 => n11943, B1 => n11952, B2 => 
                           n13595, ZN => n7827);
   U2249 : OAI22_X1 port map( A1 => n10672, A2 => n11943, B1 => n11952, B2 => 
                           n13594, ZN => n7826);
   U2250 : OAI22_X1 port map( A1 => n10665, A2 => n11943, B1 => n11952, B2 => 
                           n13593, ZN => n7825);
   U2251 : OAI22_X1 port map( A1 => n10658, A2 => n11943, B1 => n11952, B2 => 
                           n13592, ZN => n7824);
   U2252 : OAI22_X1 port map( A1 => n10651, A2 => n11943, B1 => n11953, B2 => 
                           n13591, ZN => n7823);
   U2253 : OAI22_X1 port map( A1 => n10644, A2 => n11943, B1 => n11953, B2 => 
                           n13590, ZN => n7822);
   U2254 : OAI22_X1 port map( A1 => n10637, A2 => n11943, B1 => n11953, B2 => 
                           n13589, ZN => n7821);
   U2255 : OAI22_X1 port map( A1 => n10630, A2 => n11943, B1 => n11953, B2 => 
                           n13588, ZN => n7820);
   U2256 : OAI22_X1 port map( A1 => n10847, A2 => n11933, B1 => n11934, B2 => 
                           n13587, ZN => n7819);
   U2257 : OAI22_X1 port map( A1 => n10840, A2 => n11933, B1 => n11934, B2 => 
                           n13586, ZN => n7818);
   U2258 : OAI22_X1 port map( A1 => n10833, A2 => n11933, B1 => n11934, B2 => 
                           n13585, ZN => n7817);
   U2259 : OAI22_X1 port map( A1 => n10826, A2 => n11933, B1 => n11934, B2 => 
                           n13584, ZN => n7816);
   U2260 : OAI22_X1 port map( A1 => n10819, A2 => n11933, B1 => n11935, B2 => 
                           n13583, ZN => n7815);
   U2261 : OAI22_X1 port map( A1 => n10812, A2 => n11933, B1 => n11935, B2 => 
                           n13582, ZN => n7814);
   U2262 : OAI22_X1 port map( A1 => n10805, A2 => n11933, B1 => n11935, B2 => 
                           n13581, ZN => n7813);
   U2263 : OAI22_X1 port map( A1 => n10798, A2 => n11933, B1 => n11935, B2 => 
                           n13580, ZN => n7812);
   U2264 : OAI22_X1 port map( A1 => n10791, A2 => n11932, B1 => n11936, B2 => 
                           n13579, ZN => n7811);
   U2265 : OAI22_X1 port map( A1 => n10784, A2 => n11932, B1 => n11936, B2 => 
                           n13578, ZN => n7810);
   U2266 : OAI22_X1 port map( A1 => n10777, A2 => n11932, B1 => n11936, B2 => 
                           n13577, ZN => n7809);
   U2267 : OAI22_X1 port map( A1 => n10770, A2 => n11932, B1 => n11936, B2 => 
                           n13576, ZN => n7808);
   U2268 : OAI22_X1 port map( A1 => n10763, A2 => n11932, B1 => n11937, B2 => 
                           n13575, ZN => n7807);
   U2269 : OAI22_X1 port map( A1 => n10756, A2 => n11932, B1 => n11937, B2 => 
                           n13574, ZN => n7806);
   U2270 : OAI22_X1 port map( A1 => n10749, A2 => n11932, B1 => n11937, B2 => 
                           n13573, ZN => n7805);
   U2271 : OAI22_X1 port map( A1 => n10742, A2 => n11932, B1 => n11937, B2 => 
                           n13572, ZN => n7804);
   U2272 : OAI22_X1 port map( A1 => n10735, A2 => n11932, B1 => n11938, B2 => 
                           n13571, ZN => n7803);
   U2273 : OAI22_X1 port map( A1 => n10728, A2 => n11932, B1 => n11938, B2 => 
                           n13570, ZN => n7802);
   U2274 : OAI22_X1 port map( A1 => n10721, A2 => n11932, B1 => n11938, B2 => 
                           n13569, ZN => n7801);
   U2275 : OAI22_X1 port map( A1 => n10714, A2 => n11932, B1 => n11938, B2 => 
                           n13568, ZN => n7800);
   U2276 : OAI22_X1 port map( A1 => n10707, A2 => n11931, B1 => n11939, B2 => 
                           n13567, ZN => n7799);
   U2277 : OAI22_X1 port map( A1 => n10700, A2 => n11931, B1 => n11939, B2 => 
                           n13566, ZN => n7798);
   U2278 : OAI22_X1 port map( A1 => n10693, A2 => n11931, B1 => n11939, B2 => 
                           n13565, ZN => n7797);
   U2279 : OAI22_X1 port map( A1 => n10686, A2 => n11931, B1 => n11939, B2 => 
                           n13564, ZN => n7796);
   U2280 : OAI22_X1 port map( A1 => n10679, A2 => n11931, B1 => n11940, B2 => 
                           n13563, ZN => n7795);
   U2281 : OAI22_X1 port map( A1 => n10672, A2 => n11931, B1 => n11940, B2 => 
                           n13562, ZN => n7794);
   U2282 : OAI22_X1 port map( A1 => n10665, A2 => n11931, B1 => n11940, B2 => 
                           n13561, ZN => n7793);
   U2283 : OAI22_X1 port map( A1 => n10658, A2 => n11931, B1 => n11940, B2 => 
                           n13560, ZN => n7792);
   U2284 : OAI22_X1 port map( A1 => n10651, A2 => n11931, B1 => n11941, B2 => 
                           n13559, ZN => n7791);
   U2285 : OAI22_X1 port map( A1 => n10644, A2 => n11931, B1 => n11941, B2 => 
                           n13558, ZN => n7790);
   U2286 : OAI22_X1 port map( A1 => n10637, A2 => n11931, B1 => n11941, B2 => 
                           n13557, ZN => n7789);
   U2287 : OAI22_X1 port map( A1 => n10630, A2 => n11931, B1 => n11941, B2 => 
                           n13556, ZN => n7788);
   U2288 : OAI22_X1 port map( A1 => n10847, A2 => n11897, B1 => n11898, B2 => 
                           n13491, ZN => n7723);
   U2289 : OAI22_X1 port map( A1 => n10840, A2 => n11897, B1 => n11898, B2 => 
                           n13490, ZN => n7722);
   U2290 : OAI22_X1 port map( A1 => n10833, A2 => n11897, B1 => n11898, B2 => 
                           n13489, ZN => n7721);
   U2291 : OAI22_X1 port map( A1 => n10826, A2 => n11897, B1 => n11898, B2 => 
                           n13488, ZN => n7720);
   U2292 : OAI22_X1 port map( A1 => n10819, A2 => n11897, B1 => n11899, B2 => 
                           n13487, ZN => n7719);
   U2293 : OAI22_X1 port map( A1 => n10812, A2 => n11897, B1 => n11899, B2 => 
                           n13486, ZN => n7718);
   U2294 : OAI22_X1 port map( A1 => n10805, A2 => n11897, B1 => n11899, B2 => 
                           n13485, ZN => n7717);
   U2295 : OAI22_X1 port map( A1 => n10798, A2 => n11897, B1 => n11899, B2 => 
                           n13484, ZN => n7716);
   U2296 : OAI22_X1 port map( A1 => n10791, A2 => n11896, B1 => n11900, B2 => 
                           n13483, ZN => n7715);
   U2297 : OAI22_X1 port map( A1 => n10784, A2 => n11896, B1 => n11900, B2 => 
                           n13482, ZN => n7714);
   U2298 : OAI22_X1 port map( A1 => n10777, A2 => n11896, B1 => n11900, B2 => 
                           n13481, ZN => n7713);
   U2299 : OAI22_X1 port map( A1 => n10770, A2 => n11896, B1 => n11900, B2 => 
                           n13480, ZN => n7712);
   U2300 : OAI22_X1 port map( A1 => n10763, A2 => n11896, B1 => n11901, B2 => 
                           n13479, ZN => n7711);
   U2301 : OAI22_X1 port map( A1 => n10756, A2 => n11896, B1 => n11901, B2 => 
                           n13478, ZN => n7710);
   U2302 : OAI22_X1 port map( A1 => n10749, A2 => n11896, B1 => n11901, B2 => 
                           n13477, ZN => n7709);
   U2303 : OAI22_X1 port map( A1 => n10742, A2 => n11896, B1 => n11901, B2 => 
                           n13476, ZN => n7708);
   U2304 : OAI22_X1 port map( A1 => n10735, A2 => n11896, B1 => n11902, B2 => 
                           n13475, ZN => n7707);
   U2305 : OAI22_X1 port map( A1 => n10728, A2 => n11896, B1 => n11902, B2 => 
                           n13474, ZN => n7706);
   U2306 : OAI22_X1 port map( A1 => n10721, A2 => n11896, B1 => n11902, B2 => 
                           n13473, ZN => n7705);
   U2307 : OAI22_X1 port map( A1 => n10714, A2 => n11896, B1 => n11902, B2 => 
                           n13472, ZN => n7704);
   U2308 : OAI22_X1 port map( A1 => n10707, A2 => n11895, B1 => n11903, B2 => 
                           n13471, ZN => n7703);
   U2309 : OAI22_X1 port map( A1 => n10700, A2 => n11895, B1 => n11903, B2 => 
                           n13470, ZN => n7702);
   U2310 : OAI22_X1 port map( A1 => n10693, A2 => n11895, B1 => n11903, B2 => 
                           n13469, ZN => n7701);
   U2311 : OAI22_X1 port map( A1 => n10686, A2 => n11895, B1 => n11903, B2 => 
                           n13468, ZN => n7700);
   U2312 : OAI22_X1 port map( A1 => n10679, A2 => n11895, B1 => n11904, B2 => 
                           n13467, ZN => n7699);
   U2313 : OAI22_X1 port map( A1 => n10672, A2 => n11895, B1 => n11904, B2 => 
                           n13466, ZN => n7698);
   U2314 : OAI22_X1 port map( A1 => n10665, A2 => n11895, B1 => n11904, B2 => 
                           n13465, ZN => n7697);
   U2315 : OAI22_X1 port map( A1 => n10658, A2 => n11895, B1 => n11904, B2 => 
                           n13464, ZN => n7696);
   U2316 : OAI22_X1 port map( A1 => n10651, A2 => n11895, B1 => n11905, B2 => 
                           n13463, ZN => n7695);
   U2317 : OAI22_X1 port map( A1 => n10644, A2 => n11895, B1 => n11905, B2 => 
                           n13462, ZN => n7694);
   U2318 : OAI22_X1 port map( A1 => n10637, A2 => n11895, B1 => n11905, B2 => 
                           n13461, ZN => n7693);
   U2319 : OAI22_X1 port map( A1 => n10630, A2 => n11895, B1 => n11905, B2 => 
                           n13460, ZN => n7692);
   U2320 : OAI22_X1 port map( A1 => n10847, A2 => n11873, B1 => n11874, B2 => 
                           n13459, ZN => n7659);
   U2321 : OAI22_X1 port map( A1 => n10840, A2 => n11873, B1 => n11874, B2 => 
                           n13458, ZN => n7658);
   U2322 : OAI22_X1 port map( A1 => n10833, A2 => n11873, B1 => n11874, B2 => 
                           n13457, ZN => n7657);
   U2323 : OAI22_X1 port map( A1 => n10826, A2 => n11873, B1 => n11874, B2 => 
                           n13456, ZN => n7656);
   U2324 : OAI22_X1 port map( A1 => n10819, A2 => n11873, B1 => n11875, B2 => 
                           n13455, ZN => n7655);
   U2325 : OAI22_X1 port map( A1 => n10812, A2 => n11873, B1 => n11875, B2 => 
                           n13454, ZN => n7654);
   U2326 : OAI22_X1 port map( A1 => n10805, A2 => n11873, B1 => n11875, B2 => 
                           n13453, ZN => n7653);
   U2327 : OAI22_X1 port map( A1 => n10798, A2 => n11873, B1 => n11875, B2 => 
                           n13452, ZN => n7652);
   U2328 : OAI22_X1 port map( A1 => n10791, A2 => n11872, B1 => n11876, B2 => 
                           n13451, ZN => n7651);
   U2329 : OAI22_X1 port map( A1 => n10784, A2 => n11872, B1 => n11876, B2 => 
                           n13450, ZN => n7650);
   U2330 : OAI22_X1 port map( A1 => n10777, A2 => n11872, B1 => n11876, B2 => 
                           n13449, ZN => n7649);
   U2331 : OAI22_X1 port map( A1 => n10770, A2 => n11872, B1 => n11876, B2 => 
                           n13448, ZN => n7648);
   U2332 : OAI22_X1 port map( A1 => n10763, A2 => n11872, B1 => n11877, B2 => 
                           n13447, ZN => n7647);
   U2333 : OAI22_X1 port map( A1 => n10756, A2 => n11872, B1 => n11877, B2 => 
                           n13446, ZN => n7646);
   U2334 : OAI22_X1 port map( A1 => n10749, A2 => n11872, B1 => n11877, B2 => 
                           n13445, ZN => n7645);
   U2335 : OAI22_X1 port map( A1 => n10742, A2 => n11872, B1 => n11877, B2 => 
                           n13444, ZN => n7644);
   U2336 : OAI22_X1 port map( A1 => n10735, A2 => n11872, B1 => n11878, B2 => 
                           n13443, ZN => n7643);
   U2337 : OAI22_X1 port map( A1 => n10728, A2 => n11872, B1 => n11878, B2 => 
                           n13442, ZN => n7642);
   U2338 : OAI22_X1 port map( A1 => n10721, A2 => n11872, B1 => n11878, B2 => 
                           n13441, ZN => n7641);
   U2339 : OAI22_X1 port map( A1 => n10714, A2 => n11872, B1 => n11878, B2 => 
                           n13440, ZN => n7640);
   U2340 : OAI22_X1 port map( A1 => n10707, A2 => n11871, B1 => n11879, B2 => 
                           n13439, ZN => n7639);
   U2341 : OAI22_X1 port map( A1 => n10700, A2 => n11871, B1 => n11879, B2 => 
                           n13438, ZN => n7638);
   U2342 : OAI22_X1 port map( A1 => n10693, A2 => n11871, B1 => n11879, B2 => 
                           n13437, ZN => n7637);
   U2343 : OAI22_X1 port map( A1 => n10686, A2 => n11871, B1 => n11879, B2 => 
                           n13436, ZN => n7636);
   U2344 : OAI22_X1 port map( A1 => n10679, A2 => n11871, B1 => n11880, B2 => 
                           n13435, ZN => n7635);
   U2345 : OAI22_X1 port map( A1 => n10672, A2 => n11871, B1 => n11880, B2 => 
                           n13434, ZN => n7634);
   U2346 : OAI22_X1 port map( A1 => n10665, A2 => n11871, B1 => n11880, B2 => 
                           n13433, ZN => n7633);
   U2347 : OAI22_X1 port map( A1 => n10658, A2 => n11871, B1 => n11880, B2 => 
                           n13432, ZN => n7632);
   U2348 : OAI22_X1 port map( A1 => n10651, A2 => n11871, B1 => n11881, B2 => 
                           n13431, ZN => n7631);
   U2349 : OAI22_X1 port map( A1 => n10644, A2 => n11871, B1 => n11881, B2 => 
                           n13430, ZN => n7630);
   U2350 : OAI22_X1 port map( A1 => n10637, A2 => n11871, B1 => n11881, B2 => 
                           n13429, ZN => n7629);
   U2351 : OAI22_X1 port map( A1 => n10630, A2 => n11871, B1 => n11881, B2 => 
                           n13428, ZN => n7628);
   U2352 : OAI22_X1 port map( A1 => n10847, A2 => n11849, B1 => n11850, B2 => 
                           n13427, ZN => n7595);
   U2353 : OAI22_X1 port map( A1 => n10840, A2 => n11849, B1 => n11850, B2 => 
                           n13426, ZN => n7594);
   U2354 : OAI22_X1 port map( A1 => n10833, A2 => n11849, B1 => n11850, B2 => 
                           n13425, ZN => n7593);
   U2355 : OAI22_X1 port map( A1 => n10826, A2 => n11849, B1 => n11850, B2 => 
                           n13424, ZN => n7592);
   U2356 : OAI22_X1 port map( A1 => n10819, A2 => n11849, B1 => n11851, B2 => 
                           n13423, ZN => n7591);
   U2357 : OAI22_X1 port map( A1 => n10812, A2 => n11849, B1 => n11851, B2 => 
                           n13422, ZN => n7590);
   U2358 : OAI22_X1 port map( A1 => n10805, A2 => n11849, B1 => n11851, B2 => 
                           n13421, ZN => n7589);
   U2359 : OAI22_X1 port map( A1 => n10798, A2 => n11849, B1 => n11851, B2 => 
                           n13420, ZN => n7588);
   U2360 : OAI22_X1 port map( A1 => n10791, A2 => n11848, B1 => n11852, B2 => 
                           n13419, ZN => n7587);
   U2361 : OAI22_X1 port map( A1 => n10784, A2 => n11848, B1 => n11852, B2 => 
                           n13418, ZN => n7586);
   U2362 : OAI22_X1 port map( A1 => n10777, A2 => n11848, B1 => n11852, B2 => 
                           n13417, ZN => n7585);
   U2363 : OAI22_X1 port map( A1 => n10770, A2 => n11848, B1 => n11852, B2 => 
                           n13416, ZN => n7584);
   U2364 : OAI22_X1 port map( A1 => n10763, A2 => n11848, B1 => n11853, B2 => 
                           n13415, ZN => n7583);
   U2365 : OAI22_X1 port map( A1 => n10756, A2 => n11848, B1 => n11853, B2 => 
                           n13414, ZN => n7582);
   U2366 : OAI22_X1 port map( A1 => n10749, A2 => n11848, B1 => n11853, B2 => 
                           n13413, ZN => n7581);
   U2367 : OAI22_X1 port map( A1 => n10742, A2 => n11848, B1 => n11853, B2 => 
                           n13412, ZN => n7580);
   U2368 : OAI22_X1 port map( A1 => n10735, A2 => n11848, B1 => n11854, B2 => 
                           n13411, ZN => n7579);
   U2369 : OAI22_X1 port map( A1 => n10728, A2 => n11848, B1 => n11854, B2 => 
                           n13410, ZN => n7578);
   U2370 : OAI22_X1 port map( A1 => n10721, A2 => n11848, B1 => n11854, B2 => 
                           n13409, ZN => n7577);
   U2371 : OAI22_X1 port map( A1 => n10714, A2 => n11848, B1 => n11854, B2 => 
                           n13408, ZN => n7576);
   U2372 : OAI22_X1 port map( A1 => n10707, A2 => n11847, B1 => n11855, B2 => 
                           n13407, ZN => n7575);
   U2373 : OAI22_X1 port map( A1 => n10700, A2 => n11847, B1 => n11855, B2 => 
                           n13406, ZN => n7574);
   U2374 : OAI22_X1 port map( A1 => n10693, A2 => n11847, B1 => n11855, B2 => 
                           n13405, ZN => n7573);
   U2375 : OAI22_X1 port map( A1 => n10686, A2 => n11847, B1 => n11855, B2 => 
                           n13404, ZN => n7572);
   U2376 : OAI22_X1 port map( A1 => n10679, A2 => n11847, B1 => n11856, B2 => 
                           n13403, ZN => n7571);
   U2377 : OAI22_X1 port map( A1 => n10672, A2 => n11847, B1 => n11856, B2 => 
                           n13402, ZN => n7570);
   U2378 : OAI22_X1 port map( A1 => n10665, A2 => n11847, B1 => n11856, B2 => 
                           n13401, ZN => n7569);
   U2379 : OAI22_X1 port map( A1 => n10658, A2 => n11847, B1 => n11856, B2 => 
                           n13400, ZN => n7568);
   U2380 : OAI22_X1 port map( A1 => n10651, A2 => n11847, B1 => n11857, B2 => 
                           n13399, ZN => n7567);
   U2381 : OAI22_X1 port map( A1 => n10644, A2 => n11847, B1 => n11857, B2 => 
                           n13398, ZN => n7566);
   U2382 : OAI22_X1 port map( A1 => n10637, A2 => n11847, B1 => n11857, B2 => 
                           n13397, ZN => n7565);
   U2383 : OAI22_X1 port map( A1 => n10630, A2 => n11847, B1 => n11857, B2 => 
                           n13396, ZN => n7564);
   U2384 : OAI22_X1 port map( A1 => n10848, A2 => n11693, B1 => n11694, B2 => 
                           n13203, ZN => n7179);
   U2385 : OAI22_X1 port map( A1 => n10841, A2 => n11693, B1 => n11694, B2 => 
                           n13202, ZN => n7178);
   U2386 : OAI22_X1 port map( A1 => n10834, A2 => n11693, B1 => n11694, B2 => 
                           n13201, ZN => n7177);
   U2387 : OAI22_X1 port map( A1 => n10827, A2 => n11693, B1 => n11694, B2 => 
                           n13200, ZN => n7176);
   U2388 : OAI22_X1 port map( A1 => n10820, A2 => n11693, B1 => n11695, B2 => 
                           n13199, ZN => n7175);
   U2389 : OAI22_X1 port map( A1 => n10813, A2 => n11693, B1 => n11695, B2 => 
                           n13198, ZN => n7174);
   U2390 : OAI22_X1 port map( A1 => n10806, A2 => n11693, B1 => n11695, B2 => 
                           n13197, ZN => n7173);
   U2391 : OAI22_X1 port map( A1 => n10799, A2 => n11693, B1 => n11695, B2 => 
                           n13196, ZN => n7172);
   U2392 : OAI22_X1 port map( A1 => n10792, A2 => n11692, B1 => n11696, B2 => 
                           n13195, ZN => n7171);
   U2393 : OAI22_X1 port map( A1 => n10785, A2 => n11692, B1 => n11696, B2 => 
                           n13194, ZN => n7170);
   U2394 : OAI22_X1 port map( A1 => n10778, A2 => n11692, B1 => n11696, B2 => 
                           n13193, ZN => n7169);
   U2395 : OAI22_X1 port map( A1 => n10771, A2 => n11692, B1 => n11696, B2 => 
                           n13192, ZN => n7168);
   U2396 : OAI22_X1 port map( A1 => n10764, A2 => n11692, B1 => n11697, B2 => 
                           n13191, ZN => n7167);
   U2397 : OAI22_X1 port map( A1 => n10757, A2 => n11692, B1 => n11697, B2 => 
                           n13190, ZN => n7166);
   U2398 : OAI22_X1 port map( A1 => n10750, A2 => n11692, B1 => n11697, B2 => 
                           n13189, ZN => n7165);
   U2399 : OAI22_X1 port map( A1 => n10743, A2 => n11692, B1 => n11697, B2 => 
                           n13188, ZN => n7164);
   U2400 : OAI22_X1 port map( A1 => n10736, A2 => n11692, B1 => n11698, B2 => 
                           n13187, ZN => n7163);
   U2401 : OAI22_X1 port map( A1 => n10729, A2 => n11692, B1 => n11698, B2 => 
                           n13186, ZN => n7162);
   U2402 : OAI22_X1 port map( A1 => n10722, A2 => n11692, B1 => n11698, B2 => 
                           n13185, ZN => n7161);
   U2403 : OAI22_X1 port map( A1 => n10715, A2 => n11692, B1 => n11698, B2 => 
                           n13184, ZN => n7160);
   U2404 : OAI22_X1 port map( A1 => n10708, A2 => n11691, B1 => n11699, B2 => 
                           n13183, ZN => n7159);
   U2405 : OAI22_X1 port map( A1 => n10701, A2 => n11691, B1 => n11699, B2 => 
                           n13182, ZN => n7158);
   U2406 : OAI22_X1 port map( A1 => n10694, A2 => n11691, B1 => n11699, B2 => 
                           n13181, ZN => n7157);
   U2407 : OAI22_X1 port map( A1 => n10687, A2 => n11691, B1 => n11699, B2 => 
                           n13180, ZN => n7156);
   U2408 : OAI22_X1 port map( A1 => n10680, A2 => n11691, B1 => n11700, B2 => 
                           n13179, ZN => n7155);
   U2409 : OAI22_X1 port map( A1 => n10673, A2 => n11691, B1 => n11700, B2 => 
                           n13178, ZN => n7154);
   U2410 : OAI22_X1 port map( A1 => n10666, A2 => n11691, B1 => n11700, B2 => 
                           n13177, ZN => n7153);
   U2411 : OAI22_X1 port map( A1 => n10659, A2 => n11691, B1 => n11700, B2 => 
                           n13176, ZN => n7152);
   U2412 : OAI22_X1 port map( A1 => n10652, A2 => n11691, B1 => n11701, B2 => 
                           n13175, ZN => n7151);
   U2413 : OAI22_X1 port map( A1 => n10645, A2 => n11691, B1 => n11701, B2 => 
                           n13174, ZN => n7150);
   U2414 : OAI22_X1 port map( A1 => n10638, A2 => n11691, B1 => n11701, B2 => 
                           n13173, ZN => n7149);
   U2415 : OAI22_X1 port map( A1 => n10631, A2 => n11691, B1 => n11701, B2 => 
                           n13172, ZN => n7148);
   U2416 : OAI22_X1 port map( A1 => n10848, A2 => n11681, B1 => n11682, B2 => 
                           n13171, ZN => n7147);
   U2417 : OAI22_X1 port map( A1 => n10841, A2 => n11681, B1 => n11682, B2 => 
                           n13170, ZN => n7146);
   U2418 : OAI22_X1 port map( A1 => n10834, A2 => n11681, B1 => n11682, B2 => 
                           n13169, ZN => n7145);
   U2419 : OAI22_X1 port map( A1 => n10827, A2 => n11681, B1 => n11682, B2 => 
                           n13168, ZN => n7144);
   U2420 : OAI22_X1 port map( A1 => n10820, A2 => n11681, B1 => n11683, B2 => 
                           n13167, ZN => n7143);
   U2421 : OAI22_X1 port map( A1 => n10813, A2 => n11681, B1 => n11683, B2 => 
                           n13166, ZN => n7142);
   U2422 : OAI22_X1 port map( A1 => n10806, A2 => n11681, B1 => n11683, B2 => 
                           n13165, ZN => n7141);
   U2423 : OAI22_X1 port map( A1 => n10799, A2 => n11681, B1 => n11683, B2 => 
                           n13164, ZN => n7140);
   U2424 : OAI22_X1 port map( A1 => n10792, A2 => n11680, B1 => n11684, B2 => 
                           n13163, ZN => n7139);
   U2425 : OAI22_X1 port map( A1 => n10785, A2 => n11680, B1 => n11684, B2 => 
                           n13162, ZN => n7138);
   U2426 : OAI22_X1 port map( A1 => n10778, A2 => n11680, B1 => n11684, B2 => 
                           n13161, ZN => n7137);
   U2427 : OAI22_X1 port map( A1 => n10771, A2 => n11680, B1 => n11684, B2 => 
                           n13160, ZN => n7136);
   U2428 : OAI22_X1 port map( A1 => n10764, A2 => n11680, B1 => n11685, B2 => 
                           n13159, ZN => n7135);
   U2429 : OAI22_X1 port map( A1 => n10757, A2 => n11680, B1 => n11685, B2 => 
                           n13158, ZN => n7134);
   U2430 : OAI22_X1 port map( A1 => n10750, A2 => n11680, B1 => n11685, B2 => 
                           n13157, ZN => n7133);
   U2431 : OAI22_X1 port map( A1 => n10743, A2 => n11680, B1 => n11685, B2 => 
                           n13156, ZN => n7132);
   U2432 : OAI22_X1 port map( A1 => n10736, A2 => n11680, B1 => n11686, B2 => 
                           n13155, ZN => n7131);
   U2433 : OAI22_X1 port map( A1 => n10729, A2 => n11680, B1 => n11686, B2 => 
                           n13154, ZN => n7130);
   U2434 : OAI22_X1 port map( A1 => n10722, A2 => n11680, B1 => n11686, B2 => 
                           n13153, ZN => n7129);
   U2435 : OAI22_X1 port map( A1 => n10715, A2 => n11680, B1 => n11686, B2 => 
                           n13152, ZN => n7128);
   U2436 : OAI22_X1 port map( A1 => n10708, A2 => n11679, B1 => n11687, B2 => 
                           n13151, ZN => n7127);
   U2437 : OAI22_X1 port map( A1 => n10701, A2 => n11679, B1 => n11687, B2 => 
                           n13150, ZN => n7126);
   U2438 : OAI22_X1 port map( A1 => n10694, A2 => n11679, B1 => n11687, B2 => 
                           n13149, ZN => n7125);
   U2439 : OAI22_X1 port map( A1 => n10687, A2 => n11679, B1 => n11687, B2 => 
                           n13148, ZN => n7124);
   U2440 : OAI22_X1 port map( A1 => n10680, A2 => n11679, B1 => n11688, B2 => 
                           n13147, ZN => n7123);
   U2441 : OAI22_X1 port map( A1 => n10673, A2 => n11679, B1 => n11688, B2 => 
                           n13146, ZN => n7122);
   U2442 : OAI22_X1 port map( A1 => n10666, A2 => n11679, B1 => n11688, B2 => 
                           n13145, ZN => n7121);
   U2443 : OAI22_X1 port map( A1 => n10659, A2 => n11679, B1 => n11688, B2 => 
                           n13144, ZN => n7120);
   U2444 : OAI22_X1 port map( A1 => n10652, A2 => n11679, B1 => n11689, B2 => 
                           n13143, ZN => n7119);
   U2445 : OAI22_X1 port map( A1 => n10645, A2 => n11679, B1 => n11689, B2 => 
                           n13142, ZN => n7118);
   U2446 : OAI22_X1 port map( A1 => n10638, A2 => n11679, B1 => n11689, B2 => 
                           n13141, ZN => n7117);
   U2447 : OAI22_X1 port map( A1 => n10631, A2 => n11679, B1 => n11689, B2 => 
                           n13140, ZN => n7116);
   U2448 : OAI22_X1 port map( A1 => n10848, A2 => n11669, B1 => n11670, B2 => 
                           n13139, ZN => n7115);
   U2449 : OAI22_X1 port map( A1 => n10841, A2 => n11669, B1 => n11670, B2 => 
                           n13138, ZN => n7114);
   U2450 : OAI22_X1 port map( A1 => n10834, A2 => n11669, B1 => n11670, B2 => 
                           n13137, ZN => n7113);
   U2451 : OAI22_X1 port map( A1 => n10827, A2 => n11669, B1 => n11670, B2 => 
                           n13136, ZN => n7112);
   U2452 : OAI22_X1 port map( A1 => n10820, A2 => n11669, B1 => n11671, B2 => 
                           n13135, ZN => n7111);
   U2453 : OAI22_X1 port map( A1 => n10813, A2 => n11669, B1 => n11671, B2 => 
                           n13134, ZN => n7110);
   U2454 : OAI22_X1 port map( A1 => n10806, A2 => n11669, B1 => n11671, B2 => 
                           n13133, ZN => n7109);
   U2455 : OAI22_X1 port map( A1 => n10799, A2 => n11669, B1 => n11671, B2 => 
                           n13132, ZN => n7108);
   U2456 : OAI22_X1 port map( A1 => n10792, A2 => n11668, B1 => n11672, B2 => 
                           n13131, ZN => n7107);
   U2457 : OAI22_X1 port map( A1 => n10785, A2 => n11668, B1 => n11672, B2 => 
                           n13130, ZN => n7106);
   U2458 : OAI22_X1 port map( A1 => n10778, A2 => n11668, B1 => n11672, B2 => 
                           n13129, ZN => n7105);
   U2459 : OAI22_X1 port map( A1 => n10771, A2 => n11668, B1 => n11672, B2 => 
                           n13128, ZN => n7104);
   U2460 : OAI22_X1 port map( A1 => n10764, A2 => n11668, B1 => n11673, B2 => 
                           n13127, ZN => n7103);
   U2461 : OAI22_X1 port map( A1 => n10757, A2 => n11668, B1 => n11673, B2 => 
                           n13126, ZN => n7102);
   U2462 : OAI22_X1 port map( A1 => n10750, A2 => n11668, B1 => n11673, B2 => 
                           n13125, ZN => n7101);
   U2463 : OAI22_X1 port map( A1 => n10743, A2 => n11668, B1 => n11673, B2 => 
                           n13124, ZN => n7100);
   U2464 : OAI22_X1 port map( A1 => n10736, A2 => n11668, B1 => n11674, B2 => 
                           n13123, ZN => n7099);
   U2465 : OAI22_X1 port map( A1 => n10729, A2 => n11668, B1 => n11674, B2 => 
                           n13122, ZN => n7098);
   U2466 : OAI22_X1 port map( A1 => n10722, A2 => n11668, B1 => n11674, B2 => 
                           n13121, ZN => n7097);
   U2467 : OAI22_X1 port map( A1 => n10715, A2 => n11668, B1 => n11674, B2 => 
                           n13120, ZN => n7096);
   U2468 : OAI22_X1 port map( A1 => n10708, A2 => n11667, B1 => n11675, B2 => 
                           n13119, ZN => n7095);
   U2469 : OAI22_X1 port map( A1 => n10701, A2 => n11667, B1 => n11675, B2 => 
                           n13118, ZN => n7094);
   U2470 : OAI22_X1 port map( A1 => n10694, A2 => n11667, B1 => n11675, B2 => 
                           n13117, ZN => n7093);
   U2471 : OAI22_X1 port map( A1 => n10687, A2 => n11667, B1 => n11675, B2 => 
                           n13116, ZN => n7092);
   U2472 : OAI22_X1 port map( A1 => n10680, A2 => n11667, B1 => n11676, B2 => 
                           n13115, ZN => n7091);
   U2473 : OAI22_X1 port map( A1 => n10673, A2 => n11667, B1 => n11676, B2 => 
                           n13114, ZN => n7090);
   U2474 : OAI22_X1 port map( A1 => n10666, A2 => n11667, B1 => n11676, B2 => 
                           n13113, ZN => n7089);
   U2475 : OAI22_X1 port map( A1 => n10659, A2 => n11667, B1 => n11676, B2 => 
                           n13112, ZN => n7088);
   U2476 : OAI22_X1 port map( A1 => n10652, A2 => n11667, B1 => n11677, B2 => 
                           n13111, ZN => n7087);
   U2477 : OAI22_X1 port map( A1 => n10645, A2 => n11667, B1 => n11677, B2 => 
                           n13110, ZN => n7086);
   U2478 : OAI22_X1 port map( A1 => n10638, A2 => n11667, B1 => n11677, B2 => 
                           n13109, ZN => n7085);
   U2479 : OAI22_X1 port map( A1 => n10631, A2 => n11667, B1 => n11677, B2 => 
                           n13108, ZN => n7084);
   U2480 : OAI22_X1 port map( A1 => n10640, A2 => n11475, B1 => n11485, B2 => 
                           n12787, ZN => n6573);
   U2481 : OAI22_X1 port map( A1 => n10633, A2 => n11475, B1 => n11485, B2 => 
                           n12786, ZN => n6572);
   U2482 : OAI22_X1 port map( A1 => n10647, A2 => n11439, B1 => n11449, B2 => 
                           n12785, ZN => n6478);
   U2483 : OAI22_X1 port map( A1 => n10640, A2 => n11439, B1 => n11449, B2 => 
                           n12784, ZN => n6477);
   U2484 : OAI22_X1 port map( A1 => n10633, A2 => n11439, B1 => n11449, B2 => 
                           n12783, ZN => n6476);
   U2485 : OAI22_X1 port map( A1 => n10647, A2 => n11403, B1 => n11413, B2 => 
                           n12782, ZN => n6382);
   U2486 : OAI22_X1 port map( A1 => n10640, A2 => n11403, B1 => n11413, B2 => 
                           n12781, ZN => n6381);
   U2487 : OAI22_X1 port map( A1 => n10633, A2 => n11403, B1 => n11413, B2 => 
                           n12780, ZN => n6380);
   U2488 : INV_X1 port map( A => n2478, ZN => n14517);
   U2489 : INV_X1 port map( A => n2481, ZN => n12777);
   U2490 : NAND2_X1 port map( A1 => n10625, A2 => n10626, ZN => n2487);
   U2491 : INV_X1 port map( A => n2477, ZN => n12778);
   U2492 : AOI21_X1 port map( B1 => n10625, B2 => n2478, A => n2479, ZN => 
                           n2477);
   U2493 : AOI21_X1 port map( B1 => n2480, B2 => n2481, A => n10625, ZN => 
                           n2479);
   U2494 : AOI222_X1 port map( A1 => n11064, A2 => n12979, B1 => n11061, B2 => 
                           n12915, C1 => n11058, C2 => n13043, ZN => n5639);
   U2495 : AOI222_X1 port map( A1 => n10866, A2 => n14448, B1 => n10863, B2 => 
                           n14384, C1 => n10860, C2 => n14512, ZN => n5694);
   U2496 : AOI222_X1 port map( A1 => n11328, A2 => n12979, B1 => n11325, B2 => 
                           n12915, C1 => n11322, C2 => n13043, ZN => n4206);
   U2497 : AOI222_X1 port map( A1 => n11130, A2 => n14448, B1 => n11127, B2 => 
                           n14384, C1 => n11124, C2 => n14512, ZN => n4261);
   U2498 : AOI222_X1 port map( A1 => n11064, A2 => n12978, B1 => n11061, B2 => 
                           n12914, C1 => n11058, C2 => n13042, ZN => n5598);
   U2499 : AOI222_X1 port map( A1 => n10866, A2 => n14447, B1 => n10863, B2 => 
                           n14383, C1 => n10860, C2 => n14511, ZN => n5625);
   U2500 : AOI222_X1 port map( A1 => n11328, A2 => n12978, B1 => n11325, B2 => 
                           n12914, C1 => n11322, C2 => n13042, ZN => n4165);
   U2501 : AOI222_X1 port map( A1 => n11130, A2 => n14447, B1 => n11127, B2 => 
                           n14383, C1 => n11124, C2 => n14511, ZN => n4192);
   U2502 : AOI222_X1 port map( A1 => n11064, A2 => n12977, B1 => n11061, B2 => 
                           n12913, C1 => n11058, C2 => n13041, ZN => n5557);
   U2503 : AOI222_X1 port map( A1 => n10866, A2 => n14446, B1 => n10863, B2 => 
                           n14382, C1 => n10860, C2 => n14510, ZN => n5584);
   U2504 : AOI222_X1 port map( A1 => n11328, A2 => n12977, B1 => n11325, B2 => 
                           n12913, C1 => n11322, C2 => n13041, ZN => n4124);
   U2505 : AOI222_X1 port map( A1 => n11130, A2 => n14446, B1 => n11127, B2 => 
                           n14382, C1 => n11124, C2 => n14510, ZN => n4151);
   U2506 : AOI222_X1 port map( A1 => n11064, A2 => n12976, B1 => n11061, B2 => 
                           n12912, C1 => n11058, C2 => n13040, ZN => n5516);
   U2507 : AOI222_X1 port map( A1 => n10866, A2 => n14445, B1 => n10863, B2 => 
                           n14381, C1 => n10860, C2 => n14509, ZN => n5543);
   U2508 : AOI222_X1 port map( A1 => n11328, A2 => n12976, B1 => n11325, B2 => 
                           n12912, C1 => n11322, C2 => n13040, ZN => n4083);
   U2509 : AOI222_X1 port map( A1 => n11130, A2 => n14445, B1 => n11127, B2 => 
                           n14381, C1 => n11124, C2 => n14509, ZN => n4110);
   U2510 : AOI222_X1 port map( A1 => n11064, A2 => n12975, B1 => n11061, B2 => 
                           n12911, C1 => n11058, C2 => n13039, ZN => n5475);
   U2511 : AOI222_X1 port map( A1 => n10866, A2 => n14444, B1 => n10863, B2 => 
                           n14380, C1 => n10860, C2 => n14508, ZN => n5502);
   U2512 : AOI222_X1 port map( A1 => n11328, A2 => n12975, B1 => n11325, B2 => 
                           n12911, C1 => n11322, C2 => n13039, ZN => n4042);
   U2513 : AOI222_X1 port map( A1 => n11130, A2 => n14444, B1 => n11127, B2 => 
                           n14380, C1 => n11124, C2 => n14508, ZN => n4069);
   U2514 : AOI222_X1 port map( A1 => n11064, A2 => n12974, B1 => n11061, B2 => 
                           n12910, C1 => n11058, C2 => n13038, ZN => n5434);
   U2515 : AOI222_X1 port map( A1 => n10866, A2 => n14443, B1 => n10863, B2 => 
                           n14379, C1 => n10860, C2 => n14507, ZN => n5461);
   U2516 : AOI222_X1 port map( A1 => n11328, A2 => n12974, B1 => n11325, B2 => 
                           n12910, C1 => n11322, C2 => n13038, ZN => n4001);
   U2517 : AOI222_X1 port map( A1 => n11130, A2 => n14443, B1 => n11127, B2 => 
                           n14379, C1 => n11124, C2 => n14507, ZN => n4028);
   U2518 : AOI222_X1 port map( A1 => n11064, A2 => n12973, B1 => n11061, B2 => 
                           n12909, C1 => n11058, C2 => n13037, ZN => n5393);
   U2519 : AOI222_X1 port map( A1 => n10866, A2 => n14442, B1 => n10863, B2 => 
                           n14378, C1 => n10860, C2 => n14506, ZN => n5420);
   U2520 : AOI222_X1 port map( A1 => n11328, A2 => n12973, B1 => n11325, B2 => 
                           n12909, C1 => n11322, C2 => n13037, ZN => n3960);
   U2521 : AOI222_X1 port map( A1 => n11130, A2 => n14442, B1 => n11127, B2 => 
                           n14378, C1 => n11124, C2 => n14506, ZN => n3987);
   U2522 : AOI222_X1 port map( A1 => n11064, A2 => n12972, B1 => n11061, B2 => 
                           n12908, C1 => n11058, C2 => n13036, ZN => n5352);
   U2523 : AOI222_X1 port map( A1 => n10866, A2 => n14441, B1 => n10863, B2 => 
                           n14377, C1 => n10860, C2 => n14505, ZN => n5379);
   U2524 : AOI222_X1 port map( A1 => n11328, A2 => n12972, B1 => n11325, B2 => 
                           n12908, C1 => n11322, C2 => n13036, ZN => n3919);
   U2525 : AOI222_X1 port map( A1 => n11130, A2 => n14441, B1 => n11127, B2 => 
                           n14377, C1 => n11124, C2 => n14505, ZN => n3946);
   U2526 : AOI222_X1 port map( A1 => n11064, A2 => n12971, B1 => n11061, B2 => 
                           n12907, C1 => n11058, C2 => n13035, ZN => n5311);
   U2527 : AOI222_X1 port map( A1 => n10866, A2 => n14440, B1 => n10863, B2 => 
                           n14376, C1 => n10860, C2 => n14504, ZN => n5338);
   U2528 : AOI222_X1 port map( A1 => n11328, A2 => n12971, B1 => n11325, B2 => 
                           n12907, C1 => n11322, C2 => n13035, ZN => n3878);
   U2529 : AOI222_X1 port map( A1 => n11130, A2 => n14440, B1 => n11127, B2 => 
                           n14376, C1 => n11124, C2 => n14504, ZN => n3905);
   U2530 : AOI222_X1 port map( A1 => n11064, A2 => n12970, B1 => n11061, B2 => 
                           n12906, C1 => n11058, C2 => n13034, ZN => n5270);
   U2531 : AOI222_X1 port map( A1 => n10866, A2 => n14439, B1 => n10863, B2 => 
                           n14375, C1 => n10860, C2 => n14503, ZN => n5297);
   U2532 : AOI222_X1 port map( A1 => n11328, A2 => n12970, B1 => n11325, B2 => 
                           n12906, C1 => n11322, C2 => n13034, ZN => n3837);
   U2533 : AOI222_X1 port map( A1 => n11130, A2 => n14439, B1 => n11127, B2 => 
                           n14375, C1 => n11124, C2 => n14503, ZN => n3864);
   U2534 : AOI222_X1 port map( A1 => n11064, A2 => n12969, B1 => n11061, B2 => 
                           n12905, C1 => n11058, C2 => n13033, ZN => n5229);
   U2535 : AOI222_X1 port map( A1 => n10866, A2 => n14438, B1 => n10863, B2 => 
                           n14374, C1 => n10860, C2 => n14502, ZN => n5256);
   U2536 : AOI222_X1 port map( A1 => n11328, A2 => n12969, B1 => n11325, B2 => 
                           n12905, C1 => n11322, C2 => n13033, ZN => n3796);
   U2537 : AOI222_X1 port map( A1 => n11130, A2 => n14438, B1 => n11127, B2 => 
                           n14374, C1 => n11124, C2 => n14502, ZN => n3823);
   U2538 : AOI222_X1 port map( A1 => n11064, A2 => n12968, B1 => n11061, B2 => 
                           n12904, C1 => n11058, C2 => n13032, ZN => n5188);
   U2539 : AOI222_X1 port map( A1 => n10866, A2 => n14437, B1 => n10863, B2 => 
                           n14373, C1 => n10860, C2 => n14501, ZN => n5215);
   U2540 : AOI222_X1 port map( A1 => n11328, A2 => n12968, B1 => n11325, B2 => 
                           n12904, C1 => n11322, C2 => n13032, ZN => n3755);
   U2541 : AOI222_X1 port map( A1 => n11130, A2 => n14437, B1 => n11127, B2 => 
                           n14373, C1 => n11124, C2 => n14501, ZN => n3782);
   U2542 : AOI222_X1 port map( A1 => n11065, A2 => n12967, B1 => n11062, B2 => 
                           n12903, C1 => n11059, C2 => n13031, ZN => n5147);
   U2543 : AOI222_X1 port map( A1 => n10867, A2 => n14436, B1 => n10864, B2 => 
                           n14372, C1 => n10861, C2 => n14500, ZN => n5174);
   U2544 : AOI222_X1 port map( A1 => n11329, A2 => n12967, B1 => n11326, B2 => 
                           n12903, C1 => n11323, C2 => n13031, ZN => n3714);
   U2545 : AOI222_X1 port map( A1 => n11131, A2 => n14436, B1 => n11128, B2 => 
                           n14372, C1 => n11125, C2 => n14500, ZN => n3741);
   U2546 : AOI222_X1 port map( A1 => n11065, A2 => n12966, B1 => n11062, B2 => 
                           n12902, C1 => n11059, C2 => n13030, ZN => n5106);
   U2547 : AOI222_X1 port map( A1 => n10867, A2 => n14435, B1 => n10864, B2 => 
                           n14371, C1 => n10861, C2 => n14499, ZN => n5133);
   U2548 : AOI222_X1 port map( A1 => n11329, A2 => n12966, B1 => n11326, B2 => 
                           n12902, C1 => n11323, C2 => n13030, ZN => n3673);
   U2549 : AOI222_X1 port map( A1 => n11131, A2 => n14435, B1 => n11128, B2 => 
                           n14371, C1 => n11125, C2 => n14499, ZN => n3700);
   U2550 : AOI222_X1 port map( A1 => n11065, A2 => n12965, B1 => n11062, B2 => 
                           n12901, C1 => n11059, C2 => n13029, ZN => n5065);
   U2551 : AOI222_X1 port map( A1 => n10867, A2 => n14434, B1 => n10864, B2 => 
                           n14370, C1 => n10861, C2 => n14498, ZN => n5092);
   U2552 : AOI222_X1 port map( A1 => n11329, A2 => n12965, B1 => n11326, B2 => 
                           n12901, C1 => n11323, C2 => n13029, ZN => n3632);
   U2553 : AOI222_X1 port map( A1 => n11131, A2 => n14434, B1 => n11128, B2 => 
                           n14370, C1 => n11125, C2 => n14498, ZN => n3659);
   U2554 : AOI222_X1 port map( A1 => n11065, A2 => n12964, B1 => n11062, B2 => 
                           n12900, C1 => n11059, C2 => n13028, ZN => n5024);
   U2555 : AOI222_X1 port map( A1 => n10867, A2 => n14433, B1 => n10864, B2 => 
                           n14369, C1 => n10861, C2 => n14497, ZN => n5051);
   U2556 : AOI222_X1 port map( A1 => n11329, A2 => n12964, B1 => n11326, B2 => 
                           n12900, C1 => n11323, C2 => n13028, ZN => n3591);
   U2557 : AOI222_X1 port map( A1 => n11131, A2 => n14433, B1 => n11128, B2 => 
                           n14369, C1 => n11125, C2 => n14497, ZN => n3618);
   U2558 : AOI222_X1 port map( A1 => n11065, A2 => n12963, B1 => n11062, B2 => 
                           n12899, C1 => n11059, C2 => n13027, ZN => n4983);
   U2559 : AOI222_X1 port map( A1 => n10867, A2 => n14432, B1 => n10864, B2 => 
                           n14368, C1 => n10861, C2 => n14496, ZN => n5010);
   U2560 : AOI222_X1 port map( A1 => n11329, A2 => n12963, B1 => n11326, B2 => 
                           n12899, C1 => n11323, C2 => n13027, ZN => n3550);
   U2561 : AOI222_X1 port map( A1 => n11131, A2 => n14432, B1 => n11128, B2 => 
                           n14368, C1 => n11125, C2 => n14496, ZN => n3577);
   U2562 : AOI222_X1 port map( A1 => n11065, A2 => n12962, B1 => n11062, B2 => 
                           n12898, C1 => n11059, C2 => n13026, ZN => n4942);
   U2563 : AOI222_X1 port map( A1 => n10867, A2 => n14431, B1 => n10864, B2 => 
                           n14367, C1 => n10861, C2 => n14495, ZN => n4969);
   U2564 : AOI222_X1 port map( A1 => n11329, A2 => n12962, B1 => n11326, B2 => 
                           n12898, C1 => n11323, C2 => n13026, ZN => n3509);
   U2565 : AOI222_X1 port map( A1 => n11131, A2 => n14431, B1 => n11128, B2 => 
                           n14367, C1 => n11125, C2 => n14495, ZN => n3536);
   U2566 : AOI222_X1 port map( A1 => n11065, A2 => n12961, B1 => n11062, B2 => 
                           n12897, C1 => n11059, C2 => n13025, ZN => n4901);
   U2567 : AOI222_X1 port map( A1 => n10867, A2 => n14430, B1 => n10864, B2 => 
                           n14366, C1 => n10861, C2 => n14494, ZN => n4928);
   U2568 : AOI222_X1 port map( A1 => n11329, A2 => n12961, B1 => n11326, B2 => 
                           n12897, C1 => n11323, C2 => n13025, ZN => n3468);
   U2569 : AOI222_X1 port map( A1 => n11131, A2 => n14430, B1 => n11128, B2 => 
                           n14366, C1 => n11125, C2 => n14494, ZN => n3495);
   U2570 : AOI222_X1 port map( A1 => n11065, A2 => n12960, B1 => n11062, B2 => 
                           n12896, C1 => n11059, C2 => n13024, ZN => n4860);
   U2571 : AOI222_X1 port map( A1 => n10867, A2 => n14429, B1 => n10864, B2 => 
                           n14365, C1 => n10861, C2 => n14493, ZN => n4887);
   U2572 : AOI222_X1 port map( A1 => n11329, A2 => n12960, B1 => n11326, B2 => 
                           n12896, C1 => n11323, C2 => n13024, ZN => n3427);
   U2573 : AOI222_X1 port map( A1 => n11131, A2 => n14429, B1 => n11128, B2 => 
                           n14365, C1 => n11125, C2 => n14493, ZN => n3454);
   U2574 : AOI222_X1 port map( A1 => n11065, A2 => n12959, B1 => n11062, B2 => 
                           n12895, C1 => n11059, C2 => n13023, ZN => n4819);
   U2575 : AOI222_X1 port map( A1 => n10867, A2 => n14428, B1 => n10864, B2 => 
                           n14364, C1 => n10861, C2 => n14492, ZN => n4846);
   U2576 : AOI222_X1 port map( A1 => n11329, A2 => n12959, B1 => n11326, B2 => 
                           n12895, C1 => n11323, C2 => n13023, ZN => n3386);
   U2577 : AOI222_X1 port map( A1 => n11131, A2 => n14428, B1 => n11128, B2 => 
                           n14364, C1 => n11125, C2 => n14492, ZN => n3413);
   U2578 : AOI222_X1 port map( A1 => n11065, A2 => n12958, B1 => n11062, B2 => 
                           n12894, C1 => n11059, C2 => n13022, ZN => n4778);
   U2579 : AOI222_X1 port map( A1 => n10867, A2 => n14427, B1 => n10864, B2 => 
                           n14363, C1 => n10861, C2 => n14491, ZN => n4805);
   U2580 : AOI222_X1 port map( A1 => n11329, A2 => n12958, B1 => n11326, B2 => 
                           n12894, C1 => n11323, C2 => n13022, ZN => n3345);
   U2581 : AOI222_X1 port map( A1 => n11131, A2 => n14427, B1 => n11128, B2 => 
                           n14363, C1 => n11125, C2 => n14491, ZN => n3372);
   U2582 : AOI222_X1 port map( A1 => n11065, A2 => n12957, B1 => n11062, B2 => 
                           n12893, C1 => n11059, C2 => n13021, ZN => n4737);
   U2583 : AOI222_X1 port map( A1 => n10867, A2 => n14426, B1 => n10864, B2 => 
                           n14362, C1 => n10861, C2 => n14490, ZN => n4764);
   U2584 : AOI222_X1 port map( A1 => n11329, A2 => n12957, B1 => n11326, B2 => 
                           n12893, C1 => n11323, C2 => n13021, ZN => n3304);
   U2585 : AOI222_X1 port map( A1 => n11131, A2 => n14426, B1 => n11128, B2 => 
                           n14362, C1 => n11125, C2 => n14490, ZN => n3331);
   U2586 : AOI222_X1 port map( A1 => n11065, A2 => n12956, B1 => n11062, B2 => 
                           n12892, C1 => n11059, C2 => n13020, ZN => n4696);
   U2587 : AOI222_X1 port map( A1 => n10867, A2 => n14425, B1 => n10864, B2 => 
                           n14361, C1 => n10861, C2 => n14489, ZN => n4723);
   U2588 : AOI222_X1 port map( A1 => n11329, A2 => n12956, B1 => n11326, B2 => 
                           n12892, C1 => n11323, C2 => n13020, ZN => n3263);
   U2589 : AOI222_X1 port map( A1 => n11131, A2 => n14425, B1 => n11128, B2 => 
                           n14361, C1 => n11125, C2 => n14489, ZN => n3290);
   U2590 : AOI222_X1 port map( A1 => n11066, A2 => n12955, B1 => n11063, B2 => 
                           n12891, C1 => n11060, C2 => n13019, ZN => n4655);
   U2591 : AOI222_X1 port map( A1 => n10868, A2 => n14424, B1 => n10865, B2 => 
                           n14360, C1 => n10862, C2 => n14488, ZN => n4682);
   U2592 : AOI222_X1 port map( A1 => n11330, A2 => n12955, B1 => n11327, B2 => 
                           n12891, C1 => n11324, C2 => n13019, ZN => n3222);
   U2593 : AOI222_X1 port map( A1 => n11132, A2 => n14424, B1 => n11129, B2 => 
                           n14360, C1 => n11126, C2 => n14488, ZN => n3249);
   U2594 : AOI222_X1 port map( A1 => n11066, A2 => n12954, B1 => n11063, B2 => 
                           n12890, C1 => n11060, C2 => n13018, ZN => n4614);
   U2595 : AOI222_X1 port map( A1 => n10868, A2 => n14423, B1 => n10865, B2 => 
                           n14359, C1 => n10862, C2 => n14487, ZN => n4641);
   U2596 : AOI222_X1 port map( A1 => n11330, A2 => n12954, B1 => n11327, B2 => 
                           n12890, C1 => n11324, C2 => n13018, ZN => n3181);
   U2597 : AOI222_X1 port map( A1 => n11132, A2 => n14423, B1 => n11129, B2 => 
                           n14359, C1 => n11126, C2 => n14487, ZN => n3208);
   U2598 : AOI222_X1 port map( A1 => n11066, A2 => n12953, B1 => n11063, B2 => 
                           n12889, C1 => n11060, C2 => n13017, ZN => n4573);
   U2599 : AOI222_X1 port map( A1 => n10868, A2 => n14422, B1 => n10865, B2 => 
                           n14358, C1 => n10862, C2 => n14486, ZN => n4600);
   U2600 : AOI222_X1 port map( A1 => n11330, A2 => n12953, B1 => n11327, B2 => 
                           n12889, C1 => n11324, C2 => n13017, ZN => n3140);
   U2601 : AOI222_X1 port map( A1 => n11132, A2 => n14422, B1 => n11129, B2 => 
                           n14358, C1 => n11126, C2 => n14486, ZN => n3167);
   U2602 : AOI222_X1 port map( A1 => n11066, A2 => n12952, B1 => n11063, B2 => 
                           n12888, C1 => n11060, C2 => n13016, ZN => n4532);
   U2603 : AOI222_X1 port map( A1 => n10868, A2 => n14421, B1 => n10865, B2 => 
                           n14357, C1 => n10862, C2 => n14485, ZN => n4559);
   U2604 : AOI222_X1 port map( A1 => n11330, A2 => n12952, B1 => n11327, B2 => 
                           n12888, C1 => n11324, C2 => n13016, ZN => n3099);
   U2605 : AOI222_X1 port map( A1 => n11132, A2 => n14421, B1 => n11129, B2 => 
                           n14357, C1 => n11126, C2 => n14485, ZN => n3126);
   U2606 : AOI222_X1 port map( A1 => n11066, A2 => n12951, B1 => n11063, B2 => 
                           n12887, C1 => n11060, C2 => n13015, ZN => n4491);
   U2607 : AOI222_X1 port map( A1 => n10868, A2 => n14420, B1 => n10865, B2 => 
                           n14356, C1 => n10862, C2 => n14484, ZN => n4518);
   U2608 : AOI222_X1 port map( A1 => n11330, A2 => n12951, B1 => n11327, B2 => 
                           n12887, C1 => n11324, C2 => n13015, ZN => n3058);
   U2609 : AOI222_X1 port map( A1 => n11132, A2 => n14420, B1 => n11129, B2 => 
                           n14356, C1 => n11126, C2 => n14484, ZN => n3085);
   U2610 : AOI222_X1 port map( A1 => n11066, A2 => n12950, B1 => n11063, B2 => 
                           n12886, C1 => n11060, C2 => n13014, ZN => n4450);
   U2611 : AOI222_X1 port map( A1 => n10868, A2 => n14419, B1 => n10865, B2 => 
                           n14355, C1 => n10862, C2 => n14483, ZN => n4477);
   U2612 : AOI222_X1 port map( A1 => n11330, A2 => n12950, B1 => n11327, B2 => 
                           n12886, C1 => n11324, C2 => n13014, ZN => n3017);
   U2613 : AOI222_X1 port map( A1 => n11132, A2 => n14419, B1 => n11129, B2 => 
                           n14355, C1 => n11126, C2 => n14483, ZN => n3044);
   U2614 : AOI222_X1 port map( A1 => n11066, A2 => n12949, B1 => n11063, B2 => 
                           n12885, C1 => n11060, C2 => n13013, ZN => n4409);
   U2615 : AOI222_X1 port map( A1 => n10868, A2 => n14418, B1 => n10865, B2 => 
                           n14354, C1 => n10862, C2 => n14482, ZN => n4436);
   U2616 : AOI222_X1 port map( A1 => n11330, A2 => n12949, B1 => n11327, B2 => 
                           n12885, C1 => n11324, C2 => n13013, ZN => n2976);
   U2617 : AOI222_X1 port map( A1 => n11132, A2 => n14418, B1 => n11129, B2 => 
                           n14354, C1 => n11126, C2 => n14482, ZN => n3003);
   U2618 : AOI222_X1 port map( A1 => n11066, A2 => n12948, B1 => n11063, B2 => 
                           n12884, C1 => n11060, C2 => n13012, ZN => n4280);
   U2619 : AOI222_X1 port map( A1 => n10868, A2 => n14417, B1 => n10865, B2 => 
                           n14353, C1 => n10862, C2 => n14481, ZN => n4373);
   U2620 : AOI222_X1 port map( A1 => n11330, A2 => n12948, B1 => n11327, B2 => 
                           n12884, C1 => n11324, C2 => n13012, ZN => n2748);
   U2621 : AOI222_X1 port map( A1 => n11132, A2 => n14417, B1 => n11129, B2 => 
                           n14353, C1 => n11126, C2 => n14481, ZN => n2940);
   U2622 : OAI222_X1 port map( A1 => n14042, A2 => n10910, B1 => n14074, B2 => 
                           n10907, C1 => n14010, C2 => n10904, ZN => n4687);
   U2623 : OAI222_X1 port map( A1 => n14042, A2 => n11174, B1 => n14074, B2 => 
                           n11171, C1 => n14010, C2 => n11168, ZN => n3254);
   U2624 : OAI222_X1 port map( A1 => n14041, A2 => n10910, B1 => n14073, B2 => 
                           n10907, C1 => n14009, C2 => n10904, ZN => n4646);
   U2625 : OAI222_X1 port map( A1 => n14041, A2 => n11174, B1 => n14073, B2 => 
                           n11171, C1 => n14009, C2 => n11168, ZN => n3213);
   U2626 : OAI222_X1 port map( A1 => n14040, A2 => n10910, B1 => n14072, B2 => 
                           n10907, C1 => n14008, C2 => n10904, ZN => n4605);
   U2627 : OAI222_X1 port map( A1 => n14040, A2 => n11174, B1 => n14072, B2 => 
                           n11171, C1 => n14008, C2 => n11168, ZN => n3172);
   U2628 : OAI222_X1 port map( A1 => n14039, A2 => n10910, B1 => n14071, B2 => 
                           n10907, C1 => n14007, C2 => n10904, ZN => n4564);
   U2629 : OAI222_X1 port map( A1 => n14039, A2 => n11174, B1 => n14071, B2 => 
                           n11171, C1 => n14007, C2 => n11168, ZN => n3131);
   U2630 : OAI222_X1 port map( A1 => n14038, A2 => n10910, B1 => n14070, B2 => 
                           n10907, C1 => n14006, C2 => n10904, ZN => n4523);
   U2631 : OAI222_X1 port map( A1 => n14038, A2 => n11174, B1 => n14070, B2 => 
                           n11171, C1 => n14006, C2 => n11168, ZN => n3090);
   U2632 : OAI222_X1 port map( A1 => n14037, A2 => n10910, B1 => n14069, B2 => 
                           n10907, C1 => n14005, C2 => n10904, ZN => n4482);
   U2633 : OAI222_X1 port map( A1 => n14037, A2 => n11174, B1 => n14069, B2 => 
                           n11171, C1 => n14005, C2 => n11168, ZN => n3049);
   U2634 : OAI222_X1 port map( A1 => n14036, A2 => n10910, B1 => n14068, B2 => 
                           n10907, C1 => n14004, C2 => n10904, ZN => n4441);
   U2635 : OAI222_X1 port map( A1 => n14036, A2 => n11174, B1 => n14068, B2 => 
                           n11171, C1 => n14004, C2 => n11168, ZN => n3008);
   U2636 : OAI222_X1 port map( A1 => n14066, A2 => n10908, B1 => n14098, B2 => 
                           n10905, C1 => n14034, C2 => n10902, ZN => n5699);
   U2637 : OAI222_X1 port map( A1 => n14066, A2 => n11172, B1 => n14098, B2 => 
                           n11169, C1 => n14034, C2 => n11166, ZN => n4266);
   U2638 : OAI222_X1 port map( A1 => n14065, A2 => n10908, B1 => n14097, B2 => 
                           n10905, C1 => n14033, C2 => n10902, ZN => n5630);
   U2639 : OAI222_X1 port map( A1 => n14065, A2 => n11172, B1 => n14097, B2 => 
                           n11169, C1 => n14033, C2 => n11166, ZN => n4197);
   U2640 : OAI222_X1 port map( A1 => n14064, A2 => n10908, B1 => n14096, B2 => 
                           n10905, C1 => n14032, C2 => n10902, ZN => n5589);
   U2641 : OAI222_X1 port map( A1 => n14064, A2 => n11172, B1 => n14096, B2 => 
                           n11169, C1 => n14032, C2 => n11166, ZN => n4156);
   U2642 : OAI222_X1 port map( A1 => n14063, A2 => n10908, B1 => n14095, B2 => 
                           n10905, C1 => n14031, C2 => n10902, ZN => n5548);
   U2643 : OAI222_X1 port map( A1 => n14063, A2 => n11172, B1 => n14095, B2 => 
                           n11169, C1 => n14031, C2 => n11166, ZN => n4115);
   U2644 : OAI222_X1 port map( A1 => n14062, A2 => n10908, B1 => n14094, B2 => 
                           n10905, C1 => n14030, C2 => n10902, ZN => n5507);
   U2645 : OAI222_X1 port map( A1 => n14062, A2 => n11172, B1 => n14094, B2 => 
                           n11169, C1 => n14030, C2 => n11166, ZN => n4074);
   U2646 : OAI222_X1 port map( A1 => n14061, A2 => n10908, B1 => n14093, B2 => 
                           n10905, C1 => n14029, C2 => n10902, ZN => n5466);
   U2647 : OAI222_X1 port map( A1 => n14061, A2 => n11172, B1 => n14093, B2 => 
                           n11169, C1 => n14029, C2 => n11166, ZN => n4033);
   U2648 : OAI222_X1 port map( A1 => n14060, A2 => n10908, B1 => n14092, B2 => 
                           n10905, C1 => n14028, C2 => n10902, ZN => n5425);
   U2649 : OAI222_X1 port map( A1 => n14060, A2 => n11172, B1 => n14092, B2 => 
                           n11169, C1 => n14028, C2 => n11166, ZN => n3992);
   U2650 : OAI222_X1 port map( A1 => n14059, A2 => n10908, B1 => n14091, B2 => 
                           n10905, C1 => n14027, C2 => n10902, ZN => n5384);
   U2651 : OAI222_X1 port map( A1 => n14059, A2 => n11172, B1 => n14091, B2 => 
                           n11169, C1 => n14027, C2 => n11166, ZN => n3951);
   U2652 : OAI222_X1 port map( A1 => n14058, A2 => n10908, B1 => n14090, B2 => 
                           n10905, C1 => n14026, C2 => n10902, ZN => n5343);
   U2653 : OAI222_X1 port map( A1 => n14058, A2 => n11172, B1 => n14090, B2 => 
                           n11169, C1 => n14026, C2 => n11166, ZN => n3910);
   U2654 : OAI222_X1 port map( A1 => n14057, A2 => n10908, B1 => n14089, B2 => 
                           n10905, C1 => n14025, C2 => n10902, ZN => n5302);
   U2655 : OAI222_X1 port map( A1 => n14057, A2 => n11172, B1 => n14089, B2 => 
                           n11169, C1 => n14025, C2 => n11166, ZN => n3869);
   U2656 : OAI222_X1 port map( A1 => n14056, A2 => n10908, B1 => n14088, B2 => 
                           n10905, C1 => n14024, C2 => n10902, ZN => n5261);
   U2657 : OAI222_X1 port map( A1 => n14056, A2 => n11172, B1 => n14088, B2 => 
                           n11169, C1 => n14024, C2 => n11166, ZN => n3828);
   U2658 : OAI222_X1 port map( A1 => n14055, A2 => n10908, B1 => n14087, B2 => 
                           n10905, C1 => n14023, C2 => n10902, ZN => n5220);
   U2659 : OAI222_X1 port map( A1 => n14055, A2 => n11172, B1 => n14087, B2 => 
                           n11169, C1 => n14023, C2 => n11166, ZN => n3787);
   U2660 : OAI222_X1 port map( A1 => n14054, A2 => n10909, B1 => n14086, B2 => 
                           n10906, C1 => n14022, C2 => n10903, ZN => n5179);
   U2661 : OAI222_X1 port map( A1 => n14054, A2 => n11173, B1 => n14086, B2 => 
                           n11170, C1 => n14022, C2 => n11167, ZN => n3746);
   U2662 : OAI222_X1 port map( A1 => n14053, A2 => n10909, B1 => n14085, B2 => 
                           n10906, C1 => n14021, C2 => n10903, ZN => n5138);
   U2663 : OAI222_X1 port map( A1 => n14053, A2 => n11173, B1 => n14085, B2 => 
                           n11170, C1 => n14021, C2 => n11167, ZN => n3705);
   U2664 : OAI222_X1 port map( A1 => n14052, A2 => n10909, B1 => n14084, B2 => 
                           n10906, C1 => n14020, C2 => n10903, ZN => n5097);
   U2665 : OAI222_X1 port map( A1 => n14052, A2 => n11173, B1 => n14084, B2 => 
                           n11170, C1 => n14020, C2 => n11167, ZN => n3664);
   U2666 : OAI222_X1 port map( A1 => n14051, A2 => n10909, B1 => n14083, B2 => 
                           n10906, C1 => n14019, C2 => n10903, ZN => n5056);
   U2667 : OAI222_X1 port map( A1 => n14051, A2 => n11173, B1 => n14083, B2 => 
                           n11170, C1 => n14019, C2 => n11167, ZN => n3623);
   U2668 : OAI222_X1 port map( A1 => n14050, A2 => n10909, B1 => n14082, B2 => 
                           n10906, C1 => n14018, C2 => n10903, ZN => n5015);
   U2669 : OAI222_X1 port map( A1 => n14050, A2 => n11173, B1 => n14082, B2 => 
                           n11170, C1 => n14018, C2 => n11167, ZN => n3582);
   U2670 : OAI222_X1 port map( A1 => n14049, A2 => n10909, B1 => n14081, B2 => 
                           n10906, C1 => n14017, C2 => n10903, ZN => n4974);
   U2671 : OAI222_X1 port map( A1 => n14049, A2 => n11173, B1 => n14081, B2 => 
                           n11170, C1 => n14017, C2 => n11167, ZN => n3541);
   U2672 : OAI222_X1 port map( A1 => n14048, A2 => n10909, B1 => n14080, B2 => 
                           n10906, C1 => n14016, C2 => n10903, ZN => n4933);
   U2673 : OAI222_X1 port map( A1 => n14048, A2 => n11173, B1 => n14080, B2 => 
                           n11170, C1 => n14016, C2 => n11167, ZN => n3500);
   U2674 : OAI222_X1 port map( A1 => n14047, A2 => n10909, B1 => n14079, B2 => 
                           n10906, C1 => n14015, C2 => n10903, ZN => n4892);
   U2675 : OAI222_X1 port map( A1 => n14047, A2 => n11173, B1 => n14079, B2 => 
                           n11170, C1 => n14015, C2 => n11167, ZN => n3459);
   U2676 : OAI222_X1 port map( A1 => n14046, A2 => n10909, B1 => n14078, B2 => 
                           n10906, C1 => n14014, C2 => n10903, ZN => n4851);
   U2677 : OAI222_X1 port map( A1 => n14046, A2 => n11173, B1 => n14078, B2 => 
                           n11170, C1 => n14014, C2 => n11167, ZN => n3418);
   U2678 : OAI222_X1 port map( A1 => n14045, A2 => n10909, B1 => n14077, B2 => 
                           n10906, C1 => n14013, C2 => n10903, ZN => n4810);
   U2679 : OAI222_X1 port map( A1 => n14045, A2 => n11173, B1 => n14077, B2 => 
                           n11170, C1 => n14013, C2 => n11167, ZN => n3377);
   U2680 : OAI222_X1 port map( A1 => n14044, A2 => n10909, B1 => n14076, B2 => 
                           n10906, C1 => n14012, C2 => n10903, ZN => n4769);
   U2681 : OAI222_X1 port map( A1 => n14044, A2 => n11173, B1 => n14076, B2 => 
                           n11170, C1 => n14012, C2 => n11167, ZN => n3336);
   U2682 : OAI222_X1 port map( A1 => n14043, A2 => n10909, B1 => n14075, B2 => 
                           n10906, C1 => n14011, C2 => n10903, ZN => n4728);
   U2683 : OAI222_X1 port map( A1 => n14043, A2 => n11173, B1 => n14075, B2 => 
                           n11170, C1 => n14011, C2 => n11167, ZN => n3295);
   U2684 : OAI222_X1 port map( A1 => n13147, A2 => n11009, B1 => n13179, B2 => 
                           n11006, C1 => n13115, C2 => n11003, ZN => n4671);
   U2685 : OAI222_X1 port map( A1 => n13147, A2 => n11273, B1 => n13179, B2 => 
                           n11270, C1 => n13115, C2 => n11267, ZN => n3238);
   U2686 : OAI222_X1 port map( A1 => n13146, A2 => n11009, B1 => n13178, B2 => 
                           n11006, C1 => n13114, C2 => n11003, ZN => n4630);
   U2687 : OAI222_X1 port map( A1 => n13146, A2 => n11273, B1 => n13178, B2 => 
                           n11270, C1 => n13114, C2 => n11267, ZN => n3197);
   U2688 : OAI222_X1 port map( A1 => n13145, A2 => n11009, B1 => n13177, B2 => 
                           n11006, C1 => n13113, C2 => n11003, ZN => n4589);
   U2689 : OAI222_X1 port map( A1 => n13145, A2 => n11273, B1 => n13177, B2 => 
                           n11270, C1 => n13113, C2 => n11267, ZN => n3156);
   U2690 : OAI222_X1 port map( A1 => n13144, A2 => n11009, B1 => n13176, B2 => 
                           n11006, C1 => n13112, C2 => n11003, ZN => n4548);
   U2691 : OAI222_X1 port map( A1 => n13144, A2 => n11273, B1 => n13176, B2 => 
                           n11270, C1 => n13112, C2 => n11267, ZN => n3115);
   U2692 : OAI222_X1 port map( A1 => n13143, A2 => n11009, B1 => n13175, B2 => 
                           n11006, C1 => n13111, C2 => n11003, ZN => n4507);
   U2693 : OAI222_X1 port map( A1 => n13143, A2 => n11273, B1 => n13175, B2 => 
                           n11270, C1 => n13111, C2 => n11267, ZN => n3074);
   U2694 : OAI222_X1 port map( A1 => n13142, A2 => n11009, B1 => n13174, B2 => 
                           n11006, C1 => n13110, C2 => n11003, ZN => n4466);
   U2695 : OAI222_X1 port map( A1 => n13142, A2 => n11273, B1 => n13174, B2 => 
                           n11270, C1 => n13110, C2 => n11267, ZN => n3033);
   U2696 : OAI222_X1 port map( A1 => n13141, A2 => n11009, B1 => n13173, B2 => 
                           n11006, C1 => n13109, C2 => n11003, ZN => n4425);
   U2697 : OAI222_X1 port map( A1 => n13141, A2 => n11273, B1 => n13173, B2 => 
                           n11270, C1 => n13109, C2 => n11267, ZN => n2992);
   U2698 : OAI222_X1 port map( A1 => n13140, A2 => n11009, B1 => n13172, B2 => 
                           n11006, C1 => n13108, C2 => n11003, ZN => n4331);
   U2699 : OAI222_X1 port map( A1 => n13140, A2 => n11273, B1 => n13172, B2 => 
                           n11270, C1 => n13108, C2 => n11267, ZN => n2863);
   U2700 : OAI222_X1 port map( A1 => n13171, A2 => n11007, B1 => n13203, B2 => 
                           n11004, C1 => n13139, C2 => n11001, ZN => n5677);
   U2701 : OAI222_X1 port map( A1 => n13171, A2 => n11271, B1 => n13203, B2 => 
                           n11268, C1 => n13139, C2 => n11265, ZN => n4244);
   U2702 : OAI222_X1 port map( A1 => n13170, A2 => n11007, B1 => n13202, B2 => 
                           n11004, C1 => n13138, C2 => n11001, ZN => n5614);
   U2703 : OAI222_X1 port map( A1 => n13170, A2 => n11271, B1 => n13202, B2 => 
                           n11268, C1 => n13138, C2 => n11265, ZN => n4181);
   U2704 : OAI222_X1 port map( A1 => n13169, A2 => n11007, B1 => n13201, B2 => 
                           n11004, C1 => n13137, C2 => n11001, ZN => n5573);
   U2705 : OAI222_X1 port map( A1 => n13169, A2 => n11271, B1 => n13201, B2 => 
                           n11268, C1 => n13137, C2 => n11265, ZN => n4140);
   U2706 : OAI222_X1 port map( A1 => n13168, A2 => n11007, B1 => n13200, B2 => 
                           n11004, C1 => n13136, C2 => n11001, ZN => n5532);
   U2707 : OAI222_X1 port map( A1 => n13168, A2 => n11271, B1 => n13200, B2 => 
                           n11268, C1 => n13136, C2 => n11265, ZN => n4099);
   U2708 : OAI222_X1 port map( A1 => n13167, A2 => n11007, B1 => n13199, B2 => 
                           n11004, C1 => n13135, C2 => n11001, ZN => n5491);
   U2709 : OAI222_X1 port map( A1 => n13167, A2 => n11271, B1 => n13199, B2 => 
                           n11268, C1 => n13135, C2 => n11265, ZN => n4058);
   U2710 : OAI222_X1 port map( A1 => n13166, A2 => n11007, B1 => n13198, B2 => 
                           n11004, C1 => n13134, C2 => n11001, ZN => n5450);
   U2711 : OAI222_X1 port map( A1 => n13166, A2 => n11271, B1 => n13198, B2 => 
                           n11268, C1 => n13134, C2 => n11265, ZN => n4017);
   U2712 : OAI222_X1 port map( A1 => n13165, A2 => n11007, B1 => n13197, B2 => 
                           n11004, C1 => n13133, C2 => n11001, ZN => n5409);
   U2713 : OAI222_X1 port map( A1 => n13165, A2 => n11271, B1 => n13197, B2 => 
                           n11268, C1 => n13133, C2 => n11265, ZN => n3976);
   U2714 : OAI222_X1 port map( A1 => n13164, A2 => n11007, B1 => n13196, B2 => 
                           n11004, C1 => n13132, C2 => n11001, ZN => n5368);
   U2715 : OAI222_X1 port map( A1 => n13164, A2 => n11271, B1 => n13196, B2 => 
                           n11268, C1 => n13132, C2 => n11265, ZN => n3935);
   U2716 : OAI222_X1 port map( A1 => n13163, A2 => n11007, B1 => n13195, B2 => 
                           n11004, C1 => n13131, C2 => n11001, ZN => n5327);
   U2717 : OAI222_X1 port map( A1 => n13163, A2 => n11271, B1 => n13195, B2 => 
                           n11268, C1 => n13131, C2 => n11265, ZN => n3894);
   U2718 : OAI222_X1 port map( A1 => n13162, A2 => n11007, B1 => n13194, B2 => 
                           n11004, C1 => n13130, C2 => n11001, ZN => n5286);
   U2719 : OAI222_X1 port map( A1 => n13162, A2 => n11271, B1 => n13194, B2 => 
                           n11268, C1 => n13130, C2 => n11265, ZN => n3853);
   U2720 : OAI222_X1 port map( A1 => n13161, A2 => n11007, B1 => n13193, B2 => 
                           n11004, C1 => n13129, C2 => n11001, ZN => n5245);
   U2721 : OAI222_X1 port map( A1 => n13161, A2 => n11271, B1 => n13193, B2 => 
                           n11268, C1 => n13129, C2 => n11265, ZN => n3812);
   U2722 : OAI222_X1 port map( A1 => n13160, A2 => n11007, B1 => n13192, B2 => 
                           n11004, C1 => n13128, C2 => n11001, ZN => n5204);
   U2723 : OAI222_X1 port map( A1 => n13160, A2 => n11271, B1 => n13192, B2 => 
                           n11268, C1 => n13128, C2 => n11265, ZN => n3771);
   U2724 : OAI222_X1 port map( A1 => n13159, A2 => n11008, B1 => n13191, B2 => 
                           n11005, C1 => n13127, C2 => n11002, ZN => n5163);
   U2725 : OAI222_X1 port map( A1 => n13159, A2 => n11272, B1 => n13191, B2 => 
                           n11269, C1 => n13127, C2 => n11266, ZN => n3730);
   U2726 : OAI222_X1 port map( A1 => n13158, A2 => n11008, B1 => n13190, B2 => 
                           n11005, C1 => n13126, C2 => n11002, ZN => n5122);
   U2727 : OAI222_X1 port map( A1 => n13158, A2 => n11272, B1 => n13190, B2 => 
                           n11269, C1 => n13126, C2 => n11266, ZN => n3689);
   U2728 : OAI222_X1 port map( A1 => n13157, A2 => n11008, B1 => n13189, B2 => 
                           n11005, C1 => n13125, C2 => n11002, ZN => n5081);
   U2729 : OAI222_X1 port map( A1 => n13157, A2 => n11272, B1 => n13189, B2 => 
                           n11269, C1 => n13125, C2 => n11266, ZN => n3648);
   U2730 : OAI222_X1 port map( A1 => n13156, A2 => n11008, B1 => n13188, B2 => 
                           n11005, C1 => n13124, C2 => n11002, ZN => n5040);
   U2731 : OAI222_X1 port map( A1 => n13156, A2 => n11272, B1 => n13188, B2 => 
                           n11269, C1 => n13124, C2 => n11266, ZN => n3607);
   U2732 : OAI222_X1 port map( A1 => n13155, A2 => n11008, B1 => n13187, B2 => 
                           n11005, C1 => n13123, C2 => n11002, ZN => n4999);
   U2733 : OAI222_X1 port map( A1 => n13155, A2 => n11272, B1 => n13187, B2 => 
                           n11269, C1 => n13123, C2 => n11266, ZN => n3566);
   U2734 : OAI222_X1 port map( A1 => n13154, A2 => n11008, B1 => n13186, B2 => 
                           n11005, C1 => n13122, C2 => n11002, ZN => n4958);
   U2735 : OAI222_X1 port map( A1 => n13154, A2 => n11272, B1 => n13186, B2 => 
                           n11269, C1 => n13122, C2 => n11266, ZN => n3525);
   U2736 : OAI222_X1 port map( A1 => n13153, A2 => n11008, B1 => n13185, B2 => 
                           n11005, C1 => n13121, C2 => n11002, ZN => n4917);
   U2737 : OAI222_X1 port map( A1 => n13153, A2 => n11272, B1 => n13185, B2 => 
                           n11269, C1 => n13121, C2 => n11266, ZN => n3484);
   U2738 : OAI222_X1 port map( A1 => n13152, A2 => n11008, B1 => n13184, B2 => 
                           n11005, C1 => n13120, C2 => n11002, ZN => n4876);
   U2739 : OAI222_X1 port map( A1 => n13152, A2 => n11272, B1 => n13184, B2 => 
                           n11269, C1 => n13120, C2 => n11266, ZN => n3443);
   U2740 : OAI222_X1 port map( A1 => n13151, A2 => n11008, B1 => n13183, B2 => 
                           n11005, C1 => n13119, C2 => n11002, ZN => n4835);
   U2741 : OAI222_X1 port map( A1 => n13151, A2 => n11272, B1 => n13183, B2 => 
                           n11269, C1 => n13119, C2 => n11266, ZN => n3402);
   U2742 : OAI222_X1 port map( A1 => n13150, A2 => n11008, B1 => n13182, B2 => 
                           n11005, C1 => n13118, C2 => n11002, ZN => n4794);
   U2743 : OAI222_X1 port map( A1 => n13150, A2 => n11272, B1 => n13182, B2 => 
                           n11269, C1 => n13118, C2 => n11266, ZN => n3361);
   U2744 : OAI222_X1 port map( A1 => n13149, A2 => n11008, B1 => n13181, B2 => 
                           n11005, C1 => n13117, C2 => n11002, ZN => n4753);
   U2745 : OAI222_X1 port map( A1 => n13149, A2 => n11272, B1 => n13181, B2 => 
                           n11269, C1 => n13117, C2 => n11266, ZN => n3320);
   U2746 : OAI222_X1 port map( A1 => n13148, A2 => n11008, B1 => n13180, B2 => 
                           n11005, C1 => n13116, C2 => n11002, ZN => n4712);
   U2747 : OAI222_X1 port map( A1 => n13148, A2 => n11272, B1 => n13180, B2 => 
                           n11269, C1 => n13116, C2 => n11266, ZN => n3279);
   U2748 : OAI222_X1 port map( A1 => n13467, A2 => n11024, B1 => n13403, B2 => 
                           n11021, C1 => n13435, C2 => n11018, ZN => n4667);
   U2749 : OAI222_X1 port map( A1 => n13467, A2 => n11288, B1 => n13403, B2 => 
                           n11285, C1 => n13435, C2 => n11282, ZN => n3234);
   U2750 : OAI222_X1 port map( A1 => n13466, A2 => n11024, B1 => n13402, B2 => 
                           n11021, C1 => n13434, C2 => n11018, ZN => n4626);
   U2751 : OAI222_X1 port map( A1 => n13466, A2 => n11288, B1 => n13402, B2 => 
                           n11285, C1 => n13434, C2 => n11282, ZN => n3193);
   U2752 : OAI222_X1 port map( A1 => n13465, A2 => n11024, B1 => n13401, B2 => 
                           n11021, C1 => n13433, C2 => n11018, ZN => n4585);
   U2753 : OAI222_X1 port map( A1 => n13465, A2 => n11288, B1 => n13401, B2 => 
                           n11285, C1 => n13433, C2 => n11282, ZN => n3152);
   U2754 : OAI222_X1 port map( A1 => n13464, A2 => n11024, B1 => n13400, B2 => 
                           n11021, C1 => n13432, C2 => n11018, ZN => n4544);
   U2755 : OAI222_X1 port map( A1 => n13464, A2 => n11288, B1 => n13400, B2 => 
                           n11285, C1 => n13432, C2 => n11282, ZN => n3111);
   U2756 : OAI222_X1 port map( A1 => n13463, A2 => n11024, B1 => n13399, B2 => 
                           n11021, C1 => n13431, C2 => n11018, ZN => n4503);
   U2757 : OAI222_X1 port map( A1 => n13463, A2 => n11288, B1 => n13399, B2 => 
                           n11285, C1 => n13431, C2 => n11282, ZN => n3070);
   U2758 : OAI222_X1 port map( A1 => n13462, A2 => n11024, B1 => n13398, B2 => 
                           n11021, C1 => n13430, C2 => n11018, ZN => n4462);
   U2759 : OAI222_X1 port map( A1 => n13462, A2 => n11288, B1 => n13398, B2 => 
                           n11285, C1 => n13430, C2 => n11282, ZN => n3029);
   U2760 : OAI222_X1 port map( A1 => n13461, A2 => n11024, B1 => n13397, B2 => 
                           n11021, C1 => n13429, C2 => n11018, ZN => n4421);
   U2761 : OAI222_X1 port map( A1 => n13461, A2 => n11288, B1 => n13397, B2 => 
                           n11285, C1 => n13429, C2 => n11282, ZN => n2988);
   U2762 : OAI222_X1 port map( A1 => n13460, A2 => n11024, B1 => n13396, B2 => 
                           n11021, C1 => n13428, C2 => n11018, ZN => n4314);
   U2763 : OAI222_X1 port map( A1 => n13460, A2 => n11288, B1 => n13396, B2 => 
                           n11285, C1 => n13428, C2 => n11282, ZN => n2814);
   U2764 : OAI222_X1 port map( A1 => n13491, A2 => n11022, B1 => n13427, B2 => 
                           n11019, C1 => n13459, C2 => n11016, ZN => n5670);
   U2765 : OAI222_X1 port map( A1 => n13491, A2 => n11286, B1 => n13427, B2 => 
                           n11283, C1 => n13459, C2 => n11280, ZN => n4237);
   U2766 : OAI222_X1 port map( A1 => n13490, A2 => n11022, B1 => n13426, B2 => 
                           n11019, C1 => n13458, C2 => n11016, ZN => n5610);
   U2767 : OAI222_X1 port map( A1 => n13490, A2 => n11286, B1 => n13426, B2 => 
                           n11283, C1 => n13458, C2 => n11280, ZN => n4177);
   U2768 : OAI222_X1 port map( A1 => n13489, A2 => n11022, B1 => n13425, B2 => 
                           n11019, C1 => n13457, C2 => n11016, ZN => n5569);
   U2769 : OAI222_X1 port map( A1 => n13489, A2 => n11286, B1 => n13425, B2 => 
                           n11283, C1 => n13457, C2 => n11280, ZN => n4136);
   U2770 : OAI222_X1 port map( A1 => n13488, A2 => n11022, B1 => n13424, B2 => 
                           n11019, C1 => n13456, C2 => n11016, ZN => n5528);
   U2771 : OAI222_X1 port map( A1 => n13488, A2 => n11286, B1 => n13424, B2 => 
                           n11283, C1 => n13456, C2 => n11280, ZN => n4095);
   U2772 : OAI222_X1 port map( A1 => n13487, A2 => n11022, B1 => n13423, B2 => 
                           n11019, C1 => n13455, C2 => n11016, ZN => n5487);
   U2773 : OAI222_X1 port map( A1 => n13487, A2 => n11286, B1 => n13423, B2 => 
                           n11283, C1 => n13455, C2 => n11280, ZN => n4054);
   U2774 : OAI222_X1 port map( A1 => n13486, A2 => n11022, B1 => n13422, B2 => 
                           n11019, C1 => n13454, C2 => n11016, ZN => n5446);
   U2775 : OAI222_X1 port map( A1 => n13486, A2 => n11286, B1 => n13422, B2 => 
                           n11283, C1 => n13454, C2 => n11280, ZN => n4013);
   U2776 : OAI222_X1 port map( A1 => n13485, A2 => n11022, B1 => n13421, B2 => 
                           n11019, C1 => n13453, C2 => n11016, ZN => n5405);
   U2777 : OAI222_X1 port map( A1 => n13485, A2 => n11286, B1 => n13421, B2 => 
                           n11283, C1 => n13453, C2 => n11280, ZN => n3972);
   U2778 : OAI222_X1 port map( A1 => n13484, A2 => n11022, B1 => n13420, B2 => 
                           n11019, C1 => n13452, C2 => n11016, ZN => n5364);
   U2779 : OAI222_X1 port map( A1 => n13484, A2 => n11286, B1 => n13420, B2 => 
                           n11283, C1 => n13452, C2 => n11280, ZN => n3931);
   U2780 : OAI222_X1 port map( A1 => n13483, A2 => n11022, B1 => n13419, B2 => 
                           n11019, C1 => n13451, C2 => n11016, ZN => n5323);
   U2781 : OAI222_X1 port map( A1 => n13483, A2 => n11286, B1 => n13419, B2 => 
                           n11283, C1 => n13451, C2 => n11280, ZN => n3890);
   U2782 : OAI222_X1 port map( A1 => n13482, A2 => n11022, B1 => n13418, B2 => 
                           n11019, C1 => n13450, C2 => n11016, ZN => n5282);
   U2783 : OAI222_X1 port map( A1 => n13482, A2 => n11286, B1 => n13418, B2 => 
                           n11283, C1 => n13450, C2 => n11280, ZN => n3849);
   U2784 : OAI222_X1 port map( A1 => n13481, A2 => n11022, B1 => n13417, B2 => 
                           n11019, C1 => n13449, C2 => n11016, ZN => n5241);
   U2785 : OAI222_X1 port map( A1 => n13481, A2 => n11286, B1 => n13417, B2 => 
                           n11283, C1 => n13449, C2 => n11280, ZN => n3808);
   U2786 : OAI222_X1 port map( A1 => n13480, A2 => n11022, B1 => n13416, B2 => 
                           n11019, C1 => n13448, C2 => n11016, ZN => n5200);
   U2787 : OAI222_X1 port map( A1 => n13480, A2 => n11286, B1 => n13416, B2 => 
                           n11283, C1 => n13448, C2 => n11280, ZN => n3767);
   U2788 : OAI222_X1 port map( A1 => n13479, A2 => n11023, B1 => n13415, B2 => 
                           n11020, C1 => n13447, C2 => n11017, ZN => n5159);
   U2789 : OAI222_X1 port map( A1 => n13479, A2 => n11287, B1 => n13415, B2 => 
                           n11284, C1 => n13447, C2 => n11281, ZN => n3726);
   U2790 : OAI222_X1 port map( A1 => n13478, A2 => n11023, B1 => n13414, B2 => 
                           n11020, C1 => n13446, C2 => n11017, ZN => n5118);
   U2791 : OAI222_X1 port map( A1 => n13478, A2 => n11287, B1 => n13414, B2 => 
                           n11284, C1 => n13446, C2 => n11281, ZN => n3685);
   U2792 : OAI222_X1 port map( A1 => n13477, A2 => n11023, B1 => n13413, B2 => 
                           n11020, C1 => n13445, C2 => n11017, ZN => n5077);
   U2793 : OAI222_X1 port map( A1 => n13477, A2 => n11287, B1 => n13413, B2 => 
                           n11284, C1 => n13445, C2 => n11281, ZN => n3644);
   U2794 : OAI222_X1 port map( A1 => n13476, A2 => n11023, B1 => n13412, B2 => 
                           n11020, C1 => n13444, C2 => n11017, ZN => n5036);
   U2795 : OAI222_X1 port map( A1 => n13476, A2 => n11287, B1 => n13412, B2 => 
                           n11284, C1 => n13444, C2 => n11281, ZN => n3603);
   U2796 : OAI222_X1 port map( A1 => n13475, A2 => n11023, B1 => n13411, B2 => 
                           n11020, C1 => n13443, C2 => n11017, ZN => n4995);
   U2797 : OAI222_X1 port map( A1 => n13475, A2 => n11287, B1 => n13411, B2 => 
                           n11284, C1 => n13443, C2 => n11281, ZN => n3562);
   U2798 : OAI222_X1 port map( A1 => n13474, A2 => n11023, B1 => n13410, B2 => 
                           n11020, C1 => n13442, C2 => n11017, ZN => n4954);
   U2799 : OAI222_X1 port map( A1 => n13474, A2 => n11287, B1 => n13410, B2 => 
                           n11284, C1 => n13442, C2 => n11281, ZN => n3521);
   U2800 : OAI222_X1 port map( A1 => n13473, A2 => n11023, B1 => n13409, B2 => 
                           n11020, C1 => n13441, C2 => n11017, ZN => n4913);
   U2801 : OAI222_X1 port map( A1 => n13473, A2 => n11287, B1 => n13409, B2 => 
                           n11284, C1 => n13441, C2 => n11281, ZN => n3480);
   U2802 : OAI222_X1 port map( A1 => n13472, A2 => n11023, B1 => n13408, B2 => 
                           n11020, C1 => n13440, C2 => n11017, ZN => n4872);
   U2803 : OAI222_X1 port map( A1 => n13472, A2 => n11287, B1 => n13408, B2 => 
                           n11284, C1 => n13440, C2 => n11281, ZN => n3439);
   U2804 : OAI222_X1 port map( A1 => n13471, A2 => n11023, B1 => n13407, B2 => 
                           n11020, C1 => n13439, C2 => n11017, ZN => n4831);
   U2805 : OAI222_X1 port map( A1 => n13471, A2 => n11287, B1 => n13407, B2 => 
                           n11284, C1 => n13439, C2 => n11281, ZN => n3398);
   U2806 : OAI222_X1 port map( A1 => n13470, A2 => n11023, B1 => n13406, B2 => 
                           n11020, C1 => n13438, C2 => n11017, ZN => n4790);
   U2807 : OAI222_X1 port map( A1 => n13470, A2 => n11287, B1 => n13406, B2 => 
                           n11284, C1 => n13438, C2 => n11281, ZN => n3357);
   U2808 : OAI222_X1 port map( A1 => n13469, A2 => n11023, B1 => n13405, B2 => 
                           n11020, C1 => n13437, C2 => n11017, ZN => n4749);
   U2809 : OAI222_X1 port map( A1 => n13469, A2 => n11287, B1 => n13405, B2 => 
                           n11284, C1 => n13437, C2 => n11281, ZN => n3316);
   U2810 : OAI222_X1 port map( A1 => n13468, A2 => n11023, B1 => n13404, B2 => 
                           n11020, C1 => n13436, C2 => n11017, ZN => n4708);
   U2811 : OAI222_X1 port map( A1 => n13468, A2 => n11287, B1 => n13404, B2 => 
                           n11284, C1 => n13436, C2 => n11281, ZN => n3275);
   U2812 : AOI222_X1 port map( A1 => n10857, A2 => n14320, B1 => n10854, B2 => 
                           n14352, C1 => n10851, C2 => n14416, ZN => n5693);
   U2813 : AOI222_X1 port map( A1 => n11121, A2 => n14320, B1 => n11118, B2 => 
                           n14352, C1 => n11115, C2 => n14416, ZN => n4260);
   U2814 : AOI222_X1 port map( A1 => n10857, A2 => n14319, B1 => n10854, B2 => 
                           n14351, C1 => n10851, C2 => n14415, ZN => n5624);
   U2815 : AOI222_X1 port map( A1 => n11121, A2 => n14319, B1 => n11118, B2 => 
                           n14351, C1 => n11115, C2 => n14415, ZN => n4191);
   U2816 : AOI222_X1 port map( A1 => n10857, A2 => n14318, B1 => n10854, B2 => 
                           n14350, C1 => n10851, C2 => n14414, ZN => n5583);
   U2817 : AOI222_X1 port map( A1 => n11121, A2 => n14318, B1 => n11118, B2 => 
                           n14350, C1 => n11115, C2 => n14414, ZN => n4150);
   U2818 : AOI222_X1 port map( A1 => n10857, A2 => n14317, B1 => n10854, B2 => 
                           n14349, C1 => n10851, C2 => n14413, ZN => n5542);
   U2819 : AOI222_X1 port map( A1 => n11121, A2 => n14317, B1 => n11118, B2 => 
                           n14349, C1 => n11115, C2 => n14413, ZN => n4109);
   U2820 : AOI222_X1 port map( A1 => n10857, A2 => n14316, B1 => n10854, B2 => 
                           n14348, C1 => n10851, C2 => n14412, ZN => n5501);
   U2821 : AOI222_X1 port map( A1 => n11121, A2 => n14316, B1 => n11118, B2 => 
                           n14348, C1 => n11115, C2 => n14412, ZN => n4068);
   U2822 : AOI222_X1 port map( A1 => n10857, A2 => n14315, B1 => n10854, B2 => 
                           n14347, C1 => n10851, C2 => n14411, ZN => n5460);
   U2823 : AOI222_X1 port map( A1 => n11121, A2 => n14315, B1 => n11118, B2 => 
                           n14347, C1 => n11115, C2 => n14411, ZN => n4027);
   U2824 : AOI222_X1 port map( A1 => n10857, A2 => n14314, B1 => n10854, B2 => 
                           n14346, C1 => n10851, C2 => n14410, ZN => n5419);
   U2825 : AOI222_X1 port map( A1 => n11121, A2 => n14314, B1 => n11118, B2 => 
                           n14346, C1 => n11115, C2 => n14410, ZN => n3986);
   U2826 : AOI222_X1 port map( A1 => n10857, A2 => n14313, B1 => n10854, B2 => 
                           n14345, C1 => n10851, C2 => n14409, ZN => n5378);
   U2827 : AOI222_X1 port map( A1 => n11121, A2 => n14313, B1 => n11118, B2 => 
                           n14345, C1 => n11115, C2 => n14409, ZN => n3945);
   U2828 : AOI222_X1 port map( A1 => n10857, A2 => n14312, B1 => n10854, B2 => 
                           n14344, C1 => n10851, C2 => n14408, ZN => n5337);
   U2829 : AOI222_X1 port map( A1 => n11121, A2 => n14312, B1 => n11118, B2 => 
                           n14344, C1 => n11115, C2 => n14408, ZN => n3904);
   U2830 : AOI222_X1 port map( A1 => n10857, A2 => n14311, B1 => n10854, B2 => 
                           n14343, C1 => n10851, C2 => n14407, ZN => n5296);
   U2831 : AOI222_X1 port map( A1 => n11121, A2 => n14311, B1 => n11118, B2 => 
                           n14343, C1 => n11115, C2 => n14407, ZN => n3863);
   U2832 : AOI222_X1 port map( A1 => n10857, A2 => n14310, B1 => n10854, B2 => 
                           n14342, C1 => n10851, C2 => n14406, ZN => n5255);
   U2833 : AOI222_X1 port map( A1 => n11121, A2 => n14310, B1 => n11118, B2 => 
                           n14342, C1 => n11115, C2 => n14406, ZN => n3822);
   U2834 : AOI222_X1 port map( A1 => n10857, A2 => n14309, B1 => n10854, B2 => 
                           n14341, C1 => n10851, C2 => n14405, ZN => n5214);
   U2835 : AOI222_X1 port map( A1 => n11121, A2 => n14309, B1 => n11118, B2 => 
                           n14341, C1 => n11115, C2 => n14405, ZN => n3781);
   U2836 : AOI222_X1 port map( A1 => n10858, A2 => n14308, B1 => n10855, B2 => 
                           n14340, C1 => n10852, C2 => n14404, ZN => n5173);
   U2837 : AOI222_X1 port map( A1 => n11122, A2 => n14308, B1 => n11119, B2 => 
                           n14340, C1 => n11116, C2 => n14404, ZN => n3740);
   U2838 : AOI222_X1 port map( A1 => n10858, A2 => n14307, B1 => n10855, B2 => 
                           n14339, C1 => n10852, C2 => n14403, ZN => n5132);
   U2839 : AOI222_X1 port map( A1 => n11122, A2 => n14307, B1 => n11119, B2 => 
                           n14339, C1 => n11116, C2 => n14403, ZN => n3699);
   U2840 : AOI222_X1 port map( A1 => n10858, A2 => n14306, B1 => n10855, B2 => 
                           n14338, C1 => n10852, C2 => n14402, ZN => n5091);
   U2841 : AOI222_X1 port map( A1 => n11122, A2 => n14306, B1 => n11119, B2 => 
                           n14338, C1 => n11116, C2 => n14402, ZN => n3658);
   U2842 : AOI222_X1 port map( A1 => n10858, A2 => n14305, B1 => n10855, B2 => 
                           n14337, C1 => n10852, C2 => n14401, ZN => n5050);
   U2843 : AOI222_X1 port map( A1 => n11122, A2 => n14305, B1 => n11119, B2 => 
                           n14337, C1 => n11116, C2 => n14401, ZN => n3617);
   U2844 : AOI222_X1 port map( A1 => n10858, A2 => n14304, B1 => n10855, B2 => 
                           n14336, C1 => n10852, C2 => n14400, ZN => n5009);
   U2845 : AOI222_X1 port map( A1 => n11122, A2 => n14304, B1 => n11119, B2 => 
                           n14336, C1 => n11116, C2 => n14400, ZN => n3576);
   U2846 : AOI222_X1 port map( A1 => n10858, A2 => n14303, B1 => n10855, B2 => 
                           n14335, C1 => n10852, C2 => n14399, ZN => n4968);
   U2847 : AOI222_X1 port map( A1 => n11122, A2 => n14303, B1 => n11119, B2 => 
                           n14335, C1 => n11116, C2 => n14399, ZN => n3535);
   U2848 : AOI222_X1 port map( A1 => n10858, A2 => n14302, B1 => n10855, B2 => 
                           n14334, C1 => n10852, C2 => n14398, ZN => n4927);
   U2849 : AOI222_X1 port map( A1 => n11122, A2 => n14302, B1 => n11119, B2 => 
                           n14334, C1 => n11116, C2 => n14398, ZN => n3494);
   U2850 : AOI222_X1 port map( A1 => n10858, A2 => n14301, B1 => n10855, B2 => 
                           n14333, C1 => n10852, C2 => n14397, ZN => n4886);
   U2851 : AOI222_X1 port map( A1 => n11122, A2 => n14301, B1 => n11119, B2 => 
                           n14333, C1 => n11116, C2 => n14397, ZN => n3453);
   U2852 : AOI222_X1 port map( A1 => n10858, A2 => n14300, B1 => n10855, B2 => 
                           n14332, C1 => n10852, C2 => n14396, ZN => n4845);
   U2853 : AOI222_X1 port map( A1 => n11122, A2 => n14300, B1 => n11119, B2 => 
                           n14332, C1 => n11116, C2 => n14396, ZN => n3412);
   U2854 : AOI222_X1 port map( A1 => n10858, A2 => n14299, B1 => n10855, B2 => 
                           n14331, C1 => n10852, C2 => n14395, ZN => n4804);
   U2855 : AOI222_X1 port map( A1 => n11122, A2 => n14299, B1 => n11119, B2 => 
                           n14331, C1 => n11116, C2 => n14395, ZN => n3371);
   U2856 : AOI222_X1 port map( A1 => n10858, A2 => n14298, B1 => n10855, B2 => 
                           n14330, C1 => n10852, C2 => n14394, ZN => n4763);
   U2857 : AOI222_X1 port map( A1 => n11122, A2 => n14298, B1 => n11119, B2 => 
                           n14330, C1 => n11116, C2 => n14394, ZN => n3330);
   U2858 : AOI222_X1 port map( A1 => n10858, A2 => n14297, B1 => n10855, B2 => 
                           n14329, C1 => n10852, C2 => n14393, ZN => n4722);
   U2859 : AOI222_X1 port map( A1 => n11122, A2 => n14297, B1 => n11119, B2 => 
                           n14329, C1 => n11116, C2 => n14393, ZN => n3289);
   U2860 : AOI222_X1 port map( A1 => n10859, A2 => n14296, B1 => n10856, B2 => 
                           n14328, C1 => n10853, C2 => n14392, ZN => n4681);
   U2861 : AOI222_X1 port map( A1 => n11123, A2 => n14296, B1 => n11120, B2 => 
                           n14328, C1 => n11117, C2 => n14392, ZN => n3248);
   U2862 : AOI222_X1 port map( A1 => n10859, A2 => n14295, B1 => n10856, B2 => 
                           n14327, C1 => n10853, C2 => n14391, ZN => n4640);
   U2863 : AOI222_X1 port map( A1 => n11123, A2 => n14295, B1 => n11120, B2 => 
                           n14327, C1 => n11117, C2 => n14391, ZN => n3207);
   U2864 : AOI222_X1 port map( A1 => n10859, A2 => n14294, B1 => n10856, B2 => 
                           n14326, C1 => n10853, C2 => n14390, ZN => n4599);
   U2865 : AOI222_X1 port map( A1 => n11123, A2 => n14294, B1 => n11120, B2 => 
                           n14326, C1 => n11117, C2 => n14390, ZN => n3166);
   U2866 : AOI222_X1 port map( A1 => n10859, A2 => n14293, B1 => n10856, B2 => 
                           n14325, C1 => n10853, C2 => n14389, ZN => n4558);
   U2867 : AOI222_X1 port map( A1 => n11123, A2 => n14293, B1 => n11120, B2 => 
                           n14325, C1 => n11117, C2 => n14389, ZN => n3125);
   U2868 : AOI222_X1 port map( A1 => n10859, A2 => n14292, B1 => n10856, B2 => 
                           n14324, C1 => n10853, C2 => n14388, ZN => n4517);
   U2869 : AOI222_X1 port map( A1 => n11123, A2 => n14292, B1 => n11120, B2 => 
                           n14324, C1 => n11117, C2 => n14388, ZN => n3084);
   U2870 : AOI222_X1 port map( A1 => n10859, A2 => n14291, B1 => n10856, B2 => 
                           n14323, C1 => n10853, C2 => n14387, ZN => n4476);
   U2871 : AOI222_X1 port map( A1 => n11123, A2 => n14291, B1 => n11120, B2 => 
                           n14323, C1 => n11117, C2 => n14387, ZN => n3043);
   U2872 : AOI222_X1 port map( A1 => n10859, A2 => n14290, B1 => n10856, B2 => 
                           n14322, C1 => n10853, C2 => n14386, ZN => n4435);
   U2873 : AOI222_X1 port map( A1 => n11123, A2 => n14290, B1 => n11120, B2 => 
                           n14322, C1 => n11117, C2 => n14386, ZN => n3002);
   U2874 : AOI222_X1 port map( A1 => n10859, A2 => n14289, B1 => n10856, B2 => 
                           n14321, C1 => n10853, C2 => n14385, ZN => n4372);
   U2875 : AOI222_X1 port map( A1 => n11123, A2 => n14289, B1 => n11120, B2 => 
                           n14321, C1 => n11117, C2 => n14385, ZN => n2939);
   U2876 : NOR3_X1 port map( A1 => n14514, A2 => n12769, A3 => n12771, ZN => 
                           n5706);
   U2877 : NOR3_X1 port map( A1 => n14516, A2 => n12773, A3 => n12775, ZN => 
                           n4273);
   U2878 : NOR2_X1 port map( A1 => n2597, A2 => N2173, ZN => n2615);
   U2879 : BUF_X1 port map( A => n12768, Z => n10844);
   U2880 : BUF_X1 port map( A => n12767, Z => n10837);
   U2881 : BUF_X1 port map( A => n12766, Z => n10830);
   U2882 : BUF_X1 port map( A => n12765, Z => n10823);
   U2883 : BUF_X1 port map( A => n12764, Z => n10816);
   U2884 : BUF_X1 port map( A => n12763, Z => n10809);
   U2885 : BUF_X1 port map( A => n12762, Z => n10802);
   U2886 : BUF_X1 port map( A => n12761, Z => n10795);
   U2887 : BUF_X1 port map( A => n12760, Z => n10788);
   U2888 : BUF_X1 port map( A => n12759, Z => n10781);
   U2889 : BUF_X1 port map( A => n12758, Z => n10774);
   U2890 : BUF_X1 port map( A => n12757, Z => n10767);
   U2891 : BUF_X1 port map( A => n12756, Z => n10760);
   U2892 : BUF_X1 port map( A => n12755, Z => n10753);
   U2893 : BUF_X1 port map( A => n12754, Z => n10746);
   U2894 : BUF_X1 port map( A => n12753, Z => n10739);
   U2895 : BUF_X1 port map( A => n12752, Z => n10732);
   U2896 : BUF_X1 port map( A => n12751, Z => n10725);
   U2897 : BUF_X1 port map( A => n12750, Z => n10718);
   U2898 : BUF_X1 port map( A => n12749, Z => n10711);
   U2899 : BUF_X1 port map( A => n12748, Z => n10704);
   U2900 : BUF_X1 port map( A => n12747, Z => n10697);
   U2901 : BUF_X1 port map( A => n12746, Z => n10690);
   U2902 : BUF_X1 port map( A => n12745, Z => n10683);
   U2903 : BUF_X1 port map( A => n12744, Z => n10676);
   U2904 : BUF_X1 port map( A => n12743, Z => n10669);
   U2905 : BUF_X1 port map( A => n12742, Z => n10662);
   U2906 : BUF_X1 port map( A => n12741, Z => n10655);
   U2907 : BUF_X1 port map( A => n12740, Z => n10648);
   U2908 : BUF_X1 port map( A => n12739, Z => n10641);
   U2909 : BUF_X1 port map( A => n12738, Z => n10634);
   U2910 : BUF_X1 port map( A => n12737, Z => n10627);
   U2911 : BUF_X1 port map( A => n12768, Z => n10845);
   U2912 : BUF_X1 port map( A => n12767, Z => n10838);
   U2913 : BUF_X1 port map( A => n12766, Z => n10831);
   U2914 : BUF_X1 port map( A => n12765, Z => n10824);
   U2915 : BUF_X1 port map( A => n12764, Z => n10817);
   U2916 : BUF_X1 port map( A => n12763, Z => n10810);
   U2917 : BUF_X1 port map( A => n12762, Z => n10803);
   U2918 : BUF_X1 port map( A => n12761, Z => n10796);
   U2919 : BUF_X1 port map( A => n12760, Z => n10789);
   U2920 : BUF_X1 port map( A => n12759, Z => n10782);
   U2921 : BUF_X1 port map( A => n12758, Z => n10775);
   U2922 : BUF_X1 port map( A => n12757, Z => n10768);
   U2923 : BUF_X1 port map( A => n12756, Z => n10761);
   U2924 : BUF_X1 port map( A => n12755, Z => n10754);
   U2925 : BUF_X1 port map( A => n12754, Z => n10747);
   U2926 : BUF_X1 port map( A => n12753, Z => n10740);
   U2927 : BUF_X1 port map( A => n12752, Z => n10733);
   U2928 : BUF_X1 port map( A => n12751, Z => n10726);
   U2929 : BUF_X1 port map( A => n12750, Z => n10719);
   U2930 : BUF_X1 port map( A => n12749, Z => n10712);
   U2931 : BUF_X1 port map( A => n12748, Z => n10705);
   U2932 : BUF_X1 port map( A => n12747, Z => n10698);
   U2933 : BUF_X1 port map( A => n12746, Z => n10691);
   U2934 : BUF_X1 port map( A => n12745, Z => n10684);
   U2935 : BUF_X1 port map( A => n12744, Z => n10677);
   U2936 : BUF_X1 port map( A => n12743, Z => n10670);
   U2937 : BUF_X1 port map( A => n12742, Z => n10663);
   U2938 : BUF_X1 port map( A => n12741, Z => n10656);
   U2939 : BUF_X1 port map( A => n12740, Z => n10649);
   U2940 : BUF_X1 port map( A => n12739, Z => n10642);
   U2941 : BUF_X1 port map( A => n12738, Z => n10635);
   U2942 : BUF_X1 port map( A => n12737, Z => n10628);
   U2943 : BUF_X1 port map( A => n12768, Z => n10846);
   U2944 : BUF_X1 port map( A => n12767, Z => n10839);
   U2945 : BUF_X1 port map( A => n12766, Z => n10832);
   U2946 : BUF_X1 port map( A => n12765, Z => n10825);
   U2947 : BUF_X1 port map( A => n12764, Z => n10818);
   U2948 : BUF_X1 port map( A => n12763, Z => n10811);
   U2949 : BUF_X1 port map( A => n12762, Z => n10804);
   U2950 : BUF_X1 port map( A => n12761, Z => n10797);
   U2951 : BUF_X1 port map( A => n12760, Z => n10790);
   U2952 : BUF_X1 port map( A => n12759, Z => n10783);
   U2953 : BUF_X1 port map( A => n12758, Z => n10776);
   U2954 : BUF_X1 port map( A => n12757, Z => n10769);
   U2955 : BUF_X1 port map( A => n12756, Z => n10762);
   U2956 : BUF_X1 port map( A => n12755, Z => n10755);
   U2957 : BUF_X1 port map( A => n12754, Z => n10748);
   U2958 : BUF_X1 port map( A => n12753, Z => n10741);
   U2959 : BUF_X1 port map( A => n12752, Z => n10734);
   U2960 : BUF_X1 port map( A => n12751, Z => n10727);
   U2961 : BUF_X1 port map( A => n12750, Z => n10720);
   U2962 : BUF_X1 port map( A => n12749, Z => n10713);
   U2963 : BUF_X1 port map( A => n12748, Z => n10706);
   U2964 : BUF_X1 port map( A => n12747, Z => n10699);
   U2965 : BUF_X1 port map( A => n12746, Z => n10692);
   U2966 : BUF_X1 port map( A => n12745, Z => n10685);
   U2967 : BUF_X1 port map( A => n12744, Z => n10678);
   U2968 : BUF_X1 port map( A => n12743, Z => n10671);
   U2969 : BUF_X1 port map( A => n12742, Z => n10664);
   U2970 : BUF_X1 port map( A => n12741, Z => n10657);
   U2971 : BUF_X1 port map( A => n12740, Z => n10650);
   U2972 : BUF_X1 port map( A => n12739, Z => n10643);
   U2973 : BUF_X1 port map( A => n12738, Z => n10636);
   U2974 : BUF_X1 port map( A => n12737, Z => n10629);
   U2975 : BUF_X1 port map( A => n12768, Z => n10847);
   U2976 : BUF_X1 port map( A => n12767, Z => n10840);
   U2977 : BUF_X1 port map( A => n12766, Z => n10833);
   U2978 : BUF_X1 port map( A => n12765, Z => n10826);
   U2979 : BUF_X1 port map( A => n12764, Z => n10819);
   U2980 : BUF_X1 port map( A => n12763, Z => n10812);
   U2981 : BUF_X1 port map( A => n12762, Z => n10805);
   U2982 : BUF_X1 port map( A => n12761, Z => n10798);
   U2983 : BUF_X1 port map( A => n12760, Z => n10791);
   U2984 : BUF_X1 port map( A => n12759, Z => n10784);
   U2985 : BUF_X1 port map( A => n12758, Z => n10777);
   U2986 : BUF_X1 port map( A => n12757, Z => n10770);
   U2987 : BUF_X1 port map( A => n12756, Z => n10763);
   U2988 : BUF_X1 port map( A => n12755, Z => n10756);
   U2989 : BUF_X1 port map( A => n12754, Z => n10749);
   U2990 : BUF_X1 port map( A => n12753, Z => n10742);
   U2991 : BUF_X1 port map( A => n12752, Z => n10735);
   U2992 : BUF_X1 port map( A => n12751, Z => n10728);
   U2993 : BUF_X1 port map( A => n12750, Z => n10721);
   U2994 : BUF_X1 port map( A => n12749, Z => n10714);
   U2995 : BUF_X1 port map( A => n12748, Z => n10707);
   U2996 : BUF_X1 port map( A => n12747, Z => n10700);
   U2997 : BUF_X1 port map( A => n12746, Z => n10693);
   U2998 : BUF_X1 port map( A => n12745, Z => n10686);
   U2999 : BUF_X1 port map( A => n12744, Z => n10679);
   U3000 : BUF_X1 port map( A => n12743, Z => n10672);
   U3001 : BUF_X1 port map( A => n12742, Z => n10665);
   U3002 : BUF_X1 port map( A => n12741, Z => n10658);
   U3003 : BUF_X1 port map( A => n12740, Z => n10651);
   U3004 : BUF_X1 port map( A => n12739, Z => n10644);
   U3005 : BUF_X1 port map( A => n12738, Z => n10637);
   U3006 : BUF_X1 port map( A => n12737, Z => n10630);
   U3007 : BUF_X1 port map( A => n12768, Z => n10848);
   U3008 : BUF_X1 port map( A => n12767, Z => n10841);
   U3009 : BUF_X1 port map( A => n12766, Z => n10834);
   U3010 : BUF_X1 port map( A => n12765, Z => n10827);
   U3011 : BUF_X1 port map( A => n12764, Z => n10820);
   U3012 : BUF_X1 port map( A => n12763, Z => n10813);
   U3013 : BUF_X1 port map( A => n12762, Z => n10806);
   U3014 : BUF_X1 port map( A => n12761, Z => n10799);
   U3015 : BUF_X1 port map( A => n12760, Z => n10792);
   U3016 : BUF_X1 port map( A => n12759, Z => n10785);
   U3017 : BUF_X1 port map( A => n12758, Z => n10778);
   U3018 : BUF_X1 port map( A => n12757, Z => n10771);
   U3019 : BUF_X1 port map( A => n12756, Z => n10764);
   U3020 : BUF_X1 port map( A => n12755, Z => n10757);
   U3021 : BUF_X1 port map( A => n12754, Z => n10750);
   U3022 : BUF_X1 port map( A => n12753, Z => n10743);
   U3023 : BUF_X1 port map( A => n12752, Z => n10736);
   U3024 : BUF_X1 port map( A => n12751, Z => n10729);
   U3025 : BUF_X1 port map( A => n12750, Z => n10722);
   U3026 : BUF_X1 port map( A => n12749, Z => n10715);
   U3027 : BUF_X1 port map( A => n12748, Z => n10708);
   U3028 : BUF_X1 port map( A => n12747, Z => n10701);
   U3029 : BUF_X1 port map( A => n12746, Z => n10694);
   U3030 : BUF_X1 port map( A => n12745, Z => n10687);
   U3031 : BUF_X1 port map( A => n12744, Z => n10680);
   U3032 : BUF_X1 port map( A => n12743, Z => n10673);
   U3033 : BUF_X1 port map( A => n12742, Z => n10666);
   U3034 : BUF_X1 port map( A => n12741, Z => n10659);
   U3035 : BUF_X1 port map( A => n12740, Z => n10652);
   U3036 : BUF_X1 port map( A => n12739, Z => n10645);
   U3037 : BUF_X1 port map( A => n12738, Z => n10638);
   U3038 : BUF_X1 port map( A => n12737, Z => n10631);
   U3039 : BUF_X1 port map( A => n12768, Z => n10849);
   U3040 : BUF_X1 port map( A => n12767, Z => n10842);
   U3041 : BUF_X1 port map( A => n12766, Z => n10835);
   U3042 : BUF_X1 port map( A => n12765, Z => n10828);
   U3043 : BUF_X1 port map( A => n12764, Z => n10821);
   U3044 : BUF_X1 port map( A => n12763, Z => n10814);
   U3045 : BUF_X1 port map( A => n12762, Z => n10807);
   U3046 : BUF_X1 port map( A => n12761, Z => n10800);
   U3047 : BUF_X1 port map( A => n12760, Z => n10793);
   U3048 : BUF_X1 port map( A => n12759, Z => n10786);
   U3049 : BUF_X1 port map( A => n12758, Z => n10779);
   U3050 : BUF_X1 port map( A => n12757, Z => n10772);
   U3051 : BUF_X1 port map( A => n12756, Z => n10765);
   U3052 : BUF_X1 port map( A => n12755, Z => n10758);
   U3053 : BUF_X1 port map( A => n12754, Z => n10751);
   U3054 : BUF_X1 port map( A => n12753, Z => n10744);
   U3055 : BUF_X1 port map( A => n12752, Z => n10737);
   U3056 : BUF_X1 port map( A => n12751, Z => n10730);
   U3057 : BUF_X1 port map( A => n12750, Z => n10723);
   U3058 : BUF_X1 port map( A => n12749, Z => n10716);
   U3059 : BUF_X1 port map( A => n12748, Z => n10709);
   U3060 : BUF_X1 port map( A => n12747, Z => n10702);
   U3061 : BUF_X1 port map( A => n12746, Z => n10695);
   U3062 : BUF_X1 port map( A => n12745, Z => n10688);
   U3063 : BUF_X1 port map( A => n12744, Z => n10681);
   U3064 : BUF_X1 port map( A => n12743, Z => n10674);
   U3065 : BUF_X1 port map( A => n12742, Z => n10667);
   U3066 : BUF_X1 port map( A => n12741, Z => n10660);
   U3067 : BUF_X1 port map( A => n12740, Z => n10653);
   U3068 : BUF_X1 port map( A => n12739, Z => n10646);
   U3069 : BUF_X1 port map( A => n12738, Z => n10639);
   U3070 : BUF_X1 port map( A => n12737, Z => n10632);
   U3071 : AND2_X1 port map( A1 => N2171, A2 => n2571, ZN => n2492);
   U3072 : NOR3_X1 port map( A1 => n2597, A2 => N2172, A3 => n12731, ZN => 
                           n2571);
   U3073 : INV_X1 port map( A => N2173, ZN => n12731);
   U3074 : NOR2_X1 port map( A1 => n14514, A2 => N8434, ZN => n5653);
   U3075 : NOR2_X1 port map( A1 => n14516, A2 => N8578, ZN => n4220);
   U3076 : BUF_X1 port map( A => n12768, Z => n10850);
   U3077 : BUF_X1 port map( A => n12767, Z => n10843);
   U3078 : BUF_X1 port map( A => n12766, Z => n10836);
   U3079 : BUF_X1 port map( A => n12765, Z => n10829);
   U3080 : BUF_X1 port map( A => n12764, Z => n10822);
   U3081 : BUF_X1 port map( A => n12763, Z => n10815);
   U3082 : BUF_X1 port map( A => n12762, Z => n10808);
   U3083 : BUF_X1 port map( A => n12761, Z => n10801);
   U3084 : BUF_X1 port map( A => n12760, Z => n10794);
   U3085 : BUF_X1 port map( A => n12759, Z => n10787);
   U3086 : BUF_X1 port map( A => n12758, Z => n10780);
   U3087 : BUF_X1 port map( A => n12757, Z => n10773);
   U3088 : BUF_X1 port map( A => n12756, Z => n10766);
   U3089 : BUF_X1 port map( A => n12755, Z => n10759);
   U3090 : BUF_X1 port map( A => n12754, Z => n10752);
   U3091 : BUF_X1 port map( A => n12753, Z => n10745);
   U3092 : BUF_X1 port map( A => n12752, Z => n10738);
   U3093 : BUF_X1 port map( A => n12751, Z => n10731);
   U3094 : BUF_X1 port map( A => n12750, Z => n10724);
   U3095 : BUF_X1 port map( A => n12749, Z => n10717);
   U3096 : BUF_X1 port map( A => n12748, Z => n10710);
   U3097 : BUF_X1 port map( A => n12747, Z => n10703);
   U3098 : BUF_X1 port map( A => n12746, Z => n10696);
   U3099 : BUF_X1 port map( A => n12745, Z => n10689);
   U3100 : BUF_X1 port map( A => n12744, Z => n10682);
   U3101 : BUF_X1 port map( A => n12743, Z => n10675);
   U3102 : BUF_X1 port map( A => n12742, Z => n10668);
   U3103 : BUF_X1 port map( A => n12741, Z => n10661);
   U3104 : BUF_X1 port map( A => n12740, Z => n10654);
   U3105 : BUF_X1 port map( A => n12739, Z => n10647);
   U3106 : BUF_X1 port map( A => n12738, Z => n10640);
   U3107 : BUF_X1 port map( A => n12737, Z => n10633);
   U3108 : AND2_X1 port map( A1 => n2719, A2 => n2730, ZN => n2494);
   U3109 : AND2_X1 port map( A1 => n2721, A2 => n2730, ZN => n2496);
   U3110 : AND2_X1 port map( A1 => n2723, A2 => n2730, ZN => n2498);
   U3111 : AND2_X1 port map( A1 => n2735, A2 => n2717, ZN => n2500);
   U3112 : AND2_X1 port map( A1 => n2735, A2 => n2719, ZN => n2566);
   U3113 : AND2_X1 port map( A1 => n2735, A2 => n2721, ZN => n2568);
   U3114 : AND2_X1 port map( A1 => n2735, A2 => n2723, ZN => n2570);
   U3115 : NAND2_X1 port map( A1 => N8437, A2 => n5659, ZN => n4389);
   U3116 : NAND2_X1 port map( A1 => N8581, A2 => n4226, ZN => n2956);
   U3117 : INV_X1 port map( A => N8437, ZN => n12769);
   U3118 : INV_X1 port map( A => N8581, ZN => n12773);
   U3119 : NOR2_X1 port map( A1 => n12734, A2 => N2170, ZN => n2730);
   U3120 : NOR2_X1 port map( A1 => n12735, A2 => n12736, ZN => n2717);
   U3121 : NOR2_X1 port map( A1 => n14514, A2 => n12772, ZN => n5702);
   U3122 : NOR2_X1 port map( A1 => n14516, A2 => n12776, ZN => n4269);
   U3123 : AND2_X1 port map( A1 => n5647, A2 => n5703, ZN => n5655);
   U3124 : AND2_X1 port map( A1 => n5647, A2 => n5702, ZN => n5657);
   U3125 : AND2_X1 port map( A1 => n4214, A2 => n4270, ZN => n4222);
   U3126 : AND2_X1 port map( A1 => n4214, A2 => n4269, ZN => n4224);
   U3127 : AND2_X1 port map( A1 => n5649, A2 => n5703, ZN => n5656);
   U3128 : AND2_X1 port map( A1 => n4216, A2 => n4270, ZN => n4223);
   U3129 : INV_X1 port map( A => N8435, ZN => n12771);
   U3130 : INV_X1 port map( A => N8579, ZN => n12775);
   U3131 : AND2_X1 port map( A1 => n2716, A2 => n2717, ZN => n2573);
   U3132 : AND2_X1 port map( A1 => n2716, A2 => n2719, ZN => n2576);
   U3133 : AND2_X1 port map( A1 => n2716, A2 => n2721, ZN => n2578);
   U3134 : AND2_X1 port map( A1 => n2716, A2 => n2723, ZN => n2580);
   U3135 : AND2_X1 port map( A1 => n2725, A2 => n2719, ZN => n2584);
   U3136 : AND2_X1 port map( A1 => n2725, A2 => n2721, ZN => n2586);
   U3137 : AND2_X1 port map( A1 => n2725, A2 => n2723, ZN => n2588);
   U3138 : AND2_X1 port map( A1 => n5651, A2 => n5703, ZN => n5661);
   U3139 : AND2_X1 port map( A1 => n4218, A2 => n4270, ZN => n4228);
   U3140 : NAND2_X1 port map( A1 => n5655, A2 => N8437, ZN => n4385);
   U3141 : NAND2_X1 port map( A1 => n5657, A2 => N8437, ZN => n4386);
   U3142 : NAND2_X1 port map( A1 => n5656, A2 => N8437, ZN => n4390);
   U3143 : NAND2_X1 port map( A1 => n5663, A2 => N8437, ZN => n4388);
   U3144 : NAND2_X1 port map( A1 => n5661, A2 => N8437, ZN => n4396);
   U3145 : NAND2_X1 port map( A1 => n5665, A2 => N8437, ZN => n4395);
   U3146 : NAND2_X1 port map( A1 => n4222, A2 => N8581, ZN => n2952);
   U3147 : NAND2_X1 port map( A1 => n4224, A2 => N8581, ZN => n2953);
   U3148 : NAND2_X1 port map( A1 => n4223, A2 => N8581, ZN => n2957);
   U3149 : NAND2_X1 port map( A1 => n4230, A2 => N8581, ZN => n2955);
   U3150 : NAND2_X1 port map( A1 => n4228, A2 => N8581, ZN => n2963);
   U3151 : NAND2_X1 port map( A1 => n4232, A2 => N8581, ZN => n2962);
   U3152 : NAND4_X1 port map( A1 => n5638, A2 => n5639, A3 => n5640, A4 => 
                           n5641, ZN => n5637);
   U3153 : AOI221_X1 port map( B1 => n11079, B2 => n12819, C1 => n11076, C2 => 
                           n13011, A => n5658, ZN => n5640);
   U3154 : NOR4_X1 port map( A1 => n5642, A2 => n5643, A3 => n5644, A4 => n5645
                           , ZN => n5641);
   U3155 : AOI222_X1 port map( A1 => n11055, A2 => n12851, B1 => n11052, B2 => 
                           n12883, C1 => n11049, C2 => n12947, ZN => n5638);
   U3156 : NAND4_X1 port map( A1 => n4205, A2 => n4206, A3 => n4207, A4 => 
                           n4208, ZN => n4204);
   U3157 : AOI221_X1 port map( B1 => n11343, B2 => n12819, C1 => n11340, C2 => 
                           n13011, A => n4225, ZN => n4207);
   U3158 : NOR4_X1 port map( A1 => n4209, A2 => n4210, A3 => n4211, A4 => n4212
                           , ZN => n4208);
   U3159 : AOI222_X1 port map( A1 => n11319, A2 => n12851, B1 => n11316, B2 => 
                           n12883, C1 => n11313, C2 => n12947, ZN => n4205);
   U3160 : NAND4_X1 port map( A1 => n5597, A2 => n5598, A3 => n5599, A4 => 
                           n5600, ZN => n5596);
   U3161 : AOI221_X1 port map( B1 => n11079, B2 => n12818, C1 => n11076, C2 => 
                           n13010, A => n5605, ZN => n5599);
   U3162 : NOR4_X1 port map( A1 => n5601, A2 => n5602, A3 => n5603, A4 => n5604
                           , ZN => n5600);
   U3163 : AOI222_X1 port map( A1 => n11055, A2 => n12850, B1 => n11052, B2 => 
                           n12882, C1 => n11049, C2 => n12946, ZN => n5597);
   U3164 : NAND4_X1 port map( A1 => n4164, A2 => n4165, A3 => n4166, A4 => 
                           n4167, ZN => n4163);
   U3165 : AOI221_X1 port map( B1 => n11343, B2 => n12818, C1 => n11340, C2 => 
                           n13010, A => n4172, ZN => n4166);
   U3166 : NOR4_X1 port map( A1 => n4168, A2 => n4169, A3 => n4170, A4 => n4171
                           , ZN => n4167);
   U3167 : AOI222_X1 port map( A1 => n11319, A2 => n12850, B1 => n11316, B2 => 
                           n12882, C1 => n11313, C2 => n12946, ZN => n4164);
   U3168 : NAND4_X1 port map( A1 => n5556, A2 => n5557, A3 => n5558, A4 => 
                           n5559, ZN => n5555);
   U3169 : AOI221_X1 port map( B1 => n11079, B2 => n12817, C1 => n11076, C2 => 
                           n13009, A => n5564, ZN => n5558);
   U3170 : NOR4_X1 port map( A1 => n5560, A2 => n5561, A3 => n5562, A4 => n5563
                           , ZN => n5559);
   U3171 : AOI222_X1 port map( A1 => n11055, A2 => n12849, B1 => n11052, B2 => 
                           n12881, C1 => n11049, C2 => n12945, ZN => n5556);
   U3172 : NAND4_X1 port map( A1 => n4123, A2 => n4124, A3 => n4125, A4 => 
                           n4126, ZN => n4122);
   U3173 : AOI221_X1 port map( B1 => n11343, B2 => n12817, C1 => n11340, C2 => 
                           n13009, A => n4131, ZN => n4125);
   U3174 : NOR4_X1 port map( A1 => n4127, A2 => n4128, A3 => n4129, A4 => n4130
                           , ZN => n4126);
   U3175 : AOI222_X1 port map( A1 => n11319, A2 => n12849, B1 => n11316, B2 => 
                           n12881, C1 => n11313, C2 => n12945, ZN => n4123);
   U3176 : NAND4_X1 port map( A1 => n5515, A2 => n5516, A3 => n5517, A4 => 
                           n5518, ZN => n5514);
   U3177 : AOI221_X1 port map( B1 => n11079, B2 => n12816, C1 => n11076, C2 => 
                           n13008, A => n5523, ZN => n5517);
   U3178 : NOR4_X1 port map( A1 => n5519, A2 => n5520, A3 => n5521, A4 => n5522
                           , ZN => n5518);
   U3179 : AOI222_X1 port map( A1 => n11055, A2 => n12848, B1 => n11052, B2 => 
                           n12880, C1 => n11049, C2 => n12944, ZN => n5515);
   U3180 : NAND4_X1 port map( A1 => n4082, A2 => n4083, A3 => n4084, A4 => 
                           n4085, ZN => n4081);
   U3181 : AOI221_X1 port map( B1 => n11343, B2 => n12816, C1 => n11340, C2 => 
                           n13008, A => n4090, ZN => n4084);
   U3182 : NOR4_X1 port map( A1 => n4086, A2 => n4087, A3 => n4088, A4 => n4089
                           , ZN => n4085);
   U3183 : AOI222_X1 port map( A1 => n11319, A2 => n12848, B1 => n11316, B2 => 
                           n12880, C1 => n11313, C2 => n12944, ZN => n4082);
   U3184 : NAND4_X1 port map( A1 => n5474, A2 => n5475, A3 => n5476, A4 => 
                           n5477, ZN => n5473);
   U3185 : AOI221_X1 port map( B1 => n11079, B2 => n12815, C1 => n11076, C2 => 
                           n13007, A => n5482, ZN => n5476);
   U3186 : NOR4_X1 port map( A1 => n5478, A2 => n5479, A3 => n5480, A4 => n5481
                           , ZN => n5477);
   U3187 : AOI222_X1 port map( A1 => n11055, A2 => n12847, B1 => n11052, B2 => 
                           n12879, C1 => n11049, C2 => n12943, ZN => n5474);
   U3188 : NAND4_X1 port map( A1 => n4041, A2 => n4042, A3 => n4043, A4 => 
                           n4044, ZN => n4040);
   U3189 : AOI221_X1 port map( B1 => n11343, B2 => n12815, C1 => n11340, C2 => 
                           n13007, A => n4049, ZN => n4043);
   U3190 : NOR4_X1 port map( A1 => n4045, A2 => n4046, A3 => n4047, A4 => n4048
                           , ZN => n4044);
   U3191 : AOI222_X1 port map( A1 => n11319, A2 => n12847, B1 => n11316, B2 => 
                           n12879, C1 => n11313, C2 => n12943, ZN => n4041);
   U3192 : NAND4_X1 port map( A1 => n5433, A2 => n5434, A3 => n5435, A4 => 
                           n5436, ZN => n5432);
   U3193 : AOI221_X1 port map( B1 => n11079, B2 => n12814, C1 => n11076, C2 => 
                           n13006, A => n5441, ZN => n5435);
   U3194 : NOR4_X1 port map( A1 => n5437, A2 => n5438, A3 => n5439, A4 => n5440
                           , ZN => n5436);
   U3195 : AOI222_X1 port map( A1 => n11055, A2 => n12846, B1 => n11052, B2 => 
                           n12878, C1 => n11049, C2 => n12942, ZN => n5433);
   U3196 : NAND4_X1 port map( A1 => n4000, A2 => n4001, A3 => n4002, A4 => 
                           n4003, ZN => n3999);
   U3197 : AOI221_X1 port map( B1 => n11343, B2 => n12814, C1 => n11340, C2 => 
                           n13006, A => n4008, ZN => n4002);
   U3198 : NOR4_X1 port map( A1 => n4004, A2 => n4005, A3 => n4006, A4 => n4007
                           , ZN => n4003);
   U3199 : AOI222_X1 port map( A1 => n11319, A2 => n12846, B1 => n11316, B2 => 
                           n12878, C1 => n11313, C2 => n12942, ZN => n4000);
   U3200 : NAND4_X1 port map( A1 => n5392, A2 => n5393, A3 => n5394, A4 => 
                           n5395, ZN => n5391);
   U3201 : AOI221_X1 port map( B1 => n11079, B2 => n12813, C1 => n11076, C2 => 
                           n13005, A => n5400, ZN => n5394);
   U3202 : NOR4_X1 port map( A1 => n5396, A2 => n5397, A3 => n5398, A4 => n5399
                           , ZN => n5395);
   U3203 : AOI222_X1 port map( A1 => n11055, A2 => n12845, B1 => n11052, B2 => 
                           n12877, C1 => n11049, C2 => n12941, ZN => n5392);
   U3204 : NAND4_X1 port map( A1 => n3959, A2 => n3960, A3 => n3961, A4 => 
                           n3962, ZN => n3958);
   U3205 : AOI221_X1 port map( B1 => n11343, B2 => n12813, C1 => n11340, C2 => 
                           n13005, A => n3967, ZN => n3961);
   U3206 : NOR4_X1 port map( A1 => n3963, A2 => n3964, A3 => n3965, A4 => n3966
                           , ZN => n3962);
   U3207 : AOI222_X1 port map( A1 => n11319, A2 => n12845, B1 => n11316, B2 => 
                           n12877, C1 => n11313, C2 => n12941, ZN => n3959);
   U3208 : NAND4_X1 port map( A1 => n5351, A2 => n5352, A3 => n5353, A4 => 
                           n5354, ZN => n5350);
   U3209 : AOI221_X1 port map( B1 => n11079, B2 => n12812, C1 => n11076, C2 => 
                           n13004, A => n5359, ZN => n5353);
   U3210 : NOR4_X1 port map( A1 => n5355, A2 => n5356, A3 => n5357, A4 => n5358
                           , ZN => n5354);
   U3211 : AOI222_X1 port map( A1 => n11055, A2 => n12844, B1 => n11052, B2 => 
                           n12876, C1 => n11049, C2 => n12940, ZN => n5351);
   U3212 : NAND4_X1 port map( A1 => n3918, A2 => n3919, A3 => n3920, A4 => 
                           n3921, ZN => n3917);
   U3213 : AOI221_X1 port map( B1 => n11343, B2 => n12812, C1 => n11340, C2 => 
                           n13004, A => n3926, ZN => n3920);
   U3214 : NOR4_X1 port map( A1 => n3922, A2 => n3923, A3 => n3924, A4 => n3925
                           , ZN => n3921);
   U3215 : AOI222_X1 port map( A1 => n11319, A2 => n12844, B1 => n11316, B2 => 
                           n12876, C1 => n11313, C2 => n12940, ZN => n3918);
   U3216 : NAND4_X1 port map( A1 => n5310, A2 => n5311, A3 => n5312, A4 => 
                           n5313, ZN => n5309);
   U3217 : AOI221_X1 port map( B1 => n11079, B2 => n12811, C1 => n11076, C2 => 
                           n13003, A => n5318, ZN => n5312);
   U3218 : NOR4_X1 port map( A1 => n5314, A2 => n5315, A3 => n5316, A4 => n5317
                           , ZN => n5313);
   U3219 : AOI222_X1 port map( A1 => n11055, A2 => n12843, B1 => n11052, B2 => 
                           n12875, C1 => n11049, C2 => n12939, ZN => n5310);
   U3220 : NAND4_X1 port map( A1 => n3877, A2 => n3878, A3 => n3879, A4 => 
                           n3880, ZN => n3876);
   U3221 : AOI221_X1 port map( B1 => n11343, B2 => n12811, C1 => n11340, C2 => 
                           n13003, A => n3885, ZN => n3879);
   U3222 : NOR4_X1 port map( A1 => n3881, A2 => n3882, A3 => n3883, A4 => n3884
                           , ZN => n3880);
   U3223 : AOI222_X1 port map( A1 => n11319, A2 => n12843, B1 => n11316, B2 => 
                           n12875, C1 => n11313, C2 => n12939, ZN => n3877);
   U3224 : NAND4_X1 port map( A1 => n5269, A2 => n5270, A3 => n5271, A4 => 
                           n5272, ZN => n5268);
   U3225 : AOI221_X1 port map( B1 => n11079, B2 => n12810, C1 => n11076, C2 => 
                           n13002, A => n5277, ZN => n5271);
   U3226 : NOR4_X1 port map( A1 => n5273, A2 => n5274, A3 => n5275, A4 => n5276
                           , ZN => n5272);
   U3227 : AOI222_X1 port map( A1 => n11055, A2 => n12842, B1 => n11052, B2 => 
                           n12874, C1 => n11049, C2 => n12938, ZN => n5269);
   U3228 : NAND4_X1 port map( A1 => n3836, A2 => n3837, A3 => n3838, A4 => 
                           n3839, ZN => n3835);
   U3229 : AOI221_X1 port map( B1 => n11343, B2 => n12810, C1 => n11340, C2 => 
                           n13002, A => n3844, ZN => n3838);
   U3230 : NOR4_X1 port map( A1 => n3840, A2 => n3841, A3 => n3842, A4 => n3843
                           , ZN => n3839);
   U3231 : AOI222_X1 port map( A1 => n11319, A2 => n12842, B1 => n11316, B2 => 
                           n12874, C1 => n11313, C2 => n12938, ZN => n3836);
   U3232 : NAND4_X1 port map( A1 => n5228, A2 => n5229, A3 => n5230, A4 => 
                           n5231, ZN => n5227);
   U3233 : AOI221_X1 port map( B1 => n11079, B2 => n12809, C1 => n11076, C2 => 
                           n13001, A => n5236, ZN => n5230);
   U3234 : NOR4_X1 port map( A1 => n5232, A2 => n5233, A3 => n5234, A4 => n5235
                           , ZN => n5231);
   U3235 : AOI222_X1 port map( A1 => n11055, A2 => n12841, B1 => n11052, B2 => 
                           n12873, C1 => n11049, C2 => n12937, ZN => n5228);
   U3236 : NAND4_X1 port map( A1 => n3795, A2 => n3796, A3 => n3797, A4 => 
                           n3798, ZN => n3794);
   U3237 : AOI221_X1 port map( B1 => n11343, B2 => n12809, C1 => n11340, C2 => 
                           n13001, A => n3803, ZN => n3797);
   U3238 : NOR4_X1 port map( A1 => n3799, A2 => n3800, A3 => n3801, A4 => n3802
                           , ZN => n3798);
   U3239 : AOI222_X1 port map( A1 => n11319, A2 => n12841, B1 => n11316, B2 => 
                           n12873, C1 => n11313, C2 => n12937, ZN => n3795);
   U3240 : NAND4_X1 port map( A1 => n5187, A2 => n5188, A3 => n5189, A4 => 
                           n5190, ZN => n5186);
   U3241 : AOI221_X1 port map( B1 => n11079, B2 => n12808, C1 => n11076, C2 => 
                           n13000, A => n5195, ZN => n5189);
   U3242 : NOR4_X1 port map( A1 => n5191, A2 => n5192, A3 => n5193, A4 => n5194
                           , ZN => n5190);
   U3243 : AOI222_X1 port map( A1 => n11055, A2 => n12840, B1 => n11052, B2 => 
                           n12872, C1 => n11049, C2 => n12936, ZN => n5187);
   U3244 : NAND4_X1 port map( A1 => n3754, A2 => n3755, A3 => n3756, A4 => 
                           n3757, ZN => n3753);
   U3245 : AOI221_X1 port map( B1 => n11343, B2 => n12808, C1 => n11340, C2 => 
                           n13000, A => n3762, ZN => n3756);
   U3246 : NOR4_X1 port map( A1 => n3758, A2 => n3759, A3 => n3760, A4 => n3761
                           , ZN => n3757);
   U3247 : AOI222_X1 port map( A1 => n11319, A2 => n12840, B1 => n11316, B2 => 
                           n12872, C1 => n11313, C2 => n12936, ZN => n3754);
   U3248 : NAND4_X1 port map( A1 => n5146, A2 => n5147, A3 => n5148, A4 => 
                           n5149, ZN => n5145);
   U3249 : AOI221_X1 port map( B1 => n11080, B2 => n12807, C1 => n11077, C2 => 
                           n12999, A => n5154, ZN => n5148);
   U3250 : NOR4_X1 port map( A1 => n5150, A2 => n5151, A3 => n5152, A4 => n5153
                           , ZN => n5149);
   U3251 : AOI222_X1 port map( A1 => n11056, A2 => n12839, B1 => n11053, B2 => 
                           n12871, C1 => n11050, C2 => n12935, ZN => n5146);
   U3252 : NAND4_X1 port map( A1 => n3713, A2 => n3714, A3 => n3715, A4 => 
                           n3716, ZN => n3712);
   U3253 : AOI221_X1 port map( B1 => n11344, B2 => n12807, C1 => n11341, C2 => 
                           n12999, A => n3721, ZN => n3715);
   U3254 : NOR4_X1 port map( A1 => n3717, A2 => n3718, A3 => n3719, A4 => n3720
                           , ZN => n3716);
   U3255 : AOI222_X1 port map( A1 => n11320, A2 => n12839, B1 => n11317, B2 => 
                           n12871, C1 => n11314, C2 => n12935, ZN => n3713);
   U3256 : NAND4_X1 port map( A1 => n5105, A2 => n5106, A3 => n5107, A4 => 
                           n5108, ZN => n5104);
   U3257 : AOI221_X1 port map( B1 => n11080, B2 => n12806, C1 => n11077, C2 => 
                           n12998, A => n5113, ZN => n5107);
   U3258 : NOR4_X1 port map( A1 => n5109, A2 => n5110, A3 => n5111, A4 => n5112
                           , ZN => n5108);
   U3259 : AOI222_X1 port map( A1 => n11056, A2 => n12838, B1 => n11053, B2 => 
                           n12870, C1 => n11050, C2 => n12934, ZN => n5105);
   U3260 : NAND4_X1 port map( A1 => n3672, A2 => n3673, A3 => n3674, A4 => 
                           n3675, ZN => n3671);
   U3261 : AOI221_X1 port map( B1 => n11344, B2 => n12806, C1 => n11341, C2 => 
                           n12998, A => n3680, ZN => n3674);
   U3262 : NOR4_X1 port map( A1 => n3676, A2 => n3677, A3 => n3678, A4 => n3679
                           , ZN => n3675);
   U3263 : AOI222_X1 port map( A1 => n11320, A2 => n12838, B1 => n11317, B2 => 
                           n12870, C1 => n11314, C2 => n12934, ZN => n3672);
   U3264 : NAND4_X1 port map( A1 => n5064, A2 => n5065, A3 => n5066, A4 => 
                           n5067, ZN => n5063);
   U3265 : AOI221_X1 port map( B1 => n11080, B2 => n12805, C1 => n11077, C2 => 
                           n12997, A => n5072, ZN => n5066);
   U3266 : NOR4_X1 port map( A1 => n5068, A2 => n5069, A3 => n5070, A4 => n5071
                           , ZN => n5067);
   U3267 : AOI222_X1 port map( A1 => n11056, A2 => n12837, B1 => n11053, B2 => 
                           n12869, C1 => n11050, C2 => n12933, ZN => n5064);
   U3268 : NAND4_X1 port map( A1 => n3631, A2 => n3632, A3 => n3633, A4 => 
                           n3634, ZN => n3630);
   U3269 : AOI221_X1 port map( B1 => n11344, B2 => n12805, C1 => n11341, C2 => 
                           n12997, A => n3639, ZN => n3633);
   U3270 : NOR4_X1 port map( A1 => n3635, A2 => n3636, A3 => n3637, A4 => n3638
                           , ZN => n3634);
   U3271 : AOI222_X1 port map( A1 => n11320, A2 => n12837, B1 => n11317, B2 => 
                           n12869, C1 => n11314, C2 => n12933, ZN => n3631);
   U3272 : NAND4_X1 port map( A1 => n5023, A2 => n5024, A3 => n5025, A4 => 
                           n5026, ZN => n5022);
   U3273 : AOI221_X1 port map( B1 => n11080, B2 => n12804, C1 => n11077, C2 => 
                           n12996, A => n5031, ZN => n5025);
   U3274 : NOR4_X1 port map( A1 => n5027, A2 => n5028, A3 => n5029, A4 => n5030
                           , ZN => n5026);
   U3275 : AOI222_X1 port map( A1 => n11056, A2 => n12836, B1 => n11053, B2 => 
                           n12868, C1 => n11050, C2 => n12932, ZN => n5023);
   U3276 : NAND4_X1 port map( A1 => n3590, A2 => n3591, A3 => n3592, A4 => 
                           n3593, ZN => n3589);
   U3277 : AOI221_X1 port map( B1 => n11344, B2 => n12804, C1 => n11341, C2 => 
                           n12996, A => n3598, ZN => n3592);
   U3278 : NOR4_X1 port map( A1 => n3594, A2 => n3595, A3 => n3596, A4 => n3597
                           , ZN => n3593);
   U3279 : AOI222_X1 port map( A1 => n11320, A2 => n12836, B1 => n11317, B2 => 
                           n12868, C1 => n11314, C2 => n12932, ZN => n3590);
   U3280 : NAND4_X1 port map( A1 => n4982, A2 => n4983, A3 => n4984, A4 => 
                           n4985, ZN => n4981);
   U3281 : AOI221_X1 port map( B1 => n11080, B2 => n12803, C1 => n11077, C2 => 
                           n12995, A => n4990, ZN => n4984);
   U3282 : NOR4_X1 port map( A1 => n4986, A2 => n4987, A3 => n4988, A4 => n4989
                           , ZN => n4985);
   U3283 : AOI222_X1 port map( A1 => n11056, A2 => n12835, B1 => n11053, B2 => 
                           n12867, C1 => n11050, C2 => n12931, ZN => n4982);
   U3284 : NAND4_X1 port map( A1 => n3549, A2 => n3550, A3 => n3551, A4 => 
                           n3552, ZN => n3548);
   U3285 : AOI221_X1 port map( B1 => n11344, B2 => n12803, C1 => n11341, C2 => 
                           n12995, A => n3557, ZN => n3551);
   U3286 : NOR4_X1 port map( A1 => n3553, A2 => n3554, A3 => n3555, A4 => n3556
                           , ZN => n3552);
   U3287 : AOI222_X1 port map( A1 => n11320, A2 => n12835, B1 => n11317, B2 => 
                           n12867, C1 => n11314, C2 => n12931, ZN => n3549);
   U3288 : NAND4_X1 port map( A1 => n4941, A2 => n4942, A3 => n4943, A4 => 
                           n4944, ZN => n4940);
   U3289 : AOI221_X1 port map( B1 => n11080, B2 => n12802, C1 => n11077, C2 => 
                           n12994, A => n4949, ZN => n4943);
   U3290 : NOR4_X1 port map( A1 => n4945, A2 => n4946, A3 => n4947, A4 => n4948
                           , ZN => n4944);
   U3291 : AOI222_X1 port map( A1 => n11056, A2 => n12834, B1 => n11053, B2 => 
                           n12866, C1 => n11050, C2 => n12930, ZN => n4941);
   U3292 : NAND4_X1 port map( A1 => n3508, A2 => n3509, A3 => n3510, A4 => 
                           n3511, ZN => n3507);
   U3293 : AOI221_X1 port map( B1 => n11344, B2 => n12802, C1 => n11341, C2 => 
                           n12994, A => n3516, ZN => n3510);
   U3294 : NOR4_X1 port map( A1 => n3512, A2 => n3513, A3 => n3514, A4 => n3515
                           , ZN => n3511);
   U3295 : AOI222_X1 port map( A1 => n11320, A2 => n12834, B1 => n11317, B2 => 
                           n12866, C1 => n11314, C2 => n12930, ZN => n3508);
   U3296 : NAND4_X1 port map( A1 => n4900, A2 => n4901, A3 => n4902, A4 => 
                           n4903, ZN => n4899);
   U3297 : AOI221_X1 port map( B1 => n11080, B2 => n12801, C1 => n11077, C2 => 
                           n12993, A => n4908, ZN => n4902);
   U3298 : NOR4_X1 port map( A1 => n4904, A2 => n4905, A3 => n4906, A4 => n4907
                           , ZN => n4903);
   U3299 : AOI222_X1 port map( A1 => n11056, A2 => n12833, B1 => n11053, B2 => 
                           n12865, C1 => n11050, C2 => n12929, ZN => n4900);
   U3300 : NAND4_X1 port map( A1 => n3467, A2 => n3468, A3 => n3469, A4 => 
                           n3470, ZN => n3466);
   U3301 : AOI221_X1 port map( B1 => n11344, B2 => n12801, C1 => n11341, C2 => 
                           n12993, A => n3475, ZN => n3469);
   U3302 : NOR4_X1 port map( A1 => n3471, A2 => n3472, A3 => n3473, A4 => n3474
                           , ZN => n3470);
   U3303 : AOI222_X1 port map( A1 => n11320, A2 => n12833, B1 => n11317, B2 => 
                           n12865, C1 => n11314, C2 => n12929, ZN => n3467);
   U3304 : NAND4_X1 port map( A1 => n4859, A2 => n4860, A3 => n4861, A4 => 
                           n4862, ZN => n4858);
   U3305 : AOI221_X1 port map( B1 => n11080, B2 => n12800, C1 => n11077, C2 => 
                           n12992, A => n4867, ZN => n4861);
   U3306 : NOR4_X1 port map( A1 => n4863, A2 => n4864, A3 => n4865, A4 => n4866
                           , ZN => n4862);
   U3307 : AOI222_X1 port map( A1 => n11056, A2 => n12832, B1 => n11053, B2 => 
                           n12864, C1 => n11050, C2 => n12928, ZN => n4859);
   U3308 : NAND4_X1 port map( A1 => n3426, A2 => n3427, A3 => n3428, A4 => 
                           n3429, ZN => n3425);
   U3309 : AOI221_X1 port map( B1 => n11344, B2 => n12800, C1 => n11341, C2 => 
                           n12992, A => n3434, ZN => n3428);
   U3310 : NOR4_X1 port map( A1 => n3430, A2 => n3431, A3 => n3432, A4 => n3433
                           , ZN => n3429);
   U3311 : AOI222_X1 port map( A1 => n11320, A2 => n12832, B1 => n11317, B2 => 
                           n12864, C1 => n11314, C2 => n12928, ZN => n3426);
   U3312 : NAND4_X1 port map( A1 => n4818, A2 => n4819, A3 => n4820, A4 => 
                           n4821, ZN => n4817);
   U3313 : AOI221_X1 port map( B1 => n11080, B2 => n12799, C1 => n11077, C2 => 
                           n12991, A => n4826, ZN => n4820);
   U3314 : NOR4_X1 port map( A1 => n4822, A2 => n4823, A3 => n4824, A4 => n4825
                           , ZN => n4821);
   U3315 : AOI222_X1 port map( A1 => n11056, A2 => n12831, B1 => n11053, B2 => 
                           n12863, C1 => n11050, C2 => n12927, ZN => n4818);
   U3316 : NAND4_X1 port map( A1 => n3385, A2 => n3386, A3 => n3387, A4 => 
                           n3388, ZN => n3384);
   U3317 : AOI221_X1 port map( B1 => n11344, B2 => n12799, C1 => n11341, C2 => 
                           n12991, A => n3393, ZN => n3387);
   U3318 : NOR4_X1 port map( A1 => n3389, A2 => n3390, A3 => n3391, A4 => n3392
                           , ZN => n3388);
   U3319 : AOI222_X1 port map( A1 => n11320, A2 => n12831, B1 => n11317, B2 => 
                           n12863, C1 => n11314, C2 => n12927, ZN => n3385);
   U3320 : NAND4_X1 port map( A1 => n4777, A2 => n4778, A3 => n4779, A4 => 
                           n4780, ZN => n4776);
   U3321 : AOI221_X1 port map( B1 => n11080, B2 => n12798, C1 => n11077, C2 => 
                           n12990, A => n4785, ZN => n4779);
   U3322 : NOR4_X1 port map( A1 => n4781, A2 => n4782, A3 => n4783, A4 => n4784
                           , ZN => n4780);
   U3323 : AOI222_X1 port map( A1 => n11056, A2 => n12830, B1 => n11053, B2 => 
                           n12862, C1 => n11050, C2 => n12926, ZN => n4777);
   U3324 : NAND4_X1 port map( A1 => n3344, A2 => n3345, A3 => n3346, A4 => 
                           n3347, ZN => n3343);
   U3325 : AOI221_X1 port map( B1 => n11344, B2 => n12798, C1 => n11341, C2 => 
                           n12990, A => n3352, ZN => n3346);
   U3326 : NOR4_X1 port map( A1 => n3348, A2 => n3349, A3 => n3350, A4 => n3351
                           , ZN => n3347);
   U3327 : AOI222_X1 port map( A1 => n11320, A2 => n12830, B1 => n11317, B2 => 
                           n12862, C1 => n11314, C2 => n12926, ZN => n3344);
   U3328 : NAND4_X1 port map( A1 => n4736, A2 => n4737, A3 => n4738, A4 => 
                           n4739, ZN => n4735);
   U3329 : AOI221_X1 port map( B1 => n11080, B2 => n12797, C1 => n11077, C2 => 
                           n12989, A => n4744, ZN => n4738);
   U3330 : NOR4_X1 port map( A1 => n4740, A2 => n4741, A3 => n4742, A4 => n4743
                           , ZN => n4739);
   U3331 : AOI222_X1 port map( A1 => n11056, A2 => n12829, B1 => n11053, B2 => 
                           n12861, C1 => n11050, C2 => n12925, ZN => n4736);
   U3332 : NAND4_X1 port map( A1 => n3303, A2 => n3304, A3 => n3305, A4 => 
                           n3306, ZN => n3302);
   U3333 : AOI221_X1 port map( B1 => n11344, B2 => n12797, C1 => n11341, C2 => 
                           n12989, A => n3311, ZN => n3305);
   U3334 : NOR4_X1 port map( A1 => n3307, A2 => n3308, A3 => n3309, A4 => n3310
                           , ZN => n3306);
   U3335 : AOI222_X1 port map( A1 => n11320, A2 => n12829, B1 => n11317, B2 => 
                           n12861, C1 => n11314, C2 => n12925, ZN => n3303);
   U3336 : NAND4_X1 port map( A1 => n4695, A2 => n4696, A3 => n4697, A4 => 
                           n4698, ZN => n4694);
   U3337 : AOI221_X1 port map( B1 => n11080, B2 => n12796, C1 => n11077, C2 => 
                           n12988, A => n4703, ZN => n4697);
   U3338 : NOR4_X1 port map( A1 => n4699, A2 => n4700, A3 => n4701, A4 => n4702
                           , ZN => n4698);
   U3339 : AOI222_X1 port map( A1 => n11056, A2 => n12828, B1 => n11053, B2 => 
                           n12860, C1 => n11050, C2 => n12924, ZN => n4695);
   U3340 : NAND4_X1 port map( A1 => n3262, A2 => n3263, A3 => n3264, A4 => 
                           n3265, ZN => n3261);
   U3341 : AOI221_X1 port map( B1 => n11344, B2 => n12796, C1 => n11341, C2 => 
                           n12988, A => n3270, ZN => n3264);
   U3342 : NOR4_X1 port map( A1 => n3266, A2 => n3267, A3 => n3268, A4 => n3269
                           , ZN => n3265);
   U3343 : AOI222_X1 port map( A1 => n11320, A2 => n12828, B1 => n11317, B2 => 
                           n12860, C1 => n11314, C2 => n12924, ZN => n3262);
   U3344 : NAND4_X1 port map( A1 => n4654, A2 => n4655, A3 => n4656, A4 => 
                           n4657, ZN => n4653);
   U3345 : AOI221_X1 port map( B1 => n11081, B2 => n12795, C1 => n11078, C2 => 
                           n12987, A => n4662, ZN => n4656);
   U3346 : NOR4_X1 port map( A1 => n4658, A2 => n4659, A3 => n4660, A4 => n4661
                           , ZN => n4657);
   U3347 : AOI222_X1 port map( A1 => n11057, A2 => n12827, B1 => n11054, B2 => 
                           n12859, C1 => n11051, C2 => n12923, ZN => n4654);
   U3348 : NAND4_X1 port map( A1 => n3221, A2 => n3222, A3 => n3223, A4 => 
                           n3224, ZN => n3220);
   U3349 : AOI221_X1 port map( B1 => n11345, B2 => n12795, C1 => n11342, C2 => 
                           n12987, A => n3229, ZN => n3223);
   U3350 : NOR4_X1 port map( A1 => n3225, A2 => n3226, A3 => n3227, A4 => n3228
                           , ZN => n3224);
   U3351 : AOI222_X1 port map( A1 => n11321, A2 => n12827, B1 => n11318, B2 => 
                           n12859, C1 => n11315, C2 => n12923, ZN => n3221);
   U3352 : NAND4_X1 port map( A1 => n4613, A2 => n4614, A3 => n4615, A4 => 
                           n4616, ZN => n4612);
   U3353 : AOI221_X1 port map( B1 => n11081, B2 => n12794, C1 => n11078, C2 => 
                           n12986, A => n4621, ZN => n4615);
   U3354 : NOR4_X1 port map( A1 => n4617, A2 => n4618, A3 => n4619, A4 => n4620
                           , ZN => n4616);
   U3355 : AOI222_X1 port map( A1 => n11057, A2 => n12826, B1 => n11054, B2 => 
                           n12858, C1 => n11051, C2 => n12922, ZN => n4613);
   U3356 : NAND4_X1 port map( A1 => n3180, A2 => n3181, A3 => n3182, A4 => 
                           n3183, ZN => n3179);
   U3357 : AOI221_X1 port map( B1 => n11345, B2 => n12794, C1 => n11342, C2 => 
                           n12986, A => n3188, ZN => n3182);
   U3358 : NOR4_X1 port map( A1 => n3184, A2 => n3185, A3 => n3186, A4 => n3187
                           , ZN => n3183);
   U3359 : AOI222_X1 port map( A1 => n11321, A2 => n12826, B1 => n11318, B2 => 
                           n12858, C1 => n11315, C2 => n12922, ZN => n3180);
   U3360 : NAND4_X1 port map( A1 => n4572, A2 => n4573, A3 => n4574, A4 => 
                           n4575, ZN => n4571);
   U3361 : AOI221_X1 port map( B1 => n11081, B2 => n12793, C1 => n11078, C2 => 
                           n12985, A => n4580, ZN => n4574);
   U3362 : NOR4_X1 port map( A1 => n4576, A2 => n4577, A3 => n4578, A4 => n4579
                           , ZN => n4575);
   U3363 : AOI222_X1 port map( A1 => n11057, A2 => n12825, B1 => n11054, B2 => 
                           n12857, C1 => n11051, C2 => n12921, ZN => n4572);
   U3364 : NAND4_X1 port map( A1 => n3139, A2 => n3140, A3 => n3141, A4 => 
                           n3142, ZN => n3138);
   U3365 : AOI221_X1 port map( B1 => n11345, B2 => n12793, C1 => n11342, C2 => 
                           n12985, A => n3147, ZN => n3141);
   U3366 : NOR4_X1 port map( A1 => n3143, A2 => n3144, A3 => n3145, A4 => n3146
                           , ZN => n3142);
   U3367 : AOI222_X1 port map( A1 => n11321, A2 => n12825, B1 => n11318, B2 => 
                           n12857, C1 => n11315, C2 => n12921, ZN => n3139);
   U3368 : NAND4_X1 port map( A1 => n4531, A2 => n4532, A3 => n4533, A4 => 
                           n4534, ZN => n4530);
   U3369 : AOI221_X1 port map( B1 => n11081, B2 => n12792, C1 => n11078, C2 => 
                           n12984, A => n4539, ZN => n4533);
   U3370 : NOR4_X1 port map( A1 => n4535, A2 => n4536, A3 => n4537, A4 => n4538
                           , ZN => n4534);
   U3371 : AOI222_X1 port map( A1 => n11057, A2 => n12824, B1 => n11054, B2 => 
                           n12856, C1 => n11051, C2 => n12920, ZN => n4531);
   U3372 : NAND4_X1 port map( A1 => n3098, A2 => n3099, A3 => n3100, A4 => 
                           n3101, ZN => n3097);
   U3373 : AOI221_X1 port map( B1 => n11345, B2 => n12792, C1 => n11342, C2 => 
                           n12984, A => n3106, ZN => n3100);
   U3374 : NOR4_X1 port map( A1 => n3102, A2 => n3103, A3 => n3104, A4 => n3105
                           , ZN => n3101);
   U3375 : AOI222_X1 port map( A1 => n11321, A2 => n12824, B1 => n11318, B2 => 
                           n12856, C1 => n11315, C2 => n12920, ZN => n3098);
   U3376 : NAND4_X1 port map( A1 => n4490, A2 => n4491, A3 => n4492, A4 => 
                           n4493, ZN => n4489);
   U3377 : AOI221_X1 port map( B1 => n11081, B2 => n12791, C1 => n11078, C2 => 
                           n12983, A => n4498, ZN => n4492);
   U3378 : NOR4_X1 port map( A1 => n4494, A2 => n4495, A3 => n4496, A4 => n4497
                           , ZN => n4493);
   U3379 : AOI222_X1 port map( A1 => n11057, A2 => n12823, B1 => n11054, B2 => 
                           n12855, C1 => n11051, C2 => n12919, ZN => n4490);
   U3380 : NAND4_X1 port map( A1 => n3057, A2 => n3058, A3 => n3059, A4 => 
                           n3060, ZN => n3056);
   U3381 : AOI221_X1 port map( B1 => n11345, B2 => n12791, C1 => n11342, C2 => 
                           n12983, A => n3065, ZN => n3059);
   U3382 : NOR4_X1 port map( A1 => n3061, A2 => n3062, A3 => n3063, A4 => n3064
                           , ZN => n3060);
   U3383 : AOI222_X1 port map( A1 => n11321, A2 => n12823, B1 => n11318, B2 => 
                           n12855, C1 => n11315, C2 => n12919, ZN => n3057);
   U3384 : NAND4_X1 port map( A1 => n4449, A2 => n4450, A3 => n4451, A4 => 
                           n4452, ZN => n4448);
   U3385 : AOI221_X1 port map( B1 => n11081, B2 => n12790, C1 => n11078, C2 => 
                           n12982, A => n4457, ZN => n4451);
   U3386 : NOR4_X1 port map( A1 => n4453, A2 => n4454, A3 => n4455, A4 => n4456
                           , ZN => n4452);
   U3387 : AOI222_X1 port map( A1 => n11057, A2 => n12822, B1 => n11054, B2 => 
                           n12854, C1 => n11051, C2 => n12918, ZN => n4449);
   U3388 : NAND4_X1 port map( A1 => n3016, A2 => n3017, A3 => n3018, A4 => 
                           n3019, ZN => n3015);
   U3389 : AOI221_X1 port map( B1 => n11345, B2 => n12790, C1 => n11342, C2 => 
                           n12982, A => n3024, ZN => n3018);
   U3390 : NOR4_X1 port map( A1 => n3020, A2 => n3021, A3 => n3022, A4 => n3023
                           , ZN => n3019);
   U3391 : AOI222_X1 port map( A1 => n11321, A2 => n12822, B1 => n11318, B2 => 
                           n12854, C1 => n11315, C2 => n12918, ZN => n3016);
   U3392 : NAND4_X1 port map( A1 => n4408, A2 => n4409, A3 => n4410, A4 => 
                           n4411, ZN => n4407);
   U3393 : AOI221_X1 port map( B1 => n11081, B2 => n12789, C1 => n11078, C2 => 
                           n12981, A => n4416, ZN => n4410);
   U3394 : NOR4_X1 port map( A1 => n4412, A2 => n4413, A3 => n4414, A4 => n4415
                           , ZN => n4411);
   U3395 : AOI222_X1 port map( A1 => n11057, A2 => n12821, B1 => n11054, B2 => 
                           n12853, C1 => n11051, C2 => n12917, ZN => n4408);
   U3396 : NAND4_X1 port map( A1 => n2975, A2 => n2976, A3 => n2977, A4 => 
                           n2978, ZN => n2974);
   U3397 : AOI221_X1 port map( B1 => n11345, B2 => n12789, C1 => n11342, C2 => 
                           n12981, A => n2983, ZN => n2977);
   U3398 : NOR4_X1 port map( A1 => n2979, A2 => n2980, A3 => n2981, A4 => n2982
                           , ZN => n2978);
   U3399 : AOI222_X1 port map( A1 => n11321, A2 => n12821, B1 => n11318, B2 => 
                           n12853, C1 => n11315, C2 => n12917, ZN => n2975);
   U3400 : NAND4_X1 port map( A1 => n4279, A2 => n4280, A3 => n4281, A4 => 
                           n4282, ZN => n4278);
   U3401 : AOI221_X1 port map( B1 => n11081, B2 => n12788, C1 => n11078, C2 => 
                           n12980, A => n4300, ZN => n4281);
   U3402 : NOR4_X1 port map( A1 => n4283, A2 => n4284, A3 => n4285, A4 => n4286
                           , ZN => n4282);
   U3403 : AOI222_X1 port map( A1 => n11057, A2 => n12820, B1 => n11054, B2 => 
                           n12852, C1 => n11051, C2 => n12916, ZN => n4279);
   U3404 : NAND4_X1 port map( A1 => n2747, A2 => n2748, A3 => n2749, A4 => 
                           n2750, ZN => n2746);
   U3405 : AOI221_X1 port map( B1 => n11345, B2 => n12788, C1 => n11342, C2 => 
                           n12980, A => n2800, ZN => n2749);
   U3406 : NOR4_X1 port map( A1 => n2751, A2 => n2752, A3 => n2753, A4 => n2786
                           , ZN => n2750);
   U3407 : AOI222_X1 port map( A1 => n11321, A2 => n12820, B1 => n11318, B2 => 
                           n12852, C1 => n11315, C2 => n12916, ZN => n2747);
   U3408 : AND2_X1 port map( A1 => n5650, A2 => n5703, ZN => n5659);
   U3409 : AND2_X1 port map( A1 => n4217, A2 => n4270, ZN => n4226);
   U3410 : AND2_X1 port map( A1 => n5649, A2 => n5702, ZN => n5663);
   U3411 : AND2_X1 port map( A1 => n4216, A2 => n4269, ZN => n4230);
   U3412 : AND2_X1 port map( A1 => n5651, A2 => n5702, ZN => n5665);
   U3413 : AND2_X1 port map( A1 => n4218, A2 => n4269, ZN => n4232);
   U3414 : AND2_X1 port map( A1 => n5652, A2 => n5654, ZN => n5648);
   U3415 : AND2_X1 port map( A1 => n4219, A2 => n4221, ZN => n4215);
   U3416 : AND2_X1 port map( A1 => n5702, A2 => n5650, ZN => n5660);
   U3417 : AND2_X1 port map( A1 => n4269, A2 => n4217, ZN => n4227);
   U3418 : NAND2_X1 port map( A1 => n5705, A2 => n5647, ZN => n4394);
   U3419 : NAND2_X1 port map( A1 => n4272, A2 => n4214, ZN => n2961);
   U3420 : AND2_X1 port map( A1 => n5654, A2 => n5701, ZN => n5688);
   U3421 : AND2_X1 port map( A1 => n4221, A2 => n4268, ZN => n4255);
   U3422 : NOR2_X1 port map( A1 => n12769, A2 => N8435, ZN => n5701);
   U3423 : NOR2_X1 port map( A1 => n12773, A2 => N8579, ZN => n4268);
   U3424 : AND2_X1 port map( A1 => n5675, A2 => n5654, ZN => n5676);
   U3425 : AND2_X1 port map( A1 => n4242, A2 => n4221, ZN => n4243);
   U3426 : INV_X1 port map( A => N2171, ZN => n12733);
   U3427 : NAND2_X1 port map( A1 => n5648, A2 => n5647, ZN => n4287);
   U3428 : NAND2_X1 port map( A1 => n5646, A2 => n5647, ZN => n4288);
   U3429 : NAND2_X1 port map( A1 => n5674, A2 => n5647, ZN => n4319);
   U3430 : NAND2_X1 port map( A1 => n5690, A2 => n5647, ZN => n4357);
   U3431 : NAND2_X1 port map( A1 => n5688, A2 => n5647, ZN => n4349);
   U3432 : NAND2_X1 port map( A1 => n5692, A2 => n5647, ZN => n4364);
   U3433 : NAND2_X1 port map( A1 => n4215, A2 => n4214, ZN => n2787);
   U3434 : NAND2_X1 port map( A1 => n4213, A2 => n4214, ZN => n2788);
   U3435 : NAND2_X1 port map( A1 => n4241, A2 => n4214, ZN => n2851);
   U3436 : NAND2_X1 port map( A1 => n4257, A2 => n4214, ZN => n2921);
   U3437 : NAND2_X1 port map( A1 => n4255, A2 => n4214, ZN => n2881);
   U3438 : NAND2_X1 port map( A1 => n4259, A2 => n4214, ZN => n2928);
   U3439 : BUF_X1 port map( A => N8735, Z => n12427);
   U3440 : BUF_X1 port map( A => N8702, Z => n12430);
   U3441 : BUF_X1 port map( A => N8702, Z => n12429);
   U3442 : BUF_X1 port map( A => N8735, Z => n12426);
   U3443 : NAND2_X1 port map( A1 => n5648, A2 => n5649, ZN => n4291);
   U3444 : NAND2_X1 port map( A1 => n5646, A2 => n5649, ZN => n4289);
   U3445 : NAND2_X1 port map( A1 => n5676, A2 => n5649, ZN => n4322);
   U3446 : NAND2_X1 port map( A1 => n5674, A2 => n5649, ZN => n4321);
   U3447 : NAND2_X1 port map( A1 => n5688, A2 => n5649, ZN => n4380);
   U3448 : NAND2_X1 port map( A1 => n5690, A2 => n5649, ZN => n4381);
   U3449 : NAND2_X1 port map( A1 => n4215, A2 => n4216, ZN => n2791);
   U3450 : NAND2_X1 port map( A1 => n4213, A2 => n4216, ZN => n2789);
   U3451 : NAND2_X1 port map( A1 => n4243, A2 => n4216, ZN => n2854);
   U3452 : NAND2_X1 port map( A1 => n4241, A2 => n4216, ZN => n2853);
   U3453 : NAND2_X1 port map( A1 => n4255, A2 => n4216, ZN => n2947);
   U3454 : NAND2_X1 port map( A1 => n4257, A2 => n4216, ZN => n2948);
   U3455 : INV_X1 port map( A => N8434, ZN => n12772);
   U3456 : INV_X1 port map( A => N8578, ZN => n12776);
   U3457 : BUF_X1 port map( A => N8702, Z => n12431);
   U3458 : BUF_X1 port map( A => N8735, Z => n12428);
   U3459 : NAND2_X1 port map( A1 => n5648, A2 => n5651, ZN => n4292);
   U3460 : NAND2_X1 port map( A1 => n5646, A2 => n5651, ZN => n4293);
   U3461 : NAND2_X1 port map( A1 => n5676, A2 => n5651, ZN => n4324);
   U3462 : NAND2_X1 port map( A1 => n5674, A2 => n5651, ZN => n4327);
   U3463 : NAND2_X1 port map( A1 => n5687, A2 => n5651, ZN => n4350);
   U3464 : NAND2_X1 port map( A1 => n5688, A2 => n5651, ZN => n4383);
   U3465 : NAND2_X1 port map( A1 => n4215, A2 => n4218, ZN => n2792);
   U3466 : NAND2_X1 port map( A1 => n4213, A2 => n4218, ZN => n2793);
   U3467 : NAND2_X1 port map( A1 => n4243, A2 => n4218, ZN => n2856);
   U3468 : NAND2_X1 port map( A1 => n4241, A2 => n4218, ZN => n2859);
   U3469 : NAND2_X1 port map( A1 => n4254, A2 => n4218, ZN => n2914);
   U3470 : NAND2_X1 port map( A1 => n4255, A2 => n4218, ZN => n2950);
   U3471 : NAND2_X1 port map( A1 => n5648, A2 => n5650, ZN => n4290);
   U3472 : NAND2_X1 port map( A1 => n5646, A2 => n5650, ZN => n4294);
   U3473 : NAND2_X1 port map( A1 => n5676, A2 => n5650, ZN => n4320);
   U3474 : NAND2_X1 port map( A1 => n5674, A2 => n5650, ZN => n4325);
   U3475 : NAND2_X1 port map( A1 => n5688, A2 => n5650, ZN => n4384);
   U3476 : NAND2_X1 port map( A1 => n5690, A2 => n5650, ZN => n4382);
   U3477 : NAND2_X1 port map( A1 => n4215, A2 => n4217, ZN => n2790);
   U3478 : NAND2_X1 port map( A1 => n4213, A2 => n4217, ZN => n2794);
   U3479 : NAND2_X1 port map( A1 => n4243, A2 => n4217, ZN => n2852);
   U3480 : NAND2_X1 port map( A1 => n4241, A2 => n4217, ZN => n2857);
   U3481 : NAND2_X1 port map( A1 => n4255, A2 => n4217, ZN => n2951);
   U3482 : NAND2_X1 port map( A1 => n4257, A2 => n4217, ZN => n2949);
   U3483 : AND2_X1 port map( A1 => n5660, A2 => N8437, ZN => n4391);
   U3484 : AND2_X1 port map( A1 => n4227, A2 => N8581, ZN => n2958);
   U3485 : NAND2_X1 port map( A1 => n5651, A2 => n5690, ZN => n4387);
   U3486 : NAND2_X1 port map( A1 => n4218, A2 => n4257, ZN => n2954);
   U3487 : AND3_X1 port map( A1 => n5654, A2 => n12769, A3 => n5678, ZN => 
                           n5662);
   U3488 : AND3_X1 port map( A1 => n4221, A2 => n12773, A3 => n4245, ZN => 
                           n4229);
   U3489 : AND2_X1 port map( A1 => n5689, A2 => n5654, ZN => n5692);
   U3490 : AND2_X1 port map( A1 => n4256, A2 => n4221, ZN => n4259);
   U3491 : AND2_X1 port map( A1 => n5705, A2 => n5651, ZN => n4392);
   U3492 : AND2_X1 port map( A1 => n4272, A2 => n4218, ZN => n2959);
   U3493 : AND2_X1 port map( A1 => n5687, A2 => n5647, ZN => n4369);
   U3494 : AND2_X1 port map( A1 => n5706, A2 => n5647, ZN => n4400);
   U3495 : AND2_X1 port map( A1 => n4254, A2 => n4214, ZN => n2933);
   U3496 : AND2_X1 port map( A1 => n4273, A2 => n4214, ZN => n2967);
   U3497 : AND2_X1 port map( A1 => n5664, A2 => n5649, ZN => n4304);
   U3498 : AND2_X1 port map( A1 => n4231, A2 => n4216, ZN => n2804);
   U3499 : AND2_X1 port map( A1 => n5706, A2 => n5650, ZN => n4397);
   U3500 : AND2_X1 port map( A1 => n4273, A2 => n4217, ZN => n2964);
   U3501 : AND2_X1 port map( A1 => n5664, A2 => n5651, ZN => n4329);
   U3502 : AND2_X1 port map( A1 => n5662, A2 => n5651, ZN => n4330);
   U3503 : AND2_X1 port map( A1 => n4231, A2 => n4218, ZN => n2861);
   U3504 : AND2_X1 port map( A1 => n4229, A2 => n4218, ZN => n2862);
   U3505 : AND2_X1 port map( A1 => n5662, A2 => n5650, ZN => n4299);
   U3506 : AND2_X1 port map( A1 => n5692, A2 => n5650, ZN => n4366);
   U3507 : AND2_X1 port map( A1 => n4229, A2 => n4217, ZN => n2799);
   U3508 : AND2_X1 port map( A1 => n4259, A2 => n4217, ZN => n2930);
   U3509 : AND2_X1 port map( A1 => N2170, A2 => n12734, ZN => n2725);
   U3510 : BUF_X1 port map( A => RESET, Z => n12432);
   U3511 : INV_X1 port map( A => n2740, ZN => r480_A_3_port);
   U3512 : INV_X1 port map( A => n2739, ZN => r486_A_3_port);
   U3513 : INV_X1 port map( A => n2741, ZN => r472_B_3_port);
   U3514 : AND2_X1 port map( A1 => n5705, A2 => n5649, ZN => n4401);
   U3515 : AND2_X1 port map( A1 => n5705, A2 => n5650, ZN => n4402);
   U3516 : AND2_X1 port map( A1 => n4272, A2 => n4216, ZN => n2968);
   U3517 : AND2_X1 port map( A1 => n4272, A2 => n4217, ZN => n2969);
   U3518 : AND2_X1 port map( A1 => n5664, A2 => n5647, ZN => n4305);
   U3519 : AND2_X1 port map( A1 => n5662, A2 => n5647, ZN => n4308);
   U3520 : AND2_X1 port map( A1 => n5676, A2 => n5647, ZN => n4336);
   U3521 : AND2_X1 port map( A1 => n4231, A2 => n4214, ZN => n2805);
   U3522 : AND2_X1 port map( A1 => n4229, A2 => n4214, ZN => n2808);
   U3523 : AND2_X1 port map( A1 => n4243, A2 => n4214, ZN => n2868);
   U3524 : AND2_X1 port map( A1 => n5706, A2 => n5649, ZN => n4398);
   U3525 : AND2_X1 port map( A1 => n5706, A2 => n5651, ZN => n4399);
   U3526 : AND2_X1 port map( A1 => n4273, A2 => n4216, ZN => n2965);
   U3527 : AND2_X1 port map( A1 => n4273, A2 => n4218, ZN => n2966);
   U3528 : AND2_X1 port map( A1 => n5662, A2 => n5649, ZN => n4309);
   U3529 : AND2_X1 port map( A1 => n5687, A2 => n5649, ZN => n4370);
   U3530 : AND2_X1 port map( A1 => n5692, A2 => n5649, ZN => n4371);
   U3531 : AND2_X1 port map( A1 => n4229, A2 => n4216, ZN => n2809);
   U3532 : AND2_X1 port map( A1 => n4254, A2 => n4216, ZN => n2934);
   U3533 : AND2_X1 port map( A1 => n4259, A2 => n4216, ZN => n2938);
   U3534 : AND2_X1 port map( A1 => n5692, A2 => n5651, ZN => n4367);
   U3535 : AND2_X1 port map( A1 => n4259, A2 => n4218, ZN => n2931);
   U3536 : AND2_X1 port map( A1 => n5664, A2 => n5650, ZN => n4306);
   U3537 : AND2_X1 port map( A1 => n5687, A2 => n5650, ZN => n4368);
   U3538 : AND2_X1 port map( A1 => n4231, A2 => n4217, ZN => n2806);
   U3539 : AND2_X1 port map( A1 => n4254, A2 => n4217, ZN => n2932);
   U3540 : NOR2_X1 port map( A1 => n5633, A2 => n12663, ZN => N8703);
   U3541 : NOR4_X1 port map( A1 => n5634, A2 => n5635, A3 => n5636, A4 => n5637
                           , ZN => n5633);
   U3542 : NAND4_X1 port map( A1 => n5693, A2 => n5694, A3 => n5695, A4 => 
                           n5696, ZN => n5634);
   U3543 : NAND4_X1 port map( A1 => n5679, A2 => n5680, A3 => n5681, A4 => 
                           n5682, ZN => n5635);
   U3544 : NOR2_X1 port map( A1 => n4200, A2 => n12671, ZN => N8736);
   U3545 : NOR4_X1 port map( A1 => n4201, A2 => n4202, A3 => n4203, A4 => n4204
                           , ZN => n4200);
   U3546 : NAND4_X1 port map( A1 => n4260, A2 => n4261, A3 => n4262, A4 => 
                           n4263, ZN => n4201);
   U3547 : NAND4_X1 port map( A1 => n4246, A2 => n4247, A3 => n4248, A4 => 
                           n4249, ZN => n4202);
   U3548 : NOR2_X1 port map( A1 => n5592, A2 => n12663, ZN => N8704);
   U3549 : NOR4_X1 port map( A1 => n5593, A2 => n5594, A3 => n5595, A4 => n5596
                           , ZN => n5592);
   U3550 : NAND4_X1 port map( A1 => n5624, A2 => n5625, A3 => n5626, A4 => 
                           n5627, ZN => n5593);
   U3551 : NAND4_X1 port map( A1 => n5615, A2 => n5616, A3 => n5617, A4 => 
                           n5618, ZN => n5594);
   U3552 : NOR2_X1 port map( A1 => n4159, A2 => n12671, ZN => N8737);
   U3553 : NOR4_X1 port map( A1 => n4160, A2 => n4161, A3 => n4162, A4 => n4163
                           , ZN => n4159);
   U3554 : NAND4_X1 port map( A1 => n4191, A2 => n4192, A3 => n4193, A4 => 
                           n4194, ZN => n4160);
   U3555 : NAND4_X1 port map( A1 => n4182, A2 => n4183, A3 => n4184, A4 => 
                           n4185, ZN => n4161);
   U3556 : NOR2_X1 port map( A1 => n5551, A2 => n12663, ZN => N8705);
   U3557 : NOR4_X1 port map( A1 => n5552, A2 => n5553, A3 => n5554, A4 => n5555
                           , ZN => n5551);
   U3558 : NAND4_X1 port map( A1 => n5583, A2 => n5584, A3 => n5585, A4 => 
                           n5586, ZN => n5552);
   U3559 : NAND4_X1 port map( A1 => n5574, A2 => n5575, A3 => n5576, A4 => 
                           n5577, ZN => n5553);
   U3560 : NOR2_X1 port map( A1 => n4118, A2 => n12671, ZN => N8738);
   U3561 : NOR4_X1 port map( A1 => n4119, A2 => n4120, A3 => n4121, A4 => n4122
                           , ZN => n4118);
   U3562 : NAND4_X1 port map( A1 => n4150, A2 => n4151, A3 => n4152, A4 => 
                           n4153, ZN => n4119);
   U3563 : NAND4_X1 port map( A1 => n4141, A2 => n4142, A3 => n4143, A4 => 
                           n4144, ZN => n4120);
   U3564 : NOR2_X1 port map( A1 => n5510, A2 => n12663, ZN => N8706);
   U3565 : NOR4_X1 port map( A1 => n5511, A2 => n5512, A3 => n5513, A4 => n5514
                           , ZN => n5510);
   U3566 : NAND4_X1 port map( A1 => n5542, A2 => n5543, A3 => n5544, A4 => 
                           n5545, ZN => n5511);
   U3567 : NAND4_X1 port map( A1 => n5533, A2 => n5534, A3 => n5535, A4 => 
                           n5536, ZN => n5512);
   U3568 : NOR2_X1 port map( A1 => n4077, A2 => n12672, ZN => N8739);
   U3569 : NOR4_X1 port map( A1 => n4078, A2 => n4079, A3 => n4080, A4 => n4081
                           , ZN => n4077);
   U3570 : NAND4_X1 port map( A1 => n4109, A2 => n4110, A3 => n4111, A4 => 
                           n4112, ZN => n4078);
   U3571 : NAND4_X1 port map( A1 => n4100, A2 => n4101, A3 => n4102, A4 => 
                           n4103, ZN => n4079);
   U3572 : NOR2_X1 port map( A1 => n5469, A2 => n12664, ZN => N8707);
   U3573 : NOR4_X1 port map( A1 => n5470, A2 => n5471, A3 => n5472, A4 => n5473
                           , ZN => n5469);
   U3574 : NAND4_X1 port map( A1 => n5501, A2 => n5502, A3 => n5503, A4 => 
                           n5504, ZN => n5470);
   U3575 : NAND4_X1 port map( A1 => n5492, A2 => n5493, A3 => n5494, A4 => 
                           n5495, ZN => n5471);
   U3576 : NOR2_X1 port map( A1 => n4036, A2 => n12672, ZN => N8740);
   U3577 : NOR4_X1 port map( A1 => n4037, A2 => n4038, A3 => n4039, A4 => n4040
                           , ZN => n4036);
   U3578 : NAND4_X1 port map( A1 => n4068, A2 => n4069, A3 => n4070, A4 => 
                           n4071, ZN => n4037);
   U3579 : NAND4_X1 port map( A1 => n4059, A2 => n4060, A3 => n4061, A4 => 
                           n4062, ZN => n4038);
   U3580 : NOR2_X1 port map( A1 => n5428, A2 => n12664, ZN => N8708);
   U3581 : NOR4_X1 port map( A1 => n5429, A2 => n5430, A3 => n5431, A4 => n5432
                           , ZN => n5428);
   U3582 : NAND4_X1 port map( A1 => n5460, A2 => n5461, A3 => n5462, A4 => 
                           n5463, ZN => n5429);
   U3583 : NAND4_X1 port map( A1 => n5451, A2 => n5452, A3 => n5453, A4 => 
                           n5454, ZN => n5430);
   U3584 : NOR2_X1 port map( A1 => n3995, A2 => n12672, ZN => N8741);
   U3585 : NOR4_X1 port map( A1 => n3996, A2 => n3997, A3 => n3998, A4 => n3999
                           , ZN => n3995);
   U3586 : NAND4_X1 port map( A1 => n4027, A2 => n4028, A3 => n4029, A4 => 
                           n4030, ZN => n3996);
   U3587 : NAND4_X1 port map( A1 => n4018, A2 => n4019, A3 => n4020, A4 => 
                           n4021, ZN => n3997);
   U3588 : NOR2_X1 port map( A1 => n5387, A2 => n12664, ZN => N8709);
   U3589 : NOR4_X1 port map( A1 => n5388, A2 => n5389, A3 => n5390, A4 => n5391
                           , ZN => n5387);
   U3590 : NAND4_X1 port map( A1 => n5419, A2 => n5420, A3 => n5421, A4 => 
                           n5422, ZN => n5388);
   U3591 : NAND4_X1 port map( A1 => n5410, A2 => n5411, A3 => n5412, A4 => 
                           n5413, ZN => n5389);
   U3592 : NOR2_X1 port map( A1 => n3954, A2 => n12672, ZN => N8742);
   U3593 : NOR4_X1 port map( A1 => n3955, A2 => n3956, A3 => n3957, A4 => n3958
                           , ZN => n3954);
   U3594 : NAND4_X1 port map( A1 => n3986, A2 => n3987, A3 => n3988, A4 => 
                           n3989, ZN => n3955);
   U3595 : NAND4_X1 port map( A1 => n3977, A2 => n3978, A3 => n3979, A4 => 
                           n3980, ZN => n3956);
   U3596 : NOR2_X1 port map( A1 => n5346, A2 => n12664, ZN => N8710);
   U3597 : NOR4_X1 port map( A1 => n5347, A2 => n5348, A3 => n5349, A4 => n5350
                           , ZN => n5346);
   U3598 : NAND4_X1 port map( A1 => n5378, A2 => n5379, A3 => n5380, A4 => 
                           n5381, ZN => n5347);
   U3599 : NAND4_X1 port map( A1 => n5369, A2 => n5370, A3 => n5371, A4 => 
                           n5372, ZN => n5348);
   U3600 : NOR2_X1 port map( A1 => n3913, A2 => n12673, ZN => N8743);
   U3601 : NOR4_X1 port map( A1 => n3914, A2 => n3915, A3 => n3916, A4 => n3917
                           , ZN => n3913);
   U3602 : NAND4_X1 port map( A1 => n3945, A2 => n3946, A3 => n3947, A4 => 
                           n3948, ZN => n3914);
   U3603 : NAND4_X1 port map( A1 => n3936, A2 => n3937, A3 => n3938, A4 => 
                           n3939, ZN => n3915);
   U3604 : NOR2_X1 port map( A1 => n5305, A2 => n12665, ZN => N8711);
   U3605 : NOR4_X1 port map( A1 => n5306, A2 => n5307, A3 => n5308, A4 => n5309
                           , ZN => n5305);
   U3606 : NAND4_X1 port map( A1 => n5337, A2 => n5338, A3 => n5339, A4 => 
                           n5340, ZN => n5306);
   U3607 : NAND4_X1 port map( A1 => n5328, A2 => n5329, A3 => n5330, A4 => 
                           n5331, ZN => n5307);
   U3608 : NOR2_X1 port map( A1 => n3872, A2 => n12673, ZN => N8744);
   U3609 : NOR4_X1 port map( A1 => n3873, A2 => n3874, A3 => n3875, A4 => n3876
                           , ZN => n3872);
   U3610 : NAND4_X1 port map( A1 => n3904, A2 => n3905, A3 => n3906, A4 => 
                           n3907, ZN => n3873);
   U3611 : NAND4_X1 port map( A1 => n3895, A2 => n3896, A3 => n3897, A4 => 
                           n3898, ZN => n3874);
   U3612 : NOR2_X1 port map( A1 => n5264, A2 => n12665, ZN => N8712);
   U3613 : NOR4_X1 port map( A1 => n5265, A2 => n5266, A3 => n5267, A4 => n5268
                           , ZN => n5264);
   U3614 : NAND4_X1 port map( A1 => n5296, A2 => n5297, A3 => n5298, A4 => 
                           n5299, ZN => n5265);
   U3615 : NAND4_X1 port map( A1 => n5287, A2 => n5288, A3 => n5289, A4 => 
                           n5290, ZN => n5266);
   U3616 : NOR2_X1 port map( A1 => n3831, A2 => n12673, ZN => N8745);
   U3617 : NOR4_X1 port map( A1 => n3832, A2 => n3833, A3 => n3834, A4 => n3835
                           , ZN => n3831);
   U3618 : NAND4_X1 port map( A1 => n3863, A2 => n3864, A3 => n3865, A4 => 
                           n3866, ZN => n3832);
   U3619 : NAND4_X1 port map( A1 => n3854, A2 => n3855, A3 => n3856, A4 => 
                           n3857, ZN => n3833);
   U3620 : NOR2_X1 port map( A1 => n5223, A2 => n12665, ZN => N8713);
   U3621 : NOR4_X1 port map( A1 => n5224, A2 => n5225, A3 => n5226, A4 => n5227
                           , ZN => n5223);
   U3622 : NAND4_X1 port map( A1 => n5255, A2 => n5256, A3 => n5257, A4 => 
                           n5258, ZN => n5224);
   U3623 : NAND4_X1 port map( A1 => n5246, A2 => n5247, A3 => n5248, A4 => 
                           n5249, ZN => n5225);
   U3624 : NOR2_X1 port map( A1 => n3790, A2 => n12673, ZN => N8746);
   U3625 : NOR4_X1 port map( A1 => n3791, A2 => n3792, A3 => n3793, A4 => n3794
                           , ZN => n3790);
   U3626 : NAND4_X1 port map( A1 => n3822, A2 => n3823, A3 => n3824, A4 => 
                           n3825, ZN => n3791);
   U3627 : NAND4_X1 port map( A1 => n3813, A2 => n3814, A3 => n3815, A4 => 
                           n3816, ZN => n3792);
   U3628 : NOR2_X1 port map( A1 => n5182, A2 => n12665, ZN => N8714);
   U3629 : NOR4_X1 port map( A1 => n5183, A2 => n5184, A3 => n5185, A4 => n5186
                           , ZN => n5182);
   U3630 : NAND4_X1 port map( A1 => n5214, A2 => n5215, A3 => n5216, A4 => 
                           n5217, ZN => n5183);
   U3631 : NAND4_X1 port map( A1 => n5205, A2 => n5206, A3 => n5207, A4 => 
                           n5208, ZN => n5184);
   U3632 : NOR2_X1 port map( A1 => n3749, A2 => n12674, ZN => N8747);
   U3633 : NOR4_X1 port map( A1 => n3750, A2 => n3751, A3 => n3752, A4 => n3753
                           , ZN => n3749);
   U3634 : NAND4_X1 port map( A1 => n3781, A2 => n3782, A3 => n3783, A4 => 
                           n3784, ZN => n3750);
   U3635 : NAND4_X1 port map( A1 => n3772, A2 => n3773, A3 => n3774, A4 => 
                           n3775, ZN => n3751);
   U3636 : NOR2_X1 port map( A1 => n5141, A2 => n12666, ZN => N8715);
   U3637 : NOR4_X1 port map( A1 => n5142, A2 => n5143, A3 => n5144, A4 => n5145
                           , ZN => n5141);
   U3638 : NAND4_X1 port map( A1 => n5173, A2 => n5174, A3 => n5175, A4 => 
                           n5176, ZN => n5142);
   U3639 : NAND4_X1 port map( A1 => n5164, A2 => n5165, A3 => n5166, A4 => 
                           n5167, ZN => n5143);
   U3640 : NOR2_X1 port map( A1 => n3708, A2 => n12674, ZN => N8748);
   U3641 : NOR4_X1 port map( A1 => n3709, A2 => n3710, A3 => n3711, A4 => n3712
                           , ZN => n3708);
   U3642 : NAND4_X1 port map( A1 => n3740, A2 => n3741, A3 => n3742, A4 => 
                           n3743, ZN => n3709);
   U3643 : NAND4_X1 port map( A1 => n3731, A2 => n3732, A3 => n3733, A4 => 
                           n3734, ZN => n3710);
   U3644 : NOR2_X1 port map( A1 => n5100, A2 => n12666, ZN => N8716);
   U3645 : NOR4_X1 port map( A1 => n5101, A2 => n5102, A3 => n5103, A4 => n5104
                           , ZN => n5100);
   U3646 : NAND4_X1 port map( A1 => n5132, A2 => n5133, A3 => n5134, A4 => 
                           n5135, ZN => n5101);
   U3647 : NAND4_X1 port map( A1 => n5123, A2 => n5124, A3 => n5125, A4 => 
                           n5126, ZN => n5102);
   U3648 : NOR2_X1 port map( A1 => n3667, A2 => n12674, ZN => N8749);
   U3649 : NOR4_X1 port map( A1 => n3668, A2 => n3669, A3 => n3670, A4 => n3671
                           , ZN => n3667);
   U3650 : NAND4_X1 port map( A1 => n3699, A2 => n3700, A3 => n3701, A4 => 
                           n3702, ZN => n3668);
   U3651 : NAND4_X1 port map( A1 => n3690, A2 => n3691, A3 => n3692, A4 => 
                           n3693, ZN => n3669);
   U3652 : NOR2_X1 port map( A1 => n5059, A2 => n12666, ZN => N8717);
   U3653 : NOR4_X1 port map( A1 => n5060, A2 => n5061, A3 => n5062, A4 => n5063
                           , ZN => n5059);
   U3654 : NAND4_X1 port map( A1 => n5091, A2 => n5092, A3 => n5093, A4 => 
                           n5094, ZN => n5060);
   U3655 : NAND4_X1 port map( A1 => n5082, A2 => n5083, A3 => n5084, A4 => 
                           n5085, ZN => n5061);
   U3656 : NOR2_X1 port map( A1 => n3626, A2 => n12674, ZN => N8750);
   U3657 : NOR4_X1 port map( A1 => n3627, A2 => n3628, A3 => n3629, A4 => n3630
                           , ZN => n3626);
   U3658 : NAND4_X1 port map( A1 => n3658, A2 => n3659, A3 => n3660, A4 => 
                           n3661, ZN => n3627);
   U3659 : NAND4_X1 port map( A1 => n3649, A2 => n3650, A3 => n3651, A4 => 
                           n3652, ZN => n3628);
   U3660 : NOR2_X1 port map( A1 => n5018, A2 => n12666, ZN => N8718);
   U3661 : NOR4_X1 port map( A1 => n5019, A2 => n5020, A3 => n5021, A4 => n5022
                           , ZN => n5018);
   U3662 : NAND4_X1 port map( A1 => n5050, A2 => n5051, A3 => n5052, A4 => 
                           n5053, ZN => n5019);
   U3663 : NAND4_X1 port map( A1 => n5041, A2 => n5042, A3 => n5043, A4 => 
                           n5044, ZN => n5020);
   U3664 : NOR2_X1 port map( A1 => n3585, A2 => n12675, ZN => N8751);
   U3665 : NOR4_X1 port map( A1 => n3586, A2 => n3587, A3 => n3588, A4 => n3589
                           , ZN => n3585);
   U3666 : NAND4_X1 port map( A1 => n3617, A2 => n3618, A3 => n3619, A4 => 
                           n3620, ZN => n3586);
   U3667 : NAND4_X1 port map( A1 => n3608, A2 => n3609, A3 => n3610, A4 => 
                           n3611, ZN => n3587);
   U3668 : NOR2_X1 port map( A1 => n4977, A2 => n12667, ZN => N8719);
   U3669 : NOR4_X1 port map( A1 => n4978, A2 => n4979, A3 => n4980, A4 => n4981
                           , ZN => n4977);
   U3670 : NAND4_X1 port map( A1 => n5009, A2 => n5010, A3 => n5011, A4 => 
                           n5012, ZN => n4978);
   U3671 : NAND4_X1 port map( A1 => n5000, A2 => n5001, A3 => n5002, A4 => 
                           n5003, ZN => n4979);
   U3672 : NOR2_X1 port map( A1 => n3544, A2 => n12675, ZN => N8752);
   U3673 : NOR4_X1 port map( A1 => n3545, A2 => n3546, A3 => n3547, A4 => n3548
                           , ZN => n3544);
   U3674 : NAND4_X1 port map( A1 => n3576, A2 => n3577, A3 => n3578, A4 => 
                           n3579, ZN => n3545);
   U3675 : NAND4_X1 port map( A1 => n3567, A2 => n3568, A3 => n3569, A4 => 
                           n3570, ZN => n3546);
   U3676 : NOR2_X1 port map( A1 => n4936, A2 => n12667, ZN => N8720);
   U3677 : NOR4_X1 port map( A1 => n4937, A2 => n4938, A3 => n4939, A4 => n4940
                           , ZN => n4936);
   U3678 : NAND4_X1 port map( A1 => n4968, A2 => n4969, A3 => n4970, A4 => 
                           n4971, ZN => n4937);
   U3679 : NAND4_X1 port map( A1 => n4959, A2 => n4960, A3 => n4961, A4 => 
                           n4962, ZN => n4938);
   U3680 : NOR2_X1 port map( A1 => n3503, A2 => n12675, ZN => N8753);
   U3681 : NOR4_X1 port map( A1 => n3504, A2 => n3505, A3 => n3506, A4 => n3507
                           , ZN => n3503);
   U3682 : NAND4_X1 port map( A1 => n3535, A2 => n3536, A3 => n3537, A4 => 
                           n3538, ZN => n3504);
   U3683 : NAND4_X1 port map( A1 => n3526, A2 => n3527, A3 => n3528, A4 => 
                           n3529, ZN => n3505);
   U3684 : NOR2_X1 port map( A1 => n4895, A2 => n12667, ZN => N8721);
   U3685 : NOR4_X1 port map( A1 => n4896, A2 => n4897, A3 => n4898, A4 => n4899
                           , ZN => n4895);
   U3686 : NAND4_X1 port map( A1 => n4927, A2 => n4928, A3 => n4929, A4 => 
                           n4930, ZN => n4896);
   U3687 : NAND4_X1 port map( A1 => n4918, A2 => n4919, A3 => n4920, A4 => 
                           n4921, ZN => n4897);
   U3688 : NOR2_X1 port map( A1 => n3462, A2 => n12675, ZN => N8754);
   U3689 : NOR4_X1 port map( A1 => n3463, A2 => n3464, A3 => n3465, A4 => n3466
                           , ZN => n3462);
   U3690 : NAND4_X1 port map( A1 => n3494, A2 => n3495, A3 => n3496, A4 => 
                           n3497, ZN => n3463);
   U3691 : NAND4_X1 port map( A1 => n3485, A2 => n3486, A3 => n3487, A4 => 
                           n3488, ZN => n3464);
   U3692 : NOR2_X1 port map( A1 => n4854, A2 => n12667, ZN => N8722);
   U3693 : NOR4_X1 port map( A1 => n4855, A2 => n4856, A3 => n4857, A4 => n4858
                           , ZN => n4854);
   U3694 : NAND4_X1 port map( A1 => n4886, A2 => n4887, A3 => n4888, A4 => 
                           n4889, ZN => n4855);
   U3695 : NAND4_X1 port map( A1 => n4877, A2 => n4878, A3 => n4879, A4 => 
                           n4880, ZN => n4856);
   U3696 : NOR2_X1 port map( A1 => n3421, A2 => n12676, ZN => N8755);
   U3697 : NOR4_X1 port map( A1 => n3422, A2 => n3423, A3 => n3424, A4 => n3425
                           , ZN => n3421);
   U3698 : NAND4_X1 port map( A1 => n3453, A2 => n3454, A3 => n3455, A4 => 
                           n3456, ZN => n3422);
   U3699 : NAND4_X1 port map( A1 => n3444, A2 => n3445, A3 => n3446, A4 => 
                           n3447, ZN => n3423);
   U3700 : NOR2_X1 port map( A1 => n4813, A2 => n12668, ZN => N8723);
   U3701 : NOR4_X1 port map( A1 => n4814, A2 => n4815, A3 => n4816, A4 => n4817
                           , ZN => n4813);
   U3702 : NAND4_X1 port map( A1 => n4845, A2 => n4846, A3 => n4847, A4 => 
                           n4848, ZN => n4814);
   U3703 : NAND4_X1 port map( A1 => n4836, A2 => n4837, A3 => n4838, A4 => 
                           n4839, ZN => n4815);
   U3704 : NOR2_X1 port map( A1 => n3380, A2 => n12676, ZN => N8756);
   U3705 : NOR4_X1 port map( A1 => n3381, A2 => n3382, A3 => n3383, A4 => n3384
                           , ZN => n3380);
   U3706 : NAND4_X1 port map( A1 => n3412, A2 => n3413, A3 => n3414, A4 => 
                           n3415, ZN => n3381);
   U3707 : NAND4_X1 port map( A1 => n3403, A2 => n3404, A3 => n3405, A4 => 
                           n3406, ZN => n3382);
   U3708 : NOR2_X1 port map( A1 => n4772, A2 => n12668, ZN => N8724);
   U3709 : NOR4_X1 port map( A1 => n4773, A2 => n4774, A3 => n4775, A4 => n4776
                           , ZN => n4772);
   U3710 : NAND4_X1 port map( A1 => n4804, A2 => n4805, A3 => n4806, A4 => 
                           n4807, ZN => n4773);
   U3711 : NAND4_X1 port map( A1 => n4795, A2 => n4796, A3 => n4797, A4 => 
                           n4798, ZN => n4774);
   U3712 : NOR2_X1 port map( A1 => n3339, A2 => n12676, ZN => N8757);
   U3713 : NOR4_X1 port map( A1 => n3340, A2 => n3341, A3 => n3342, A4 => n3343
                           , ZN => n3339);
   U3714 : NAND4_X1 port map( A1 => n3371, A2 => n3372, A3 => n3373, A4 => 
                           n3374, ZN => n3340);
   U3715 : NAND4_X1 port map( A1 => n3362, A2 => n3363, A3 => n3364, A4 => 
                           n3365, ZN => n3341);
   U3716 : NOR2_X1 port map( A1 => n4731, A2 => n12668, ZN => N8725);
   U3717 : NOR4_X1 port map( A1 => n4732, A2 => n4733, A3 => n4734, A4 => n4735
                           , ZN => n4731);
   U3718 : NAND4_X1 port map( A1 => n4763, A2 => n4764, A3 => n4765, A4 => 
                           n4766, ZN => n4732);
   U3719 : NAND4_X1 port map( A1 => n4754, A2 => n4755, A3 => n4756, A4 => 
                           n4757, ZN => n4733);
   U3720 : NOR2_X1 port map( A1 => n3298, A2 => n12676, ZN => N8758);
   U3721 : NOR4_X1 port map( A1 => n3299, A2 => n3300, A3 => n3301, A4 => n3302
                           , ZN => n3298);
   U3722 : NAND4_X1 port map( A1 => n3330, A2 => n3331, A3 => n3332, A4 => 
                           n3333, ZN => n3299);
   U3723 : NAND4_X1 port map( A1 => n3321, A2 => n3322, A3 => n3323, A4 => 
                           n3324, ZN => n3300);
   U3724 : NOR2_X1 port map( A1 => n4690, A2 => n12668, ZN => N8726);
   U3725 : NOR4_X1 port map( A1 => n4691, A2 => n4692, A3 => n4693, A4 => n4694
                           , ZN => n4690);
   U3726 : NAND4_X1 port map( A1 => n4722, A2 => n4723, A3 => n4724, A4 => 
                           n4725, ZN => n4691);
   U3727 : NAND4_X1 port map( A1 => n4713, A2 => n4714, A3 => n4715, A4 => 
                           n4716, ZN => n4692);
   U3728 : NOR2_X1 port map( A1 => n3257, A2 => n12677, ZN => N8759);
   U3729 : NOR4_X1 port map( A1 => n3258, A2 => n3259, A3 => n3260, A4 => n3261
                           , ZN => n3257);
   U3730 : NAND4_X1 port map( A1 => n3289, A2 => n3290, A3 => n3291, A4 => 
                           n3292, ZN => n3258);
   U3731 : NAND4_X1 port map( A1 => n3280, A2 => n3281, A3 => n3282, A4 => 
                           n3283, ZN => n3259);
   U3732 : NOR2_X1 port map( A1 => n4649, A2 => n12669, ZN => N8727);
   U3733 : NOR4_X1 port map( A1 => n4650, A2 => n4651, A3 => n4652, A4 => n4653
                           , ZN => n4649);
   U3734 : NAND4_X1 port map( A1 => n4681, A2 => n4682, A3 => n4683, A4 => 
                           n4684, ZN => n4650);
   U3735 : NAND4_X1 port map( A1 => n4672, A2 => n4673, A3 => n4674, A4 => 
                           n4675, ZN => n4651);
   U3736 : NOR2_X1 port map( A1 => n3216, A2 => n12677, ZN => N8760);
   U3737 : NOR4_X1 port map( A1 => n3217, A2 => n3218, A3 => n3219, A4 => n3220
                           , ZN => n3216);
   U3738 : NAND4_X1 port map( A1 => n3248, A2 => n3249, A3 => n3250, A4 => 
                           n3251, ZN => n3217);
   U3739 : NAND4_X1 port map( A1 => n3239, A2 => n3240, A3 => n3241, A4 => 
                           n3242, ZN => n3218);
   U3740 : NOR2_X1 port map( A1 => n4608, A2 => n12669, ZN => N8728);
   U3741 : NOR4_X1 port map( A1 => n4609, A2 => n4610, A3 => n4611, A4 => n4612
                           , ZN => n4608);
   U3742 : NAND4_X1 port map( A1 => n4640, A2 => n4641, A3 => n4642, A4 => 
                           n4643, ZN => n4609);
   U3743 : NAND4_X1 port map( A1 => n4631, A2 => n4632, A3 => n4633, A4 => 
                           n4634, ZN => n4610);
   U3744 : NOR2_X1 port map( A1 => n3175, A2 => n12677, ZN => N8761);
   U3745 : NOR4_X1 port map( A1 => n3176, A2 => n3177, A3 => n3178, A4 => n3179
                           , ZN => n3175);
   U3746 : NAND4_X1 port map( A1 => n3207, A2 => n3208, A3 => n3209, A4 => 
                           n3210, ZN => n3176);
   U3747 : NAND4_X1 port map( A1 => n3198, A2 => n3199, A3 => n3200, A4 => 
                           n3201, ZN => n3177);
   U3748 : NOR2_X1 port map( A1 => n4567, A2 => n12669, ZN => N8729);
   U3749 : NOR4_X1 port map( A1 => n4568, A2 => n4569, A3 => n4570, A4 => n4571
                           , ZN => n4567);
   U3750 : NAND4_X1 port map( A1 => n4599, A2 => n4600, A3 => n4601, A4 => 
                           n4602, ZN => n4568);
   U3751 : NAND4_X1 port map( A1 => n4590, A2 => n4591, A3 => n4592, A4 => 
                           n4593, ZN => n4569);
   U3752 : NOR2_X1 port map( A1 => n3134, A2 => n12677, ZN => N8762);
   U3753 : NOR4_X1 port map( A1 => n3135, A2 => n3136, A3 => n3137, A4 => n3138
                           , ZN => n3134);
   U3754 : NAND4_X1 port map( A1 => n3166, A2 => n3167, A3 => n3168, A4 => 
                           n3169, ZN => n3135);
   U3755 : NAND4_X1 port map( A1 => n3157, A2 => n3158, A3 => n3159, A4 => 
                           n3160, ZN => n3136);
   U3756 : NOR2_X1 port map( A1 => n4526, A2 => n12669, ZN => N8730);
   U3757 : NOR4_X1 port map( A1 => n4527, A2 => n4528, A3 => n4529, A4 => n4530
                           , ZN => n4526);
   U3758 : NAND4_X1 port map( A1 => n4558, A2 => n4559, A3 => n4560, A4 => 
                           n4561, ZN => n4527);
   U3759 : NAND4_X1 port map( A1 => n4549, A2 => n4550, A3 => n4551, A4 => 
                           n4552, ZN => n4528);
   U3760 : NOR2_X1 port map( A1 => n3093, A2 => n12678, ZN => N8763);
   U3761 : NOR4_X1 port map( A1 => n3094, A2 => n3095, A3 => n3096, A4 => n3097
                           , ZN => n3093);
   U3762 : NAND4_X1 port map( A1 => n3125, A2 => n3126, A3 => n3127, A4 => 
                           n3128, ZN => n3094);
   U3763 : NAND4_X1 port map( A1 => n3116, A2 => n3117, A3 => n3118, A4 => 
                           n3119, ZN => n3095);
   U3764 : NOR2_X1 port map( A1 => n4485, A2 => n12670, ZN => N8731);
   U3765 : NOR4_X1 port map( A1 => n4486, A2 => n4487, A3 => n4488, A4 => n4489
                           , ZN => n4485);
   U3766 : NAND4_X1 port map( A1 => n4517, A2 => n4518, A3 => n4519, A4 => 
                           n4520, ZN => n4486);
   U3767 : NAND4_X1 port map( A1 => n4508, A2 => n4509, A3 => n4510, A4 => 
                           n4511, ZN => n4487);
   U3768 : NOR2_X1 port map( A1 => n3052, A2 => n12678, ZN => N8764);
   U3769 : NOR4_X1 port map( A1 => n3053, A2 => n3054, A3 => n3055, A4 => n3056
                           , ZN => n3052);
   U3770 : NAND4_X1 port map( A1 => n3084, A2 => n3085, A3 => n3086, A4 => 
                           n3087, ZN => n3053);
   U3771 : NAND4_X1 port map( A1 => n3075, A2 => n3076, A3 => n3077, A4 => 
                           n3078, ZN => n3054);
   U3772 : NOR2_X1 port map( A1 => n4444, A2 => n12670, ZN => N8732);
   U3773 : NOR4_X1 port map( A1 => n4445, A2 => n4446, A3 => n4447, A4 => n4448
                           , ZN => n4444);
   U3774 : NAND4_X1 port map( A1 => n4476, A2 => n4477, A3 => n4478, A4 => 
                           n4479, ZN => n4445);
   U3775 : NAND4_X1 port map( A1 => n4467, A2 => n4468, A3 => n4469, A4 => 
                           n4470, ZN => n4446);
   U3776 : NOR2_X1 port map( A1 => n3011, A2 => n12678, ZN => N8765);
   U3777 : NOR4_X1 port map( A1 => n3012, A2 => n3013, A3 => n3014, A4 => n3015
                           , ZN => n3011);
   U3778 : NAND4_X1 port map( A1 => n3043, A2 => n3044, A3 => n3045, A4 => 
                           n3046, ZN => n3012);
   U3779 : NAND4_X1 port map( A1 => n3034, A2 => n3035, A3 => n3036, A4 => 
                           n3037, ZN => n3013);
   U3780 : NOR2_X1 port map( A1 => n4403, A2 => n12670, ZN => N8733);
   U3781 : NOR4_X1 port map( A1 => n4404, A2 => n4405, A3 => n4406, A4 => n4407
                           , ZN => n4403);
   U3782 : NAND4_X1 port map( A1 => n4435, A2 => n4436, A3 => n4437, A4 => 
                           n4438, ZN => n4404);
   U3783 : NAND4_X1 port map( A1 => n4426, A2 => n4427, A3 => n4428, A4 => 
                           n4429, ZN => n4405);
   U3784 : NOR2_X1 port map( A1 => n2970, A2 => n12678, ZN => N8766);
   U3785 : NOR4_X1 port map( A1 => n2971, A2 => n2972, A3 => n2973, A4 => n2974
                           , ZN => n2970);
   U3786 : NAND4_X1 port map( A1 => n3002, A2 => n3003, A3 => n3004, A4 => 
                           n3005, ZN => n2971);
   U3787 : NAND4_X1 port map( A1 => n2993, A2 => n2994, A3 => n2995, A4 => 
                           n2996, ZN => n2972);
   U3788 : NOR2_X1 port map( A1 => n4274, A2 => n12670, ZN => N8734);
   U3789 : NOR4_X1 port map( A1 => n4275, A2 => n4276, A3 => n4277, A4 => n4278
                           , ZN => n4274);
   U3790 : NAND4_X1 port map( A1 => n4372, A2 => n4373, A3 => n4374, A4 => 
                           n4375, ZN => n4275);
   U3791 : NAND4_X1 port map( A1 => n4341, A2 => n4342, A3 => n4343, A4 => 
                           n4344, ZN => n4276);
   U3792 : NOR2_X1 port map( A1 => n2742, A2 => n12671, ZN => N8767);
   U3793 : NOR4_X1 port map( A1 => n2743, A2 => n2744, A3 => n2745, A4 => n2746
                           , ZN => n2742);
   U3794 : NAND4_X1 port map( A1 => n2939, A2 => n2940, A3 => n2941, A4 => 
                           n2942, ZN => n2743);
   U3795 : NAND4_X1 port map( A1 => n2873, A2 => n2874, A3 => n2875, A4 => 
                           n2876, ZN => n2744);
   U3796 : OAI222_X1 port map( A1 => n12779, A2 => n2481, B1 => n2482, B2 => 
                           n2480, C1 => n2936, C2 => n14517, ZN => n9133);
   U3797 : INV_X1 port map( A => n2482, ZN => n12779);
   U3798 : XNOR2_X1 port map( A => n10626, B => n2937, ZN => n2482);
   U3799 : OAI21_X1 port map( B1 => RETRN, B2 => CALL, A => ENABLE, ZN => n2478
                           );
   U3800 : OR3_X1 port map( A1 => n10626, A2 => n2935, A3 => n10625, ZN => 
                           n2489);
   U3801 : OAI221_X1 port map( B1 => n2483, B2 => n2484, C1 => n2935, C2 => 
                           n2485, A => n2486, ZN => n9132);
   U3802 : NAND2_X1 port map( A1 => RETRN, A2 => n14517, ZN => n2484);
   U3803 : NAND4_X1 port map( A1 => n12777, A2 => n2935, A3 => n10626, A4 => 
                           n10625, ZN => n2486);
   U3804 : AOI211_X1 port map( C1 => n12777, C2 => n2487, A => n2478, B => 
                           n2488, ZN => n2485);
   U3805 : OAI22_X1 port map( A1 => n10844, A2 => n12317, B1 => n10511, B2 => 
                           n12318, ZN => n8843);
   U3806 : OAI22_X1 port map( A1 => n10837, A2 => n12317, B1 => n10479, B2 => 
                           n12318, ZN => n8842);
   U3807 : OAI22_X1 port map( A1 => n10830, A2 => n12317, B1 => n10447, B2 => 
                           n12318, ZN => n8841);
   U3808 : OAI22_X1 port map( A1 => n10823, A2 => n12317, B1 => n10415, B2 => 
                           n12318, ZN => n8840);
   U3809 : OAI22_X1 port map( A1 => n10816, A2 => n12317, B1 => n10380, B2 => 
                           n12319, ZN => n8839);
   U3810 : OAI22_X1 port map( A1 => n10809, A2 => n12317, B1 => n10348, B2 => 
                           n12319, ZN => n8838);
   U3811 : OAI22_X1 port map( A1 => n10802, A2 => n12317, B1 => n10316, B2 => 
                           n12319, ZN => n8837);
   U3812 : OAI22_X1 port map( A1 => n10795, A2 => n12317, B1 => n10281, B2 => 
                           n12319, ZN => n8836);
   U3813 : OAI22_X1 port map( A1 => n10788, A2 => n12316, B1 => n10249, B2 => 
                           n12320, ZN => n8835);
   U3814 : OAI22_X1 port map( A1 => n10781, A2 => n12316, B1 => n10217, B2 => 
                           n12320, ZN => n8834);
   U3815 : OAI22_X1 port map( A1 => n10774, A2 => n12316, B1 => n10183, B2 => 
                           n12320, ZN => n8833);
   U3816 : OAI22_X1 port map( A1 => n10767, A2 => n12316, B1 => n10151, B2 => 
                           n12320, ZN => n8832);
   U3817 : OAI22_X1 port map( A1 => n10760, A2 => n12316, B1 => n10119, B2 => 
                           n12321, ZN => n8831);
   U3818 : OAI22_X1 port map( A1 => n10753, A2 => n12316, B1 => n10087, B2 => 
                           n12321, ZN => n8830);
   U3819 : OAI22_X1 port map( A1 => n10746, A2 => n12316, B1 => n10055, B2 => 
                           n12321, ZN => n8829);
   U3820 : OAI22_X1 port map( A1 => n10739, A2 => n12316, B1 => n10023, B2 => 
                           n12321, ZN => n8828);
   U3821 : OAI22_X1 port map( A1 => n10732, A2 => n12316, B1 => n9661, B2 => 
                           n12322, ZN => n8827);
   U3822 : OAI22_X1 port map( A1 => n10725, A2 => n12316, B1 => n9629, B2 => 
                           n12322, ZN => n8826);
   U3823 : OAI22_X1 port map( A1 => n10718, A2 => n12316, B1 => n9597, B2 => 
                           n12322, ZN => n8825);
   U3824 : OAI22_X1 port map( A1 => n10711, A2 => n12316, B1 => n9263, B2 => 
                           n12322, ZN => n8824);
   U3825 : OAI22_X1 port map( A1 => n10704, A2 => n12315, B1 => n9199, B2 => 
                           n12323, ZN => n8823);
   U3826 : OAI22_X1 port map( A1 => n10697, A2 => n12315, B1 => n9167, B2 => 
                           n12323, ZN => n8822);
   U3827 : OAI22_X1 port map( A1 => n10690, A2 => n12315, B1 => n9135, B2 => 
                           n12323, ZN => n8821);
   U3828 : OAI22_X1 port map( A1 => n10683, A2 => n12315, B1 => n6000, B2 => 
                           n12323, ZN => n8820);
   U3829 : OAI22_X1 port map( A1 => n10676, A2 => n12315, B1 => n5936, B2 => 
                           n12324, ZN => n8819);
   U3830 : OAI22_X1 port map( A1 => n10669, A2 => n12315, B1 => n5904, B2 => 
                           n12324, ZN => n8818);
   U3831 : OAI22_X1 port map( A1 => n10662, A2 => n12315, B1 => n5872, B2 => 
                           n12324, ZN => n8817);
   U3832 : OAI22_X1 port map( A1 => n10655, A2 => n12315, B1 => n5840, B2 => 
                           n12324, ZN => n8816);
   U3833 : OAI22_X1 port map( A1 => n10648, A2 => n12315, B1 => n5808, B2 => 
                           n12325, ZN => n8815);
   U3834 : OAI22_X1 port map( A1 => n10641, A2 => n12315, B1 => n5776, B2 => 
                           n12325, ZN => n8814);
   U3835 : OAI22_X1 port map( A1 => n10634, A2 => n12315, B1 => n5744, B2 => 
                           n12325, ZN => n8813);
   U3836 : OAI22_X1 port map( A1 => n10627, A2 => n12315, B1 => n5712, B2 => 
                           n12325, ZN => n8812);
   U3837 : OAI22_X1 port map( A1 => n10628, A2 => n12267, B1 => n996, B2 => 
                           n12270, ZN => n8684);
   U3838 : OAI22_X1 port map( A1 => n10628, A2 => n12231, B1 => n997, B2 => 
                           n12234, ZN => n8588);
   U3839 : OAI22_X1 port map( A1 => n10628, A2 => n12195, B1 => n998, B2 => 
                           n12198, ZN => n8492);
   U3840 : OAI22_X1 port map( A1 => n10846, A2 => n12089, B1 => n10516, B2 => 
                           n12090, ZN => n8235);
   U3841 : OAI22_X1 port map( A1 => n10839, A2 => n12089, B1 => n10484, B2 => 
                           n12090, ZN => n8234);
   U3842 : OAI22_X1 port map( A1 => n10832, A2 => n12089, B1 => n10452, B2 => 
                           n12090, ZN => n8233);
   U3843 : OAI22_X1 port map( A1 => n10825, A2 => n12089, B1 => n10420, B2 => 
                           n12090, ZN => n8232);
   U3844 : OAI22_X1 port map( A1 => n10818, A2 => n12089, B1 => n10385, B2 => 
                           n12091, ZN => n8231);
   U3845 : OAI22_X1 port map( A1 => n10811, A2 => n12089, B1 => n10353, B2 => 
                           n12091, ZN => n8230);
   U3846 : OAI22_X1 port map( A1 => n10804, A2 => n12089, B1 => n10321, B2 => 
                           n12091, ZN => n8229);
   U3847 : OAI22_X1 port map( A1 => n10797, A2 => n12089, B1 => n10286, B2 => 
                           n12091, ZN => n8228);
   U3848 : OAI22_X1 port map( A1 => n10790, A2 => n12088, B1 => n10254, B2 => 
                           n12092, ZN => n8227);
   U3849 : OAI22_X1 port map( A1 => n10783, A2 => n12088, B1 => n10222, B2 => 
                           n12092, ZN => n8226);
   U3850 : OAI22_X1 port map( A1 => n10776, A2 => n12088, B1 => n10188, B2 => 
                           n12092, ZN => n8225);
   U3851 : OAI22_X1 port map( A1 => n10769, A2 => n12088, B1 => n10156, B2 => 
                           n12092, ZN => n8224);
   U3852 : OAI22_X1 port map( A1 => n10762, A2 => n12088, B1 => n10124, B2 => 
                           n12093, ZN => n8223);
   U3853 : OAI22_X1 port map( A1 => n10755, A2 => n12088, B1 => n10092, B2 => 
                           n12093, ZN => n8222);
   U3854 : OAI22_X1 port map( A1 => n10748, A2 => n12088, B1 => n10060, B2 => 
                           n12093, ZN => n8221);
   U3855 : OAI22_X1 port map( A1 => n10741, A2 => n12088, B1 => n10028, B2 => 
                           n12093, ZN => n8220);
   U3856 : OAI22_X1 port map( A1 => n10734, A2 => n12088, B1 => n9698, B2 => 
                           n12094, ZN => n8219);
   U3857 : OAI22_X1 port map( A1 => n10727, A2 => n12088, B1 => n9634, B2 => 
                           n12094, ZN => n8218);
   U3858 : OAI22_X1 port map( A1 => n10720, A2 => n12088, B1 => n9602, B2 => 
                           n12094, ZN => n8217);
   U3859 : OAI22_X1 port map( A1 => n10713, A2 => n12088, B1 => n9570, B2 => 
                           n12094, ZN => n8216);
   U3860 : OAI22_X1 port map( A1 => n10706, A2 => n12087, B1 => n9204, B2 => 
                           n12095, ZN => n8215);
   U3861 : OAI22_X1 port map( A1 => n10699, A2 => n12087, B1 => n9172, B2 => 
                           n12095, ZN => n8214);
   U3862 : OAI22_X1 port map( A1 => n10692, A2 => n12087, B1 => n9140, B2 => 
                           n12095, ZN => n8213);
   U3863 : OAI22_X1 port map( A1 => n10685, A2 => n12087, B1 => n6005, B2 => 
                           n12095, ZN => n8212);
   U3864 : OAI22_X1 port map( A1 => n10678, A2 => n12087, B1 => n5941, B2 => 
                           n12096, ZN => n8211);
   U3865 : OAI22_X1 port map( A1 => n10671, A2 => n12087, B1 => n5909, B2 => 
                           n12096, ZN => n8210);
   U3866 : OAI22_X1 port map( A1 => n10664, A2 => n12087, B1 => n5877, B2 => 
                           n12096, ZN => n8209);
   U3867 : OAI22_X1 port map( A1 => n10657, A2 => n12087, B1 => n5845, B2 => 
                           n12096, ZN => n8208);
   U3868 : OAI22_X1 port map( A1 => n10650, A2 => n12087, B1 => n5813, B2 => 
                           n12097, ZN => n8207);
   U3869 : OAI22_X1 port map( A1 => n10643, A2 => n12087, B1 => n5781, B2 => 
                           n12097, ZN => n8206);
   U3870 : OAI22_X1 port map( A1 => n10636, A2 => n12087, B1 => n5749, B2 => 
                           n12097, ZN => n8205);
   U3871 : OAI22_X1 port map( A1 => n10629, A2 => n12087, B1 => n5717, B2 => 
                           n12097, ZN => n8204);
   U3872 : OAI22_X1 port map( A1 => n10846, A2 => n12053, B1 => n10519, B2 => 
                           n12054, ZN => n8139);
   U3873 : OAI22_X1 port map( A1 => n10839, A2 => n12053, B1 => n10487, B2 => 
                           n12054, ZN => n8138);
   U3874 : OAI22_X1 port map( A1 => n10832, A2 => n12053, B1 => n10455, B2 => 
                           n12054, ZN => n8137);
   U3875 : OAI22_X1 port map( A1 => n10825, A2 => n12053, B1 => n10423, B2 => 
                           n12054, ZN => n8136);
   U3876 : OAI22_X1 port map( A1 => n10818, A2 => n12053, B1 => n10388, B2 => 
                           n12055, ZN => n8135);
   U3877 : OAI22_X1 port map( A1 => n10811, A2 => n12053, B1 => n10356, B2 => 
                           n12055, ZN => n8134);
   U3878 : OAI22_X1 port map( A1 => n10804, A2 => n12053, B1 => n10324, B2 => 
                           n12055, ZN => n8133);
   U3879 : OAI22_X1 port map( A1 => n10797, A2 => n12053, B1 => n10289, B2 => 
                           n12055, ZN => n8132);
   U3880 : OAI22_X1 port map( A1 => n10790, A2 => n12052, B1 => n10257, B2 => 
                           n12056, ZN => n8131);
   U3881 : OAI22_X1 port map( A1 => n10783, A2 => n12052, B1 => n10225, B2 => 
                           n12056, ZN => n8130);
   U3882 : OAI22_X1 port map( A1 => n10776, A2 => n12052, B1 => n10191, B2 => 
                           n12056, ZN => n8129);
   U3883 : OAI22_X1 port map( A1 => n10769, A2 => n12052, B1 => n10159, B2 => 
                           n12056, ZN => n8128);
   U3884 : OAI22_X1 port map( A1 => n10762, A2 => n12052, B1 => n10127, B2 => 
                           n12057, ZN => n8127);
   U3885 : OAI22_X1 port map( A1 => n10755, A2 => n12052, B1 => n10095, B2 => 
                           n12057, ZN => n8126);
   U3886 : OAI22_X1 port map( A1 => n10748, A2 => n12052, B1 => n10063, B2 => 
                           n12057, ZN => n8125);
   U3887 : OAI22_X1 port map( A1 => n10741, A2 => n12052, B1 => n10031, B2 => 
                           n12057, ZN => n8124);
   U3888 : OAI22_X1 port map( A1 => n10734, A2 => n12052, B1 => n9701, B2 => 
                           n12058, ZN => n8123);
   U3889 : OAI22_X1 port map( A1 => n10727, A2 => n12052, B1 => n9637, B2 => 
                           n12058, ZN => n8122);
   U3890 : OAI22_X1 port map( A1 => n10720, A2 => n12052, B1 => n9605, B2 => 
                           n12058, ZN => n8121);
   U3891 : OAI22_X1 port map( A1 => n10713, A2 => n12052, B1 => n9573, B2 => 
                           n12058, ZN => n8120);
   U3892 : OAI22_X1 port map( A1 => n10706, A2 => n12051, B1 => n9207, B2 => 
                           n12059, ZN => n8119);
   U3893 : OAI22_X1 port map( A1 => n10699, A2 => n12051, B1 => n9175, B2 => 
                           n12059, ZN => n8118);
   U3894 : OAI22_X1 port map( A1 => n10692, A2 => n12051, B1 => n9143, B2 => 
                           n12059, ZN => n8117);
   U3895 : OAI22_X1 port map( A1 => n10685, A2 => n12051, B1 => n6008, B2 => 
                           n12059, ZN => n8116);
   U3896 : OAI22_X1 port map( A1 => n10678, A2 => n12051, B1 => n5944, B2 => 
                           n12060, ZN => n8115);
   U3897 : OAI22_X1 port map( A1 => n10671, A2 => n12051, B1 => n5912, B2 => 
                           n12060, ZN => n8114);
   U3898 : OAI22_X1 port map( A1 => n10664, A2 => n12051, B1 => n5880, B2 => 
                           n12060, ZN => n8113);
   U3899 : OAI22_X1 port map( A1 => n10657, A2 => n12051, B1 => n5848, B2 => 
                           n12060, ZN => n8112);
   U3900 : OAI22_X1 port map( A1 => n10650, A2 => n12051, B1 => n5816, B2 => 
                           n12061, ZN => n8111);
   U3901 : OAI22_X1 port map( A1 => n10643, A2 => n12051, B1 => n5784, B2 => 
                           n12061, ZN => n8110);
   U3902 : OAI22_X1 port map( A1 => n10636, A2 => n12051, B1 => n5752, B2 => 
                           n12061, ZN => n8109);
   U3903 : OAI22_X1 port map( A1 => n10629, A2 => n12051, B1 => n5720, B2 => 
                           n12061, ZN => n8108);
   U3904 : OAI22_X1 port map( A1 => n10847, A2 => n11825, B1 => n10524, B2 => 
                           n11826, ZN => n7531);
   U3905 : OAI22_X1 port map( A1 => n10840, A2 => n11825, B1 => n10492, B2 => 
                           n11826, ZN => n7530);
   U3906 : OAI22_X1 port map( A1 => n10833, A2 => n11825, B1 => n10460, B2 => 
                           n11826, ZN => n7529);
   U3907 : OAI22_X1 port map( A1 => n10826, A2 => n11825, B1 => n10428, B2 => 
                           n11826, ZN => n7528);
   U3908 : OAI22_X1 port map( A1 => n10819, A2 => n11825, B1 => n10393, B2 => 
                           n11827, ZN => n7527);
   U3909 : OAI22_X1 port map( A1 => n10812, A2 => n11825, B1 => n10361, B2 => 
                           n11827, ZN => n7526);
   U3910 : OAI22_X1 port map( A1 => n10805, A2 => n11825, B1 => n10329, B2 => 
                           n11827, ZN => n7525);
   U3911 : OAI22_X1 port map( A1 => n10798, A2 => n11825, B1 => n10294, B2 => 
                           n11827, ZN => n7524);
   U3912 : OAI22_X1 port map( A1 => n10791, A2 => n11824, B1 => n10262, B2 => 
                           n11828, ZN => n7523);
   U3913 : OAI22_X1 port map( A1 => n10784, A2 => n11824, B1 => n10230, B2 => 
                           n11828, ZN => n7522);
   U3914 : OAI22_X1 port map( A1 => n10777, A2 => n11824, B1 => n10196, B2 => 
                           n11828, ZN => n7521);
   U3915 : OAI22_X1 port map( A1 => n10770, A2 => n11824, B1 => n10164, B2 => 
                           n11828, ZN => n7520);
   U3916 : OAI22_X1 port map( A1 => n10763, A2 => n11824, B1 => n10132, B2 => 
                           n11829, ZN => n7519);
   U3917 : OAI22_X1 port map( A1 => n10756, A2 => n11824, B1 => n10100, B2 => 
                           n11829, ZN => n7518);
   U3918 : OAI22_X1 port map( A1 => n10749, A2 => n11824, B1 => n10068, B2 => 
                           n11829, ZN => n7517);
   U3919 : OAI22_X1 port map( A1 => n10742, A2 => n11824, B1 => n10036, B2 => 
                           n11829, ZN => n7516);
   U3920 : OAI22_X1 port map( A1 => n10735, A2 => n11824, B1 => n10004, B2 => 
                           n11830, ZN => n7515);
   U3921 : OAI22_X1 port map( A1 => n10728, A2 => n11824, B1 => n9642, B2 => 
                           n11830, ZN => n7514);
   U3922 : OAI22_X1 port map( A1 => n10721, A2 => n11824, B1 => n9610, B2 => 
                           n11830, ZN => n7513);
   U3923 : OAI22_X1 port map( A1 => n10714, A2 => n11824, B1 => n9578, B2 => 
                           n11830, ZN => n7512);
   U3924 : OAI22_X1 port map( A1 => n10707, A2 => n11823, B1 => n9212, B2 => 
                           n11831, ZN => n7511);
   U3925 : OAI22_X1 port map( A1 => n10700, A2 => n11823, B1 => n9180, B2 => 
                           n11831, ZN => n7510);
   U3926 : OAI22_X1 port map( A1 => n10693, A2 => n11823, B1 => n9148, B2 => 
                           n11831, ZN => n7509);
   U3927 : OAI22_X1 port map( A1 => n10686, A2 => n11823, B1 => n6044, B2 => 
                           n11831, ZN => n7508);
   U3928 : OAI22_X1 port map( A1 => n10679, A2 => n11823, B1 => n5981, B2 => 
                           n11832, ZN => n7507);
   U3929 : OAI22_X1 port map( A1 => n10672, A2 => n11823, B1 => n5917, B2 => 
                           n11832, ZN => n7506);
   U3930 : OAI22_X1 port map( A1 => n10665, A2 => n11823, B1 => n5885, B2 => 
                           n11832, ZN => n7505);
   U3931 : OAI22_X1 port map( A1 => n10658, A2 => n11823, B1 => n5853, B2 => 
                           n11832, ZN => n7504);
   U3932 : OAI22_X1 port map( A1 => n10651, A2 => n11823, B1 => n5821, B2 => 
                           n11833, ZN => n7503);
   U3933 : OAI22_X1 port map( A1 => n10644, A2 => n11823, B1 => n5789, B2 => 
                           n11833, ZN => n7502);
   U3934 : OAI22_X1 port map( A1 => n10637, A2 => n11823, B1 => n5757, B2 => 
                           n11833, ZN => n7501);
   U3935 : OAI22_X1 port map( A1 => n10630, A2 => n11823, B1 => n5725, B2 => 
                           n11833, ZN => n7500);
   U3936 : OAI22_X1 port map( A1 => n10848, A2 => n11789, B1 => n10527, B2 => 
                           n11790, ZN => n7435);
   U3937 : OAI22_X1 port map( A1 => n10841, A2 => n11789, B1 => n10495, B2 => 
                           n11790, ZN => n7434);
   U3938 : OAI22_X1 port map( A1 => n10834, A2 => n11789, B1 => n10463, B2 => 
                           n11790, ZN => n7433);
   U3939 : OAI22_X1 port map( A1 => n10827, A2 => n11789, B1 => n10431, B2 => 
                           n11790, ZN => n7432);
   U3940 : OAI22_X1 port map( A1 => n10820, A2 => n11789, B1 => n10396, B2 => 
                           n11791, ZN => n7431);
   U3941 : OAI22_X1 port map( A1 => n10813, A2 => n11789, B1 => n10364, B2 => 
                           n11791, ZN => n7430);
   U3942 : OAI22_X1 port map( A1 => n10806, A2 => n11789, B1 => n10332, B2 => 
                           n11791, ZN => n7429);
   U3943 : OAI22_X1 port map( A1 => n10799, A2 => n11789, B1 => n10297, B2 => 
                           n11791, ZN => n7428);
   U3944 : OAI22_X1 port map( A1 => n10792, A2 => n11788, B1 => n10265, B2 => 
                           n11792, ZN => n7427);
   U3945 : OAI22_X1 port map( A1 => n10785, A2 => n11788, B1 => n10233, B2 => 
                           n11792, ZN => n7426);
   U3946 : OAI22_X1 port map( A1 => n10778, A2 => n11788, B1 => n10199, B2 => 
                           n11792, ZN => n7425);
   U3947 : OAI22_X1 port map( A1 => n10771, A2 => n11788, B1 => n10167, B2 => 
                           n11792, ZN => n7424);
   U3948 : OAI22_X1 port map( A1 => n10764, A2 => n11788, B1 => n10135, B2 => 
                           n11793, ZN => n7423);
   U3949 : OAI22_X1 port map( A1 => n10757, A2 => n11788, B1 => n10103, B2 => 
                           n11793, ZN => n7422);
   U3950 : OAI22_X1 port map( A1 => n10750, A2 => n11788, B1 => n10071, B2 => 
                           n11793, ZN => n7421);
   U3951 : OAI22_X1 port map( A1 => n10743, A2 => n11788, B1 => n10039, B2 => 
                           n11793, ZN => n7420);
   U3952 : OAI22_X1 port map( A1 => n10736, A2 => n11788, B1 => n10007, B2 => 
                           n11794, ZN => n7419);
   U3953 : OAI22_X1 port map( A1 => n10729, A2 => n11788, B1 => n9645, B2 => 
                           n11794, ZN => n7418);
   U3954 : OAI22_X1 port map( A1 => n10722, A2 => n11788, B1 => n9613, B2 => 
                           n11794, ZN => n7417);
   U3955 : OAI22_X1 port map( A1 => n10715, A2 => n11788, B1 => n9581, B2 => 
                           n11794, ZN => n7416);
   U3956 : OAI22_X1 port map( A1 => n10708, A2 => n11787, B1 => n9215, B2 => 
                           n11795, ZN => n7415);
   U3957 : OAI22_X1 port map( A1 => n10701, A2 => n11787, B1 => n9183, B2 => 
                           n11795, ZN => n7414);
   U3958 : OAI22_X1 port map( A1 => n10694, A2 => n11787, B1 => n9151, B2 => 
                           n11795, ZN => n7413);
   U3959 : OAI22_X1 port map( A1 => n10687, A2 => n11787, B1 => n6301, B2 => 
                           n11795, ZN => n7412);
   U3960 : OAI22_X1 port map( A1 => n10680, A2 => n11787, B1 => n5984, B2 => 
                           n11796, ZN => n7411);
   U3961 : OAI22_X1 port map( A1 => n10673, A2 => n11787, B1 => n5920, B2 => 
                           n11796, ZN => n7410);
   U3962 : OAI22_X1 port map( A1 => n10666, A2 => n11787, B1 => n5888, B2 => 
                           n11796, ZN => n7409);
   U3963 : OAI22_X1 port map( A1 => n10659, A2 => n11787, B1 => n5856, B2 => 
                           n11796, ZN => n7408);
   U3964 : OAI22_X1 port map( A1 => n10652, A2 => n11787, B1 => n5824, B2 => 
                           n11797, ZN => n7407);
   U3965 : OAI22_X1 port map( A1 => n10645, A2 => n11787, B1 => n5792, B2 => 
                           n11797, ZN => n7406);
   U3966 : OAI22_X1 port map( A1 => n10638, A2 => n11787, B1 => n5760, B2 => 
                           n11797, ZN => n7405);
   U3967 : OAI22_X1 port map( A1 => n10631, A2 => n11787, B1 => n5728, B2 => 
                           n11797, ZN => n7404);
   U3968 : OAI22_X1 port map( A1 => n10849, A2 => n11525, B1 => n10535, B2 => 
                           n11526, ZN => n6731);
   U3969 : OAI22_X1 port map( A1 => n10842, A2 => n11525, B1 => n10503, B2 => 
                           n11526, ZN => n6730);
   U3970 : OAI22_X1 port map( A1 => n10835, A2 => n11525, B1 => n10471, B2 => 
                           n11526, ZN => n6729);
   U3971 : OAI22_X1 port map( A1 => n10828, A2 => n11525, B1 => n10439, B2 => 
                           n11526, ZN => n6728);
   U3972 : OAI22_X1 port map( A1 => n10821, A2 => n11525, B1 => n10407, B2 => 
                           n11527, ZN => n6727);
   U3973 : OAI22_X1 port map( A1 => n10814, A2 => n11525, B1 => n10372, B2 => 
                           n11527, ZN => n6726);
   U3974 : OAI22_X1 port map( A1 => n10807, A2 => n11525, B1 => n10340, B2 => 
                           n11527, ZN => n6725);
   U3975 : OAI22_X1 port map( A1 => n10800, A2 => n11525, B1 => n10308, B2 => 
                           n11527, ZN => n6724);
   U3976 : OAI22_X1 port map( A1 => n10793, A2 => n11524, B1 => n10273, B2 => 
                           n11528, ZN => n6723);
   U3977 : OAI22_X1 port map( A1 => n10786, A2 => n11524, B1 => n10241, B2 => 
                           n11528, ZN => n6722);
   U3978 : OAI22_X1 port map( A1 => n10779, A2 => n11524, B1 => n10209, B2 => 
                           n11528, ZN => n6721);
   U3979 : OAI22_X1 port map( A1 => n10772, A2 => n11524, B1 => n10175, B2 => 
                           n11528, ZN => n6720);
   U3980 : OAI22_X1 port map( A1 => n10765, A2 => n11524, B1 => n10143, B2 => 
                           n11529, ZN => n6719);
   U3981 : OAI22_X1 port map( A1 => n10758, A2 => n11524, B1 => n10111, B2 => 
                           n11529, ZN => n6718);
   U3982 : OAI22_X1 port map( A1 => n10751, A2 => n11524, B1 => n10079, B2 => 
                           n11529, ZN => n6717);
   U3983 : OAI22_X1 port map( A1 => n10744, A2 => n11524, B1 => n10047, B2 => 
                           n11529, ZN => n6716);
   U3984 : OAI22_X1 port map( A1 => n10737, A2 => n11524, B1 => n10015, B2 => 
                           n11530, ZN => n6715);
   U3985 : OAI22_X1 port map( A1 => n10730, A2 => n11524, B1 => n9653, B2 => 
                           n11530, ZN => n6714);
   U3986 : OAI22_X1 port map( A1 => n10723, A2 => n11524, B1 => n9621, B2 => 
                           n11530, ZN => n6713);
   U3987 : OAI22_X1 port map( A1 => n10716, A2 => n11524, B1 => n9589, B2 => 
                           n11530, ZN => n6712);
   U3988 : OAI22_X1 port map( A1 => n10709, A2 => n11523, B1 => n9255, B2 => 
                           n11531, ZN => n6711);
   U3989 : OAI22_X1 port map( A1 => n10702, A2 => n11523, B1 => n9191, B2 => 
                           n11531, ZN => n6710);
   U3990 : OAI22_X1 port map( A1 => n10695, A2 => n11523, B1 => n9159, B2 => 
                           n11531, ZN => n6709);
   U3991 : OAI22_X1 port map( A1 => n10688, A2 => n11523, B1 => n6309, B2 => 
                           n11531, ZN => n6708);
   U3992 : OAI22_X1 port map( A1 => n10681, A2 => n11523, B1 => n5992, B2 => 
                           n11532, ZN => n6707);
   U3993 : OAI22_X1 port map( A1 => n10674, A2 => n11523, B1 => n5928, B2 => 
                           n11532, ZN => n6706);
   U3994 : OAI22_X1 port map( A1 => n10667, A2 => n11523, B1 => n5896, B2 => 
                           n11532, ZN => n6705);
   U3995 : OAI22_X1 port map( A1 => n10660, A2 => n11523, B1 => n5864, B2 => 
                           n11532, ZN => n6704);
   U3996 : OAI22_X1 port map( A1 => n10653, A2 => n11523, B1 => n5832, B2 => 
                           n11533, ZN => n6703);
   U3997 : OAI22_X1 port map( A1 => n10646, A2 => n11523, B1 => n5800, B2 => 
                           n11533, ZN => n6702);
   U3998 : OAI22_X1 port map( A1 => n10639, A2 => n11523, B1 => n5768, B2 => 
                           n11533, ZN => n6701);
   U3999 : OAI22_X1 port map( A1 => n10632, A2 => n11523, B1 => n5736, B2 => 
                           n11533, ZN => n6700);
   U4000 : OAI22_X1 port map( A1 => n10850, A2 => n11477, B1 => n1409, B2 => 
                           n11478, ZN => n6603);
   U4001 : OAI22_X1 port map( A1 => n10843, A2 => n11477, B1 => n1397, B2 => 
                           n11478, ZN => n6602);
   U4002 : OAI22_X1 port map( A1 => n10836, A2 => n11477, B1 => n1385, B2 => 
                           n11478, ZN => n6601);
   U4003 : OAI22_X1 port map( A1 => n10829, A2 => n11477, B1 => n1341, B2 => 
                           n11478, ZN => n6600);
   U4004 : OAI22_X1 port map( A1 => n10822, A2 => n11477, B1 => n1329, B2 => 
                           n11479, ZN => n6599);
   U4005 : OAI22_X1 port map( A1 => n10815, A2 => n11477, B1 => n1317, B2 => 
                           n11479, ZN => n6598);
   U4006 : OAI22_X1 port map( A1 => n10808, A2 => n11477, B1 => n1305, B2 => 
                           n11479, ZN => n6597);
   U4007 : OAI22_X1 port map( A1 => n10801, A2 => n11477, B1 => n1293, B2 => 
                           n11479, ZN => n6596);
   U4008 : OAI22_X1 port map( A1 => n10794, A2 => n11476, B1 => n1281, B2 => 
                           n11480, ZN => n6595);
   U4009 : OAI22_X1 port map( A1 => n10787, A2 => n11476, B1 => n1269, B2 => 
                           n11480, ZN => n6594);
   U4010 : OAI22_X1 port map( A1 => n10780, A2 => n11476, B1 => n1257, B2 => 
                           n11480, ZN => n6593);
   U4011 : OAI22_X1 port map( A1 => n10773, A2 => n11476, B1 => n1245, B2 => 
                           n11480, ZN => n6592);
   U4012 : OAI22_X1 port map( A1 => n10766, A2 => n11476, B1 => n1233, B2 => 
                           n11481, ZN => n6591);
   U4013 : OAI22_X1 port map( A1 => n10759, A2 => n11476, B1 => n1221, B2 => 
                           n11481, ZN => n6590);
   U4014 : OAI22_X1 port map( A1 => n10752, A2 => n11476, B1 => n1209, B2 => 
                           n11481, ZN => n6589);
   U4015 : OAI22_X1 port map( A1 => n10745, A2 => n11476, B1 => n1197, B2 => 
                           n11481, ZN => n6588);
   U4016 : OAI22_X1 port map( A1 => n10738, A2 => n11476, B1 => n1185, B2 => 
                           n11482, ZN => n6587);
   U4017 : OAI22_X1 port map( A1 => n10731, A2 => n11476, B1 => n1173, B2 => 
                           n11482, ZN => n6586);
   U4018 : OAI22_X1 port map( A1 => n10724, A2 => n11476, B1 => n1161, B2 => 
                           n11482, ZN => n6585);
   U4019 : OAI22_X1 port map( A1 => n10717, A2 => n11476, B1 => n1149, B2 => 
                           n11482, ZN => n6584);
   U4020 : OAI22_X1 port map( A1 => n10710, A2 => n11475, B1 => n1137, B2 => 
                           n11483, ZN => n6583);
   U4021 : OAI22_X1 port map( A1 => n10703, A2 => n11475, B1 => n1125, B2 => 
                           n11483, ZN => n6582);
   U4022 : OAI22_X1 port map( A1 => n10696, A2 => n11475, B1 => n1113, B2 => 
                           n11483, ZN => n6581);
   U4023 : OAI22_X1 port map( A1 => n10689, A2 => n11475, B1 => n1101, B2 => 
                           n11483, ZN => n6580);
   U4024 : OAI22_X1 port map( A1 => n10682, A2 => n11475, B1 => n1089, B2 => 
                           n11484, ZN => n6579);
   U4025 : OAI22_X1 port map( A1 => n10675, A2 => n11475, B1 => n1077, B2 => 
                           n11484, ZN => n6578);
   U4026 : OAI22_X1 port map( A1 => n10668, A2 => n11475, B1 => n1065, B2 => 
                           n11484, ZN => n6577);
   U4027 : OAI22_X1 port map( A1 => n10661, A2 => n11475, B1 => n1053, B2 => 
                           n11484, ZN => n6576);
   U4028 : OAI22_X1 port map( A1 => n10654, A2 => n11475, B1 => n1041, B2 => 
                           n11485, ZN => n6575);
   U4029 : OAI22_X1 port map( A1 => n10647, A2 => n11475, B1 => n1029, B2 => 
                           n11485, ZN => n6574);
   U4030 : OAI22_X1 port map( A1 => n10850, A2 => n11441, B1 => n1442, B2 => 
                           n11442, ZN => n6507);
   U4031 : OAI22_X1 port map( A1 => n10843, A2 => n11441, B1 => n1398, B2 => 
                           n11442, ZN => n6506);
   U4032 : OAI22_X1 port map( A1 => n10836, A2 => n11441, B1 => n1386, B2 => 
                           n11442, ZN => n6505);
   U4033 : OAI22_X1 port map( A1 => n10829, A2 => n11441, B1 => n1342, B2 => 
                           n11442, ZN => n6504);
   U4034 : OAI22_X1 port map( A1 => n10822, A2 => n11441, B1 => n1330, B2 => 
                           n11443, ZN => n6503);
   U4035 : OAI22_X1 port map( A1 => n10815, A2 => n11441, B1 => n1318, B2 => 
                           n11443, ZN => n6502);
   U4036 : OAI22_X1 port map( A1 => n10808, A2 => n11441, B1 => n1306, B2 => 
                           n11443, ZN => n6501);
   U4037 : OAI22_X1 port map( A1 => n10801, A2 => n11441, B1 => n1294, B2 => 
                           n11443, ZN => n6500);
   U4038 : OAI22_X1 port map( A1 => n10794, A2 => n11440, B1 => n1282, B2 => 
                           n11444, ZN => n6499);
   U4039 : OAI22_X1 port map( A1 => n10787, A2 => n11440, B1 => n1270, B2 => 
                           n11444, ZN => n6498);
   U4040 : OAI22_X1 port map( A1 => n10780, A2 => n11440, B1 => n1258, B2 => 
                           n11444, ZN => n6497);
   U4041 : OAI22_X1 port map( A1 => n10773, A2 => n11440, B1 => n1246, B2 => 
                           n11444, ZN => n6496);
   U4042 : OAI22_X1 port map( A1 => n10766, A2 => n11440, B1 => n1234, B2 => 
                           n11445, ZN => n6495);
   U4043 : OAI22_X1 port map( A1 => n10759, A2 => n11440, B1 => n1222, B2 => 
                           n11445, ZN => n6494);
   U4044 : OAI22_X1 port map( A1 => n10752, A2 => n11440, B1 => n1210, B2 => 
                           n11445, ZN => n6493);
   U4045 : OAI22_X1 port map( A1 => n10745, A2 => n11440, B1 => n1198, B2 => 
                           n11445, ZN => n6492);
   U4046 : OAI22_X1 port map( A1 => n10738, A2 => n11440, B1 => n1186, B2 => 
                           n11446, ZN => n6491);
   U4047 : OAI22_X1 port map( A1 => n10731, A2 => n11440, B1 => n1174, B2 => 
                           n11446, ZN => n6490);
   U4048 : OAI22_X1 port map( A1 => n10724, A2 => n11440, B1 => n1162, B2 => 
                           n11446, ZN => n6489);
   U4049 : OAI22_X1 port map( A1 => n10717, A2 => n11440, B1 => n1150, B2 => 
                           n11446, ZN => n6488);
   U4050 : OAI22_X1 port map( A1 => n10710, A2 => n11439, B1 => n1138, B2 => 
                           n11447, ZN => n6487);
   U4051 : OAI22_X1 port map( A1 => n10703, A2 => n11439, B1 => n1126, B2 => 
                           n11447, ZN => n6486);
   U4052 : OAI22_X1 port map( A1 => n10696, A2 => n11439, B1 => n1114, B2 => 
                           n11447, ZN => n6485);
   U4053 : OAI22_X1 port map( A1 => n10689, A2 => n11439, B1 => n1102, B2 => 
                           n11447, ZN => n6484);
   U4054 : OAI22_X1 port map( A1 => n10682, A2 => n11439, B1 => n1090, B2 => 
                           n11448, ZN => n6483);
   U4055 : OAI22_X1 port map( A1 => n10675, A2 => n11439, B1 => n1078, B2 => 
                           n11448, ZN => n6482);
   U4056 : OAI22_X1 port map( A1 => n10668, A2 => n11439, B1 => n1066, B2 => 
                           n11448, ZN => n6481);
   U4057 : OAI22_X1 port map( A1 => n10661, A2 => n11439, B1 => n1054, B2 => 
                           n11448, ZN => n6480);
   U4058 : OAI22_X1 port map( A1 => n10654, A2 => n11439, B1 => n1042, B2 => 
                           n11449, ZN => n6479);
   U4059 : OAI22_X1 port map( A1 => n10850, A2 => n11405, B1 => n1443, B2 => 
                           n11406, ZN => n6411);
   U4060 : OAI22_X1 port map( A1 => n10843, A2 => n11405, B1 => n1399, B2 => 
                           n11406, ZN => n6410);
   U4061 : OAI22_X1 port map( A1 => n10836, A2 => n11405, B1 => n1387, B2 => 
                           n11406, ZN => n6409);
   U4062 : OAI22_X1 port map( A1 => n10829, A2 => n11405, B1 => n1343, B2 => 
                           n11406, ZN => n6408);
   U4063 : OAI22_X1 port map( A1 => n10822, A2 => n11405, B1 => n1331, B2 => 
                           n11407, ZN => n6407);
   U4064 : OAI22_X1 port map( A1 => n10815, A2 => n11405, B1 => n1319, B2 => 
                           n11407, ZN => n6406);
   U4065 : OAI22_X1 port map( A1 => n10808, A2 => n11405, B1 => n1307, B2 => 
                           n11407, ZN => n6405);
   U4066 : OAI22_X1 port map( A1 => n10801, A2 => n11405, B1 => n1295, B2 => 
                           n11407, ZN => n6404);
   U4067 : OAI22_X1 port map( A1 => n10794, A2 => n11404, B1 => n1283, B2 => 
                           n11408, ZN => n6403);
   U4068 : OAI22_X1 port map( A1 => n10787, A2 => n11404, B1 => n1271, B2 => 
                           n11408, ZN => n6402);
   U4069 : OAI22_X1 port map( A1 => n10780, A2 => n11404, B1 => n1259, B2 => 
                           n11408, ZN => n6401);
   U4070 : OAI22_X1 port map( A1 => n10773, A2 => n11404, B1 => n1247, B2 => 
                           n11408, ZN => n6400);
   U4071 : OAI22_X1 port map( A1 => n10766, A2 => n11404, B1 => n1235, B2 => 
                           n11409, ZN => n6399);
   U4072 : OAI22_X1 port map( A1 => n10759, A2 => n11404, B1 => n1223, B2 => 
                           n11409, ZN => n6398);
   U4073 : OAI22_X1 port map( A1 => n10752, A2 => n11404, B1 => n1211, B2 => 
                           n11409, ZN => n6397);
   U4074 : OAI22_X1 port map( A1 => n10745, A2 => n11404, B1 => n1199, B2 => 
                           n11409, ZN => n6396);
   U4075 : OAI22_X1 port map( A1 => n10738, A2 => n11404, B1 => n1187, B2 => 
                           n11410, ZN => n6395);
   U4076 : OAI22_X1 port map( A1 => n10731, A2 => n11404, B1 => n1175, B2 => 
                           n11410, ZN => n6394);
   U4077 : OAI22_X1 port map( A1 => n10724, A2 => n11404, B1 => n1163, B2 => 
                           n11410, ZN => n6393);
   U4078 : OAI22_X1 port map( A1 => n10717, A2 => n11404, B1 => n1151, B2 => 
                           n11410, ZN => n6392);
   U4079 : OAI22_X1 port map( A1 => n10710, A2 => n11403, B1 => n1139, B2 => 
                           n11411, ZN => n6391);
   U4080 : OAI22_X1 port map( A1 => n10703, A2 => n11403, B1 => n1127, B2 => 
                           n11411, ZN => n6390);
   U4081 : OAI22_X1 port map( A1 => n10696, A2 => n11403, B1 => n1115, B2 => 
                           n11411, ZN => n6389);
   U4082 : OAI22_X1 port map( A1 => n10689, A2 => n11403, B1 => n1103, B2 => 
                           n11411, ZN => n6388);
   U4083 : OAI22_X1 port map( A1 => n10682, A2 => n11403, B1 => n1091, B2 => 
                           n11412, ZN => n6387);
   U4084 : OAI22_X1 port map( A1 => n10675, A2 => n11403, B1 => n1079, B2 => 
                           n11412, ZN => n6386);
   U4085 : OAI22_X1 port map( A1 => n10668, A2 => n11403, B1 => n1067, B2 => 
                           n11412, ZN => n6385);
   U4086 : OAI22_X1 port map( A1 => n10661, A2 => n11403, B1 => n1055, B2 => 
                           n11412, ZN => n6384);
   U4087 : OAI22_X1 port map( A1 => n10654, A2 => n11403, B1 => n1043, B2 => 
                           n11413, ZN => n6383);
   U4088 : OAI22_X1 port map( A1 => n10844, A2 => n12329, B1 => n10509, B2 => 
                           n12330, ZN => n8875);
   U4089 : OAI22_X1 port map( A1 => n10837, A2 => n12329, B1 => n10477, B2 => 
                           n12330, ZN => n8874);
   U4090 : OAI22_X1 port map( A1 => n10830, A2 => n12329, B1 => n10445, B2 => 
                           n12330, ZN => n8873);
   U4091 : OAI22_X1 port map( A1 => n10823, A2 => n12329, B1 => n10413, B2 => 
                           n12330, ZN => n8872);
   U4092 : OAI22_X1 port map( A1 => n10816, A2 => n12329, B1 => n10378, B2 => 
                           n12331, ZN => n8871);
   U4093 : OAI22_X1 port map( A1 => n10809, A2 => n12329, B1 => n10346, B2 => 
                           n12331, ZN => n8870);
   U4094 : OAI22_X1 port map( A1 => n10802, A2 => n12329, B1 => n10314, B2 => 
                           n12331, ZN => n8869);
   U4095 : OAI22_X1 port map( A1 => n10795, A2 => n12329, B1 => n10279, B2 => 
                           n12331, ZN => n8868);
   U4096 : OAI22_X1 port map( A1 => n10788, A2 => n12328, B1 => n10247, B2 => 
                           n12332, ZN => n8867);
   U4097 : OAI22_X1 port map( A1 => n10781, A2 => n12328, B1 => n10215, B2 => 
                           n12332, ZN => n8866);
   U4098 : OAI22_X1 port map( A1 => n10774, A2 => n12328, B1 => n10181, B2 => 
                           n12332, ZN => n8865);
   U4099 : OAI22_X1 port map( A1 => n10767, A2 => n12328, B1 => n10149, B2 => 
                           n12332, ZN => n8864);
   U4100 : OAI22_X1 port map( A1 => n10760, A2 => n12328, B1 => n10117, B2 => 
                           n12333, ZN => n8863);
   U4101 : OAI22_X1 port map( A1 => n10753, A2 => n12328, B1 => n10085, B2 => 
                           n12333, ZN => n8862);
   U4102 : OAI22_X1 port map( A1 => n10746, A2 => n12328, B1 => n10053, B2 => 
                           n12333, ZN => n8861);
   U4103 : OAI22_X1 port map( A1 => n10739, A2 => n12328, B1 => n10021, B2 => 
                           n12333, ZN => n8860);
   U4104 : OAI22_X1 port map( A1 => n10732, A2 => n12328, B1 => n9659, B2 => 
                           n12334, ZN => n8859);
   U4105 : OAI22_X1 port map( A1 => n10725, A2 => n12328, B1 => n9627, B2 => 
                           n12334, ZN => n8858);
   U4106 : OAI22_X1 port map( A1 => n10718, A2 => n12328, B1 => n9595, B2 => 
                           n12334, ZN => n8857);
   U4107 : OAI22_X1 port map( A1 => n10711, A2 => n12328, B1 => n9261, B2 => 
                           n12334, ZN => n8856);
   U4108 : OAI22_X1 port map( A1 => n10704, A2 => n12327, B1 => n9197, B2 => 
                           n12335, ZN => n8855);
   U4109 : OAI22_X1 port map( A1 => n10697, A2 => n12327, B1 => n9165, B2 => 
                           n12335, ZN => n8854);
   U4110 : OAI22_X1 port map( A1 => n10690, A2 => n12327, B1 => n6315, B2 => 
                           n12335, ZN => n8853);
   U4111 : OAI22_X1 port map( A1 => n10683, A2 => n12327, B1 => n5998, B2 => 
                           n12335, ZN => n8852);
   U4112 : OAI22_X1 port map( A1 => n10676, A2 => n12327, B1 => n5934, B2 => 
                           n12336, ZN => n8851);
   U4113 : OAI22_X1 port map( A1 => n10669, A2 => n12327, B1 => n5902, B2 => 
                           n12336, ZN => n8850);
   U4114 : OAI22_X1 port map( A1 => n10662, A2 => n12327, B1 => n5870, B2 => 
                           n12336, ZN => n8849);
   U4115 : OAI22_X1 port map( A1 => n10655, A2 => n12327, B1 => n5838, B2 => 
                           n12336, ZN => n8848);
   U4116 : OAI22_X1 port map( A1 => n10648, A2 => n12327, B1 => n5806, B2 => 
                           n12337, ZN => n8847);
   U4117 : OAI22_X1 port map( A1 => n10641, A2 => n12327, B1 => n5774, B2 => 
                           n12337, ZN => n8846);
   U4118 : OAI22_X1 port map( A1 => n10634, A2 => n12327, B1 => n5742, B2 => 
                           n12337, ZN => n8845);
   U4119 : OAI22_X1 port map( A1 => n10627, A2 => n12327, B1 => n5710, B2 => 
                           n12337, ZN => n8844);
   U4120 : OAI22_X1 port map( A1 => n10846, A2 => n12101, B1 => n10514, B2 => 
                           n12102, ZN => n8267);
   U4121 : OAI22_X1 port map( A1 => n10839, A2 => n12101, B1 => n10482, B2 => 
                           n12102, ZN => n8266);
   U4122 : OAI22_X1 port map( A1 => n10832, A2 => n12101, B1 => n10450, B2 => 
                           n12102, ZN => n8265);
   U4123 : OAI22_X1 port map( A1 => n10825, A2 => n12101, B1 => n10418, B2 => 
                           n12102, ZN => n8264);
   U4124 : OAI22_X1 port map( A1 => n10818, A2 => n12101, B1 => n10383, B2 => 
                           n12103, ZN => n8263);
   U4125 : OAI22_X1 port map( A1 => n10811, A2 => n12101, B1 => n10351, B2 => 
                           n12103, ZN => n8262);
   U4126 : OAI22_X1 port map( A1 => n10804, A2 => n12101, B1 => n10319, B2 => 
                           n12103, ZN => n8261);
   U4127 : OAI22_X1 port map( A1 => n10797, A2 => n12101, B1 => n10284, B2 => 
                           n12103, ZN => n8260);
   U4128 : OAI22_X1 port map( A1 => n10790, A2 => n12100, B1 => n10252, B2 => 
                           n12104, ZN => n8259);
   U4129 : OAI22_X1 port map( A1 => n10783, A2 => n12100, B1 => n10220, B2 => 
                           n12104, ZN => n8258);
   U4130 : OAI22_X1 port map( A1 => n10776, A2 => n12100, B1 => n10186, B2 => 
                           n12104, ZN => n8257);
   U4131 : OAI22_X1 port map( A1 => n10769, A2 => n12100, B1 => n10154, B2 => 
                           n12104, ZN => n8256);
   U4132 : OAI22_X1 port map( A1 => n10762, A2 => n12100, B1 => n10122, B2 => 
                           n12105, ZN => n8255);
   U4133 : OAI22_X1 port map( A1 => n10755, A2 => n12100, B1 => n10090, B2 => 
                           n12105, ZN => n8254);
   U4134 : OAI22_X1 port map( A1 => n10748, A2 => n12100, B1 => n10058, B2 => 
                           n12105, ZN => n8253);
   U4135 : OAI22_X1 port map( A1 => n10741, A2 => n12100, B1 => n10026, B2 => 
                           n12105, ZN => n8252);
   U4136 : OAI22_X1 port map( A1 => n10734, A2 => n12100, B1 => n9696, B2 => 
                           n12106, ZN => n8251);
   U4137 : OAI22_X1 port map( A1 => n10727, A2 => n12100, B1 => n9632, B2 => 
                           n12106, ZN => n8250);
   U4138 : OAI22_X1 port map( A1 => n10720, A2 => n12100, B1 => n9600, B2 => 
                           n12106, ZN => n8249);
   U4139 : OAI22_X1 port map( A1 => n10713, A2 => n12100, B1 => n9568, B2 => 
                           n12106, ZN => n8248);
   U4140 : OAI22_X1 port map( A1 => n10706, A2 => n12099, B1 => n9202, B2 => 
                           n12107, ZN => n8247);
   U4141 : OAI22_X1 port map( A1 => n10699, A2 => n12099, B1 => n9170, B2 => 
                           n12107, ZN => n8246);
   U4142 : OAI22_X1 port map( A1 => n10692, A2 => n12099, B1 => n9138, B2 => 
                           n12107, ZN => n8245);
   U4143 : OAI22_X1 port map( A1 => n10685, A2 => n12099, B1 => n6003, B2 => 
                           n12107, ZN => n8244);
   U4144 : OAI22_X1 port map( A1 => n10678, A2 => n12099, B1 => n5939, B2 => 
                           n12108, ZN => n8243);
   U4145 : OAI22_X1 port map( A1 => n10671, A2 => n12099, B1 => n5907, B2 => 
                           n12108, ZN => n8242);
   U4146 : OAI22_X1 port map( A1 => n10664, A2 => n12099, B1 => n5875, B2 => 
                           n12108, ZN => n8241);
   U4147 : OAI22_X1 port map( A1 => n10657, A2 => n12099, B1 => n5843, B2 => 
                           n12108, ZN => n8240);
   U4148 : OAI22_X1 port map( A1 => n10650, A2 => n12099, B1 => n5811, B2 => 
                           n12109, ZN => n8239);
   U4149 : OAI22_X1 port map( A1 => n10643, A2 => n12099, B1 => n5779, B2 => 
                           n12109, ZN => n8238);
   U4150 : OAI22_X1 port map( A1 => n10636, A2 => n12099, B1 => n5747, B2 => 
                           n12109, ZN => n8237);
   U4151 : OAI22_X1 port map( A1 => n10629, A2 => n12099, B1 => n5715, B2 => 
                           n12109, ZN => n8236);
   U4152 : OAI22_X1 port map( A1 => n10846, A2 => n12065, B1 => n10517, B2 => 
                           n12066, ZN => n8171);
   U4153 : OAI22_X1 port map( A1 => n10839, A2 => n12065, B1 => n10485, B2 => 
                           n12066, ZN => n8170);
   U4154 : OAI22_X1 port map( A1 => n10832, A2 => n12065, B1 => n10453, B2 => 
                           n12066, ZN => n8169);
   U4155 : OAI22_X1 port map( A1 => n10825, A2 => n12065, B1 => n10421, B2 => 
                           n12066, ZN => n8168);
   U4156 : OAI22_X1 port map( A1 => n10818, A2 => n12065, B1 => n10386, B2 => 
                           n12067, ZN => n8167);
   U4157 : OAI22_X1 port map( A1 => n10811, A2 => n12065, B1 => n10354, B2 => 
                           n12067, ZN => n8166);
   U4158 : OAI22_X1 port map( A1 => n10804, A2 => n12065, B1 => n10322, B2 => 
                           n12067, ZN => n8165);
   U4159 : OAI22_X1 port map( A1 => n10797, A2 => n12065, B1 => n10287, B2 => 
                           n12067, ZN => n8164);
   U4160 : OAI22_X1 port map( A1 => n10790, A2 => n12064, B1 => n10255, B2 => 
                           n12068, ZN => n8163);
   U4161 : OAI22_X1 port map( A1 => n10783, A2 => n12064, B1 => n10223, B2 => 
                           n12068, ZN => n8162);
   U4162 : OAI22_X1 port map( A1 => n10776, A2 => n12064, B1 => n10189, B2 => 
                           n12068, ZN => n8161);
   U4163 : OAI22_X1 port map( A1 => n10769, A2 => n12064, B1 => n10157, B2 => 
                           n12068, ZN => n8160);
   U4164 : OAI22_X1 port map( A1 => n10762, A2 => n12064, B1 => n10125, B2 => 
                           n12069, ZN => n8159);
   U4165 : OAI22_X1 port map( A1 => n10755, A2 => n12064, B1 => n10093, B2 => 
                           n12069, ZN => n8158);
   U4166 : OAI22_X1 port map( A1 => n10748, A2 => n12064, B1 => n10061, B2 => 
                           n12069, ZN => n8157);
   U4167 : OAI22_X1 port map( A1 => n10741, A2 => n12064, B1 => n10029, B2 => 
                           n12069, ZN => n8156);
   U4168 : OAI22_X1 port map( A1 => n10734, A2 => n12064, B1 => n9699, B2 => 
                           n12070, ZN => n8155);
   U4169 : OAI22_X1 port map( A1 => n10727, A2 => n12064, B1 => n9635, B2 => 
                           n12070, ZN => n8154);
   U4170 : OAI22_X1 port map( A1 => n10720, A2 => n12064, B1 => n9603, B2 => 
                           n12070, ZN => n8153);
   U4171 : OAI22_X1 port map( A1 => n10713, A2 => n12064, B1 => n9571, B2 => 
                           n12070, ZN => n8152);
   U4172 : OAI22_X1 port map( A1 => n10706, A2 => n12063, B1 => n9205, B2 => 
                           n12071, ZN => n8151);
   U4173 : OAI22_X1 port map( A1 => n10699, A2 => n12063, B1 => n9173, B2 => 
                           n12071, ZN => n8150);
   U4174 : OAI22_X1 port map( A1 => n10692, A2 => n12063, B1 => n9141, B2 => 
                           n12071, ZN => n8149);
   U4175 : OAI22_X1 port map( A1 => n10685, A2 => n12063, B1 => n6006, B2 => 
                           n12071, ZN => n8148);
   U4176 : OAI22_X1 port map( A1 => n10678, A2 => n12063, B1 => n5942, B2 => 
                           n12072, ZN => n8147);
   U4177 : OAI22_X1 port map( A1 => n10671, A2 => n12063, B1 => n5910, B2 => 
                           n12072, ZN => n8146);
   U4178 : OAI22_X1 port map( A1 => n10664, A2 => n12063, B1 => n5878, B2 => 
                           n12072, ZN => n8145);
   U4179 : OAI22_X1 port map( A1 => n10657, A2 => n12063, B1 => n5846, B2 => 
                           n12072, ZN => n8144);
   U4180 : OAI22_X1 port map( A1 => n10650, A2 => n12063, B1 => n5814, B2 => 
                           n12073, ZN => n8143);
   U4181 : OAI22_X1 port map( A1 => n10643, A2 => n12063, B1 => n5782, B2 => 
                           n12073, ZN => n8142);
   U4182 : OAI22_X1 port map( A1 => n10636, A2 => n12063, B1 => n5750, B2 => 
                           n12073, ZN => n8141);
   U4183 : OAI22_X1 port map( A1 => n10629, A2 => n12063, B1 => n5718, B2 => 
                           n12073, ZN => n8140);
   U4184 : OAI22_X1 port map( A1 => n10847, A2 => n11837, B1 => n10522, B2 => 
                           n11838, ZN => n7563);
   U4185 : OAI22_X1 port map( A1 => n10840, A2 => n11837, B1 => n10490, B2 => 
                           n11838, ZN => n7562);
   U4186 : OAI22_X1 port map( A1 => n10833, A2 => n11837, B1 => n10458, B2 => 
                           n11838, ZN => n7561);
   U4187 : OAI22_X1 port map( A1 => n10826, A2 => n11837, B1 => n10426, B2 => 
                           n11838, ZN => n7560);
   U4188 : OAI22_X1 port map( A1 => n10819, A2 => n11837, B1 => n10391, B2 => 
                           n11839, ZN => n7559);
   U4189 : OAI22_X1 port map( A1 => n10812, A2 => n11837, B1 => n10359, B2 => 
                           n11839, ZN => n7558);
   U4190 : OAI22_X1 port map( A1 => n10805, A2 => n11837, B1 => n10327, B2 => 
                           n11839, ZN => n7557);
   U4191 : OAI22_X1 port map( A1 => n10798, A2 => n11837, B1 => n10292, B2 => 
                           n11839, ZN => n7556);
   U4192 : OAI22_X1 port map( A1 => n10791, A2 => n11836, B1 => n10260, B2 => 
                           n11840, ZN => n7555);
   U4193 : OAI22_X1 port map( A1 => n10784, A2 => n11836, B1 => n10228, B2 => 
                           n11840, ZN => n7554);
   U4194 : OAI22_X1 port map( A1 => n10777, A2 => n11836, B1 => n10194, B2 => 
                           n11840, ZN => n7553);
   U4195 : OAI22_X1 port map( A1 => n10770, A2 => n11836, B1 => n10162, B2 => 
                           n11840, ZN => n7552);
   U4196 : OAI22_X1 port map( A1 => n10763, A2 => n11836, B1 => n10130, B2 => 
                           n11841, ZN => n7551);
   U4197 : OAI22_X1 port map( A1 => n10756, A2 => n11836, B1 => n10098, B2 => 
                           n11841, ZN => n7550);
   U4198 : OAI22_X1 port map( A1 => n10749, A2 => n11836, B1 => n10066, B2 => 
                           n11841, ZN => n7549);
   U4199 : OAI22_X1 port map( A1 => n10742, A2 => n11836, B1 => n10034, B2 => 
                           n11841, ZN => n7548);
   U4200 : OAI22_X1 port map( A1 => n10735, A2 => n11836, B1 => n10002, B2 => 
                           n11842, ZN => n7547);
   U4201 : OAI22_X1 port map( A1 => n10728, A2 => n11836, B1 => n9640, B2 => 
                           n11842, ZN => n7546);
   U4202 : OAI22_X1 port map( A1 => n10721, A2 => n11836, B1 => n9608, B2 => 
                           n11842, ZN => n7545);
   U4203 : OAI22_X1 port map( A1 => n10714, A2 => n11836, B1 => n9576, B2 => 
                           n11842, ZN => n7544);
   U4204 : OAI22_X1 port map( A1 => n10707, A2 => n11835, B1 => n9210, B2 => 
                           n11843, ZN => n7543);
   U4205 : OAI22_X1 port map( A1 => n10700, A2 => n11835, B1 => n9178, B2 => 
                           n11843, ZN => n7542);
   U4206 : OAI22_X1 port map( A1 => n10693, A2 => n11835, B1 => n9146, B2 => 
                           n11843, ZN => n7541);
   U4207 : OAI22_X1 port map( A1 => n10686, A2 => n11835, B1 => n6011, B2 => 
                           n11843, ZN => n7540);
   U4208 : OAI22_X1 port map( A1 => n10679, A2 => n11835, B1 => n5947, B2 => 
                           n11844, ZN => n7539);
   U4209 : OAI22_X1 port map( A1 => n10672, A2 => n11835, B1 => n5915, B2 => 
                           n11844, ZN => n7538);
   U4210 : OAI22_X1 port map( A1 => n10665, A2 => n11835, B1 => n5883, B2 => 
                           n11844, ZN => n7537);
   U4211 : OAI22_X1 port map( A1 => n10658, A2 => n11835, B1 => n5851, B2 => 
                           n11844, ZN => n7536);
   U4212 : OAI22_X1 port map( A1 => n10651, A2 => n11835, B1 => n5819, B2 => 
                           n11845, ZN => n7535);
   U4213 : OAI22_X1 port map( A1 => n10644, A2 => n11835, B1 => n5787, B2 => 
                           n11845, ZN => n7534);
   U4214 : OAI22_X1 port map( A1 => n10637, A2 => n11835, B1 => n5755, B2 => 
                           n11845, ZN => n7533);
   U4215 : OAI22_X1 port map( A1 => n10630, A2 => n11835, B1 => n5723, B2 => 
                           n11845, ZN => n7532);
   U4216 : OAI22_X1 port map( A1 => n10848, A2 => n11801, B1 => n10525, B2 => 
                           n11802, ZN => n7467);
   U4217 : OAI22_X1 port map( A1 => n10841, A2 => n11801, B1 => n10493, B2 => 
                           n11802, ZN => n7466);
   U4218 : OAI22_X1 port map( A1 => n10834, A2 => n11801, B1 => n10461, B2 => 
                           n11802, ZN => n7465);
   U4219 : OAI22_X1 port map( A1 => n10827, A2 => n11801, B1 => n10429, B2 => 
                           n11802, ZN => n7464);
   U4220 : OAI22_X1 port map( A1 => n10820, A2 => n11801, B1 => n10394, B2 => 
                           n11803, ZN => n7463);
   U4221 : OAI22_X1 port map( A1 => n10813, A2 => n11801, B1 => n10362, B2 => 
                           n11803, ZN => n7462);
   U4222 : OAI22_X1 port map( A1 => n10806, A2 => n11801, B1 => n10330, B2 => 
                           n11803, ZN => n7461);
   U4223 : OAI22_X1 port map( A1 => n10799, A2 => n11801, B1 => n10295, B2 => 
                           n11803, ZN => n7460);
   U4224 : OAI22_X1 port map( A1 => n10792, A2 => n11800, B1 => n10263, B2 => 
                           n11804, ZN => n7459);
   U4225 : OAI22_X1 port map( A1 => n10785, A2 => n11800, B1 => n10231, B2 => 
                           n11804, ZN => n7458);
   U4226 : OAI22_X1 port map( A1 => n10778, A2 => n11800, B1 => n10197, B2 => 
                           n11804, ZN => n7457);
   U4227 : OAI22_X1 port map( A1 => n10771, A2 => n11800, B1 => n10165, B2 => 
                           n11804, ZN => n7456);
   U4228 : OAI22_X1 port map( A1 => n10764, A2 => n11800, B1 => n10133, B2 => 
                           n11805, ZN => n7455);
   U4229 : OAI22_X1 port map( A1 => n10757, A2 => n11800, B1 => n10101, B2 => 
                           n11805, ZN => n7454);
   U4230 : OAI22_X1 port map( A1 => n10750, A2 => n11800, B1 => n10069, B2 => 
                           n11805, ZN => n7453);
   U4231 : OAI22_X1 port map( A1 => n10743, A2 => n11800, B1 => n10037, B2 => 
                           n11805, ZN => n7452);
   U4232 : OAI22_X1 port map( A1 => n10736, A2 => n11800, B1 => n10005, B2 => 
                           n11806, ZN => n7451);
   U4233 : OAI22_X1 port map( A1 => n10729, A2 => n11800, B1 => n9643, B2 => 
                           n11806, ZN => n7450);
   U4234 : OAI22_X1 port map( A1 => n10722, A2 => n11800, B1 => n9611, B2 => 
                           n11806, ZN => n7449);
   U4235 : OAI22_X1 port map( A1 => n10715, A2 => n11800, B1 => n9579, B2 => 
                           n11806, ZN => n7448);
   U4236 : OAI22_X1 port map( A1 => n10708, A2 => n11799, B1 => n9213, B2 => 
                           n11807, ZN => n7447);
   U4237 : OAI22_X1 port map( A1 => n10701, A2 => n11799, B1 => n9181, B2 => 
                           n11807, ZN => n7446);
   U4238 : OAI22_X1 port map( A1 => n10694, A2 => n11799, B1 => n9149, B2 => 
                           n11807, ZN => n7445);
   U4239 : OAI22_X1 port map( A1 => n10687, A2 => n11799, B1 => n6140, B2 => 
                           n11807, ZN => n7444);
   U4240 : OAI22_X1 port map( A1 => n10680, A2 => n11799, B1 => n5982, B2 => 
                           n11808, ZN => n7443);
   U4241 : OAI22_X1 port map( A1 => n10673, A2 => n11799, B1 => n5918, B2 => 
                           n11808, ZN => n7442);
   U4242 : OAI22_X1 port map( A1 => n10666, A2 => n11799, B1 => n5886, B2 => 
                           n11808, ZN => n7441);
   U4243 : OAI22_X1 port map( A1 => n10659, A2 => n11799, B1 => n5854, B2 => 
                           n11808, ZN => n7440);
   U4244 : OAI22_X1 port map( A1 => n10652, A2 => n11799, B1 => n5822, B2 => 
                           n11809, ZN => n7439);
   U4245 : OAI22_X1 port map( A1 => n10645, A2 => n11799, B1 => n5790, B2 => 
                           n11809, ZN => n7438);
   U4246 : OAI22_X1 port map( A1 => n10638, A2 => n11799, B1 => n5758, B2 => 
                           n11809, ZN => n7437);
   U4247 : OAI22_X1 port map( A1 => n10631, A2 => n11799, B1 => n5726, B2 => 
                           n11809, ZN => n7436);
   U4248 : OAI22_X1 port map( A1 => n10849, A2 => n11537, B1 => n10533, B2 => 
                           n11538, ZN => n6763);
   U4249 : OAI22_X1 port map( A1 => n10842, A2 => n11537, B1 => n10501, B2 => 
                           n11538, ZN => n6762);
   U4250 : OAI22_X1 port map( A1 => n10835, A2 => n11537, B1 => n10469, B2 => 
                           n11538, ZN => n6761);
   U4251 : OAI22_X1 port map( A1 => n10828, A2 => n11537, B1 => n10437, B2 => 
                           n11538, ZN => n6760);
   U4252 : OAI22_X1 port map( A1 => n10821, A2 => n11537, B1 => n10405, B2 => 
                           n11539, ZN => n6759);
   U4253 : OAI22_X1 port map( A1 => n10814, A2 => n11537, B1 => n10370, B2 => 
                           n11539, ZN => n6758);
   U4254 : OAI22_X1 port map( A1 => n10807, A2 => n11537, B1 => n10338, B2 => 
                           n11539, ZN => n6757);
   U4255 : OAI22_X1 port map( A1 => n10800, A2 => n11537, B1 => n10306, B2 => 
                           n11539, ZN => n6756);
   U4256 : OAI22_X1 port map( A1 => n10793, A2 => n11536, B1 => n10271, B2 => 
                           n11540, ZN => n6755);
   U4257 : OAI22_X1 port map( A1 => n10786, A2 => n11536, B1 => n10239, B2 => 
                           n11540, ZN => n6754);
   U4258 : OAI22_X1 port map( A1 => n10779, A2 => n11536, B1 => n10205, B2 => 
                           n11540, ZN => n6753);
   U4259 : OAI22_X1 port map( A1 => n10772, A2 => n11536, B1 => n10173, B2 => 
                           n11540, ZN => n6752);
   U4260 : OAI22_X1 port map( A1 => n10765, A2 => n11536, B1 => n10141, B2 => 
                           n11541, ZN => n6751);
   U4261 : OAI22_X1 port map( A1 => n10758, A2 => n11536, B1 => n10109, B2 => 
                           n11541, ZN => n6750);
   U4262 : OAI22_X1 port map( A1 => n10751, A2 => n11536, B1 => n10077, B2 => 
                           n11541, ZN => n6749);
   U4263 : OAI22_X1 port map( A1 => n10744, A2 => n11536, B1 => n10045, B2 => 
                           n11541, ZN => n6748);
   U4264 : OAI22_X1 port map( A1 => n10737, A2 => n11536, B1 => n10013, B2 => 
                           n11542, ZN => n6747);
   U4265 : OAI22_X1 port map( A1 => n10730, A2 => n11536, B1 => n9651, B2 => 
                           n11542, ZN => n6746);
   U4266 : OAI22_X1 port map( A1 => n10723, A2 => n11536, B1 => n9619, B2 => 
                           n11542, ZN => n6745);
   U4267 : OAI22_X1 port map( A1 => n10716, A2 => n11536, B1 => n9587, B2 => 
                           n11542, ZN => n6744);
   U4268 : OAI22_X1 port map( A1 => n10709, A2 => n11535, B1 => n9253, B2 => 
                           n11543, ZN => n6743);
   U4269 : OAI22_X1 port map( A1 => n10702, A2 => n11535, B1 => n9189, B2 => 
                           n11543, ZN => n6742);
   U4270 : OAI22_X1 port map( A1 => n10695, A2 => n11535, B1 => n9157, B2 => 
                           n11543, ZN => n6741);
   U4271 : OAI22_X1 port map( A1 => n10688, A2 => n11535, B1 => n6307, B2 => 
                           n11543, ZN => n6740);
   U4272 : OAI22_X1 port map( A1 => n10681, A2 => n11535, B1 => n5990, B2 => 
                           n11544, ZN => n6739);
   U4273 : OAI22_X1 port map( A1 => n10674, A2 => n11535, B1 => n5926, B2 => 
                           n11544, ZN => n6738);
   U4274 : OAI22_X1 port map( A1 => n10667, A2 => n11535, B1 => n5894, B2 => 
                           n11544, ZN => n6737);
   U4275 : OAI22_X1 port map( A1 => n10660, A2 => n11535, B1 => n5862, B2 => 
                           n11544, ZN => n6736);
   U4276 : OAI22_X1 port map( A1 => n10653, A2 => n11535, B1 => n5830, B2 => 
                           n11545, ZN => n6735);
   U4277 : OAI22_X1 port map( A1 => n10646, A2 => n11535, B1 => n5798, B2 => 
                           n11545, ZN => n6734);
   U4278 : OAI22_X1 port map( A1 => n10639, A2 => n11535, B1 => n5766, B2 => 
                           n11545, ZN => n6733);
   U4279 : OAI22_X1 port map( A1 => n10632, A2 => n11535, B1 => n5734, B2 => 
                           n11545, ZN => n6732);
   U4280 : OAI22_X1 port map( A1 => n10849, A2 => n11501, B1 => n1859, B2 => 
                           n11502, ZN => n6667);
   U4281 : OAI22_X1 port map( A1 => n10842, A2 => n11501, B1 => n1855, B2 => 
                           n11502, ZN => n6666);
   U4282 : OAI22_X1 port map( A1 => n10835, A2 => n11501, B1 => n1851, B2 => 
                           n11502, ZN => n6665);
   U4283 : OAI22_X1 port map( A1 => n10828, A2 => n11501, B1 => n1847, B2 => 
                           n11502, ZN => n6664);
   U4284 : OAI22_X1 port map( A1 => n10821, A2 => n11501, B1 => n1843, B2 => 
                           n11503, ZN => n6663);
   U4285 : OAI22_X1 port map( A1 => n10814, A2 => n11501, B1 => n1839, B2 => 
                           n11503, ZN => n6662);
   U4286 : OAI22_X1 port map( A1 => n10807, A2 => n11501, B1 => n1835, B2 => 
                           n11503, ZN => n6661);
   U4287 : OAI22_X1 port map( A1 => n10800, A2 => n11501, B1 => n1831, B2 => 
                           n11503, ZN => n6660);
   U4288 : OAI22_X1 port map( A1 => n10793, A2 => n11500, B1 => n1827, B2 => 
                           n11504, ZN => n6659);
   U4289 : OAI22_X1 port map( A1 => n10786, A2 => n11500, B1 => n1823, B2 => 
                           n11504, ZN => n6658);
   U4290 : OAI22_X1 port map( A1 => n10779, A2 => n11500, B1 => n1819, B2 => 
                           n11504, ZN => n6657);
   U4291 : OAI22_X1 port map( A1 => n10772, A2 => n11500, B1 => n1815, B2 => 
                           n11504, ZN => n6656);
   U4292 : OAI22_X1 port map( A1 => n10765, A2 => n11500, B1 => n1811, B2 => 
                           n11505, ZN => n6655);
   U4293 : OAI22_X1 port map( A1 => n10758, A2 => n11500, B1 => n1807, B2 => 
                           n11505, ZN => n6654);
   U4294 : OAI22_X1 port map( A1 => n10751, A2 => n11500, B1 => n1803, B2 => 
                           n11505, ZN => n6653);
   U4295 : OAI22_X1 port map( A1 => n10744, A2 => n11500, B1 => n1799, B2 => 
                           n11505, ZN => n6652);
   U4296 : OAI22_X1 port map( A1 => n10737, A2 => n11500, B1 => n1795, B2 => 
                           n11506, ZN => n6651);
   U4297 : OAI22_X1 port map( A1 => n10730, A2 => n11500, B1 => n1791, B2 => 
                           n11506, ZN => n6650);
   U4298 : OAI22_X1 port map( A1 => n10723, A2 => n11500, B1 => n1787, B2 => 
                           n11506, ZN => n6649);
   U4299 : OAI22_X1 port map( A1 => n10716, A2 => n11500, B1 => n1783, B2 => 
                           n11506, ZN => n6648);
   U4300 : OAI22_X1 port map( A1 => n10709, A2 => n11499, B1 => n1779, B2 => 
                           n11507, ZN => n6647);
   U4301 : OAI22_X1 port map( A1 => n10702, A2 => n11499, B1 => n1775, B2 => 
                           n11507, ZN => n6646);
   U4302 : OAI22_X1 port map( A1 => n10695, A2 => n11499, B1 => n1771, B2 => 
                           n11507, ZN => n6645);
   U4303 : OAI22_X1 port map( A1 => n10688, A2 => n11499, B1 => n1767, B2 => 
                           n11507, ZN => n6644);
   U4304 : OAI22_X1 port map( A1 => n10681, A2 => n11499, B1 => n1763, B2 => 
                           n11508, ZN => n6643);
   U4305 : OAI22_X1 port map( A1 => n10674, A2 => n11499, B1 => n1759, B2 => 
                           n11508, ZN => n6642);
   U4306 : OAI22_X1 port map( A1 => n10667, A2 => n11499, B1 => n1755, B2 => 
                           n11508, ZN => n6641);
   U4307 : OAI22_X1 port map( A1 => n10660, A2 => n11499, B1 => n1751, B2 => 
                           n11508, ZN => n6640);
   U4308 : OAI22_X1 port map( A1 => n10653, A2 => n11499, B1 => n1747, B2 => 
                           n11509, ZN => n6639);
   U4309 : OAI22_X1 port map( A1 => n10646, A2 => n11499, B1 => n1743, B2 => 
                           n11509, ZN => n6638);
   U4310 : OAI22_X1 port map( A1 => n10639, A2 => n11499, B1 => n1739, B2 => 
                           n11509, ZN => n6637);
   U4311 : OAI22_X1 port map( A1 => n10632, A2 => n11499, B1 => n1735, B2 => 
                           n11509, ZN => n6636);
   U4312 : OAI22_X1 port map( A1 => n10850, A2 => n11465, B1 => n513, B2 => 
                           n11466, ZN => n6571);
   U4313 : OAI22_X1 port map( A1 => n10843, A2 => n11465, B1 => n501, B2 => 
                           n11466, ZN => n6570);
   U4314 : OAI22_X1 port map( A1 => n10836, A2 => n11465, B1 => n489, B2 => 
                           n11466, ZN => n6569);
   U4315 : OAI22_X1 port map( A1 => n10829, A2 => n11465, B1 => n477, B2 => 
                           n11466, ZN => n6568);
   U4316 : OAI22_X1 port map( A1 => n10822, A2 => n11465, B1 => n465, B2 => 
                           n11467, ZN => n6567);
   U4317 : OAI22_X1 port map( A1 => n10815, A2 => n11465, B1 => n453, B2 => 
                           n11467, ZN => n6566);
   U4318 : OAI22_X1 port map( A1 => n10808, A2 => n11465, B1 => n441, B2 => 
                           n11467, ZN => n6565);
   U4319 : OAI22_X1 port map( A1 => n10801, A2 => n11465, B1 => n429, B2 => 
                           n11467, ZN => n6564);
   U4320 : OAI22_X1 port map( A1 => n10794, A2 => n11464, B1 => n417, B2 => 
                           n11468, ZN => n6563);
   U4321 : OAI22_X1 port map( A1 => n10787, A2 => n11464, B1 => n405, B2 => 
                           n11468, ZN => n6562);
   U4322 : OAI22_X1 port map( A1 => n10780, A2 => n11464, B1 => n393, B2 => 
                           n11468, ZN => n6561);
   U4323 : OAI22_X1 port map( A1 => n10773, A2 => n11464, B1 => n381, B2 => 
                           n11468, ZN => n6560);
   U4324 : OAI22_X1 port map( A1 => n10766, A2 => n11464, B1 => n369, B2 => 
                           n11469, ZN => n6559);
   U4325 : OAI22_X1 port map( A1 => n10759, A2 => n11464, B1 => n357, B2 => 
                           n11469, ZN => n6558);
   U4326 : OAI22_X1 port map( A1 => n10752, A2 => n11464, B1 => n345, B2 => 
                           n11469, ZN => n6557);
   U4327 : OAI22_X1 port map( A1 => n10745, A2 => n11464, B1 => n333, B2 => 
                           n11469, ZN => n6556);
   U4328 : OAI22_X1 port map( A1 => n10738, A2 => n11464, B1 => n321, B2 => 
                           n11470, ZN => n6555);
   U4329 : OAI22_X1 port map( A1 => n10731, A2 => n11464, B1 => n309, B2 => 
                           n11470, ZN => n6554);
   U4330 : OAI22_X1 port map( A1 => n10724, A2 => n11464, B1 => n297, B2 => 
                           n11470, ZN => n6553);
   U4331 : OAI22_X1 port map( A1 => n10717, A2 => n11464, B1 => n285, B2 => 
                           n11470, ZN => n6552);
   U4332 : OAI22_X1 port map( A1 => n10710, A2 => n11463, B1 => n273, B2 => 
                           n11471, ZN => n6551);
   U4333 : OAI22_X1 port map( A1 => n10703, A2 => n11463, B1 => n261, B2 => 
                           n11471, ZN => n6550);
   U4334 : OAI22_X1 port map( A1 => n10696, A2 => n11463, B1 => n249, B2 => 
                           n11471, ZN => n6549);
   U4335 : OAI22_X1 port map( A1 => n10689, A2 => n11463, B1 => n237, B2 => 
                           n11471, ZN => n6548);
   U4336 : OAI22_X1 port map( A1 => n10682, A2 => n11463, B1 => n225, B2 => 
                           n11472, ZN => n6547);
   U4337 : OAI22_X1 port map( A1 => n10675, A2 => n11463, B1 => n213, B2 => 
                           n11472, ZN => n6546);
   U4338 : OAI22_X1 port map( A1 => n10668, A2 => n11463, B1 => n201, B2 => 
                           n11472, ZN => n6545);
   U4339 : OAI22_X1 port map( A1 => n10661, A2 => n11463, B1 => n189, B2 => 
                           n11472, ZN => n6544);
   U4340 : OAI22_X1 port map( A1 => n10654, A2 => n11463, B1 => n177, B2 => 
                           n11473, ZN => n6543);
   U4341 : OAI22_X1 port map( A1 => n10647, A2 => n11463, B1 => n165, B2 => 
                           n11473, ZN => n6542);
   U4342 : OAI22_X1 port map( A1 => n10640, A2 => n11463, B1 => n153, B2 => 
                           n11473, ZN => n6541);
   U4343 : OAI22_X1 port map( A1 => n10633, A2 => n11463, B1 => n141, B2 => 
                           n11473, ZN => n6540);
   U4344 : OAI22_X1 port map( A1 => n10850, A2 => n11429, B1 => n514, B2 => 
                           n11430, ZN => n6475);
   U4345 : OAI22_X1 port map( A1 => n10843, A2 => n11429, B1 => n502, B2 => 
                           n11430, ZN => n6474);
   U4346 : OAI22_X1 port map( A1 => n10836, A2 => n11429, B1 => n490, B2 => 
                           n11430, ZN => n6473);
   U4347 : OAI22_X1 port map( A1 => n10829, A2 => n11429, B1 => n478, B2 => 
                           n11430, ZN => n6472);
   U4348 : OAI22_X1 port map( A1 => n10822, A2 => n11429, B1 => n466, B2 => 
                           n11431, ZN => n6471);
   U4349 : OAI22_X1 port map( A1 => n10815, A2 => n11429, B1 => n454, B2 => 
                           n11431, ZN => n6470);
   U4350 : OAI22_X1 port map( A1 => n10808, A2 => n11429, B1 => n442, B2 => 
                           n11431, ZN => n6469);
   U4351 : OAI22_X1 port map( A1 => n10801, A2 => n11429, B1 => n430, B2 => 
                           n11431, ZN => n6468);
   U4352 : OAI22_X1 port map( A1 => n10794, A2 => n11428, B1 => n418, B2 => 
                           n11432, ZN => n6467);
   U4353 : OAI22_X1 port map( A1 => n10787, A2 => n11428, B1 => n406, B2 => 
                           n11432, ZN => n6466);
   U4354 : OAI22_X1 port map( A1 => n10780, A2 => n11428, B1 => n394, B2 => 
                           n11432, ZN => n6465);
   U4355 : OAI22_X1 port map( A1 => n10773, A2 => n11428, B1 => n382, B2 => 
                           n11432, ZN => n6464);
   U4356 : OAI22_X1 port map( A1 => n10766, A2 => n11428, B1 => n370, B2 => 
                           n11433, ZN => n6463);
   U4357 : OAI22_X1 port map( A1 => n10759, A2 => n11428, B1 => n358, B2 => 
                           n11433, ZN => n6462);
   U4358 : OAI22_X1 port map( A1 => n10752, A2 => n11428, B1 => n346, B2 => 
                           n11433, ZN => n6461);
   U4360 : OAI22_X1 port map( A1 => n10745, A2 => n11428, B1 => n334, B2 => 
                           n11433, ZN => n6460);
   U4361 : OAI22_X1 port map( A1 => n10738, A2 => n11428, B1 => n322, B2 => 
                           n11434, ZN => n6459);
   U4362 : OAI22_X1 port map( A1 => n10731, A2 => n11428, B1 => n310, B2 => 
                           n11434, ZN => n6458);
   U4363 : OAI22_X1 port map( A1 => n10724, A2 => n11428, B1 => n298, B2 => 
                           n11434, ZN => n6457);
   U4364 : OAI22_X1 port map( A1 => n10717, A2 => n11428, B1 => n286, B2 => 
                           n11434, ZN => n6456);
   U4365 : OAI22_X1 port map( A1 => n10710, A2 => n11427, B1 => n274, B2 => 
                           n11435, ZN => n6455);
   U4366 : OAI22_X1 port map( A1 => n10703, A2 => n11427, B1 => n262, B2 => 
                           n11435, ZN => n6454);
   U4367 : OAI22_X1 port map( A1 => n10696, A2 => n11427, B1 => n250, B2 => 
                           n11435, ZN => n6453);
   U4368 : OAI22_X1 port map( A1 => n10689, A2 => n11427, B1 => n238, B2 => 
                           n11435, ZN => n6452);
   U4369 : OAI22_X1 port map( A1 => n10682, A2 => n11427, B1 => n226, B2 => 
                           n11436, ZN => n6451);
   U4370 : OAI22_X1 port map( A1 => n10675, A2 => n11427, B1 => n214, B2 => 
                           n11436, ZN => n6450);
   U4371 : OAI22_X1 port map( A1 => n10668, A2 => n11427, B1 => n202, B2 => 
                           n11436, ZN => n6449);
   U4372 : OAI22_X1 port map( A1 => n10661, A2 => n11427, B1 => n190, B2 => 
                           n11436, ZN => n6448);
   U4373 : OAI22_X1 port map( A1 => n10654, A2 => n11427, B1 => n178, B2 => 
                           n11437, ZN => n6447);
   U4374 : OAI22_X1 port map( A1 => n10647, A2 => n11427, B1 => n166, B2 => 
                           n11437, ZN => n6446);
   U4375 : OAI22_X1 port map( A1 => n10640, A2 => n11427, B1 => n154, B2 => 
                           n11437, ZN => n6445);
   U4376 : OAI22_X1 port map( A1 => n10633, A2 => n11427, B1 => n142, B2 => 
                           n11437, ZN => n6444);
   U4377 : OAI22_X1 port map( A1 => n10844, A2 => n12340, B1 => n10510, B2 => 
                           n12341, ZN => n8907);
   U4378 : OAI22_X1 port map( A1 => n10837, A2 => n12339, B1 => n10478, B2 => 
                           n12341, ZN => n8906);
   U4379 : OAI22_X1 port map( A1 => n10830, A2 => n12340, B1 => n10446, B2 => 
                           n12341, ZN => n8905);
   U4380 : OAI22_X1 port map( A1 => n10823, A2 => n12339, B1 => n10414, B2 => 
                           n12341, ZN => n8904);
   U4381 : OAI22_X1 port map( A1 => n10816, A2 => n12340, B1 => n10379, B2 => 
                           n12342, ZN => n8903);
   U4382 : OAI22_X1 port map( A1 => n10809, A2 => n12339, B1 => n10347, B2 => 
                           n12342, ZN => n8902);
   U4383 : OAI22_X1 port map( A1 => n10802, A2 => n12340, B1 => n10315, B2 => 
                           n12342, ZN => n8901);
   U4384 : OAI22_X1 port map( A1 => n10795, A2 => n12339, B1 => n10280, B2 => 
                           n12342, ZN => n8900);
   U4385 : OAI22_X1 port map( A1 => n10788, A2 => n12340, B1 => n10248, B2 => 
                           n12343, ZN => n8899);
   U4386 : OAI22_X1 port map( A1 => n10781, A2 => n12340, B1 => n10216, B2 => 
                           n12343, ZN => n8898);
   U4387 : OAI22_X1 port map( A1 => n10774, A2 => n12340, B1 => n10182, B2 => 
                           n12343, ZN => n8897);
   U4388 : OAI22_X1 port map( A1 => n10767, A2 => n12340, B1 => n10150, B2 => 
                           n12343, ZN => n8896);
   U4389 : OAI22_X1 port map( A1 => n10760, A2 => n12340, B1 => n10118, B2 => 
                           n12344, ZN => n8895);
   U4390 : OAI22_X1 port map( A1 => n10753, A2 => n12340, B1 => n10086, B2 => 
                           n12344, ZN => n8894);
   U4391 : OAI22_X1 port map( A1 => n10746, A2 => n12340, B1 => n10054, B2 => 
                           n12344, ZN => n8893);
   U4392 : OAI22_X1 port map( A1 => n10739, A2 => n12340, B1 => n10022, B2 => 
                           n12344, ZN => n8892);
   U4393 : OAI22_X1 port map( A1 => n10732, A2 => n12340, B1 => n9660, B2 => 
                           n12345, ZN => n8891);
   U4394 : OAI22_X1 port map( A1 => n10725, A2 => n12340, B1 => n9628, B2 => 
                           n12345, ZN => n8890);
   U4395 : OAI22_X1 port map( A1 => n10718, A2 => n12340, B1 => n9596, B2 => 
                           n12345, ZN => n8889);
   U4396 : OAI22_X1 port map( A1 => n10711, A2 => n12340, B1 => n9262, B2 => 
                           n12345, ZN => n8888);
   U4397 : OAI22_X1 port map( A1 => n10704, A2 => n12339, B1 => n9198, B2 => 
                           n12346, ZN => n8887);
   U4398 : OAI22_X1 port map( A1 => n10697, A2 => n12339, B1 => n9166, B2 => 
                           n12346, ZN => n8886);
   U4399 : OAI22_X1 port map( A1 => n10690, A2 => n12339, B1 => n9134, B2 => 
                           n12346, ZN => n8885);
   U4400 : OAI22_X1 port map( A1 => n10683, A2 => n12339, B1 => n5999, B2 => 
                           n12346, ZN => n8884);
   U4401 : OAI22_X1 port map( A1 => n10676, A2 => n12339, B1 => n5935, B2 => 
                           n12347, ZN => n8883);
   U4402 : OAI22_X1 port map( A1 => n10669, A2 => n12339, B1 => n5903, B2 => 
                           n12347, ZN => n8882);
   U4403 : OAI22_X1 port map( A1 => n10662, A2 => n12339, B1 => n5871, B2 => 
                           n12347, ZN => n8881);
   U4404 : OAI22_X1 port map( A1 => n10655, A2 => n12339, B1 => n5839, B2 => 
                           n12347, ZN => n8880);
   U4405 : OAI22_X1 port map( A1 => n10648, A2 => n12339, B1 => n5807, B2 => 
                           n12348, ZN => n8879);
   U4406 : OAI22_X1 port map( A1 => n10641, A2 => n12339, B1 => n5775, B2 => 
                           n12348, ZN => n8878);
   U4407 : OAI22_X1 port map( A1 => n10634, A2 => n12339, B1 => n5743, B2 => 
                           n12348, ZN => n8877);
   U4408 : OAI22_X1 port map( A1 => n10627, A2 => n12339, B1 => n5711, B2 => 
                           n12348, ZN => n8876);
   U4409 : OAI22_X1 port map( A1 => n10844, A2 => n12281, B1 => n992, B2 => 
                           n12282, ZN => n8747_port);
   U4410 : OAI22_X1 port map( A1 => n10837, A2 => n12281, B1 => n988, B2 => 
                           n12282, ZN => n8746_port);
   U4411 : OAI22_X1 port map( A1 => n10830, A2 => n12281, B1 => n984, B2 => 
                           n12282, ZN => n8745_port);
   U4412 : OAI22_X1 port map( A1 => n10823, A2 => n12281, B1 => n980, B2 => 
                           n12282, ZN => n8744_port);
   U4413 : OAI22_X1 port map( A1 => n10816, A2 => n12281, B1 => n976, B2 => 
                           n12283, ZN => n8743_port);
   U4414 : OAI22_X1 port map( A1 => n10809, A2 => n12281, B1 => n972, B2 => 
                           n12283, ZN => n8742_port);
   U4415 : OAI22_X1 port map( A1 => n10802, A2 => n12281, B1 => n968, B2 => 
                           n12283, ZN => n8741_port);
   U4416 : OAI22_X1 port map( A1 => n10795, A2 => n12281, B1 => n964, B2 => 
                           n12283, ZN => n8740_port);
   U4417 : OAI22_X1 port map( A1 => n10788, A2 => n12280, B1 => n960, B2 => 
                           n12284, ZN => n8739_port);
   U4418 : OAI22_X1 port map( A1 => n10781, A2 => n12280, B1 => n956, B2 => 
                           n12284, ZN => n8738_port);
   U4419 : OAI22_X1 port map( A1 => n10774, A2 => n12280, B1 => n952, B2 => 
                           n12284, ZN => n8737_port);
   U4420 : OAI22_X1 port map( A1 => n10767, A2 => n12280, B1 => n948, B2 => 
                           n12284, ZN => n8736_port);
   U4421 : OAI22_X1 port map( A1 => n10760, A2 => n12280, B1 => n944, B2 => 
                           n12285, ZN => n8735_port);
   U4422 : OAI22_X1 port map( A1 => n10753, A2 => n12280, B1 => n940, B2 => 
                           n12285, ZN => n8734_port);
   U4423 : OAI22_X1 port map( A1 => n10746, A2 => n12280, B1 => n936, B2 => 
                           n12285, ZN => n8733_port);
   U4424 : OAI22_X1 port map( A1 => n10739, A2 => n12280, B1 => n932, B2 => 
                           n12285, ZN => n8732_port);
   U4425 : OAI22_X1 port map( A1 => n10732, A2 => n12280, B1 => n928, B2 => 
                           n12286, ZN => n8731_port);
   U4426 : OAI22_X1 port map( A1 => n10725, A2 => n12280, B1 => n924, B2 => 
                           n12286, ZN => n8730_port);
   U4427 : OAI22_X1 port map( A1 => n10718, A2 => n12280, B1 => n920, B2 => 
                           n12286, ZN => n8729_port);
   U4428 : OAI22_X1 port map( A1 => n10711, A2 => n12280, B1 => n916, B2 => 
                           n12286, ZN => n8728_port);
   U4429 : OAI22_X1 port map( A1 => n10704, A2 => n12279, B1 => n912, B2 => 
                           n12287, ZN => n8727_port);
   U4430 : OAI22_X1 port map( A1 => n10697, A2 => n12279, B1 => n908, B2 => 
                           n12287, ZN => n8726_port);
   U4431 : OAI22_X1 port map( A1 => n10690, A2 => n12279, B1 => n904, B2 => 
                           n12287, ZN => n8725_port);
   U4432 : OAI22_X1 port map( A1 => n10683, A2 => n12279, B1 => n900, B2 => 
                           n12287, ZN => n8724_port);
   U4433 : OAI22_X1 port map( A1 => n10676, A2 => n12279, B1 => n896, B2 => 
                           n12288, ZN => n8723_port);
   U4434 : OAI22_X1 port map( A1 => n10669, A2 => n12279, B1 => n892, B2 => 
                           n12288, ZN => n8722_port);
   U4435 : OAI22_X1 port map( A1 => n10662, A2 => n12279, B1 => n888, B2 => 
                           n12288, ZN => n8721_port);
   U4436 : OAI22_X1 port map( A1 => n10655, A2 => n12279, B1 => n884, B2 => 
                           n12288, ZN => n8720_port);
   U4437 : OAI22_X1 port map( A1 => n10648, A2 => n12279, B1 => n880, B2 => 
                           n12289, ZN => n8719_port);
   U4438 : OAI22_X1 port map( A1 => n10641, A2 => n12279, B1 => n876, B2 => 
                           n12289, ZN => n8718_port);
   U4439 : OAI22_X1 port map( A1 => n10634, A2 => n12279, B1 => n872, B2 => 
                           n12289, ZN => n8717_port);
   U4440 : OAI22_X1 port map( A1 => n10627, A2 => n12279, B1 => n868, B2 => 
                           n12289, ZN => n8716_port);
   U4441 : OAI22_X1 port map( A1 => n10845, A2 => n12125, B1 => n10515, B2 => 
                           n12126, ZN => n8331);
   U4442 : OAI22_X1 port map( A1 => n10838, A2 => n12125, B1 => n10483, B2 => 
                           n12126, ZN => n8330);
   U4443 : OAI22_X1 port map( A1 => n10831, A2 => n12125, B1 => n10451, B2 => 
                           n12126, ZN => n8329);
   U4444 : OAI22_X1 port map( A1 => n10824, A2 => n12125, B1 => n10419, B2 => 
                           n12126, ZN => n8328);
   U4445 : OAI22_X1 port map( A1 => n10817, A2 => n12125, B1 => n10384, B2 => 
                           n12127, ZN => n8327);
   U4446 : OAI22_X1 port map( A1 => n10810, A2 => n12125, B1 => n10352, B2 => 
                           n12127, ZN => n8326);
   U4447 : OAI22_X1 port map( A1 => n10803, A2 => n12125, B1 => n10320, B2 => 
                           n12127, ZN => n8325);
   U4448 : OAI22_X1 port map( A1 => n10796, A2 => n12125, B1 => n10285, B2 => 
                           n12127, ZN => n8324);
   U4449 : OAI22_X1 port map( A1 => n10789, A2 => n12124, B1 => n10253, B2 => 
                           n12128, ZN => n8323);
   U4450 : OAI22_X1 port map( A1 => n10782, A2 => n12124, B1 => n10221, B2 => 
                           n12128, ZN => n8322);
   U4451 : OAI22_X1 port map( A1 => n10775, A2 => n12124, B1 => n10187, B2 => 
                           n12128, ZN => n8321);
   U4452 : OAI22_X1 port map( A1 => n10768, A2 => n12124, B1 => n10155, B2 => 
                           n12128, ZN => n8320);
   U4453 : OAI22_X1 port map( A1 => n10761, A2 => n12124, B1 => n10123, B2 => 
                           n12129, ZN => n8319);
   U4454 : OAI22_X1 port map( A1 => n10754, A2 => n12124, B1 => n10091, B2 => 
                           n12129, ZN => n8318);
   U4455 : OAI22_X1 port map( A1 => n10747, A2 => n12124, B1 => n10059, B2 => 
                           n12129, ZN => n8317);
   U4456 : OAI22_X1 port map( A1 => n10740, A2 => n12124, B1 => n10027, B2 => 
                           n12129, ZN => n8316);
   U4457 : OAI22_X1 port map( A1 => n10733, A2 => n12124, B1 => n9697, B2 => 
                           n12130, ZN => n8315);
   U4458 : OAI22_X1 port map( A1 => n10726, A2 => n12124, B1 => n9633, B2 => 
                           n12130, ZN => n8314);
   U4459 : OAI22_X1 port map( A1 => n10719, A2 => n12124, B1 => n9601, B2 => 
                           n12130, ZN => n8313);
   U4460 : OAI22_X1 port map( A1 => n10712, A2 => n12124, B1 => n9569, B2 => 
                           n12130, ZN => n8312);
   U4461 : OAI22_X1 port map( A1 => n10705, A2 => n12123, B1 => n9203, B2 => 
                           n12131, ZN => n8311);
   U4462 : OAI22_X1 port map( A1 => n10698, A2 => n12123, B1 => n9171, B2 => 
                           n12131, ZN => n8310);
   U4463 : OAI22_X1 port map( A1 => n10691, A2 => n12123, B1 => n9139, B2 => 
                           n12131, ZN => n8309);
   U4464 : OAI22_X1 port map( A1 => n10684, A2 => n12123, B1 => n6004, B2 => 
                           n12131, ZN => n8308);
   U4465 : OAI22_X1 port map( A1 => n10677, A2 => n12123, B1 => n5940, B2 => 
                           n12132, ZN => n8307);
   U4466 : OAI22_X1 port map( A1 => n10670, A2 => n12123, B1 => n5908, B2 => 
                           n12132, ZN => n8306);
   U4467 : OAI22_X1 port map( A1 => n10663, A2 => n12123, B1 => n5876, B2 => 
                           n12132, ZN => n8305);
   U4468 : OAI22_X1 port map( A1 => n10656, A2 => n12123, B1 => n5844, B2 => 
                           n12132, ZN => n8304);
   U4469 : OAI22_X1 port map( A1 => n10649, A2 => n12123, B1 => n5812, B2 => 
                           n12133, ZN => n8303);
   U4470 : OAI22_X1 port map( A1 => n10642, A2 => n12123, B1 => n5780, B2 => 
                           n12133, ZN => n8302);
   U4471 : OAI22_X1 port map( A1 => n10635, A2 => n12123, B1 => n5748, B2 => 
                           n12133, ZN => n8301);
   U4472 : OAI22_X1 port map( A1 => n10628, A2 => n12123, B1 => n5716, B2 => 
                           n12133, ZN => n8300);
   U4473 : OAI22_X1 port map( A1 => n10846, A2 => n12077, B1 => n10518, B2 => 
                           n12078, ZN => n8203);
   U4474 : OAI22_X1 port map( A1 => n10839, A2 => n12077, B1 => n10486, B2 => 
                           n12078, ZN => n8202);
   U4475 : OAI22_X1 port map( A1 => n10832, A2 => n12077, B1 => n10454, B2 => 
                           n12078, ZN => n8201);
   U4476 : OAI22_X1 port map( A1 => n10825, A2 => n12077, B1 => n10422, B2 => 
                           n12078, ZN => n8200);
   U4477 : OAI22_X1 port map( A1 => n10818, A2 => n12077, B1 => n10387, B2 => 
                           n12079, ZN => n8199);
   U4478 : OAI22_X1 port map( A1 => n10811, A2 => n12077, B1 => n10355, B2 => 
                           n12079, ZN => n8198);
   U4479 : OAI22_X1 port map( A1 => n10804, A2 => n12077, B1 => n10323, B2 => 
                           n12079, ZN => n8197);
   U4480 : OAI22_X1 port map( A1 => n10797, A2 => n12077, B1 => n10288, B2 => 
                           n12079, ZN => n8196);
   U4481 : OAI22_X1 port map( A1 => n10790, A2 => n12076, B1 => n10256, B2 => 
                           n12080, ZN => n8195);
   U4482 : OAI22_X1 port map( A1 => n10783, A2 => n12076, B1 => n10224, B2 => 
                           n12080, ZN => n8194);
   U4483 : OAI22_X1 port map( A1 => n10776, A2 => n12076, B1 => n10190, B2 => 
                           n12080, ZN => n8193);
   U4484 : OAI22_X1 port map( A1 => n10769, A2 => n12076, B1 => n10158, B2 => 
                           n12080, ZN => n8192);
   U4485 : OAI22_X1 port map( A1 => n10762, A2 => n12076, B1 => n10126, B2 => 
                           n12081, ZN => n8191);
   U4486 : OAI22_X1 port map( A1 => n10755, A2 => n12076, B1 => n10094, B2 => 
                           n12081, ZN => n8190);
   U4487 : OAI22_X1 port map( A1 => n10748, A2 => n12076, B1 => n10062, B2 => 
                           n12081, ZN => n8189);
   U4488 : OAI22_X1 port map( A1 => n10741, A2 => n12076, B1 => n10030, B2 => 
                           n12081, ZN => n8188);
   U4489 : OAI22_X1 port map( A1 => n10734, A2 => n12076, B1 => n9700, B2 => 
                           n12082, ZN => n8187);
   U4490 : OAI22_X1 port map( A1 => n10727, A2 => n12076, B1 => n9636, B2 => 
                           n12082, ZN => n8186);
   U4491 : OAI22_X1 port map( A1 => n10720, A2 => n12076, B1 => n9604, B2 => 
                           n12082, ZN => n8185);
   U4492 : OAI22_X1 port map( A1 => n10713, A2 => n12076, B1 => n9572, B2 => 
                           n12082, ZN => n8184);
   U4493 : OAI22_X1 port map( A1 => n10706, A2 => n12075, B1 => n9206, B2 => 
                           n12083, ZN => n8183);
   U4494 : OAI22_X1 port map( A1 => n10699, A2 => n12075, B1 => n9174, B2 => 
                           n12083, ZN => n8182);
   U4495 : OAI22_X1 port map( A1 => n10692, A2 => n12075, B1 => n9142, B2 => 
                           n12083, ZN => n8181);
   U4496 : OAI22_X1 port map( A1 => n10685, A2 => n12075, B1 => n6007, B2 => 
                           n12083, ZN => n8180);
   U4497 : OAI22_X1 port map( A1 => n10678, A2 => n12075, B1 => n5943, B2 => 
                           n12084, ZN => n8179);
   U4498 : OAI22_X1 port map( A1 => n10671, A2 => n12075, B1 => n5911, B2 => 
                           n12084, ZN => n8178);
   U4499 : OAI22_X1 port map( A1 => n10664, A2 => n12075, B1 => n5879, B2 => 
                           n12084, ZN => n8177);
   U4500 : OAI22_X1 port map( A1 => n10657, A2 => n12075, B1 => n5847, B2 => 
                           n12084, ZN => n8176);
   U4501 : OAI22_X1 port map( A1 => n10650, A2 => n12075, B1 => n5815, B2 => 
                           n12085, ZN => n8175);
   U4502 : OAI22_X1 port map( A1 => n10643, A2 => n12075, B1 => n5783, B2 => 
                           n12085, ZN => n8174);
   U4503 : OAI22_X1 port map( A1 => n10636, A2 => n12075, B1 => n5751, B2 => 
                           n12085, ZN => n8173);
   U4504 : OAI22_X1 port map( A1 => n10629, A2 => n12075, B1 => n5719, B2 => 
                           n12085, ZN => n8172);
   U4505 : OAI22_X1 port map( A1 => n10847, A2 => n11861, B1 => n10523, B2 => 
                           n11862, ZN => n7627);
   U4506 : OAI22_X1 port map( A1 => n10840, A2 => n11861, B1 => n10491, B2 => 
                           n11862, ZN => n7626);
   U4507 : OAI22_X1 port map( A1 => n10833, A2 => n11861, B1 => n10459, B2 => 
                           n11862, ZN => n7625);
   U4508 : OAI22_X1 port map( A1 => n10826, A2 => n11861, B1 => n10427, B2 => 
                           n11862, ZN => n7624);
   U4509 : OAI22_X1 port map( A1 => n10819, A2 => n11861, B1 => n10392, B2 => 
                           n11863, ZN => n7623);
   U4510 : OAI22_X1 port map( A1 => n10812, A2 => n11861, B1 => n10360, B2 => 
                           n11863, ZN => n7622);
   U4511 : OAI22_X1 port map( A1 => n10805, A2 => n11861, B1 => n10328, B2 => 
                           n11863, ZN => n7621);
   U4512 : OAI22_X1 port map( A1 => n10798, A2 => n11861, B1 => n10293, B2 => 
                           n11863, ZN => n7620);
   U4513 : OAI22_X1 port map( A1 => n10791, A2 => n11860, B1 => n10261, B2 => 
                           n11864, ZN => n7619);
   U4514 : OAI22_X1 port map( A1 => n10784, A2 => n11860, B1 => n10229, B2 => 
                           n11864, ZN => n7618);
   U4515 : OAI22_X1 port map( A1 => n10777, A2 => n11860, B1 => n10195, B2 => 
                           n11864, ZN => n7617);
   U4516 : OAI22_X1 port map( A1 => n10770, A2 => n11860, B1 => n10163, B2 => 
                           n11864, ZN => n7616);
   U4517 : OAI22_X1 port map( A1 => n10763, A2 => n11860, B1 => n10131, B2 => 
                           n11865, ZN => n7615);
   U4518 : OAI22_X1 port map( A1 => n10756, A2 => n11860, B1 => n10099, B2 => 
                           n11865, ZN => n7614);
   U4519 : OAI22_X1 port map( A1 => n10749, A2 => n11860, B1 => n10067, B2 => 
                           n11865, ZN => n7613);
   U4520 : OAI22_X1 port map( A1 => n10742, A2 => n11860, B1 => n10035, B2 => 
                           n11865, ZN => n7612);
   U4521 : OAI22_X1 port map( A1 => n10735, A2 => n11860, B1 => n10003, B2 => 
                           n11866, ZN => n7611);
   U4522 : OAI22_X1 port map( A1 => n10728, A2 => n11860, B1 => n9641, B2 => 
                           n11866, ZN => n7610);
   U4523 : OAI22_X1 port map( A1 => n10721, A2 => n11860, B1 => n9609, B2 => 
                           n11866, ZN => n7609);
   U4524 : OAI22_X1 port map( A1 => n10714, A2 => n11860, B1 => n9577, B2 => 
                           n11866, ZN => n7608);
   U4525 : OAI22_X1 port map( A1 => n10707, A2 => n11859, B1 => n9211, B2 => 
                           n11867, ZN => n7607);
   U4526 : OAI22_X1 port map( A1 => n10700, A2 => n11859, B1 => n9179, B2 => 
                           n11867, ZN => n7606);
   U4527 : OAI22_X1 port map( A1 => n10693, A2 => n11859, B1 => n9147, B2 => 
                           n11867, ZN => n7605);
   U4528 : OAI22_X1 port map( A1 => n10686, A2 => n11859, B1 => n6012, B2 => 
                           n11867, ZN => n7604);
   U4529 : OAI22_X1 port map( A1 => n10679, A2 => n11859, B1 => n5948, B2 => 
                           n11868, ZN => n7603);
   U4530 : OAI22_X1 port map( A1 => n10672, A2 => n11859, B1 => n5916, B2 => 
                           n11868, ZN => n7602);
   U4531 : OAI22_X1 port map( A1 => n10665, A2 => n11859, B1 => n5884, B2 => 
                           n11868, ZN => n7601);
   U4532 : OAI22_X1 port map( A1 => n10658, A2 => n11859, B1 => n5852, B2 => 
                           n11868, ZN => n7600);
   U4533 : OAI22_X1 port map( A1 => n10651, A2 => n11859, B1 => n5820, B2 => 
                           n11869, ZN => n7599);
   U4534 : OAI22_X1 port map( A1 => n10644, A2 => n11859, B1 => n5788, B2 => 
                           n11869, ZN => n7598);
   U4535 : OAI22_X1 port map( A1 => n10637, A2 => n11859, B1 => n5756, B2 => 
                           n11869, ZN => n7597);
   U4536 : OAI22_X1 port map( A1 => n10630, A2 => n11859, B1 => n5724, B2 => 
                           n11869, ZN => n7596);
   U4537 : OAI22_X1 port map( A1 => n10847, A2 => n11813, B1 => n10526, B2 => 
                           n11814, ZN => n7499);
   U4538 : OAI22_X1 port map( A1 => n10840, A2 => n11813, B1 => n10494, B2 => 
                           n11814, ZN => n7498);
   U4539 : OAI22_X1 port map( A1 => n10833, A2 => n11813, B1 => n10462, B2 => 
                           n11814, ZN => n7497);
   U4540 : OAI22_X1 port map( A1 => n10826, A2 => n11813, B1 => n10430, B2 => 
                           n11814, ZN => n7496);
   U4541 : OAI22_X1 port map( A1 => n10819, A2 => n11813, B1 => n10395, B2 => 
                           n11815, ZN => n7495);
   U4542 : OAI22_X1 port map( A1 => n10812, A2 => n11813, B1 => n10363, B2 => 
                           n11815, ZN => n7494);
   U4543 : OAI22_X1 port map( A1 => n10805, A2 => n11813, B1 => n10331, B2 => 
                           n11815, ZN => n7493);
   U4544 : OAI22_X1 port map( A1 => n10798, A2 => n11813, B1 => n10296, B2 => 
                           n11815, ZN => n7492);
   U4545 : OAI22_X1 port map( A1 => n10791, A2 => n11812, B1 => n10264, B2 => 
                           n11816, ZN => n7491);
   U4546 : OAI22_X1 port map( A1 => n10784, A2 => n11812, B1 => n10232, B2 => 
                           n11816, ZN => n7490);
   U4547 : OAI22_X1 port map( A1 => n10777, A2 => n11812, B1 => n10198, B2 => 
                           n11816, ZN => n7489);
   U4548 : OAI22_X1 port map( A1 => n10770, A2 => n11812, B1 => n10166, B2 => 
                           n11816, ZN => n7488);
   U4549 : OAI22_X1 port map( A1 => n10763, A2 => n11812, B1 => n10134, B2 => 
                           n11817, ZN => n7487);
   U4550 : OAI22_X1 port map( A1 => n10756, A2 => n11812, B1 => n10102, B2 => 
                           n11817, ZN => n7486);
   U4551 : OAI22_X1 port map( A1 => n10749, A2 => n11812, B1 => n10070, B2 => 
                           n11817, ZN => n7485);
   U4552 : OAI22_X1 port map( A1 => n10742, A2 => n11812, B1 => n10038, B2 => 
                           n11817, ZN => n7484);
   U4553 : OAI22_X1 port map( A1 => n10735, A2 => n11812, B1 => n10006, B2 => 
                           n11818, ZN => n7483);
   U4554 : OAI22_X1 port map( A1 => n10728, A2 => n11812, B1 => n9644, B2 => 
                           n11818, ZN => n7482);
   U4555 : OAI22_X1 port map( A1 => n10721, A2 => n11812, B1 => n9612, B2 => 
                           n11818, ZN => n7481);
   U4556 : OAI22_X1 port map( A1 => n10714, A2 => n11812, B1 => n9580, B2 => 
                           n11818, ZN => n7480);
   U4557 : OAI22_X1 port map( A1 => n10707, A2 => n11811, B1 => n9214, B2 => 
                           n11819, ZN => n7479);
   U4558 : OAI22_X1 port map( A1 => n10700, A2 => n11811, B1 => n9182, B2 => 
                           n11819, ZN => n7478);
   U4559 : OAI22_X1 port map( A1 => n10693, A2 => n11811, B1 => n9150, B2 => 
                           n11819, ZN => n7477);
   U4560 : OAI22_X1 port map( A1 => n10686, A2 => n11811, B1 => n6236, B2 => 
                           n11819, ZN => n7476);
   U4561 : OAI22_X1 port map( A1 => n10679, A2 => n11811, B1 => n5983, B2 => 
                           n11820, ZN => n7475);
   U4562 : OAI22_X1 port map( A1 => n10672, A2 => n11811, B1 => n5919, B2 => 
                           n11820, ZN => n7474);
   U4563 : OAI22_X1 port map( A1 => n10665, A2 => n11811, B1 => n5887, B2 => 
                           n11820, ZN => n7473);
   U4564 : OAI22_X1 port map( A1 => n10658, A2 => n11811, B1 => n5855, B2 => 
                           n11820, ZN => n7472);
   U4565 : OAI22_X1 port map( A1 => n10651, A2 => n11811, B1 => n5823, B2 => 
                           n11821, ZN => n7471);
   U4566 : OAI22_X1 port map( A1 => n10644, A2 => n11811, B1 => n5791, B2 => 
                           n11821, ZN => n7470);
   U4567 : OAI22_X1 port map( A1 => n10637, A2 => n11811, B1 => n5759, B2 => 
                           n11821, ZN => n7469);
   U4568 : OAI22_X1 port map( A1 => n10630, A2 => n11811, B1 => n5727, B2 => 
                           n11821, ZN => n7468);
   U4569 : OAI22_X1 port map( A1 => n10849, A2 => n11549, B1 => n10534, B2 => 
                           n11550, ZN => n6795);
   U4570 : OAI22_X1 port map( A1 => n10842, A2 => n11549, B1 => n10502, B2 => 
                           n11550, ZN => n6794);
   U4571 : OAI22_X1 port map( A1 => n10835, A2 => n11549, B1 => n10470, B2 => 
                           n11550, ZN => n6793);
   U4572 : OAI22_X1 port map( A1 => n10828, A2 => n11549, B1 => n10438, B2 => 
                           n11550, ZN => n6792);
   U4573 : OAI22_X1 port map( A1 => n10821, A2 => n11549, B1 => n10406, B2 => 
                           n11551, ZN => n6791);
   U4574 : OAI22_X1 port map( A1 => n10814, A2 => n11549, B1 => n10371, B2 => 
                           n11551, ZN => n6790);
   U4575 : OAI22_X1 port map( A1 => n10807, A2 => n11549, B1 => n10339, B2 => 
                           n11551, ZN => n6789);
   U4576 : OAI22_X1 port map( A1 => n10800, A2 => n11549, B1 => n10307, B2 => 
                           n11551, ZN => n6788);
   U4577 : OAI22_X1 port map( A1 => n10793, A2 => n11548, B1 => n10272, B2 => 
                           n11552, ZN => n6787);
   U4578 : OAI22_X1 port map( A1 => n10786, A2 => n11548, B1 => n10240, B2 => 
                           n11552, ZN => n6786);
   U4579 : OAI22_X1 port map( A1 => n10779, A2 => n11548, B1 => n10208, B2 => 
                           n11552, ZN => n6785);
   U4580 : OAI22_X1 port map( A1 => n10772, A2 => n11548, B1 => n10174, B2 => 
                           n11552, ZN => n6784);
   U4581 : OAI22_X1 port map( A1 => n10765, A2 => n11548, B1 => n10142, B2 => 
                           n11553, ZN => n6783);
   U4582 : OAI22_X1 port map( A1 => n10758, A2 => n11548, B1 => n10110, B2 => 
                           n11553, ZN => n6782);
   U4583 : OAI22_X1 port map( A1 => n10751, A2 => n11548, B1 => n10078, B2 => 
                           n11553, ZN => n6781);
   U4584 : OAI22_X1 port map( A1 => n10744, A2 => n11548, B1 => n10046, B2 => 
                           n11553, ZN => n6780);
   U4585 : OAI22_X1 port map( A1 => n10737, A2 => n11548, B1 => n10014, B2 => 
                           n11554, ZN => n6779);
   U4586 : OAI22_X1 port map( A1 => n10730, A2 => n11548, B1 => n9652, B2 => 
                           n11554, ZN => n6778);
   U4587 : OAI22_X1 port map( A1 => n10723, A2 => n11548, B1 => n9620, B2 => 
                           n11554, ZN => n6777);
   U4588 : OAI22_X1 port map( A1 => n10716, A2 => n11548, B1 => n9588, B2 => 
                           n11554, ZN => n6776);
   U4589 : OAI22_X1 port map( A1 => n10709, A2 => n11547, B1 => n9254, B2 => 
                           n11555, ZN => n6775);
   U4590 : OAI22_X1 port map( A1 => n10702, A2 => n11547, B1 => n9190, B2 => 
                           n11555, ZN => n6774);
   U4591 : OAI22_X1 port map( A1 => n10695, A2 => n11547, B1 => n9158, B2 => 
                           n11555, ZN => n6773);
   U4592 : OAI22_X1 port map( A1 => n10688, A2 => n11547, B1 => n6308, B2 => 
                           n11555, ZN => n6772);
   U4593 : OAI22_X1 port map( A1 => n10681, A2 => n11547, B1 => n5991, B2 => 
                           n11556, ZN => n6771);
   U4594 : OAI22_X1 port map( A1 => n10674, A2 => n11547, B1 => n5927, B2 => 
                           n11556, ZN => n6770);
   U4595 : OAI22_X1 port map( A1 => n10667, A2 => n11547, B1 => n5895, B2 => 
                           n11556, ZN => n6769);
   U4596 : OAI22_X1 port map( A1 => n10660, A2 => n11547, B1 => n5863, B2 => 
                           n11556, ZN => n6768);
   U4597 : OAI22_X1 port map( A1 => n10653, A2 => n11547, B1 => n5831, B2 => 
                           n11557, ZN => n6767);
   U4598 : OAI22_X1 port map( A1 => n10646, A2 => n11547, B1 => n5799, B2 => 
                           n11557, ZN => n6766);
   U4599 : OAI22_X1 port map( A1 => n10639, A2 => n11547, B1 => n5767, B2 => 
                           n11557, ZN => n6765);
   U4600 : OAI22_X1 port map( A1 => n10632, A2 => n11547, B1 => n5735, B2 => 
                           n11557, ZN => n6764);
   U4601 : OAI22_X1 port map( A1 => n10850, A2 => n11489, B1 => n995, B2 => 
                           n11490, ZN => n6635);
   U4602 : OAI22_X1 port map( A1 => n10843, A2 => n11489, B1 => n991, B2 => 
                           n11490, ZN => n6634);
   U4603 : OAI22_X1 port map( A1 => n10836, A2 => n11489, B1 => n987, B2 => 
                           n11490, ZN => n6633);
   U4604 : OAI22_X1 port map( A1 => n10829, A2 => n11489, B1 => n983, B2 => 
                           n11490, ZN => n6632);
   U4605 : OAI22_X1 port map( A1 => n10822, A2 => n11489, B1 => n979, B2 => 
                           n11491, ZN => n6631);
   U4606 : OAI22_X1 port map( A1 => n10815, A2 => n11489, B1 => n975, B2 => 
                           n11491, ZN => n6630);
   U4607 : OAI22_X1 port map( A1 => n10808, A2 => n11489, B1 => n971, B2 => 
                           n11491, ZN => n6629);
   U4608 : OAI22_X1 port map( A1 => n10801, A2 => n11489, B1 => n967, B2 => 
                           n11491, ZN => n6628);
   U4609 : OAI22_X1 port map( A1 => n10794, A2 => n11488, B1 => n963, B2 => 
                           n11492, ZN => n6627);
   U4610 : OAI22_X1 port map( A1 => n10787, A2 => n11488, B1 => n959, B2 => 
                           n11492, ZN => n6626);
   U4611 : OAI22_X1 port map( A1 => n10780, A2 => n11488, B1 => n955, B2 => 
                           n11492, ZN => n6625);
   U4612 : OAI22_X1 port map( A1 => n10773, A2 => n11488, B1 => n951, B2 => 
                           n11492, ZN => n6624);
   U4613 : OAI22_X1 port map( A1 => n10766, A2 => n11488, B1 => n947, B2 => 
                           n11493, ZN => n6623);
   U4614 : OAI22_X1 port map( A1 => n10759, A2 => n11488, B1 => n943, B2 => 
                           n11493, ZN => n6622);
   U4615 : OAI22_X1 port map( A1 => n10752, A2 => n11488, B1 => n939, B2 => 
                           n11493, ZN => n6621);
   U4616 : OAI22_X1 port map( A1 => n10745, A2 => n11488, B1 => n935, B2 => 
                           n11493, ZN => n6620);
   U4617 : OAI22_X1 port map( A1 => n10738, A2 => n11488, B1 => n931, B2 => 
                           n11494, ZN => n6619);
   U4618 : OAI22_X1 port map( A1 => n10731, A2 => n11488, B1 => n927, B2 => 
                           n11494, ZN => n6618);
   U4619 : OAI22_X1 port map( A1 => n10724, A2 => n11488, B1 => n923, B2 => 
                           n11494, ZN => n6617);
   U4620 : OAI22_X1 port map( A1 => n10717, A2 => n11488, B1 => n919, B2 => 
                           n11494, ZN => n6616);
   U4621 : OAI22_X1 port map( A1 => n10710, A2 => n11487, B1 => n915, B2 => 
                           n11495, ZN => n6615);
   U4622 : OAI22_X1 port map( A1 => n10703, A2 => n11487, B1 => n911, B2 => 
                           n11495, ZN => n6614);
   U4623 : OAI22_X1 port map( A1 => n10696, A2 => n11487, B1 => n907, B2 => 
                           n11495, ZN => n6613);
   U4624 : OAI22_X1 port map( A1 => n10689, A2 => n11487, B1 => n903, B2 => 
                           n11495, ZN => n6612);
   U4625 : OAI22_X1 port map( A1 => n10682, A2 => n11487, B1 => n899, B2 => 
                           n11496, ZN => n6611);
   U4626 : OAI22_X1 port map( A1 => n10675, A2 => n11487, B1 => n895, B2 => 
                           n11496, ZN => n6610);
   U4627 : OAI22_X1 port map( A1 => n10668, A2 => n11487, B1 => n891, B2 => 
                           n11496, ZN => n6609);
   U4628 : OAI22_X1 port map( A1 => n10661, A2 => n11487, B1 => n887, B2 => 
                           n11496, ZN => n6608);
   U4629 : OAI22_X1 port map( A1 => n10654, A2 => n11487, B1 => n883, B2 => 
                           n11497, ZN => n6607);
   U4630 : OAI22_X1 port map( A1 => n10647, A2 => n11487, B1 => n879, B2 => 
                           n11497, ZN => n6606);
   U4631 : OAI22_X1 port map( A1 => n10640, A2 => n11487, B1 => n875, B2 => 
                           n11497, ZN => n6605);
   U4632 : OAI22_X1 port map( A1 => n10633, A2 => n11487, B1 => n871, B2 => 
                           n11497, ZN => n6604);
   U4633 : OAI22_X1 port map( A1 => n10850, A2 => n11453, B1 => n2337, B2 => 
                           n11454, ZN => n6539);
   U4634 : OAI22_X1 port map( A1 => n10843, A2 => n11453, B1 => n2325, B2 => 
                           n11454, ZN => n6538);
   U4635 : OAI22_X1 port map( A1 => n10836, A2 => n11453, B1 => n2313, B2 => 
                           n11454, ZN => n6537);
   U4636 : OAI22_X1 port map( A1 => n10829, A2 => n11453, B1 => n2301, B2 => 
                           n11454, ZN => n6536);
   U4637 : OAI22_X1 port map( A1 => n10822, A2 => n11453, B1 => n2289, B2 => 
                           n11455, ZN => n6535);
   U4638 : OAI22_X1 port map( A1 => n10815, A2 => n11453, B1 => n2277, B2 => 
                           n11455, ZN => n6534);
   U4639 : OAI22_X1 port map( A1 => n10808, A2 => n11453, B1 => n2265, B2 => 
                           n11455, ZN => n6533);
   U4640 : OAI22_X1 port map( A1 => n10801, A2 => n11453, B1 => n2253, B2 => 
                           n11455, ZN => n6532);
   U4641 : OAI22_X1 port map( A1 => n10794, A2 => n11452, B1 => n2241, B2 => 
                           n11456, ZN => n6531);
   U4642 : OAI22_X1 port map( A1 => n10787, A2 => n11452, B1 => n2229, B2 => 
                           n11456, ZN => n6530);
   U4643 : OAI22_X1 port map( A1 => n10780, A2 => n11452, B1 => n2217, B2 => 
                           n11456, ZN => n6529);
   U4644 : OAI22_X1 port map( A1 => n10773, A2 => n11452, B1 => n2173_port, B2 
                           => n11456, ZN => n6528);
   U4645 : OAI22_X1 port map( A1 => n10766, A2 => n11452, B1 => n2161, B2 => 
                           n11457, ZN => n6527);
   U4646 : OAI22_X1 port map( A1 => n10759, A2 => n11452, B1 => n2149, B2 => 
                           n11457, ZN => n6526);
   U4647 : OAI22_X1 port map( A1 => n10752, A2 => n11452, B1 => n2105, B2 => 
                           n11457, ZN => n6525);
   U4648 : OAI22_X1 port map( A1 => n10745, A2 => n11452, B1 => n2093, B2 => 
                           n11457, ZN => n6524);
   U4649 : OAI22_X1 port map( A1 => n10738, A2 => n11452, B1 => n2049, B2 => 
                           n11458, ZN => n6523);
   U4650 : OAI22_X1 port map( A1 => n10731, A2 => n11452, B1 => n2037, B2 => 
                           n11458, ZN => n6522);
   U4651 : OAI22_X1 port map( A1 => n10724, A2 => n11452, B1 => n2025, B2 => 
                           n11458, ZN => n6521);
   U4652 : OAI22_X1 port map( A1 => n10717, A2 => n11452, B1 => n2013, B2 => 
                           n11458, ZN => n6520);
   U4653 : OAI22_X1 port map( A1 => n10710, A2 => n11451, B1 => n2001, B2 => 
                           n11459, ZN => n6519);
   U4654 : OAI22_X1 port map( A1 => n10703, A2 => n11451, B1 => n1989, B2 => 
                           n11459, ZN => n6518);
   U4655 : OAI22_X1 port map( A1 => n10696, A2 => n11451, B1 => n1977, B2 => 
                           n11459, ZN => n6517);
   U4656 : OAI22_X1 port map( A1 => n10689, A2 => n11451, B1 => n1965, B2 => 
                           n11459, ZN => n6516);
   U4657 : OAI22_X1 port map( A1 => n10682, A2 => n11451, B1 => n1953, B2 => 
                           n11460, ZN => n6515);
   U4658 : OAI22_X1 port map( A1 => n10675, A2 => n11451, B1 => n1941, B2 => 
                           n11460, ZN => n6514);
   U4659 : OAI22_X1 port map( A1 => n10668, A2 => n11451, B1 => n1929, B2 => 
                           n11460, ZN => n6513);
   U4660 : OAI22_X1 port map( A1 => n10661, A2 => n11451, B1 => n1917, B2 => 
                           n11460, ZN => n6512);
   U4661 : OAI22_X1 port map( A1 => n10654, A2 => n11451, B1 => n1905, B2 => 
                           n11461, ZN => n6511);
   U4662 : OAI22_X1 port map( A1 => n10647, A2 => n11451, B1 => n1893, B2 => 
                           n11461, ZN => n6510);
   U4663 : OAI22_X1 port map( A1 => n10640, A2 => n11451, B1 => n1881, B2 => 
                           n11461, ZN => n6509);
   U4664 : OAI22_X1 port map( A1 => n10633, A2 => n11451, B1 => n1869, B2 => 
                           n11461, ZN => n6508);
   U4665 : OAI22_X1 port map( A1 => n10850, A2 => n11417, B1 => n2338, B2 => 
                           n11418, ZN => n6443);
   U4666 : OAI22_X1 port map( A1 => n10843, A2 => n11417, B1 => n2326, B2 => 
                           n11418, ZN => n6442);
   U4667 : OAI22_X1 port map( A1 => n10836, A2 => n11417, B1 => n2314, B2 => 
                           n11418, ZN => n6441);
   U4668 : OAI22_X1 port map( A1 => n10829, A2 => n11417, B1 => n2302, B2 => 
                           n11418, ZN => n6440);
   U4669 : OAI22_X1 port map( A1 => n10822, A2 => n11417, B1 => n2290, B2 => 
                           n11419, ZN => n6439);
   U4670 : OAI22_X1 port map( A1 => n10815, A2 => n11417, B1 => n2278, B2 => 
                           n11419, ZN => n6438);
   U4671 : OAI22_X1 port map( A1 => n10808, A2 => n11417, B1 => n2266, B2 => 
                           n11419, ZN => n6437);
   U4672 : OAI22_X1 port map( A1 => n10801, A2 => n11417, B1 => n2254, B2 => 
                           n11419, ZN => n6436);
   U4673 : OAI22_X1 port map( A1 => n10794, A2 => n11416, B1 => n2242, B2 => 
                           n11420, ZN => n6435);
   U4674 : OAI22_X1 port map( A1 => n10787, A2 => n11416, B1 => n2230, B2 => 
                           n11420, ZN => n6434);
   U4675 : OAI22_X1 port map( A1 => n10780, A2 => n11416, B1 => n2218, B2 => 
                           n11420, ZN => n6433);
   U4676 : OAI22_X1 port map( A1 => n10773, A2 => n11416, B1 => n2174, B2 => 
                           n11420, ZN => n6432);
   U4677 : OAI22_X1 port map( A1 => n10766, A2 => n11416, B1 => n2162, B2 => 
                           n11421, ZN => n6431);
   U4678 : OAI22_X1 port map( A1 => n10759, A2 => n11416, B1 => n2150, B2 => 
                           n11421, ZN => n6430);
   U4679 : OAI22_X1 port map( A1 => n10752, A2 => n11416, B1 => n2106, B2 => 
                           n11421, ZN => n6429);
   U4680 : OAI22_X1 port map( A1 => n10745, A2 => n11416, B1 => n2094, B2 => 
                           n11421, ZN => n6428);
   U4681 : OAI22_X1 port map( A1 => n10738, A2 => n11416, B1 => n2082, B2 => 
                           n11422, ZN => n6427);
   U4682 : OAI22_X1 port map( A1 => n10731, A2 => n11416, B1 => n2038, B2 => 
                           n11422, ZN => n6426);
   U4683 : OAI22_X1 port map( A1 => n10724, A2 => n11416, B1 => n2026, B2 => 
                           n11422, ZN => n6425);
   U4684 : OAI22_X1 port map( A1 => n10717, A2 => n11416, B1 => n2014, B2 => 
                           n11422, ZN => n6424);
   U4685 : OAI22_X1 port map( A1 => n10710, A2 => n11415, B1 => n2002, B2 => 
                           n11423, ZN => n6423);
   U4686 : OAI22_X1 port map( A1 => n10703, A2 => n11415, B1 => n1990, B2 => 
                           n11423, ZN => n6422);
   U4687 : OAI22_X1 port map( A1 => n10696, A2 => n11415, B1 => n1978, B2 => 
                           n11423, ZN => n6421);
   U4688 : OAI22_X1 port map( A1 => n10689, A2 => n11415, B1 => n1966, B2 => 
                           n11423, ZN => n6420);
   U4689 : OAI22_X1 port map( A1 => n10682, A2 => n11415, B1 => n1954, B2 => 
                           n11424, ZN => n6419);
   U4690 : OAI22_X1 port map( A1 => n10675, A2 => n11415, B1 => n1942, B2 => 
                           n11424, ZN => n6418);
   U4691 : OAI22_X1 port map( A1 => n10668, A2 => n11415, B1 => n1930, B2 => 
                           n11424, ZN => n6417);
   U4692 : OAI22_X1 port map( A1 => n10661, A2 => n11415, B1 => n1918, B2 => 
                           n11424, ZN => n6416);
   U4693 : OAI22_X1 port map( A1 => n10654, A2 => n11415, B1 => n1906, B2 => 
                           n11425, ZN => n6415);
   U4694 : OAI22_X1 port map( A1 => n10647, A2 => n11415, B1 => n1894, B2 => 
                           n11425, ZN => n6414);
   U4695 : OAI22_X1 port map( A1 => n10640, A2 => n11415, B1 => n1882, B2 => 
                           n11425, ZN => n6413);
   U4696 : OAI22_X1 port map( A1 => n10633, A2 => n11415, B1 => n1870, B2 => 
                           n11425, ZN => n6412);
   U4697 : OAI22_X1 port map( A1 => n10846, A2 => n12041, B1 => n10520, B2 => 
                           n12042, ZN => n8107);
   U4698 : OAI22_X1 port map( A1 => n10839, A2 => n12041, B1 => n10488, B2 => 
                           n12042, ZN => n8106);
   U4699 : OAI22_X1 port map( A1 => n10832, A2 => n12041, B1 => n10456, B2 => 
                           n12042, ZN => n8105);
   U4700 : OAI22_X1 port map( A1 => n10825, A2 => n12041, B1 => n10424, B2 => 
                           n12042, ZN => n8104);
   U4701 : OAI22_X1 port map( A1 => n10818, A2 => n12041, B1 => n10389, B2 => 
                           n12043, ZN => n8103);
   U4702 : OAI22_X1 port map( A1 => n10811, A2 => n12041, B1 => n10357, B2 => 
                           n12043, ZN => n8102);
   U4703 : OAI22_X1 port map( A1 => n10804, A2 => n12041, B1 => n10325, B2 => 
                           n12043, ZN => n8101);
   U4704 : OAI22_X1 port map( A1 => n10797, A2 => n12041, B1 => n10290, B2 => 
                           n12043, ZN => n8100);
   U4705 : OAI22_X1 port map( A1 => n10790, A2 => n12040, B1 => n10258, B2 => 
                           n12044, ZN => n8099);
   U4706 : OAI22_X1 port map( A1 => n10783, A2 => n12040, B1 => n10226, B2 => 
                           n12044, ZN => n8098);
   U4707 : OAI22_X1 port map( A1 => n10776, A2 => n12040, B1 => n10192, B2 => 
                           n12044, ZN => n8097);
   U4708 : OAI22_X1 port map( A1 => n10769, A2 => n12040, B1 => n10160, B2 => 
                           n12044, ZN => n8096);
   U4709 : OAI22_X1 port map( A1 => n10762, A2 => n12040, B1 => n10128, B2 => 
                           n12045, ZN => n8095);
   U4710 : OAI22_X1 port map( A1 => n10755, A2 => n12040, B1 => n10096, B2 => 
                           n12045, ZN => n8094);
   U4711 : OAI22_X1 port map( A1 => n10748, A2 => n12040, B1 => n10064, B2 => 
                           n12045, ZN => n8093);
   U4712 : OAI22_X1 port map( A1 => n10741, A2 => n12040, B1 => n10032, B2 => 
                           n12045, ZN => n8092);
   U4713 : OAI22_X1 port map( A1 => n10734, A2 => n12040, B1 => n10000, B2 => 
                           n12046, ZN => n8091);
   U4714 : OAI22_X1 port map( A1 => n10727, A2 => n12040, B1 => n9638, B2 => 
                           n12046, ZN => n8090);
   U4715 : OAI22_X1 port map( A1 => n10720, A2 => n12040, B1 => n9606, B2 => 
                           n12046, ZN => n8089);
   U4716 : OAI22_X1 port map( A1 => n10713, A2 => n12040, B1 => n9574, B2 => 
                           n12046, ZN => n8088);
   U4717 : OAI22_X1 port map( A1 => n10706, A2 => n12039, B1 => n9208, B2 => 
                           n12047, ZN => n8087);
   U4718 : OAI22_X1 port map( A1 => n10699, A2 => n12039, B1 => n9176, B2 => 
                           n12047, ZN => n8086);
   U4719 : OAI22_X1 port map( A1 => n10692, A2 => n12039, B1 => n9144, B2 => 
                           n12047, ZN => n8085);
   U4720 : OAI22_X1 port map( A1 => n10685, A2 => n12039, B1 => n6009, B2 => 
                           n12047, ZN => n8084);
   U4721 : OAI22_X1 port map( A1 => n10678, A2 => n12039, B1 => n5945, B2 => 
                           n12048, ZN => n8083);
   U4722 : OAI22_X1 port map( A1 => n10671, A2 => n12039, B1 => n5913, B2 => 
                           n12048, ZN => n8082);
   U4723 : OAI22_X1 port map( A1 => n10664, A2 => n12039, B1 => n5881, B2 => 
                           n12048, ZN => n8081);
   U4724 : OAI22_X1 port map( A1 => n10657, A2 => n12039, B1 => n5849, B2 => 
                           n12048, ZN => n8080);
   U4725 : OAI22_X1 port map( A1 => n10650, A2 => n12039, B1 => n5817, B2 => 
                           n12049, ZN => n8079);
   U4726 : OAI22_X1 port map( A1 => n10643, A2 => n12039, B1 => n5785, B2 => 
                           n12049, ZN => n8078);
   U4727 : OAI22_X1 port map( A1 => n10636, A2 => n12039, B1 => n5753, B2 => 
                           n12049, ZN => n8077);
   U4728 : OAI22_X1 port map( A1 => n10629, A2 => n12039, B1 => n5721, B2 => 
                           n12049, ZN => n8076);
   U4729 : OAI22_X1 port map( A1 => n10848, A2 => n11777, B1 => n10528, B2 => 
                           n11778, ZN => n7403);
   U4730 : OAI22_X1 port map( A1 => n10841, A2 => n11777, B1 => n10496, B2 => 
                           n11778, ZN => n7402);
   U4731 : OAI22_X1 port map( A1 => n10834, A2 => n11777, B1 => n10464, B2 => 
                           n11778, ZN => n7401);
   U4732 : OAI22_X1 port map( A1 => n10827, A2 => n11777, B1 => n10432, B2 => 
                           n11778, ZN => n7400);
   U4733 : OAI22_X1 port map( A1 => n10820, A2 => n11777, B1 => n10400, B2 => 
                           n11779, ZN => n7399);
   U4734 : OAI22_X1 port map( A1 => n10813, A2 => n11777, B1 => n10365, B2 => 
                           n11779, ZN => n7398);
   U4735 : OAI22_X1 port map( A1 => n10806, A2 => n11777, B1 => n10333, B2 => 
                           n11779, ZN => n7397);
   U4736 : OAI22_X1 port map( A1 => n10799, A2 => n11777, B1 => n10298, B2 => 
                           n11779, ZN => n7396);
   U4737 : OAI22_X1 port map( A1 => n10792, A2 => n11776, B1 => n10266, B2 => 
                           n11780, ZN => n7395);
   U4738 : OAI22_X1 port map( A1 => n10785, A2 => n11776, B1 => n10234, B2 => 
                           n11780, ZN => n7394);
   U4739 : OAI22_X1 port map( A1 => n10778, A2 => n11776, B1 => n10200, B2 => 
                           n11780, ZN => n7393);
   U4740 : OAI22_X1 port map( A1 => n10771, A2 => n11776, B1 => n10168, B2 => 
                           n11780, ZN => n7392);
   U4741 : OAI22_X1 port map( A1 => n10764, A2 => n11776, B1 => n10136, B2 => 
                           n11781, ZN => n7391);
   U4742 : OAI22_X1 port map( A1 => n10757, A2 => n11776, B1 => n10104, B2 => 
                           n11781, ZN => n7390);
   U4743 : OAI22_X1 port map( A1 => n10750, A2 => n11776, B1 => n10072, B2 => 
                           n11781, ZN => n7389);
   U4744 : OAI22_X1 port map( A1 => n10743, A2 => n11776, B1 => n10040, B2 => 
                           n11781, ZN => n7388);
   U4745 : OAI22_X1 port map( A1 => n10736, A2 => n11776, B1 => n10008, B2 => 
                           n11782, ZN => n7387);
   U4746 : OAI22_X1 port map( A1 => n10729, A2 => n11776, B1 => n9646, B2 => 
                           n11782, ZN => n7386);
   U4747 : OAI22_X1 port map( A1 => n10722, A2 => n11776, B1 => n9614, B2 => 
                           n11782, ZN => n7385);
   U4748 : OAI22_X1 port map( A1 => n10715, A2 => n11776, B1 => n9582, B2 => 
                           n11782, ZN => n7384);
   U4749 : OAI22_X1 port map( A1 => n10708, A2 => n11775, B1 => n9248, B2 => 
                           n11783, ZN => n7383);
   U4750 : OAI22_X1 port map( A1 => n10701, A2 => n11775, B1 => n9184, B2 => 
                           n11783, ZN => n7382);
   U4751 : OAI22_X1 port map( A1 => n10694, A2 => n11775, B1 => n9152, B2 => 
                           n11783, ZN => n7381);
   U4752 : OAI22_X1 port map( A1 => n10687, A2 => n11775, B1 => n6302, B2 => 
                           n11783, ZN => n7380);
   U4753 : OAI22_X1 port map( A1 => n10680, A2 => n11775, B1 => n5985, B2 => 
                           n11784, ZN => n7379);
   U4754 : OAI22_X1 port map( A1 => n10673, A2 => n11775, B1 => n5921, B2 => 
                           n11784, ZN => n7378);
   U4755 : OAI22_X1 port map( A1 => n10666, A2 => n11775, B1 => n5889, B2 => 
                           n11784, ZN => n7377);
   U4756 : OAI22_X1 port map( A1 => n10659, A2 => n11775, B1 => n5857, B2 => 
                           n11784, ZN => n7376);
   U4757 : OAI22_X1 port map( A1 => n10652, A2 => n11775, B1 => n5825, B2 => 
                           n11785, ZN => n7375);
   U4758 : OAI22_X1 port map( A1 => n10645, A2 => n11775, B1 => n5793, B2 => 
                           n11785, ZN => n7374);
   U4759 : OAI22_X1 port map( A1 => n10638, A2 => n11775, B1 => n5761, B2 => 
                           n11785, ZN => n7373);
   U4760 : OAI22_X1 port map( A1 => n10631, A2 => n11775, B1 => n5729, B2 => 
                           n11785, ZN => n7372);
   U4761 : OAI22_X1 port map( A1 => n10850, A2 => n11393, B1 => n515, B2 => 
                           n11394, ZN => n6379);
   U4762 : OAI22_X1 port map( A1 => n10843, A2 => n11393, B1 => n503, B2 => 
                           n11394, ZN => n6378);
   U4763 : OAI22_X1 port map( A1 => n10836, A2 => n11393, B1 => n491, B2 => 
                           n11394, ZN => n6377);
   U4764 : OAI22_X1 port map( A1 => n10829, A2 => n11393, B1 => n479, B2 => 
                           n11394, ZN => n6376);
   U4765 : OAI22_X1 port map( A1 => n10822, A2 => n11393, B1 => n467, B2 => 
                           n11395, ZN => n6375);
   U4766 : OAI22_X1 port map( A1 => n10815, A2 => n11393, B1 => n455, B2 => 
                           n11395, ZN => n6374);
   U4767 : OAI22_X1 port map( A1 => n10808, A2 => n11393, B1 => n443, B2 => 
                           n11395, ZN => n6373);
   U4768 : OAI22_X1 port map( A1 => n10801, A2 => n11393, B1 => n431, B2 => 
                           n11395, ZN => n6372);
   U4769 : OAI22_X1 port map( A1 => n10794, A2 => n11392, B1 => n419, B2 => 
                           n11396, ZN => n6371);
   U4770 : OAI22_X1 port map( A1 => n10787, A2 => n11392, B1 => n407, B2 => 
                           n11396, ZN => n6370);
   U4771 : OAI22_X1 port map( A1 => n10780, A2 => n11392, B1 => n395, B2 => 
                           n11396, ZN => n6369);
   U4772 : OAI22_X1 port map( A1 => n10773, A2 => n11392, B1 => n383, B2 => 
                           n11396, ZN => n6368);
   U4773 : OAI22_X1 port map( A1 => n10766, A2 => n11392, B1 => n371, B2 => 
                           n11397, ZN => n6367);
   U4774 : OAI22_X1 port map( A1 => n10759, A2 => n11392, B1 => n359, B2 => 
                           n11397, ZN => n6366);
   U4775 : OAI22_X1 port map( A1 => n10752, A2 => n11392, B1 => n347, B2 => 
                           n11397, ZN => n6365);
   U4776 : OAI22_X1 port map( A1 => n10745, A2 => n11392, B1 => n335, B2 => 
                           n11397, ZN => n6364);
   U4777 : OAI22_X1 port map( A1 => n10738, A2 => n11392, B1 => n323, B2 => 
                           n11398, ZN => n6363);
   U4778 : OAI22_X1 port map( A1 => n10731, A2 => n11392, B1 => n311, B2 => 
                           n11398, ZN => n6362);
   U4779 : OAI22_X1 port map( A1 => n10724, A2 => n11392, B1 => n299, B2 => 
                           n11398, ZN => n6361);
   U4780 : OAI22_X1 port map( A1 => n10717, A2 => n11392, B1 => n287, B2 => 
                           n11398, ZN => n6360);
   U4781 : OAI22_X1 port map( A1 => n10710, A2 => n11391, B1 => n275, B2 => 
                           n11399, ZN => n6359);
   U4782 : OAI22_X1 port map( A1 => n10703, A2 => n11391, B1 => n263, B2 => 
                           n11399, ZN => n6358);
   U4783 : OAI22_X1 port map( A1 => n10696, A2 => n11391, B1 => n251, B2 => 
                           n11399, ZN => n6357);
   U4784 : OAI22_X1 port map( A1 => n10689, A2 => n11391, B1 => n239, B2 => 
                           n11399, ZN => n6356);
   U4785 : OAI22_X1 port map( A1 => n10682, A2 => n11391, B1 => n227, B2 => 
                           n11400, ZN => n6355);
   U4786 : OAI22_X1 port map( A1 => n10675, A2 => n11391, B1 => n215, B2 => 
                           n11400, ZN => n6354);
   U4787 : OAI22_X1 port map( A1 => n10668, A2 => n11391, B1 => n203, B2 => 
                           n11400, ZN => n6353);
   U4788 : OAI22_X1 port map( A1 => n10661, A2 => n11391, B1 => n191, B2 => 
                           n11400, ZN => n6352);
   U4789 : OAI22_X1 port map( A1 => n10654, A2 => n11391, B1 => n179, B2 => 
                           n11401, ZN => n6351);
   U4790 : OAI22_X1 port map( A1 => n10647, A2 => n11391, B1 => n167, B2 => 
                           n11401, ZN => n6350);
   U4791 : OAI22_X1 port map( A1 => n10640, A2 => n11391, B1 => n155, B2 => 
                           n11401, ZN => n6349);
   U4792 : OAI22_X1 port map( A1 => n10633, A2 => n11391, B1 => n143, B2 => 
                           n11401, ZN => n6348);
   U4793 : OAI22_X1 port map( A1 => n10845, A2 => n12149, B1 => n10521, B2 => 
                           n12150, ZN => n8395);
   U4794 : OAI22_X1 port map( A1 => n10838, A2 => n12149, B1 => n10489, B2 => 
                           n12150, ZN => n8394);
   U4795 : OAI22_X1 port map( A1 => n10831, A2 => n12149, B1 => n10457, B2 => 
                           n12150, ZN => n8393);
   U4796 : OAI22_X1 port map( A1 => n10824, A2 => n12149, B1 => n10425, B2 => 
                           n12150, ZN => n8392);
   U4797 : OAI22_X1 port map( A1 => n10817, A2 => n12149, B1 => n10390, B2 => 
                           n12151, ZN => n8391);
   U4798 : OAI22_X1 port map( A1 => n10810, A2 => n12149, B1 => n10358, B2 => 
                           n12151, ZN => n8390);
   U4799 : OAI22_X1 port map( A1 => n10803, A2 => n12149, B1 => n10326, B2 => 
                           n12151, ZN => n8389);
   U4800 : OAI22_X1 port map( A1 => n10796, A2 => n12149, B1 => n10291, B2 => 
                           n12151, ZN => n8388);
   U4801 : OAI22_X1 port map( A1 => n10789, A2 => n12148, B1 => n10259, B2 => 
                           n12152, ZN => n8387);
   U4802 : OAI22_X1 port map( A1 => n10782, A2 => n12148, B1 => n10227, B2 => 
                           n12152, ZN => n8386);
   U4803 : OAI22_X1 port map( A1 => n10775, A2 => n12148, B1 => n10193, B2 => 
                           n12152, ZN => n8385);
   U4804 : OAI22_X1 port map( A1 => n10768, A2 => n12148, B1 => n10161, B2 => 
                           n12152, ZN => n8384);
   U4805 : OAI22_X1 port map( A1 => n10761, A2 => n12148, B1 => n10129, B2 => 
                           n12153, ZN => n8383);
   U4806 : OAI22_X1 port map( A1 => n10754, A2 => n12148, B1 => n10097, B2 => 
                           n12153, ZN => n8382);
   U4807 : OAI22_X1 port map( A1 => n10747, A2 => n12148, B1 => n10065, B2 => 
                           n12153, ZN => n8381);
   U4808 : OAI22_X1 port map( A1 => n10740, A2 => n12148, B1 => n10033, B2 => 
                           n12153, ZN => n8380);
   U4809 : OAI22_X1 port map( A1 => n10733, A2 => n12148, B1 => n10001, B2 => 
                           n12154, ZN => n8379);
   U4810 : OAI22_X1 port map( A1 => n10726, A2 => n12148, B1 => n9639, B2 => 
                           n12154, ZN => n8378);
   U4811 : OAI22_X1 port map( A1 => n10719, A2 => n12148, B1 => n9607, B2 => 
                           n12154, ZN => n8377);
   U4812 : OAI22_X1 port map( A1 => n10712, A2 => n12148, B1 => n9575, B2 => 
                           n12154, ZN => n8376);
   U4813 : OAI22_X1 port map( A1 => n10705, A2 => n12147, B1 => n9209, B2 => 
                           n12155, ZN => n8375);
   U4814 : OAI22_X1 port map( A1 => n10698, A2 => n12147, B1 => n9177, B2 => 
                           n12155, ZN => n8374);
   U4815 : OAI22_X1 port map( A1 => n10691, A2 => n12147, B1 => n9145, B2 => 
                           n12155, ZN => n8373);
   U4816 : OAI22_X1 port map( A1 => n10684, A2 => n12147, B1 => n6010, B2 => 
                           n12155, ZN => n8372);
   U4817 : OAI22_X1 port map( A1 => n10677, A2 => n12147, B1 => n5946, B2 => 
                           n12156, ZN => n8371);
   U4818 : OAI22_X1 port map( A1 => n10670, A2 => n12147, B1 => n5914, B2 => 
                           n12156, ZN => n8370);
   U4819 : OAI22_X1 port map( A1 => n10663, A2 => n12147, B1 => n5882, B2 => 
                           n12156, ZN => n8369);
   U4820 : OAI22_X1 port map( A1 => n10656, A2 => n12147, B1 => n5850, B2 => 
                           n12156, ZN => n8368);
   U4821 : OAI22_X1 port map( A1 => n10649, A2 => n12147, B1 => n5818, B2 => 
                           n12157, ZN => n8367);
   U4822 : OAI22_X1 port map( A1 => n10642, A2 => n12147, B1 => n5786, B2 => 
                           n12157, ZN => n8366);
   U4823 : OAI22_X1 port map( A1 => n10635, A2 => n12147, B1 => n5754, B2 => 
                           n12157, ZN => n8365);
   U4824 : OAI22_X1 port map( A1 => n10628, A2 => n12147, B1 => n5722, B2 => 
                           n12157, ZN => n8364);
   U4825 : OAI22_X1 port map( A1 => n10847, A2 => n11885, B1 => n10529, B2 => 
                           n11886, ZN => n7691);
   U4826 : OAI22_X1 port map( A1 => n10840, A2 => n11885, B1 => n10497, B2 => 
                           n11886, ZN => n7690);
   U4827 : OAI22_X1 port map( A1 => n10833, A2 => n11885, B1 => n10465, B2 => 
                           n11886, ZN => n7689);
   U4828 : OAI22_X1 port map( A1 => n10826, A2 => n11885, B1 => n10433, B2 => 
                           n11886, ZN => n7688);
   U4829 : OAI22_X1 port map( A1 => n10819, A2 => n11885, B1 => n10401, B2 => 
                           n11887, ZN => n7687);
   U4830 : OAI22_X1 port map( A1 => n10812, A2 => n11885, B1 => n10366, B2 => 
                           n11887, ZN => n7686);
   U4831 : OAI22_X1 port map( A1 => n10805, A2 => n11885, B1 => n10334, B2 => 
                           n11887, ZN => n7685);
   U4832 : OAI22_X1 port map( A1 => n10798, A2 => n11885, B1 => n10299, B2 => 
                           n11887, ZN => n7684);
   U4833 : OAI22_X1 port map( A1 => n10791, A2 => n11884, B1 => n10267, B2 => 
                           n11888, ZN => n7683);
   U4834 : OAI22_X1 port map( A1 => n10784, A2 => n11884, B1 => n10235, B2 => 
                           n11888, ZN => n7682);
   U4835 : OAI22_X1 port map( A1 => n10777, A2 => n11884, B1 => n10201, B2 => 
                           n11888, ZN => n7681);
   U4836 : OAI22_X1 port map( A1 => n10770, A2 => n11884, B1 => n10169, B2 => 
                           n11888, ZN => n7680);
   U4837 : OAI22_X1 port map( A1 => n10763, A2 => n11884, B1 => n10137, B2 => 
                           n11889, ZN => n7679);
   U4838 : OAI22_X1 port map( A1 => n10756, A2 => n11884, B1 => n10105, B2 => 
                           n11889, ZN => n7678);
   U4839 : OAI22_X1 port map( A1 => n10749, A2 => n11884, B1 => n10073, B2 => 
                           n11889, ZN => n7677);
   U4840 : OAI22_X1 port map( A1 => n10742, A2 => n11884, B1 => n10041, B2 => 
                           n11889, ZN => n7676);
   U4841 : OAI22_X1 port map( A1 => n10735, A2 => n11884, B1 => n10009, B2 => 
                           n11890, ZN => n7675);
   U4842 : OAI22_X1 port map( A1 => n10728, A2 => n11884, B1 => n9647, B2 => 
                           n11890, ZN => n7674);
   U4843 : OAI22_X1 port map( A1 => n10721, A2 => n11884, B1 => n9615, B2 => 
                           n11890, ZN => n7673);
   U4844 : OAI22_X1 port map( A1 => n10714, A2 => n11884, B1 => n9583, B2 => 
                           n11890, ZN => n7672);
   U4845 : OAI22_X1 port map( A1 => n10707, A2 => n11883, B1 => n9249, B2 => 
                           n11891, ZN => n7671);
   U4846 : OAI22_X1 port map( A1 => n10700, A2 => n11883, B1 => n9185, B2 => 
                           n11891, ZN => n7670);
   U4847 : OAI22_X1 port map( A1 => n10693, A2 => n11883, B1 => n9153, B2 => 
                           n11891, ZN => n7669);
   U4848 : OAI22_X1 port map( A1 => n10686, A2 => n11883, B1 => n6303, B2 => 
                           n11891, ZN => n7668);
   U4849 : OAI22_X1 port map( A1 => n10679, A2 => n11883, B1 => n5986, B2 => 
                           n11892, ZN => n7667);
   U4850 : OAI22_X1 port map( A1 => n10672, A2 => n11883, B1 => n5922, B2 => 
                           n11892, ZN => n7666);
   U4851 : OAI22_X1 port map( A1 => n10665, A2 => n11883, B1 => n5890, B2 => 
                           n11892, ZN => n7665);
   U4852 : OAI22_X1 port map( A1 => n10658, A2 => n11883, B1 => n5858, B2 => 
                           n11892, ZN => n7664);
   U4853 : OAI22_X1 port map( A1 => n10651, A2 => n11883, B1 => n5826, B2 => 
                           n11893, ZN => n7663);
   U4854 : OAI22_X1 port map( A1 => n10644, A2 => n11883, B1 => n5794, B2 => 
                           n11893, ZN => n7662);
   U4855 : OAI22_X1 port map( A1 => n10637, A2 => n11883, B1 => n5762, B2 => 
                           n11893, ZN => n7661);
   U4856 : OAI22_X1 port map( A1 => n10630, A2 => n11883, B1 => n5730, B2 => 
                           n11893, ZN => n7660);
   U4857 : OAI22_X1 port map( A1 => n10850, A2 => n11381, B1 => n2339, B2 => 
                           n11382, ZN => n6347);
   U4858 : OAI22_X1 port map( A1 => n10843, A2 => n11381, B1 => n2327, B2 => 
                           n11382, ZN => n6346);
   U4859 : OAI22_X1 port map( A1 => n10836, A2 => n11381, B1 => n2315, B2 => 
                           n11382, ZN => n6345);
   U4860 : OAI22_X1 port map( A1 => n10829, A2 => n11381, B1 => n2303, B2 => 
                           n11382, ZN => n6344);
   U4861 : OAI22_X1 port map( A1 => n10822, A2 => n11381, B1 => n2291, B2 => 
                           n11383, ZN => n6343);
   U4862 : OAI22_X1 port map( A1 => n10815, A2 => n11381, B1 => n2279, B2 => 
                           n11383, ZN => n6342);
   U4863 : OAI22_X1 port map( A1 => n10808, A2 => n11381, B1 => n2267, B2 => 
                           n11383, ZN => n6341);
   U4864 : OAI22_X1 port map( A1 => n10801, A2 => n11381, B1 => n2255, B2 => 
                           n11383, ZN => n6340);
   U4865 : OAI22_X1 port map( A1 => n10794, A2 => n11380, B1 => n2243, B2 => 
                           n11384, ZN => n6339);
   U4866 : OAI22_X1 port map( A1 => n10787, A2 => n11380, B1 => n2231, B2 => 
                           n11384, ZN => n6338);
   U4867 : OAI22_X1 port map( A1 => n10780, A2 => n11380, B1 => n2219, B2 => 
                           n11384, ZN => n6337);
   U4868 : OAI22_X1 port map( A1 => n10773, A2 => n11380, B1 => n2175, B2 => 
                           n11384, ZN => n6336);
   U4869 : OAI22_X1 port map( A1 => n10766, A2 => n11380, B1 => n2163, B2 => 
                           n11385, ZN => n6335);
   U4870 : OAI22_X1 port map( A1 => n10759, A2 => n11380, B1 => n2151, B2 => 
                           n11385, ZN => n6334);
   U4871 : OAI22_X1 port map( A1 => n10752, A2 => n11380, B1 => n2107, B2 => 
                           n11385, ZN => n6333);
   U4872 : OAI22_X1 port map( A1 => n10745, A2 => n11380, B1 => n2095, B2 => 
                           n11385, ZN => n6332);
   U4873 : OAI22_X1 port map( A1 => n10738, A2 => n11380, B1 => n2083, B2 => 
                           n11386, ZN => n6331);
   U4874 : OAI22_X1 port map( A1 => n10731, A2 => n11380, B1 => n2039, B2 => 
                           n11386, ZN => n6330);
   U4875 : OAI22_X1 port map( A1 => n10724, A2 => n11380, B1 => n2027, B2 => 
                           n11386, ZN => n6329);
   U4876 : OAI22_X1 port map( A1 => n10717, A2 => n11380, B1 => n2015, B2 => 
                           n11386, ZN => n6328);
   U4877 : OAI22_X1 port map( A1 => n10710, A2 => n11379, B1 => n2003, B2 => 
                           n11387, ZN => n6327);
   U4878 : OAI22_X1 port map( A1 => n10703, A2 => n11379, B1 => n1991, B2 => 
                           n11387, ZN => n6326);
   U4879 : OAI22_X1 port map( A1 => n10696, A2 => n11379, B1 => n1979, B2 => 
                           n11387, ZN => n6325);
   U4880 : OAI22_X1 port map( A1 => n10689, A2 => n11379, B1 => n1967, B2 => 
                           n11387, ZN => n6324);
   U4881 : OAI22_X1 port map( A1 => n10682, A2 => n11379, B1 => n1955, B2 => 
                           n11388, ZN => n6323);
   U4882 : OAI22_X1 port map( A1 => n10675, A2 => n11379, B1 => n1943, B2 => 
                           n11388, ZN => n6322);
   U4883 : OAI22_X1 port map( A1 => n10668, A2 => n11379, B1 => n1931, B2 => 
                           n11388, ZN => n6321);
   U4884 : OAI22_X1 port map( A1 => n10661, A2 => n11379, B1 => n1919, B2 => 
                           n11388, ZN => n6320);
   U4885 : OAI22_X1 port map( A1 => n10654, A2 => n11379, B1 => n1907, B2 => 
                           n11389, ZN => n6319);
   U4886 : OAI22_X1 port map( A1 => n10647, A2 => n11379, B1 => n1895, B2 => 
                           n11389, ZN => n6318);
   U4887 : OAI22_X1 port map( A1 => n10640, A2 => n11379, B1 => n1883, B2 => 
                           n11389, ZN => n6317);
   U4888 : OAI22_X1 port map( A1 => n10633, A2 => n11379, B1 => n1871, B2 => 
                           n11389, ZN => n6316);
   U4889 : OAI22_X1 port map( A1 => n10844, A2 => n12406, B1 => n10513, B2 => 
                           n12407, ZN => n9099);
   U4890 : OAI22_X1 port map( A1 => n10837, A2 => n12405, B1 => n10481, B2 => 
                           n12407, ZN => n9098);
   U4891 : OAI22_X1 port map( A1 => n10830, A2 => n12406, B1 => n10449, B2 => 
                           n12407, ZN => n9097);
   U4892 : OAI22_X1 port map( A1 => n10823, A2 => n12405, B1 => n10417, B2 => 
                           n12407, ZN => n9096);
   U4893 : OAI22_X1 port map( A1 => n10816, A2 => n12406, B1 => n10382, B2 => 
                           n12408, ZN => n9095);
   U4894 : OAI22_X1 port map( A1 => n10809, A2 => n12405, B1 => n10350, B2 => 
                           n12408, ZN => n9094);
   U4895 : OAI22_X1 port map( A1 => n10802, A2 => n12406, B1 => n10318, B2 => 
                           n12408, ZN => n9093);
   U4896 : OAI22_X1 port map( A1 => n10795, A2 => n12405, B1 => n10283, B2 => 
                           n12408, ZN => n9092);
   U4897 : OAI22_X1 port map( A1 => n10788, A2 => n12406, B1 => n10251, B2 => 
                           n12409, ZN => n9091);
   U4898 : OAI22_X1 port map( A1 => n10781, A2 => n12406, B1 => n10219, B2 => 
                           n12409, ZN => n9090);
   U4899 : OAI22_X1 port map( A1 => n10774, A2 => n12406, B1 => n10185, B2 => 
                           n12409, ZN => n9089);
   U4900 : OAI22_X1 port map( A1 => n10767, A2 => n12406, B1 => n10153, B2 => 
                           n12409, ZN => n9088);
   U4901 : OAI22_X1 port map( A1 => n10760, A2 => n12406, B1 => n10121, B2 => 
                           n12410, ZN => n9087);
   U4902 : OAI22_X1 port map( A1 => n10753, A2 => n12406, B1 => n10089, B2 => 
                           n12410, ZN => n9086);
   U4903 : OAI22_X1 port map( A1 => n10746, A2 => n12406, B1 => n10057, B2 => 
                           n12410, ZN => n9085);
   U4904 : OAI22_X1 port map( A1 => n10739, A2 => n12406, B1 => n10025, B2 => 
                           n12410, ZN => n9084);
   U4905 : OAI22_X1 port map( A1 => n10732, A2 => n12406, B1 => n9663, B2 => 
                           n12411, ZN => n9083);
   U4906 : OAI22_X1 port map( A1 => n10725, A2 => n12406, B1 => n9631, B2 => 
                           n12411, ZN => n9082);
   U4907 : OAI22_X1 port map( A1 => n10718, A2 => n12406, B1 => n9599, B2 => 
                           n12411, ZN => n9081);
   U4908 : OAI22_X1 port map( A1 => n10711, A2 => n12406, B1 => n9311, B2 => 
                           n12411, ZN => n9080);
   U4909 : OAI22_X1 port map( A1 => n10704, A2 => n12405, B1 => n9201, B2 => 
                           n12412, ZN => n9079);
   U4910 : OAI22_X1 port map( A1 => n10697, A2 => n12405, B1 => n9169, B2 => 
                           n12412, ZN => n9078);
   U4911 : OAI22_X1 port map( A1 => n10690, A2 => n12405, B1 => n9137, B2 => 
                           n12412, ZN => n9077);
   U4912 : OAI22_X1 port map( A1 => n10683, A2 => n12405, B1 => n6002, B2 => 
                           n12412, ZN => n9076);
   U4913 : OAI22_X1 port map( A1 => n10676, A2 => n12405, B1 => n5938, B2 => 
                           n12413, ZN => n9075);
   U4914 : OAI22_X1 port map( A1 => n10669, A2 => n12405, B1 => n5906, B2 => 
                           n12413, ZN => n9074);
   U4915 : OAI22_X1 port map( A1 => n10662, A2 => n12405, B1 => n5874, B2 => 
                           n12413, ZN => n9073);
   U4916 : OAI22_X1 port map( A1 => n10655, A2 => n12405, B1 => n5842, B2 => 
                           n12413, ZN => n9072);
   U4917 : OAI22_X1 port map( A1 => n10648, A2 => n12405, B1 => n5810, B2 => 
                           n12414, ZN => n9071);
   U4918 : OAI22_X1 port map( A1 => n10641, A2 => n12405, B1 => n5778, B2 => 
                           n12414, ZN => n9070);
   U4919 : OAI22_X1 port map( A1 => n10634, A2 => n12405, B1 => n5746, B2 => 
                           n12414, ZN => n9069);
   U4920 : OAI22_X1 port map( A1 => n10627, A2 => n12405, B1 => n5714, B2 => 
                           n12414, ZN => n9068);
   U4921 : OAI22_X1 port map( A1 => n10844, A2 => n12395, B1 => n2849, B2 => 
                           n12396, ZN => n9067);
   U4922 : OAI22_X1 port map( A1 => n10837, A2 => n12394, B1 => n2848, B2 => 
                           n12396, ZN => n9066);
   U4923 : OAI22_X1 port map( A1 => n10830, A2 => n12395, B1 => n2847, B2 => 
                           n12396, ZN => n9065);
   U4924 : OAI22_X1 port map( A1 => n10823, A2 => n12394, B1 => n2846, B2 => 
                           n12396, ZN => n9064);
   U4925 : OAI22_X1 port map( A1 => n10816, A2 => n12395, B1 => n2845, B2 => 
                           n12397, ZN => n9063);
   U4926 : OAI22_X1 port map( A1 => n10809, A2 => n12394, B1 => n2844, B2 => 
                           n12397, ZN => n9062);
   U4927 : OAI22_X1 port map( A1 => n10802, A2 => n12395, B1 => n2843, B2 => 
                           n12397, ZN => n9061);
   U4928 : OAI22_X1 port map( A1 => n10795, A2 => n12394, B1 => n2842, B2 => 
                           n12397, ZN => n9060);
   U4929 : OAI22_X1 port map( A1 => n10788, A2 => n12395, B1 => n2841, B2 => 
                           n12398, ZN => n9059);
   U4930 : OAI22_X1 port map( A1 => n10781, A2 => n12395, B1 => n2840, B2 => 
                           n12398, ZN => n9058);
   U4931 : OAI22_X1 port map( A1 => n10774, A2 => n12395, B1 => n2839, B2 => 
                           n12398, ZN => n9057);
   U4932 : OAI22_X1 port map( A1 => n10767, A2 => n12395, B1 => n2838, B2 => 
                           n12398, ZN => n9056);
   U4933 : OAI22_X1 port map( A1 => n10760, A2 => n12395, B1 => n2837, B2 => 
                           n12399, ZN => n9055);
   U4934 : OAI22_X1 port map( A1 => n10753, A2 => n12395, B1 => n2836, B2 => 
                           n12399, ZN => n9054);
   U4935 : OAI22_X1 port map( A1 => n10746, A2 => n12395, B1 => n2835, B2 => 
                           n12399, ZN => n9053);
   U4936 : OAI22_X1 port map( A1 => n10739, A2 => n12395, B1 => n2834, B2 => 
                           n12399, ZN => n9052);
   U4937 : OAI22_X1 port map( A1 => n10732, A2 => n12395, B1 => n2833, B2 => 
                           n12400, ZN => n9051);
   U4938 : OAI22_X1 port map( A1 => n10725, A2 => n12395, B1 => n2832, B2 => 
                           n12400, ZN => n9050);
   U4939 : OAI22_X1 port map( A1 => n10718, A2 => n12395, B1 => n2831, B2 => 
                           n12400, ZN => n9049);
   U4940 : OAI22_X1 port map( A1 => n10711, A2 => n12395, B1 => n2830, B2 => 
                           n12400, ZN => n9048);
   U4941 : OAI22_X1 port map( A1 => n10704, A2 => n12394, B1 => n2829, B2 => 
                           n12401, ZN => n9047);
   U4942 : OAI22_X1 port map( A1 => n10697, A2 => n12394, B1 => n2828, B2 => 
                           n12401, ZN => n9046);
   U4943 : OAI22_X1 port map( A1 => n10690, A2 => n12394, B1 => n2827, B2 => 
                           n12401, ZN => n9045);
   U4944 : OAI22_X1 port map( A1 => n10683, A2 => n12394, B1 => n2826, B2 => 
                           n12401, ZN => n9044);
   U4945 : OAI22_X1 port map( A1 => n10676, A2 => n12394, B1 => n2825, B2 => 
                           n12402, ZN => n9043);
   U4946 : OAI22_X1 port map( A1 => n10669, A2 => n12394, B1 => n2824, B2 => 
                           n12402, ZN => n9042);
   U4947 : OAI22_X1 port map( A1 => n10662, A2 => n12394, B1 => n2823, B2 => 
                           n12402, ZN => n9041);
   U4948 : OAI22_X1 port map( A1 => n10655, A2 => n12394, B1 => n2822, B2 => 
                           n12402, ZN => n9040);
   U4949 : OAI22_X1 port map( A1 => n10648, A2 => n12394, B1 => n2821, B2 => 
                           n12403, ZN => n9039);
   U4950 : OAI22_X1 port map( A1 => n10641, A2 => n12394, B1 => n2820, B2 => 
                           n12403, ZN => n9038);
   U4951 : OAI22_X1 port map( A1 => n10634, A2 => n12394, B1 => n2819, B2 => 
                           n12403, ZN => n9037);
   U4952 : OAI22_X1 port map( A1 => n10627, A2 => n12394, B1 => n2818, B2 => 
                           n12403, ZN => n9036);
   U4953 : OAI22_X1 port map( A1 => n10844, A2 => n12384, B1 => n10507, B2 => 
                           n12385, ZN => n9035);
   U4954 : OAI22_X1 port map( A1 => n10837, A2 => n12383, B1 => n10475, B2 => 
                           n12385, ZN => n9034);
   U4955 : OAI22_X1 port map( A1 => n10830, A2 => n12384, B1 => n10443, B2 => 
                           n12385, ZN => n9033);
   U4956 : OAI22_X1 port map( A1 => n10823, A2 => n12383, B1 => n10411, B2 => 
                           n12385, ZN => n9032);
   U4957 : OAI22_X1 port map( A1 => n10816, A2 => n12384, B1 => n10376, B2 => 
                           n12386, ZN => n9031);
   U4958 : OAI22_X1 port map( A1 => n10809, A2 => n12383, B1 => n10344, B2 => 
                           n12386, ZN => n9030);
   U4959 : OAI22_X1 port map( A1 => n10802, A2 => n12384, B1 => n10312, B2 => 
                           n12386, ZN => n9029);
   U4960 : OAI22_X1 port map( A1 => n10795, A2 => n12383, B1 => n10277, B2 => 
                           n12386, ZN => n9028);
   U4961 : OAI22_X1 port map( A1 => n10788, A2 => n12384, B1 => n10245, B2 => 
                           n12387, ZN => n9027);
   U4962 : OAI22_X1 port map( A1 => n10781, A2 => n12384, B1 => n10213, B2 => 
                           n12387, ZN => n9026);
   U4963 : OAI22_X1 port map( A1 => n10774, A2 => n12384, B1 => n10179, B2 => 
                           n12387, ZN => n9025);
   U4964 : OAI22_X1 port map( A1 => n10767, A2 => n12384, B1 => n10147, B2 => 
                           n12387, ZN => n9024);
   U4965 : OAI22_X1 port map( A1 => n10760, A2 => n12384, B1 => n10115, B2 => 
                           n12388, ZN => n9023);
   U4966 : OAI22_X1 port map( A1 => n10753, A2 => n12384, B1 => n10083, B2 => 
                           n12388, ZN => n9022);
   U4967 : OAI22_X1 port map( A1 => n10746, A2 => n12384, B1 => n10051, B2 => 
                           n12388, ZN => n9021);
   U4968 : OAI22_X1 port map( A1 => n10739, A2 => n12384, B1 => n10019, B2 => 
                           n12388, ZN => n9020);
   U4969 : OAI22_X1 port map( A1 => n10732, A2 => n12384, B1 => n9657, B2 => 
                           n12389, ZN => n9019);
   U4970 : OAI22_X1 port map( A1 => n10725, A2 => n12384, B1 => n9625, B2 => 
                           n12389, ZN => n9018);
   U4971 : OAI22_X1 port map( A1 => n10718, A2 => n12384, B1 => n9593, B2 => 
                           n12389, ZN => n9017);
   U4972 : OAI22_X1 port map( A1 => n10711, A2 => n12384, B1 => n9259, B2 => 
                           n12389, ZN => n9016);
   U4973 : OAI22_X1 port map( A1 => n10704, A2 => n12383, B1 => n9195, B2 => 
                           n12390, ZN => n9015);
   U4974 : OAI22_X1 port map( A1 => n10697, A2 => n12383, B1 => n9163, B2 => 
                           n12390, ZN => n9014);
   U4975 : OAI22_X1 port map( A1 => n10690, A2 => n12383, B1 => n6313, B2 => 
                           n12390, ZN => n9013);
   U4976 : OAI22_X1 port map( A1 => n10683, A2 => n12383, B1 => n5996, B2 => 
                           n12390, ZN => n9012);
   U4977 : OAI22_X1 port map( A1 => n10676, A2 => n12383, B1 => n5932, B2 => 
                           n12391, ZN => n9011);
   U4978 : OAI22_X1 port map( A1 => n10669, A2 => n12383, B1 => n5900, B2 => 
                           n12391, ZN => n9010);
   U4979 : OAI22_X1 port map( A1 => n10662, A2 => n12383, B1 => n5868, B2 => 
                           n12391, ZN => n9009);
   U4980 : OAI22_X1 port map( A1 => n10655, A2 => n12383, B1 => n5836, B2 => 
                           n12391, ZN => n9008);
   U4981 : OAI22_X1 port map( A1 => n10648, A2 => n12383, B1 => n5804, B2 => 
                           n12392, ZN => n9007);
   U4982 : OAI22_X1 port map( A1 => n10641, A2 => n12383, B1 => n5772, B2 => 
                           n12392, ZN => n9006);
   U4983 : OAI22_X1 port map( A1 => n10634, A2 => n12383, B1 => n5740, B2 => 
                           n12392, ZN => n9005);
   U4984 : OAI22_X1 port map( A1 => n10627, A2 => n12383, B1 => n5708, B2 => 
                           n12392, ZN => n9004);
   U4985 : OAI22_X1 port map( A1 => n10844, A2 => n12373, B1 => n2785, B2 => 
                           n12374, ZN => n9003);
   U4986 : OAI22_X1 port map( A1 => n10837, A2 => n12372, B1 => n2784, B2 => 
                           n12374, ZN => n9002);
   U4987 : OAI22_X1 port map( A1 => n10830, A2 => n12373, B1 => n2783, B2 => 
                           n12374, ZN => n9001);
   U4988 : OAI22_X1 port map( A1 => n10823, A2 => n12372, B1 => n2782, B2 => 
                           n12374, ZN => n9000);
   U4989 : OAI22_X1 port map( A1 => n10816, A2 => n12373, B1 => n2781, B2 => 
                           n12375, ZN => n8999);
   U4990 : OAI22_X1 port map( A1 => n10809, A2 => n12372, B1 => n2780, B2 => 
                           n12375, ZN => n8998);
   U4991 : OAI22_X1 port map( A1 => n10802, A2 => n12373, B1 => n2779, B2 => 
                           n12375, ZN => n8997);
   U4992 : OAI22_X1 port map( A1 => n10795, A2 => n12372, B1 => n2778, B2 => 
                           n12375, ZN => n8996);
   U4993 : OAI22_X1 port map( A1 => n10788, A2 => n12373, B1 => n2777, B2 => 
                           n12376, ZN => n8995);
   U4994 : OAI22_X1 port map( A1 => n10781, A2 => n12373, B1 => n2776, B2 => 
                           n12376, ZN => n8994);
   U4995 : OAI22_X1 port map( A1 => n10774, A2 => n12373, B1 => n2775, B2 => 
                           n12376, ZN => n8993);
   U4996 : OAI22_X1 port map( A1 => n10767, A2 => n12373, B1 => n2774, B2 => 
                           n12376, ZN => n8992);
   U4997 : OAI22_X1 port map( A1 => n10760, A2 => n12373, B1 => n2773, B2 => 
                           n12377, ZN => n8991);
   U4998 : OAI22_X1 port map( A1 => n10753, A2 => n12373, B1 => n2772, B2 => 
                           n12377, ZN => n8990);
   U4999 : OAI22_X1 port map( A1 => n10746, A2 => n12373, B1 => n2771, B2 => 
                           n12377, ZN => n8989);
   U5000 : OAI22_X1 port map( A1 => n10739, A2 => n12373, B1 => n2770, B2 => 
                           n12377, ZN => n8988);
   U5001 : OAI22_X1 port map( A1 => n10732, A2 => n12373, B1 => n2769, B2 => 
                           n12378, ZN => n8987);
   U5002 : OAI22_X1 port map( A1 => n10725, A2 => n12373, B1 => n2768, B2 => 
                           n12378, ZN => n8986);
   U5003 : OAI22_X1 port map( A1 => n10718, A2 => n12373, B1 => n2767, B2 => 
                           n12378, ZN => n8985);
   U5004 : OAI22_X1 port map( A1 => n10711, A2 => n12373, B1 => n2766, B2 => 
                           n12378, ZN => n8984);
   U5005 : OAI22_X1 port map( A1 => n10704, A2 => n12372, B1 => n2765, B2 => 
                           n12379, ZN => n8983);
   U5006 : OAI22_X1 port map( A1 => n10697, A2 => n12372, B1 => n2764, B2 => 
                           n12379, ZN => n8982);
   U5007 : OAI22_X1 port map( A1 => n10690, A2 => n12372, B1 => n2763, B2 => 
                           n12379, ZN => n8981);
   U5008 : OAI22_X1 port map( A1 => n10683, A2 => n12372, B1 => n2762, B2 => 
                           n12379, ZN => n8980);
   U5009 : OAI22_X1 port map( A1 => n10676, A2 => n12372, B1 => n2761, B2 => 
                           n12380, ZN => n8979);
   U5010 : OAI22_X1 port map( A1 => n10669, A2 => n12372, B1 => n2760, B2 => 
                           n12380, ZN => n8978);
   U5011 : OAI22_X1 port map( A1 => n10662, A2 => n12372, B1 => n2759, B2 => 
                           n12380, ZN => n8977);
   U5012 : OAI22_X1 port map( A1 => n10655, A2 => n12372, B1 => n2758, B2 => 
                           n12380, ZN => n8976);
   U5013 : OAI22_X1 port map( A1 => n10648, A2 => n12372, B1 => n2757, B2 => 
                           n12381, ZN => n8975);
   U5014 : OAI22_X1 port map( A1 => n10641, A2 => n12372, B1 => n2756, B2 => 
                           n12381, ZN => n8974);
   U5015 : OAI22_X1 port map( A1 => n10634, A2 => n12372, B1 => n2755, B2 => 
                           n12381, ZN => n8973);
   U5016 : OAI22_X1 port map( A1 => n10627, A2 => n12372, B1 => n2754, B2 => 
                           n12381, ZN => n8972);
   U5017 : OAI22_X1 port map( A1 => n10844, A2 => n12362, B1 => n10506, B2 => 
                           n12363, ZN => n8971);
   U5018 : OAI22_X1 port map( A1 => n10837, A2 => n12361, B1 => n10474, B2 => 
                           n12363, ZN => n8970);
   U5019 : OAI22_X1 port map( A1 => n10830, A2 => n12362, B1 => n10442, B2 => 
                           n12363, ZN => n8969);
   U5020 : OAI22_X1 port map( A1 => n10823, A2 => n12361, B1 => n10410, B2 => 
                           n12363, ZN => n8968);
   U5021 : OAI22_X1 port map( A1 => n10816, A2 => n12362, B1 => n10375, B2 => 
                           n12364, ZN => n8967);
   U5022 : OAI22_X1 port map( A1 => n10809, A2 => n12361, B1 => n10343, B2 => 
                           n12364, ZN => n8966);
   U5023 : OAI22_X1 port map( A1 => n10802, A2 => n12362, B1 => n10311, B2 => 
                           n12364, ZN => n8965);
   U5024 : OAI22_X1 port map( A1 => n10795, A2 => n12361, B1 => n10276, B2 => 
                           n12364, ZN => n8964);
   U5025 : OAI22_X1 port map( A1 => n10788, A2 => n12362, B1 => n10244, B2 => 
                           n12365, ZN => n8963);
   U5026 : OAI22_X1 port map( A1 => n10781, A2 => n12362, B1 => n10212, B2 => 
                           n12365, ZN => n8962);
   U5027 : OAI22_X1 port map( A1 => n10774, A2 => n12362, B1 => n10178, B2 => 
                           n12365, ZN => n8961);
   U5028 : OAI22_X1 port map( A1 => n10767, A2 => n12362, B1 => n10146, B2 => 
                           n12365, ZN => n8960);
   U5029 : OAI22_X1 port map( A1 => n10760, A2 => n12362, B1 => n10114, B2 => 
                           n12366, ZN => n8959);
   U5030 : OAI22_X1 port map( A1 => n10753, A2 => n12362, B1 => n10082, B2 => 
                           n12366, ZN => n8958);
   U5031 : OAI22_X1 port map( A1 => n10746, A2 => n12362, B1 => n10050, B2 => 
                           n12366, ZN => n8957);
   U5032 : OAI22_X1 port map( A1 => n10739, A2 => n12362, B1 => n10018, B2 => 
                           n12366, ZN => n8956);
   U5033 : OAI22_X1 port map( A1 => n10732, A2 => n12362, B1 => n9656, B2 => 
                           n12367, ZN => n8955);
   U5034 : OAI22_X1 port map( A1 => n10725, A2 => n12362, B1 => n9624, B2 => 
                           n12367, ZN => n8954);
   U5035 : OAI22_X1 port map( A1 => n10718, A2 => n12362, B1 => n9592, B2 => 
                           n12367, ZN => n8953);
   U5036 : OAI22_X1 port map( A1 => n10711, A2 => n12362, B1 => n9258, B2 => 
                           n12367, ZN => n8952);
   U5037 : OAI22_X1 port map( A1 => n10704, A2 => n12361, B1 => n9194, B2 => 
                           n12368, ZN => n8951);
   U5038 : OAI22_X1 port map( A1 => n10697, A2 => n12361, B1 => n9162, B2 => 
                           n12368, ZN => n8950);
   U5039 : OAI22_X1 port map( A1 => n10690, A2 => n12361, B1 => n6312, B2 => 
                           n12368, ZN => n8949);
   U5040 : OAI22_X1 port map( A1 => n10683, A2 => n12361, B1 => n5995, B2 => 
                           n12368, ZN => n8948);
   U5041 : OAI22_X1 port map( A1 => n10676, A2 => n12361, B1 => n5931, B2 => 
                           n12369, ZN => n8947);
   U5042 : OAI22_X1 port map( A1 => n10669, A2 => n12361, B1 => n5899, B2 => 
                           n12369, ZN => n8946);
   U5043 : OAI22_X1 port map( A1 => n10662, A2 => n12361, B1 => n5867, B2 => 
                           n12369, ZN => n8945);
   U5044 : OAI22_X1 port map( A1 => n10655, A2 => n12361, B1 => n5835, B2 => 
                           n12369, ZN => n8944);
   U5045 : OAI22_X1 port map( A1 => n10648, A2 => n12361, B1 => n5803, B2 => 
                           n12370, ZN => n8943);
   U5046 : OAI22_X1 port map( A1 => n10641, A2 => n12361, B1 => n5771, B2 => 
                           n12370, ZN => n8942);
   U5047 : OAI22_X1 port map( A1 => n10634, A2 => n12361, B1 => n5739, B2 => 
                           n12370, ZN => n8941);
   U5048 : OAI22_X1 port map( A1 => n10627, A2 => n12361, B1 => n5707, B2 => 
                           n12370, ZN => n8940);
   U5049 : OAI22_X1 port map( A1 => n10844, A2 => n12351, B1 => n10508, B2 => 
                           n12352, ZN => n8939);
   U5050 : OAI22_X1 port map( A1 => n10837, A2 => n12350, B1 => n10476, B2 => 
                           n12352, ZN => n8938);
   U5051 : OAI22_X1 port map( A1 => n10830, A2 => n12351, B1 => n10444, B2 => 
                           n12352, ZN => n8937);
   U5052 : OAI22_X1 port map( A1 => n10823, A2 => n12350, B1 => n10412, B2 => 
                           n12352, ZN => n8936);
   U5053 : OAI22_X1 port map( A1 => n10816, A2 => n12351, B1 => n10377, B2 => 
                           n12353, ZN => n8935);
   U5054 : OAI22_X1 port map( A1 => n10809, A2 => n12350, B1 => n10345, B2 => 
                           n12353, ZN => n8934);
   U5055 : OAI22_X1 port map( A1 => n10802, A2 => n12351, B1 => n10313, B2 => 
                           n12353, ZN => n8933);
   U5056 : OAI22_X1 port map( A1 => n10795, A2 => n12350, B1 => n10278, B2 => 
                           n12353, ZN => n8932);
   U5057 : OAI22_X1 port map( A1 => n10788, A2 => n12351, B1 => n10246, B2 => 
                           n12354, ZN => n8931);
   U5058 : OAI22_X1 port map( A1 => n10781, A2 => n12351, B1 => n10214, B2 => 
                           n12354, ZN => n8930);
   U5059 : OAI22_X1 port map( A1 => n10774, A2 => n12351, B1 => n10180, B2 => 
                           n12354, ZN => n8929);
   U5060 : OAI22_X1 port map( A1 => n10767, A2 => n12351, B1 => n10148, B2 => 
                           n12354, ZN => n8928);
   U5061 : OAI22_X1 port map( A1 => n10760, A2 => n12351, B1 => n10116, B2 => 
                           n12355, ZN => n8927);
   U5062 : OAI22_X1 port map( A1 => n10753, A2 => n12351, B1 => n10084, B2 => 
                           n12355, ZN => n8926);
   U5063 : OAI22_X1 port map( A1 => n10746, A2 => n12351, B1 => n10052, B2 => 
                           n12355, ZN => n8925);
   U5064 : OAI22_X1 port map( A1 => n10739, A2 => n12351, B1 => n10020, B2 => 
                           n12355, ZN => n8924);
   U5065 : OAI22_X1 port map( A1 => n10732, A2 => n12351, B1 => n9658, B2 => 
                           n12356, ZN => n8923);
   U5066 : OAI22_X1 port map( A1 => n10725, A2 => n12351, B1 => n9626, B2 => 
                           n12356, ZN => n8922);
   U5067 : OAI22_X1 port map( A1 => n10718, A2 => n12351, B1 => n9594, B2 => 
                           n12356, ZN => n8921);
   U5068 : OAI22_X1 port map( A1 => n10711, A2 => n12351, B1 => n9260, B2 => 
                           n12356, ZN => n8920);
   U5069 : OAI22_X1 port map( A1 => n10704, A2 => n12350, B1 => n9196, B2 => 
                           n12357, ZN => n8919);
   U5070 : OAI22_X1 port map( A1 => n10697, A2 => n12350, B1 => n9164, B2 => 
                           n12357, ZN => n8918);
   U5071 : OAI22_X1 port map( A1 => n10690, A2 => n12350, B1 => n6314, B2 => 
                           n12357, ZN => n8917);
   U5072 : OAI22_X1 port map( A1 => n10683, A2 => n12350, B1 => n5997, B2 => 
                           n12357, ZN => n8916);
   U5073 : OAI22_X1 port map( A1 => n10676, A2 => n12350, B1 => n5933, B2 => 
                           n12358, ZN => n8915);
   U5074 : OAI22_X1 port map( A1 => n10669, A2 => n12350, B1 => n5901, B2 => 
                           n12358, ZN => n8914);
   U5075 : OAI22_X1 port map( A1 => n10662, A2 => n12350, B1 => n5869, B2 => 
                           n12358, ZN => n8913);
   U5076 : OAI22_X1 port map( A1 => n10655, A2 => n12350, B1 => n5837, B2 => 
                           n12358, ZN => n8912);
   U5077 : OAI22_X1 port map( A1 => n10648, A2 => n12350, B1 => n5805, B2 => 
                           n12359, ZN => n8911);
   U5078 : OAI22_X1 port map( A1 => n10641, A2 => n12350, B1 => n5773, B2 => 
                           n12359, ZN => n8910);
   U5079 : OAI22_X1 port map( A1 => n10634, A2 => n12350, B1 => n5741, B2 => 
                           n12359, ZN => n8909);
   U5080 : OAI22_X1 port map( A1 => n10627, A2 => n12350, B1 => n5709, B2 => 
                           n12359, ZN => n8908);
   U5081 : OAI22_X1 port map( A1 => n10844, A2 => n12305, B1 => n10512, B2 => 
                           n12306, ZN => n8811);
   U5082 : OAI22_X1 port map( A1 => n10837, A2 => n12305, B1 => n10480, B2 => 
                           n12306, ZN => n8810);
   U5083 : OAI22_X1 port map( A1 => n10830, A2 => n12305, B1 => n10448, B2 => 
                           n12306, ZN => n8809);
   U5084 : OAI22_X1 port map( A1 => n10823, A2 => n12305, B1 => n10416, B2 => 
                           n12306, ZN => n8808);
   U5085 : OAI22_X1 port map( A1 => n10816, A2 => n12305, B1 => n10381, B2 => 
                           n12307, ZN => n8807);
   U5086 : OAI22_X1 port map( A1 => n10809, A2 => n12305, B1 => n10349, B2 => 
                           n12307, ZN => n8806);
   U5087 : OAI22_X1 port map( A1 => n10802, A2 => n12305, B1 => n10317, B2 => 
                           n12307, ZN => n8805);
   U5088 : OAI22_X1 port map( A1 => n10795, A2 => n12305, B1 => n10282, B2 => 
                           n12307, ZN => n8804);
   U5089 : OAI22_X1 port map( A1 => n10788, A2 => n12304, B1 => n10250, B2 => 
                           n12308, ZN => n8803);
   U5090 : OAI22_X1 port map( A1 => n10781, A2 => n12304, B1 => n10218, B2 => 
                           n12308, ZN => n8802);
   U5091 : OAI22_X1 port map( A1 => n10774, A2 => n12304, B1 => n10184, B2 => 
                           n12308, ZN => n8801);
   U5092 : OAI22_X1 port map( A1 => n10767, A2 => n12304, B1 => n10152, B2 => 
                           n12308, ZN => n8800);
   U5093 : OAI22_X1 port map( A1 => n10760, A2 => n12304, B1 => n10120, B2 => 
                           n12309, ZN => n8799);
   U5094 : OAI22_X1 port map( A1 => n10753, A2 => n12304, B1 => n10088, B2 => 
                           n12309, ZN => n8798);
   U5095 : OAI22_X1 port map( A1 => n10746, A2 => n12304, B1 => n10056, B2 => 
                           n12309, ZN => n8797);
   U5096 : OAI22_X1 port map( A1 => n10739, A2 => n12304, B1 => n10024, B2 => 
                           n12309, ZN => n8796);
   U5097 : OAI22_X1 port map( A1 => n10732, A2 => n12304, B1 => n9662, B2 => 
                           n12310, ZN => n8795);
   U5098 : OAI22_X1 port map( A1 => n10725, A2 => n12304, B1 => n9630, B2 => 
                           n12310, ZN => n8794);
   U5099 : OAI22_X1 port map( A1 => n10718, A2 => n12304, B1 => n9598, B2 => 
                           n12310, ZN => n8793);
   U5100 : OAI22_X1 port map( A1 => n10711, A2 => n12304, B1 => n9264, B2 => 
                           n12310, ZN => n8792);
   U5101 : OAI22_X1 port map( A1 => n10704, A2 => n12303, B1 => n9200, B2 => 
                           n12311, ZN => n8791);
   U5102 : OAI22_X1 port map( A1 => n10697, A2 => n12303, B1 => n9168, B2 => 
                           n12311, ZN => n8790);
   U5103 : OAI22_X1 port map( A1 => n10690, A2 => n12303, B1 => n9136, B2 => 
                           n12311, ZN => n8789);
   U5104 : OAI22_X1 port map( A1 => n10683, A2 => n12303, B1 => n6001, B2 => 
                           n12311, ZN => n8788);
   U5105 : OAI22_X1 port map( A1 => n10676, A2 => n12303, B1 => n5937, B2 => 
                           n12312, ZN => n8787);
   U5106 : OAI22_X1 port map( A1 => n10669, A2 => n12303, B1 => n5905, B2 => 
                           n12312, ZN => n8786);
   U5107 : OAI22_X1 port map( A1 => n10662, A2 => n12303, B1 => n5873, B2 => 
                           n12312, ZN => n8785);
   U5108 : OAI22_X1 port map( A1 => n10655, A2 => n12303, B1 => n5841, B2 => 
                           n12312, ZN => n8784);
   U5109 : OAI22_X1 port map( A1 => n10648, A2 => n12303, B1 => n5809, B2 => 
                           n12313, ZN => n8783);
   U5110 : OAI22_X1 port map( A1 => n10641, A2 => n12303, B1 => n5777, B2 => 
                           n12313, ZN => n8782);
   U5111 : OAI22_X1 port map( A1 => n10634, A2 => n12303, B1 => n5745, B2 => 
                           n12313, ZN => n8781);
   U5112 : OAI22_X1 port map( A1 => n10627, A2 => n12303, B1 => n5713, B2 => 
                           n12313, ZN => n8780);
   U5113 : OAI22_X1 port map( A1 => n10846, A2 => n12017, B1 => n993, B2 => 
                           n12018, ZN => n8043);
   U5114 : OAI22_X1 port map( A1 => n10839, A2 => n12017, B1 => n989, B2 => 
                           n12018, ZN => n8042);
   U5115 : OAI22_X1 port map( A1 => n10832, A2 => n12017, B1 => n985, B2 => 
                           n12018, ZN => n8041);
   U5116 : OAI22_X1 port map( A1 => n10825, A2 => n12017, B1 => n981, B2 => 
                           n12018, ZN => n8040);
   U5117 : OAI22_X1 port map( A1 => n10818, A2 => n12017, B1 => n977, B2 => 
                           n12019, ZN => n8039);
   U5118 : OAI22_X1 port map( A1 => n10811, A2 => n12017, B1 => n973, B2 => 
                           n12019, ZN => n8038);
   U5119 : OAI22_X1 port map( A1 => n10804, A2 => n12017, B1 => n969, B2 => 
                           n12019, ZN => n8037);
   U5120 : OAI22_X1 port map( A1 => n10797, A2 => n12017, B1 => n965, B2 => 
                           n12019, ZN => n8036);
   U5121 : OAI22_X1 port map( A1 => n10790, A2 => n12016, B1 => n961, B2 => 
                           n12020, ZN => n8035);
   U5122 : OAI22_X1 port map( A1 => n10783, A2 => n12016, B1 => n957, B2 => 
                           n12020, ZN => n8034);
   U5123 : OAI22_X1 port map( A1 => n10776, A2 => n12016, B1 => n953, B2 => 
                           n12020, ZN => n8033);
   U5124 : OAI22_X1 port map( A1 => n10769, A2 => n12016, B1 => n949, B2 => 
                           n12020, ZN => n8032);
   U5125 : OAI22_X1 port map( A1 => n10762, A2 => n12016, B1 => n945, B2 => 
                           n12021, ZN => n8031);
   U5126 : OAI22_X1 port map( A1 => n10755, A2 => n12016, B1 => n941, B2 => 
                           n12021, ZN => n8030);
   U5127 : OAI22_X1 port map( A1 => n10748, A2 => n12016, B1 => n937, B2 => 
                           n12021, ZN => n8029);
   U5128 : OAI22_X1 port map( A1 => n10741, A2 => n12016, B1 => n933, B2 => 
                           n12021, ZN => n8028);
   U5129 : OAI22_X1 port map( A1 => n10734, A2 => n12016, B1 => n929, B2 => 
                           n12022, ZN => n8027);
   U5130 : OAI22_X1 port map( A1 => n10629, A2 => n12003, B1 => n999, B2 => 
                           n12006, ZN => n7980);
   U5131 : OAI22_X1 port map( A1 => n10848, A2 => n11753, B1 => n994, B2 => 
                           n11754, ZN => n7339);
   U5132 : OAI22_X1 port map( A1 => n10841, A2 => n11753, B1 => n990, B2 => 
                           n11754, ZN => n7338);
   U5133 : OAI22_X1 port map( A1 => n10834, A2 => n11753, B1 => n986, B2 => 
                           n11754, ZN => n7337);
   U5134 : OAI22_X1 port map( A1 => n10827, A2 => n11753, B1 => n982, B2 => 
                           n11754, ZN => n7336);
   U5135 : OAI22_X1 port map( A1 => n10820, A2 => n11753, B1 => n978, B2 => 
                           n11755, ZN => n7335);
   U5136 : OAI22_X1 port map( A1 => n10813, A2 => n11753, B1 => n974, B2 => 
                           n11755, ZN => n7334);
   U5137 : OAI22_X1 port map( A1 => n10737, A2 => n11644, B1 => n2048, B2 => 
                           n11646, ZN => n7035);
   U5138 : OAI22_X1 port map( A1 => n10730, A2 => n11644, B1 => n2036, B2 => 
                           n11646, ZN => n7034);
   U5139 : OAI22_X1 port map( A1 => n10723, A2 => n11644, B1 => n2024, B2 => 
                           n11646, ZN => n7033);
   U5140 : OAI22_X1 port map( A1 => n10716, A2 => n11644, B1 => n2012, B2 => 
                           n11646, ZN => n7032);
   U5141 : OAI22_X1 port map( A1 => n10709, A2 => n11643, B1 => n2000, B2 => 
                           n11647, ZN => n7031);
   U5142 : OAI22_X1 port map( A1 => n10702, A2 => n11643, B1 => n1988, B2 => 
                           n11647, ZN => n7030);
   U5143 : OAI22_X1 port map( A1 => n10695, A2 => n11643, B1 => n1976, B2 => 
                           n11647, ZN => n7029);
   U5144 : OAI22_X1 port map( A1 => n10688, A2 => n11643, B1 => n1964, B2 => 
                           n11647, ZN => n7028);
   U5145 : OAI22_X1 port map( A1 => n10681, A2 => n11643, B1 => n1952, B2 => 
                           n11648, ZN => n7027);
   U5146 : OAI22_X1 port map( A1 => n10674, A2 => n11643, B1 => n1940, B2 => 
                           n11648, ZN => n7026);
   U5147 : OAI22_X1 port map( A1 => n10667, A2 => n11643, B1 => n1928, B2 => 
                           n11648, ZN => n7025);
   U5148 : OAI22_X1 port map( A1 => n10660, A2 => n11643, B1 => n1916, B2 => 
                           n11648, ZN => n7024);
   U5149 : OAI22_X1 port map( A1 => n10653, A2 => n11643, B1 => n1904, B2 => 
                           n11649, ZN => n7023);
   U5150 : OAI22_X1 port map( A1 => n10646, A2 => n11643, B1 => n1892, B2 => 
                           n11649, ZN => n7022);
   U5151 : OAI22_X1 port map( A1 => n10639, A2 => n11643, B1 => n1880, B2 => 
                           n11649, ZN => n7021);
   U5152 : OAI22_X1 port map( A1 => n10632, A2 => n11643, B1 => n1868, B2 => 
                           n11649, ZN => n7020);
   U5153 : OAI22_X1 port map( A1 => n10849, A2 => n11633, B1 => n801, B2 => 
                           n11634, ZN => n7019);
   U5154 : OAI22_X1 port map( A1 => n10842, A2 => n11633, B1 => n800, B2 => 
                           n11634, ZN => n7018);
   U5155 : OAI22_X1 port map( A1 => n10835, A2 => n11633, B1 => n799, B2 => 
                           n11634, ZN => n7017);
   U5156 : OAI22_X1 port map( A1 => n10828, A2 => n11633, B1 => n798, B2 => 
                           n11634, ZN => n7016);
   U5157 : OAI22_X1 port map( A1 => n10821, A2 => n11633, B1 => n797, B2 => 
                           n11635, ZN => n7015);
   U5158 : OAI22_X1 port map( A1 => n10814, A2 => n11633, B1 => n796, B2 => 
                           n11635, ZN => n7014);
   U5159 : OAI22_X1 port map( A1 => n10807, A2 => n11633, B1 => n795, B2 => 
                           n11635, ZN => n7013);
   U5160 : OAI22_X1 port map( A1 => n10800, A2 => n11633, B1 => n794, B2 => 
                           n11635, ZN => n7012);
   U5161 : OAI22_X1 port map( A1 => n10793, A2 => n11632, B1 => n793, B2 => 
                           n11636, ZN => n7011);
   U5162 : OAI22_X1 port map( A1 => n10786, A2 => n11632, B1 => n792, B2 => 
                           n11636, ZN => n7010);
   U5163 : OAI22_X1 port map( A1 => n10779, A2 => n11632, B1 => n791, B2 => 
                           n11636, ZN => n7009);
   U5164 : OAI22_X1 port map( A1 => n10772, A2 => n11632, B1 => n790, B2 => 
                           n11636, ZN => n7008);
   U5165 : OAI22_X1 port map( A1 => n10765, A2 => n11632, B1 => n789, B2 => 
                           n11637, ZN => n7007);
   U5166 : OAI22_X1 port map( A1 => n10758, A2 => n11632, B1 => n788, B2 => 
                           n11637, ZN => n7006);
   U5167 : OAI22_X1 port map( A1 => n10751, A2 => n11632, B1 => n787, B2 => 
                           n11637, ZN => n7005);
   U5168 : OAI22_X1 port map( A1 => n10744, A2 => n11632, B1 => n786, B2 => 
                           n11637, ZN => n7004);
   U5169 : OAI22_X1 port map( A1 => n10737, A2 => n11632, B1 => n785, B2 => 
                           n11638, ZN => n7003);
   U5170 : OAI22_X1 port map( A1 => n10730, A2 => n11632, B1 => n784, B2 => 
                           n11638, ZN => n7002);
   U5171 : OAI22_X1 port map( A1 => n10723, A2 => n11632, B1 => n783, B2 => 
                           n11638, ZN => n7001);
   U5172 : OAI22_X1 port map( A1 => n10716, A2 => n11632, B1 => n782, B2 => 
                           n11638, ZN => n7000);
   U5173 : OAI22_X1 port map( A1 => n10709, A2 => n11631, B1 => n781, B2 => 
                           n11639, ZN => n6999);
   U5174 : OAI22_X1 port map( A1 => n10702, A2 => n11631, B1 => n780, B2 => 
                           n11639, ZN => n6998);
   U5175 : OAI22_X1 port map( A1 => n10695, A2 => n11631, B1 => n779, B2 => 
                           n11639, ZN => n6997);
   U5176 : OAI22_X1 port map( A1 => n10688, A2 => n11631, B1 => n778, B2 => 
                           n11639, ZN => n6996);
   U5177 : OAI22_X1 port map( A1 => n10681, A2 => n11631, B1 => n777, B2 => 
                           n11640, ZN => n6995);
   U5178 : OAI22_X1 port map( A1 => n10674, A2 => n11631, B1 => n776, B2 => 
                           n11640, ZN => n6994);
   U5179 : OAI22_X1 port map( A1 => n10667, A2 => n11631, B1 => n775, B2 => 
                           n11640, ZN => n6993);
   U5180 : OAI22_X1 port map( A1 => n10660, A2 => n11631, B1 => n774, B2 => 
                           n11640, ZN => n6992);
   U5181 : OAI22_X1 port map( A1 => n10653, A2 => n11631, B1 => n773, B2 => 
                           n11641, ZN => n6991);
   U5182 : OAI22_X1 port map( A1 => n10646, A2 => n11631, B1 => n772, B2 => 
                           n11641, ZN => n6990);
   U5183 : OAI22_X1 port map( A1 => n10639, A2 => n11631, B1 => n771, B2 => 
                           n11641, ZN => n6989);
   U5184 : OAI22_X1 port map( A1 => n10632, A2 => n11631, B1 => n770, B2 => 
                           n11641, ZN => n6988);
   U5185 : OAI22_X1 port map( A1 => n10849, A2 => n11621, B1 => n10537, B2 => 
                           n11622, ZN => n6987);
   U5186 : OAI22_X1 port map( A1 => n10842, A2 => n11621, B1 => n10505, B2 => 
                           n11622, ZN => n6986);
   U5187 : OAI22_X1 port map( A1 => n10835, A2 => n11621, B1 => n10473, B2 => 
                           n11622, ZN => n6985);
   U5188 : OAI22_X1 port map( A1 => n10828, A2 => n11621, B1 => n10441, B2 => 
                           n11622, ZN => n6984);
   U5189 : OAI22_X1 port map( A1 => n10821, A2 => n11621, B1 => n10409, B2 => 
                           n11623, ZN => n6983);
   U5190 : OAI22_X1 port map( A1 => n10814, A2 => n11621, B1 => n10374, B2 => 
                           n11623, ZN => n6982);
   U5191 : OAI22_X1 port map( A1 => n10807, A2 => n11621, B1 => n10342, B2 => 
                           n11623, ZN => n6981);
   U5192 : OAI22_X1 port map( A1 => n10800, A2 => n11621, B1 => n10310, B2 => 
                           n11623, ZN => n6980);
   U5193 : OAI22_X1 port map( A1 => n10793, A2 => n11620, B1 => n10275, B2 => 
                           n11624, ZN => n6979);
   U5194 : OAI22_X1 port map( A1 => n10786, A2 => n11620, B1 => n10243, B2 => 
                           n11624, ZN => n6978);
   U5195 : OAI22_X1 port map( A1 => n10779, A2 => n11620, B1 => n10211, B2 => 
                           n11624, ZN => n6977);
   U5196 : OAI22_X1 port map( A1 => n10772, A2 => n11620, B1 => n10177, B2 => 
                           n11624, ZN => n6976);
   U5197 : OAI22_X1 port map( A1 => n10765, A2 => n11620, B1 => n10145, B2 => 
                           n11625, ZN => n6975);
   U5198 : OAI22_X1 port map( A1 => n10758, A2 => n11620, B1 => n10113, B2 => 
                           n11625, ZN => n6974);
   U5199 : OAI22_X1 port map( A1 => n10751, A2 => n11620, B1 => n10081, B2 => 
                           n11625, ZN => n6973);
   U5200 : OAI22_X1 port map( A1 => n10744, A2 => n11620, B1 => n10049, B2 => 
                           n11625, ZN => n6972);
   U5201 : OAI22_X1 port map( A1 => n10737, A2 => n11620, B1 => n10017, B2 => 
                           n11626, ZN => n6971);
   U5202 : OAI22_X1 port map( A1 => n10730, A2 => n11620, B1 => n9655, B2 => 
                           n11626, ZN => n6970);
   U5203 : OAI22_X1 port map( A1 => n10723, A2 => n11620, B1 => n9623, B2 => 
                           n11626, ZN => n6969);
   U5204 : OAI22_X1 port map( A1 => n10716, A2 => n11620, B1 => n9591, B2 => 
                           n11626, ZN => n6968);
   U5205 : OAI22_X1 port map( A1 => n10709, A2 => n11619, B1 => n9257, B2 => 
                           n11627, ZN => n6967);
   U5206 : OAI22_X1 port map( A1 => n10702, A2 => n11619, B1 => n9193, B2 => 
                           n11627, ZN => n6966);
   U5207 : OAI22_X1 port map( A1 => n10695, A2 => n11619, B1 => n9161, B2 => 
                           n11627, ZN => n6965);
   U5208 : OAI22_X1 port map( A1 => n10688, A2 => n11619, B1 => n6311, B2 => 
                           n11627, ZN => n6964);
   U5209 : OAI22_X1 port map( A1 => n10681, A2 => n11619, B1 => n5994, B2 => 
                           n11628, ZN => n6963);
   U5210 : OAI22_X1 port map( A1 => n10674, A2 => n11619, B1 => n5930, B2 => 
                           n11628, ZN => n6962);
   U5211 : OAI22_X1 port map( A1 => n10667, A2 => n11619, B1 => n5898, B2 => 
                           n11628, ZN => n6961);
   U5212 : OAI22_X1 port map( A1 => n10660, A2 => n11619, B1 => n5866, B2 => 
                           n11628, ZN => n6960);
   U5213 : OAI22_X1 port map( A1 => n10653, A2 => n11619, B1 => n5834, B2 => 
                           n11629, ZN => n6959);
   U5214 : OAI22_X1 port map( A1 => n10646, A2 => n11619, B1 => n5802, B2 => 
                           n11629, ZN => n6958);
   U5215 : OAI22_X1 port map( A1 => n10639, A2 => n11619, B1 => n5770, B2 => 
                           n11629, ZN => n6957);
   U5216 : OAI22_X1 port map( A1 => n10632, A2 => n11619, B1 => n5738, B2 => 
                           n11629, ZN => n6956);
   U5217 : OAI22_X1 port map( A1 => n10849, A2 => n11609, B1 => n737, B2 => 
                           n11610, ZN => n6955);
   U5218 : OAI22_X1 port map( A1 => n10842, A2 => n11609, B1 => n736, B2 => 
                           n11610, ZN => n6954);
   U5219 : OAI22_X1 port map( A1 => n10835, A2 => n11609, B1 => n735, B2 => 
                           n11610, ZN => n6953);
   U5220 : OAI22_X1 port map( A1 => n10828, A2 => n11609, B1 => n734, B2 => 
                           n11610, ZN => n6952);
   U5221 : OAI22_X1 port map( A1 => n10821, A2 => n11609, B1 => n733, B2 => 
                           n11611, ZN => n6951);
   U5222 : OAI22_X1 port map( A1 => n10814, A2 => n11609, B1 => n732, B2 => 
                           n11611, ZN => n6950);
   U5223 : OAI22_X1 port map( A1 => n10807, A2 => n11609, B1 => n731, B2 => 
                           n11611, ZN => n6949);
   U5224 : OAI22_X1 port map( A1 => n10800, A2 => n11609, B1 => n730, B2 => 
                           n11611, ZN => n6948);
   U5225 : OAI22_X1 port map( A1 => n10793, A2 => n11608, B1 => n729, B2 => 
                           n11612, ZN => n6947);
   U5226 : OAI22_X1 port map( A1 => n10786, A2 => n11608, B1 => n728, B2 => 
                           n11612, ZN => n6946);
   U5227 : OAI22_X1 port map( A1 => n10779, A2 => n11608, B1 => n727, B2 => 
                           n11612, ZN => n6945);
   U5228 : OAI22_X1 port map( A1 => n10772, A2 => n11608, B1 => n726, B2 => 
                           n11612, ZN => n6944);
   U5229 : OAI22_X1 port map( A1 => n10765, A2 => n11608, B1 => n725, B2 => 
                           n11613, ZN => n6943);
   U5230 : OAI22_X1 port map( A1 => n10758, A2 => n11608, B1 => n724, B2 => 
                           n11613, ZN => n6942);
   U5231 : OAI22_X1 port map( A1 => n10751, A2 => n11608, B1 => n723, B2 => 
                           n11613, ZN => n6941);
   U5232 : OAI22_X1 port map( A1 => n10744, A2 => n11608, B1 => n722, B2 => 
                           n11613, ZN => n6940);
   U5233 : OAI22_X1 port map( A1 => n10737, A2 => n11608, B1 => n721, B2 => 
                           n11614, ZN => n6939);
   U5234 : OAI22_X1 port map( A1 => n10730, A2 => n11608, B1 => n720, B2 => 
                           n11614, ZN => n6938);
   U5235 : OAI22_X1 port map( A1 => n10723, A2 => n11608, B1 => n719, B2 => 
                           n11614, ZN => n6937);
   U5236 : OAI22_X1 port map( A1 => n10716, A2 => n11608, B1 => n718, B2 => 
                           n11614, ZN => n6936);
   U5237 : OAI22_X1 port map( A1 => n10709, A2 => n11607, B1 => n717, B2 => 
                           n11615, ZN => n6935);
   U5238 : OAI22_X1 port map( A1 => n10702, A2 => n11607, B1 => n716, B2 => 
                           n11615, ZN => n6934);
   U5239 : OAI22_X1 port map( A1 => n10695, A2 => n11607, B1 => n715, B2 => 
                           n11615, ZN => n6933);
   U5240 : OAI22_X1 port map( A1 => n10688, A2 => n11607, B1 => n714, B2 => 
                           n11615, ZN => n6932);
   U5241 : OAI22_X1 port map( A1 => n10681, A2 => n11607, B1 => n713, B2 => 
                           n11616, ZN => n6931);
   U5242 : OAI22_X1 port map( A1 => n10674, A2 => n11607, B1 => n712, B2 => 
                           n11616, ZN => n6930);
   U5243 : OAI22_X1 port map( A1 => n10667, A2 => n11607, B1 => n711, B2 => 
                           n11616, ZN => n6929);
   U5244 : OAI22_X1 port map( A1 => n10660, A2 => n11607, B1 => n710, B2 => 
                           n11616, ZN => n6928);
   U5245 : OAI22_X1 port map( A1 => n10653, A2 => n11607, B1 => n709, B2 => 
                           n11617, ZN => n6927);
   U5246 : OAI22_X1 port map( A1 => n10646, A2 => n11607, B1 => n708, B2 => 
                           n11617, ZN => n6926);
   U5247 : OAI22_X1 port map( A1 => n10639, A2 => n11607, B1 => n707, B2 => 
                           n11617, ZN => n6925);
   U5248 : OAI22_X1 port map( A1 => n10632, A2 => n11607, B1 => n706, B2 => 
                           n11617, ZN => n6924);
   U5249 : OAI22_X1 port map( A1 => n10849, A2 => n11597, B1 => n10531, B2 => 
                           n11598, ZN => n6923);
   U5250 : OAI22_X1 port map( A1 => n10842, A2 => n11597, B1 => n10499, B2 => 
                           n11598, ZN => n6922);
   U5251 : OAI22_X1 port map( A1 => n10835, A2 => n11597, B1 => n10467, B2 => 
                           n11598, ZN => n6921);
   U5252 : OAI22_X1 port map( A1 => n10828, A2 => n11597, B1 => n10435, B2 => 
                           n11598, ZN => n6920);
   U5253 : OAI22_X1 port map( A1 => n10821, A2 => n11597, B1 => n10403, B2 => 
                           n11599, ZN => n6919);
   U5254 : OAI22_X1 port map( A1 => n10814, A2 => n11597, B1 => n10368, B2 => 
                           n11599, ZN => n6918);
   U5255 : OAI22_X1 port map( A1 => n10807, A2 => n11597, B1 => n10336, B2 => 
                           n11599, ZN => n6917);
   U5256 : OAI22_X1 port map( A1 => n10800, A2 => n11597, B1 => n10304, B2 => 
                           n11599, ZN => n6916);
   U5257 : OAI22_X1 port map( A1 => n10793, A2 => n11596, B1 => n10269, B2 => 
                           n11600, ZN => n6915);
   U5258 : OAI22_X1 port map( A1 => n10786, A2 => n11596, B1 => n10237, B2 => 
                           n11600, ZN => n6914);
   U5259 : OAI22_X1 port map( A1 => n10779, A2 => n11596, B1 => n10203, B2 => 
                           n11600, ZN => n6913);
   U5260 : OAI22_X1 port map( A1 => n10772, A2 => n11596, B1 => n10171, B2 => 
                           n11600, ZN => n6912);
   U5261 : OAI22_X1 port map( A1 => n10765, A2 => n11596, B1 => n10139, B2 => 
                           n11601, ZN => n6911);
   U5262 : OAI22_X1 port map( A1 => n10758, A2 => n11596, B1 => n10107, B2 => 
                           n11601, ZN => n6910);
   U5263 : OAI22_X1 port map( A1 => n10751, A2 => n11596, B1 => n10075, B2 => 
                           n11601, ZN => n6909);
   U5264 : OAI22_X1 port map( A1 => n10744, A2 => n11596, B1 => n10043, B2 => 
                           n11601, ZN => n6908);
   U5265 : OAI22_X1 port map( A1 => n10737, A2 => n11596, B1 => n10011, B2 => 
                           n11602, ZN => n6907);
   U5266 : OAI22_X1 port map( A1 => n10730, A2 => n11596, B1 => n9649, B2 => 
                           n11602, ZN => n6906);
   U5267 : OAI22_X1 port map( A1 => n10723, A2 => n11596, B1 => n9617, B2 => 
                           n11602, ZN => n6905);
   U5268 : OAI22_X1 port map( A1 => n10716, A2 => n11596, B1 => n9585, B2 => 
                           n11602, ZN => n6904);
   U5269 : OAI22_X1 port map( A1 => n10709, A2 => n11595, B1 => n9251, B2 => 
                           n11603, ZN => n6903);
   U5270 : OAI22_X1 port map( A1 => n10702, A2 => n11595, B1 => n9187, B2 => 
                           n11603, ZN => n6902);
   U5271 : OAI22_X1 port map( A1 => n10695, A2 => n11595, B1 => n9155, B2 => 
                           n11603, ZN => n6901);
   U5272 : OAI22_X1 port map( A1 => n10688, A2 => n11595, B1 => n6305, B2 => 
                           n11603, ZN => n6900);
   U5273 : OAI22_X1 port map( A1 => n10681, A2 => n11595, B1 => n5988, B2 => 
                           n11604, ZN => n6899);
   U5274 : OAI22_X1 port map( A1 => n10674, A2 => n11595, B1 => n5924, B2 => 
                           n11604, ZN => n6898);
   U5275 : OAI22_X1 port map( A1 => n10667, A2 => n11595, B1 => n5892, B2 => 
                           n11604, ZN => n6897);
   U5276 : OAI22_X1 port map( A1 => n10660, A2 => n11595, B1 => n5860, B2 => 
                           n11604, ZN => n6896);
   U5277 : OAI22_X1 port map( A1 => n10653, A2 => n11595, B1 => n5828, B2 => 
                           n11605, ZN => n6895);
   U5278 : OAI22_X1 port map( A1 => n10646, A2 => n11595, B1 => n5796, B2 => 
                           n11605, ZN => n6894);
   U5279 : OAI22_X1 port map( A1 => n10639, A2 => n11595, B1 => n5764, B2 => 
                           n11605, ZN => n6893);
   U5280 : OAI22_X1 port map( A1 => n10632, A2 => n11595, B1 => n5732, B2 => 
                           n11605, ZN => n6892);
   U5281 : OAI22_X1 port map( A1 => n10849, A2 => n11585, B1 => n673, B2 => 
                           n11586, ZN => n6891);
   U5282 : OAI22_X1 port map( A1 => n10842, A2 => n11585, B1 => n672, B2 => 
                           n11586, ZN => n6890);
   U5283 : OAI22_X1 port map( A1 => n10835, A2 => n11585, B1 => n671, B2 => 
                           n11586, ZN => n6889);
   U5284 : OAI22_X1 port map( A1 => n10828, A2 => n11585, B1 => n670, B2 => 
                           n11586, ZN => n6888);
   U5285 : OAI22_X1 port map( A1 => n10821, A2 => n11585, B1 => n669, B2 => 
                           n11587, ZN => n6887);
   U5286 : OAI22_X1 port map( A1 => n10814, A2 => n11585, B1 => n668, B2 => 
                           n11587, ZN => n6886);
   U5287 : OAI22_X1 port map( A1 => n10807, A2 => n11585, B1 => n667, B2 => 
                           n11587, ZN => n6885);
   U5288 : OAI22_X1 port map( A1 => n10800, A2 => n11585, B1 => n666, B2 => 
                           n11587, ZN => n6884);
   U5289 : OAI22_X1 port map( A1 => n10793, A2 => n11584, B1 => n665, B2 => 
                           n11588, ZN => n6883);
   U5290 : OAI22_X1 port map( A1 => n10786, A2 => n11584, B1 => n664, B2 => 
                           n11588, ZN => n6882);
   U5291 : OAI22_X1 port map( A1 => n10779, A2 => n11584, B1 => n663, B2 => 
                           n11588, ZN => n6881);
   U5292 : OAI22_X1 port map( A1 => n10772, A2 => n11584, B1 => n662, B2 => 
                           n11588, ZN => n6880);
   U5293 : OAI22_X1 port map( A1 => n10765, A2 => n11584, B1 => n661, B2 => 
                           n11589, ZN => n6879);
   U5294 : OAI22_X1 port map( A1 => n10758, A2 => n11584, B1 => n660, B2 => 
                           n11589, ZN => n6878);
   U5295 : OAI22_X1 port map( A1 => n10751, A2 => n11584, B1 => n659, B2 => 
                           n11589, ZN => n6877);
   U5296 : OAI22_X1 port map( A1 => n10744, A2 => n11584, B1 => n658, B2 => 
                           n11589, ZN => n6876);
   U5297 : OAI22_X1 port map( A1 => n10737, A2 => n11584, B1 => n657, B2 => 
                           n11590, ZN => n6875);
   U5298 : OAI22_X1 port map( A1 => n10730, A2 => n11584, B1 => n656, B2 => 
                           n11590, ZN => n6874);
   U5299 : OAI22_X1 port map( A1 => n10723, A2 => n11584, B1 => n655, B2 => 
                           n11590, ZN => n6873);
   U5300 : OAI22_X1 port map( A1 => n10716, A2 => n11584, B1 => n654, B2 => 
                           n11590, ZN => n6872);
   U5301 : OAI22_X1 port map( A1 => n10709, A2 => n11583, B1 => n653, B2 => 
                           n11591, ZN => n6871);
   U5302 : OAI22_X1 port map( A1 => n10702, A2 => n11583, B1 => n652, B2 => 
                           n11591, ZN => n6870);
   U5303 : OAI22_X1 port map( A1 => n10695, A2 => n11583, B1 => n651, B2 => 
                           n11591, ZN => n6869);
   U5304 : OAI22_X1 port map( A1 => n10688, A2 => n11583, B1 => n650, B2 => 
                           n11591, ZN => n6868);
   U5305 : OAI22_X1 port map( A1 => n10681, A2 => n11583, B1 => n649, B2 => 
                           n11592, ZN => n6867);
   U5306 : OAI22_X1 port map( A1 => n10674, A2 => n11583, B1 => n648, B2 => 
                           n11592, ZN => n6866);
   U5307 : OAI22_X1 port map( A1 => n10667, A2 => n11583, B1 => n647, B2 => 
                           n11592, ZN => n6865);
   U5308 : OAI22_X1 port map( A1 => n10660, A2 => n11583, B1 => n646, B2 => 
                           n11592, ZN => n6864);
   U5309 : OAI22_X1 port map( A1 => n10653, A2 => n11583, B1 => n645, B2 => 
                           n11593, ZN => n6863);
   U5310 : OAI22_X1 port map( A1 => n10646, A2 => n11583, B1 => n644, B2 => 
                           n11593, ZN => n6862);
   U5311 : OAI22_X1 port map( A1 => n10639, A2 => n11583, B1 => n643, B2 => 
                           n11593, ZN => n6861);
   U5312 : OAI22_X1 port map( A1 => n10632, A2 => n11583, B1 => n642, B2 => 
                           n11593, ZN => n6860);
   U5313 : OAI22_X1 port map( A1 => n10849, A2 => n11573, B1 => n10530, B2 => 
                           n11574, ZN => n6859);
   U5314 : OAI22_X1 port map( A1 => n10842, A2 => n11573, B1 => n10498, B2 => 
                           n11574, ZN => n6858);
   U5315 : OAI22_X1 port map( A1 => n10835, A2 => n11573, B1 => n10466, B2 => 
                           n11574, ZN => n6857);
   U5316 : OAI22_X1 port map( A1 => n10828, A2 => n11573, B1 => n10434, B2 => 
                           n11574, ZN => n6856);
   U5317 : OAI22_X1 port map( A1 => n10821, A2 => n11573, B1 => n10402, B2 => 
                           n11575, ZN => n6855);
   U5318 : OAI22_X1 port map( A1 => n10814, A2 => n11573, B1 => n10367, B2 => 
                           n11575, ZN => n6854);
   U5319 : OAI22_X1 port map( A1 => n10807, A2 => n11573, B1 => n10335, B2 => 
                           n11575, ZN => n6853);
   U5320 : OAI22_X1 port map( A1 => n10800, A2 => n11573, B1 => n10300, B2 => 
                           n11575, ZN => n6852);
   U5321 : OAI22_X1 port map( A1 => n10793, A2 => n11572, B1 => n10268, B2 => 
                           n11576, ZN => n6851);
   U5322 : OAI22_X1 port map( A1 => n10786, A2 => n11572, B1 => n10236, B2 => 
                           n11576, ZN => n6850);
   U5323 : OAI22_X1 port map( A1 => n10779, A2 => n11572, B1 => n10202, B2 => 
                           n11576, ZN => n6849);
   U5324 : OAI22_X1 port map( A1 => n10772, A2 => n11572, B1 => n10170, B2 => 
                           n11576, ZN => n6848);
   U5325 : OAI22_X1 port map( A1 => n10765, A2 => n11572, B1 => n10138, B2 => 
                           n11577, ZN => n6847);
   U5326 : OAI22_X1 port map( A1 => n10758, A2 => n11572, B1 => n10106, B2 => 
                           n11577, ZN => n6846);
   U5327 : OAI22_X1 port map( A1 => n10751, A2 => n11572, B1 => n10074, B2 => 
                           n11577, ZN => n6845);
   U5328 : OAI22_X1 port map( A1 => n10744, A2 => n11572, B1 => n10042, B2 => 
                           n11577, ZN => n6844);
   U5329 : OAI22_X1 port map( A1 => n10737, A2 => n11572, B1 => n10010, B2 => 
                           n11578, ZN => n6843);
   U5330 : OAI22_X1 port map( A1 => n10730, A2 => n11572, B1 => n9648, B2 => 
                           n11578, ZN => n6842);
   U5331 : OAI22_X1 port map( A1 => n10723, A2 => n11572, B1 => n9616, B2 => 
                           n11578, ZN => n6841);
   U5332 : OAI22_X1 port map( A1 => n10716, A2 => n11572, B1 => n9584, B2 => 
                           n11578, ZN => n6840);
   U5333 : OAI22_X1 port map( A1 => n10709, A2 => n11571, B1 => n9250, B2 => 
                           n11579, ZN => n6839);
   U5334 : OAI22_X1 port map( A1 => n10702, A2 => n11571, B1 => n9186, B2 => 
                           n11579, ZN => n6838);
   U5335 : OAI22_X1 port map( A1 => n10695, A2 => n11571, B1 => n9154, B2 => 
                           n11579, ZN => n6837);
   U5336 : OAI22_X1 port map( A1 => n10688, A2 => n11571, B1 => n6304, B2 => 
                           n11579, ZN => n6836);
   U5337 : OAI22_X1 port map( A1 => n10681, A2 => n11571, B1 => n5987, B2 => 
                           n11580, ZN => n6835);
   U5338 : OAI22_X1 port map( A1 => n10674, A2 => n11571, B1 => n5923, B2 => 
                           n11580, ZN => n6834);
   U5339 : OAI22_X1 port map( A1 => n10667, A2 => n11571, B1 => n5891, B2 => 
                           n11580, ZN => n6833);
   U5340 : OAI22_X1 port map( A1 => n10660, A2 => n11571, B1 => n5859, B2 => 
                           n11580, ZN => n6832);
   U5341 : OAI22_X1 port map( A1 => n10653, A2 => n11571, B1 => n5827, B2 => 
                           n11581, ZN => n6831);
   U5342 : OAI22_X1 port map( A1 => n10646, A2 => n11571, B1 => n5795, B2 => 
                           n11581, ZN => n6830);
   U5343 : OAI22_X1 port map( A1 => n10639, A2 => n11571, B1 => n5763, B2 => 
                           n11581, ZN => n6829);
   U5344 : OAI22_X1 port map( A1 => n10632, A2 => n11571, B1 => n5731, B2 => 
                           n11581, ZN => n6828);
   U5345 : OAI22_X1 port map( A1 => n10849, A2 => n11561, B1 => n10532, B2 => 
                           n11562, ZN => n6827);
   U5346 : OAI22_X1 port map( A1 => n10842, A2 => n11561, B1 => n10500, B2 => 
                           n11562, ZN => n6826);
   U5347 : OAI22_X1 port map( A1 => n10835, A2 => n11561, B1 => n10468, B2 => 
                           n11562, ZN => n6825);
   U5348 : OAI22_X1 port map( A1 => n10828, A2 => n11561, B1 => n10436, B2 => 
                           n11562, ZN => n6824);
   U5349 : OAI22_X1 port map( A1 => n10821, A2 => n11561, B1 => n10404, B2 => 
                           n11563, ZN => n6823);
   U5350 : OAI22_X1 port map( A1 => n10814, A2 => n11561, B1 => n10369, B2 => 
                           n11563, ZN => n6822);
   U5351 : OAI22_X1 port map( A1 => n10807, A2 => n11561, B1 => n10337, B2 => 
                           n11563, ZN => n6821);
   U5352 : OAI22_X1 port map( A1 => n10800, A2 => n11561, B1 => n10305, B2 => 
                           n11563, ZN => n6820);
   U5353 : OAI22_X1 port map( A1 => n10793, A2 => n11560, B1 => n10270, B2 => 
                           n11564, ZN => n6819);
   U5354 : OAI22_X1 port map( A1 => n10786, A2 => n11560, B1 => n10238, B2 => 
                           n11564, ZN => n6818);
   U5355 : OAI22_X1 port map( A1 => n10779, A2 => n11560, B1 => n10204, B2 => 
                           n11564, ZN => n6817);
   U5356 : OAI22_X1 port map( A1 => n10772, A2 => n11560, B1 => n10172, B2 => 
                           n11564, ZN => n6816);
   U5357 : OAI22_X1 port map( A1 => n10765, A2 => n11560, B1 => n10140, B2 => 
                           n11565, ZN => n6815);
   U5358 : OAI22_X1 port map( A1 => n10758, A2 => n11560, B1 => n10108, B2 => 
                           n11565, ZN => n6814);
   U5359 : OAI22_X1 port map( A1 => n10751, A2 => n11560, B1 => n10076, B2 => 
                           n11565, ZN => n6813);
   U5360 : OAI22_X1 port map( A1 => n10744, A2 => n11560, B1 => n10044, B2 => 
                           n11565, ZN => n6812);
   U5361 : OAI22_X1 port map( A1 => n10737, A2 => n11560, B1 => n10012, B2 => 
                           n11566, ZN => n6811);
   U5362 : OAI22_X1 port map( A1 => n10730, A2 => n11560, B1 => n9650, B2 => 
                           n11566, ZN => n6810);
   U5363 : OAI22_X1 port map( A1 => n10723, A2 => n11560, B1 => n9618, B2 => 
                           n11566, ZN => n6809);
   U5364 : OAI22_X1 port map( A1 => n10716, A2 => n11560, B1 => n9586, B2 => 
                           n11566, ZN => n6808);
   U5365 : OAI22_X1 port map( A1 => n10709, A2 => n11559, B1 => n9252, B2 => 
                           n11567, ZN => n6807);
   U5366 : OAI22_X1 port map( A1 => n10702, A2 => n11559, B1 => n9188, B2 => 
                           n11567, ZN => n6806);
   U5367 : OAI22_X1 port map( A1 => n10695, A2 => n11559, B1 => n9156, B2 => 
                           n11567, ZN => n6805);
   U5368 : OAI22_X1 port map( A1 => n10688, A2 => n11559, B1 => n6306, B2 => 
                           n11567, ZN => n6804);
   U5369 : OAI22_X1 port map( A1 => n10681, A2 => n11559, B1 => n5989, B2 => 
                           n11568, ZN => n6803);
   U5370 : OAI22_X1 port map( A1 => n10674, A2 => n11559, B1 => n5925, B2 => 
                           n11568, ZN => n6802);
   U5371 : OAI22_X1 port map( A1 => n10667, A2 => n11559, B1 => n5893, B2 => 
                           n11568, ZN => n6801);
   U5372 : OAI22_X1 port map( A1 => n10660, A2 => n11559, B1 => n5861, B2 => 
                           n11568, ZN => n6800);
   U5373 : OAI22_X1 port map( A1 => n10653, A2 => n11559, B1 => n5829, B2 => 
                           n11569, ZN => n6799);
   U5374 : OAI22_X1 port map( A1 => n10646, A2 => n11559, B1 => n5797, B2 => 
                           n11569, ZN => n6798);
   U5375 : OAI22_X1 port map( A1 => n10639, A2 => n11559, B1 => n5765, B2 => 
                           n11569, ZN => n6797);
   U5376 : OAI22_X1 port map( A1 => n10632, A2 => n11559, B1 => n5733, B2 => 
                           n11569, ZN => n6796);
   U5377 : OAI22_X1 port map( A1 => n10849, A2 => n11513, B1 => n10536, B2 => 
                           n11514, ZN => n6699);
   U5378 : OAI22_X1 port map( A1 => n10842, A2 => n11513, B1 => n10504, B2 => 
                           n11514, ZN => n6698);
   U5379 : OAI22_X1 port map( A1 => n10835, A2 => n11513, B1 => n10472, B2 => 
                           n11514, ZN => n6697);
   U5380 : OAI22_X1 port map( A1 => n10828, A2 => n11513, B1 => n10440, B2 => 
                           n11514, ZN => n6696);
   U5381 : OAI22_X1 port map( A1 => n10821, A2 => n11513, B1 => n10408, B2 => 
                           n11515, ZN => n6695);
   U5382 : OAI22_X1 port map( A1 => n10814, A2 => n11513, B1 => n10373, B2 => 
                           n11515, ZN => n6694);
   U5383 : OAI22_X1 port map( A1 => n10807, A2 => n11513, B1 => n10341, B2 => 
                           n11515, ZN => n6693);
   U5384 : OAI22_X1 port map( A1 => n10800, A2 => n11513, B1 => n10309, B2 => 
                           n11515, ZN => n6692);
   U5385 : OAI22_X1 port map( A1 => n10793, A2 => n11512, B1 => n10274, B2 => 
                           n11516, ZN => n6691);
   U5386 : OAI22_X1 port map( A1 => n10786, A2 => n11512, B1 => n10242, B2 => 
                           n11516, ZN => n6690);
   U5387 : OAI22_X1 port map( A1 => n10779, A2 => n11512, B1 => n10210, B2 => 
                           n11516, ZN => n6689);
   U5388 : OAI22_X1 port map( A1 => n10772, A2 => n11512, B1 => n10176, B2 => 
                           n11516, ZN => n6688);
   U5389 : OAI22_X1 port map( A1 => n10765, A2 => n11512, B1 => n10144, B2 => 
                           n11517, ZN => n6687);
   U5390 : OAI22_X1 port map( A1 => n10758, A2 => n11512, B1 => n10112, B2 => 
                           n11517, ZN => n6686);
   U5391 : OAI22_X1 port map( A1 => n10751, A2 => n11512, B1 => n10080, B2 => 
                           n11517, ZN => n6685);
   U5392 : OAI22_X1 port map( A1 => n10744, A2 => n11512, B1 => n10048, B2 => 
                           n11517, ZN => n6684);
   U5393 : OAI22_X1 port map( A1 => n10737, A2 => n11512, B1 => n10016, B2 => 
                           n11518, ZN => n6683);
   U5394 : OAI22_X1 port map( A1 => n10730, A2 => n11512, B1 => n9654, B2 => 
                           n11518, ZN => n6682);
   U5395 : OAI22_X1 port map( A1 => n10723, A2 => n11512, B1 => n9622, B2 => 
                           n11518, ZN => n6681);
   U5396 : OAI22_X1 port map( A1 => n10716, A2 => n11512, B1 => n9590, B2 => 
                           n11518, ZN => n6680);
   U5397 : OAI22_X1 port map( A1 => n10709, A2 => n11511, B1 => n9256, B2 => 
                           n11519, ZN => n6679);
   U5398 : OAI22_X1 port map( A1 => n10702, A2 => n11511, B1 => n9192, B2 => 
                           n11519, ZN => n6678);
   U5399 : OAI22_X1 port map( A1 => n10695, A2 => n11511, B1 => n9160, B2 => 
                           n11519, ZN => n6677);
   U5400 : OAI22_X1 port map( A1 => n10688, A2 => n11511, B1 => n6310, B2 => 
                           n11519, ZN => n6676);
   U5401 : OAI22_X1 port map( A1 => n10681, A2 => n11511, B1 => n5993, B2 => 
                           n11520, ZN => n6675);
   U5402 : OAI22_X1 port map( A1 => n10674, A2 => n11511, B1 => n5929, B2 => 
                           n11520, ZN => n6674);
   U5403 : OAI22_X1 port map( A1 => n10667, A2 => n11511, B1 => n5897, B2 => 
                           n11520, ZN => n6673);
   U5404 : OAI22_X1 port map( A1 => n10660, A2 => n11511, B1 => n5865, B2 => 
                           n11520, ZN => n6672);
   U5405 : OAI22_X1 port map( A1 => n10653, A2 => n11511, B1 => n5833, B2 => 
                           n11521, ZN => n6671);
   U5406 : OAI22_X1 port map( A1 => n10646, A2 => n11511, B1 => n5801, B2 => 
                           n11521, ZN => n6670);
   U5407 : OAI22_X1 port map( A1 => n10639, A2 => n11511, B1 => n5769, B2 => 
                           n11521, ZN => n6669);
   U5408 : OAI22_X1 port map( A1 => n10632, A2 => n11511, B1 => n5737, B2 => 
                           n11521, ZN => n6668);
   U5409 : OAI22_X1 port map( A1 => n10846, A2 => n12029, B1 => n12030, B2 => 
                           n13843, ZN => n8075);
   U5410 : OAI22_X1 port map( A1 => n10839, A2 => n12029, B1 => n12030, B2 => 
                           n13842, ZN => n8074);
   U5411 : OAI22_X1 port map( A1 => n10832, A2 => n12029, B1 => n12030, B2 => 
                           n13841, ZN => n8073);
   U5412 : OAI22_X1 port map( A1 => n10825, A2 => n12029, B1 => n12030, B2 => 
                           n13840, ZN => n8072);
   U5413 : OAI22_X1 port map( A1 => n10818, A2 => n12029, B1 => n12031, B2 => 
                           n13839, ZN => n8071);
   U5414 : OAI22_X1 port map( A1 => n10811, A2 => n12029, B1 => n12031, B2 => 
                           n13838, ZN => n8070);
   U5415 : OAI22_X1 port map( A1 => n10804, A2 => n12029, B1 => n12031, B2 => 
                           n13837, ZN => n8069);
   U5416 : OAI22_X1 port map( A1 => n10797, A2 => n12029, B1 => n12031, B2 => 
                           n13836, ZN => n8068);
   U5417 : OAI22_X1 port map( A1 => n10790, A2 => n12028, B1 => n12032, B2 => 
                           n13835, ZN => n8067);
   U5418 : OAI22_X1 port map( A1 => n10783, A2 => n12028, B1 => n12032, B2 => 
                           n13834, ZN => n8066);
   U5419 : OAI22_X1 port map( A1 => n10776, A2 => n12028, B1 => n12032, B2 => 
                           n13833, ZN => n8065);
   U5420 : OAI22_X1 port map( A1 => n10769, A2 => n12028, B1 => n12032, B2 => 
                           n13832, ZN => n8064);
   U5421 : OAI22_X1 port map( A1 => n10762, A2 => n12028, B1 => n12033, B2 => 
                           n13831, ZN => n8063);
   U5422 : OAI22_X1 port map( A1 => n10755, A2 => n12028, B1 => n12033, B2 => 
                           n13830, ZN => n8062);
   U5423 : OAI22_X1 port map( A1 => n10748, A2 => n12028, B1 => n12033, B2 => 
                           n13829, ZN => n8061);
   U5424 : OAI22_X1 port map( A1 => n10741, A2 => n12028, B1 => n12033, B2 => 
                           n13828, ZN => n8060);
   U5425 : OAI22_X1 port map( A1 => n10734, A2 => n12028, B1 => n12034, B2 => 
                           n13827, ZN => n8059);
   U5426 : OAI22_X1 port map( A1 => n10727, A2 => n12028, B1 => n12034, B2 => 
                           n13826, ZN => n8058);
   U5427 : OAI22_X1 port map( A1 => n10720, A2 => n12028, B1 => n12034, B2 => 
                           n13825, ZN => n8057);
   U5428 : OAI22_X1 port map( A1 => n10713, A2 => n12028, B1 => n12034, B2 => 
                           n13824, ZN => n8056);
   U5429 : OAI22_X1 port map( A1 => n10706, A2 => n12027, B1 => n12035, B2 => 
                           n13823, ZN => n8055);
   U5430 : OAI22_X1 port map( A1 => n10699, A2 => n12027, B1 => n12035, B2 => 
                           n13822, ZN => n8054);
   U5431 : OAI22_X1 port map( A1 => n10692, A2 => n12027, B1 => n12035, B2 => 
                           n13821, ZN => n8053);
   U5432 : OAI22_X1 port map( A1 => n10685, A2 => n12027, B1 => n12035, B2 => 
                           n13820, ZN => n8052);
   U5433 : OAI22_X1 port map( A1 => n10678, A2 => n12027, B1 => n12036, B2 => 
                           n13819, ZN => n8051);
   U5434 : OAI22_X1 port map( A1 => n10671, A2 => n12027, B1 => n12036, B2 => 
                           n13818, ZN => n8050);
   U5435 : OAI22_X1 port map( A1 => n10664, A2 => n12027, B1 => n12036, B2 => 
                           n13817, ZN => n8049);
   U5436 : OAI22_X1 port map( A1 => n10657, A2 => n12027, B1 => n12036, B2 => 
                           n13816, ZN => n8048);
   U5437 : OAI22_X1 port map( A1 => n10650, A2 => n12027, B1 => n12037, B2 => 
                           n13815, ZN => n8047);
   U5438 : OAI22_X1 port map( A1 => n10643, A2 => n12027, B1 => n12037, B2 => 
                           n13814, ZN => n8046);
   U5439 : OAI22_X1 port map( A1 => n10636, A2 => n12027, B1 => n12037, B2 => 
                           n13813, ZN => n8045);
   U5440 : OAI22_X1 port map( A1 => n10629, A2 => n12027, B1 => n12037, B2 => 
                           n13812, ZN => n8044);
   U5441 : OAI22_X1 port map( A1 => n10727, A2 => n12016, B1 => n12022, B2 => 
                           n13794, ZN => n8026);
   U5442 : OAI22_X1 port map( A1 => n10720, A2 => n12016, B1 => n12022, B2 => 
                           n13793, ZN => n8025);
   U5443 : OAI22_X1 port map( A1 => n10713, A2 => n12016, B1 => n12022, B2 => 
                           n13792, ZN => n8024);
   U5444 : OAI22_X1 port map( A1 => n10706, A2 => n12015, B1 => n12023, B2 => 
                           n13791, ZN => n8023);
   U5445 : OAI22_X1 port map( A1 => n10699, A2 => n12015, B1 => n12023, B2 => 
                           n13790, ZN => n8022);
   U5446 : OAI22_X1 port map( A1 => n10692, A2 => n12015, B1 => n12023, B2 => 
                           n13789, ZN => n8021);
   U5447 : OAI22_X1 port map( A1 => n10685, A2 => n12015, B1 => n12023, B2 => 
                           n13788, ZN => n8020);
   U5448 : OAI22_X1 port map( A1 => n10678, A2 => n12015, B1 => n12024, B2 => 
                           n13787, ZN => n8019);
   U5449 : OAI22_X1 port map( A1 => n10671, A2 => n12015, B1 => n12024, B2 => 
                           n13786, ZN => n8018);
   U5450 : OAI22_X1 port map( A1 => n10664, A2 => n12015, B1 => n12024, B2 => 
                           n13785, ZN => n8017);
   U5451 : OAI22_X1 port map( A1 => n10657, A2 => n12015, B1 => n12024, B2 => 
                           n13784, ZN => n8016);
   U5452 : OAI22_X1 port map( A1 => n10650, A2 => n12015, B1 => n12025, B2 => 
                           n13783, ZN => n8015);
   U5453 : OAI22_X1 port map( A1 => n10643, A2 => n12015, B1 => n12025, B2 => 
                           n13782, ZN => n8014);
   U5454 : OAI22_X1 port map( A1 => n10636, A2 => n12015, B1 => n12025, B2 => 
                           n13781, ZN => n8013);
   U5455 : OAI22_X1 port map( A1 => n10629, A2 => n12015, B1 => n12025, B2 => 
                           n13780, ZN => n8012);
   U5456 : OAI22_X1 port map( A1 => n10846, A2 => n12005, B1 => n12010, B2 => 
                           n13779, ZN => n8011);
   U5457 : OAI22_X1 port map( A1 => n10839, A2 => n12005, B1 => n12006, B2 => 
                           n13778, ZN => n8010);
   U5458 : OAI22_X1 port map( A1 => n10832, A2 => n12005, B1 => n12006, B2 => 
                           n13777, ZN => n8009);
   U5459 : OAI22_X1 port map( A1 => n10825, A2 => n12005, B1 => n12006, B2 => 
                           n13776, ZN => n8008);
   U5460 : OAI22_X1 port map( A1 => n10818, A2 => n12005, B1 => n12007, B2 => 
                           n13775, ZN => n8007);
   U5461 : OAI22_X1 port map( A1 => n10811, A2 => n12005, B1 => n12007, B2 => 
                           n13774, ZN => n8006);
   U5462 : OAI22_X1 port map( A1 => n10804, A2 => n12005, B1 => n12007, B2 => 
                           n13773, ZN => n8005);
   U5463 : OAI22_X1 port map( A1 => n10797, A2 => n12005, B1 => n12007, B2 => 
                           n13772, ZN => n8004);
   U5464 : OAI22_X1 port map( A1 => n10790, A2 => n12004, B1 => n12008, B2 => 
                           n13771, ZN => n8003);
   U5465 : OAI22_X1 port map( A1 => n10783, A2 => n12004, B1 => n12008, B2 => 
                           n13770, ZN => n8002);
   U5466 : OAI22_X1 port map( A1 => n10776, A2 => n12004, B1 => n12008, B2 => 
                           n13769, ZN => n8001);
   U5467 : OAI22_X1 port map( A1 => n10769, A2 => n12004, B1 => n12008, B2 => 
                           n13768, ZN => n8000);
   U5468 : OAI22_X1 port map( A1 => n10762, A2 => n12004, B1 => n12009, B2 => 
                           n13767, ZN => n7999);
   U5469 : OAI22_X1 port map( A1 => n10755, A2 => n12004, B1 => n12009, B2 => 
                           n13766, ZN => n7998);
   U5470 : OAI22_X1 port map( A1 => n10748, A2 => n12004, B1 => n12009, B2 => 
                           n13765, ZN => n7997);
   U5471 : OAI22_X1 port map( A1 => n10741, A2 => n12004, B1 => n12009, B2 => 
                           n13764, ZN => n7996);
   U5472 : OAI22_X1 port map( A1 => n10734, A2 => n12004, B1 => n12010, B2 => 
                           n13763, ZN => n7995);
   U5473 : OAI22_X1 port map( A1 => n10727, A2 => n12004, B1 => n12010, B2 => 
                           n13762, ZN => n7994);
   U5474 : OAI22_X1 port map( A1 => n10720, A2 => n12004, B1 => n12010, B2 => 
                           n13761, ZN => n7993);
   U5475 : OAI22_X1 port map( A1 => n10713, A2 => n12004, B1 => n12011, B2 => 
                           n13760, ZN => n7992);
   U5476 : OAI22_X1 port map( A1 => n10706, A2 => n12003, B1 => n12011, B2 => 
                           n13759, ZN => n7991);
   U5477 : OAI22_X1 port map( A1 => n10699, A2 => n12003, B1 => n12011, B2 => 
                           n13758, ZN => n7990);
   U5478 : OAI22_X1 port map( A1 => n10692, A2 => n12003, B1 => n12011, B2 => 
                           n13757, ZN => n7989);
   U5479 : OAI22_X1 port map( A1 => n10685, A2 => n12003, B1 => n12012, B2 => 
                           n13756, ZN => n7988);
   U5480 : OAI22_X1 port map( A1 => n10678, A2 => n12003, B1 => n12012, B2 => 
                           n13755, ZN => n7987);
   U5481 : OAI22_X1 port map( A1 => n10671, A2 => n12003, B1 => n12012, B2 => 
                           n13754, ZN => n7986);
   U5482 : OAI22_X1 port map( A1 => n10664, A2 => n12003, B1 => n12012, B2 => 
                           n13753, ZN => n7985);
   U5483 : OAI22_X1 port map( A1 => n10657, A2 => n12003, B1 => n12013, B2 => 
                           n13752, ZN => n7984);
   U5484 : OAI22_X1 port map( A1 => n10650, A2 => n12003, B1 => n12013, B2 => 
                           n13751, ZN => n7983);
   U5485 : OAI22_X1 port map( A1 => n10643, A2 => n12003, B1 => n12013, B2 => 
                           n13750, ZN => n7982);
   U5486 : OAI22_X1 port map( A1 => n10636, A2 => n12003, B1 => n12013, B2 => 
                           n13749, ZN => n7981);
   U5487 : OAI22_X1 port map( A1 => n10846, A2 => n11993, B1 => n11994, B2 => 
                           n13747, ZN => n7979);
   U5488 : OAI22_X1 port map( A1 => n10839, A2 => n11993, B1 => n11994, B2 => 
                           n13746, ZN => n7978);
   U5489 : OAI22_X1 port map( A1 => n10832, A2 => n11993, B1 => n11994, B2 => 
                           n13745, ZN => n7977);
   U5490 : OAI22_X1 port map( A1 => n10825, A2 => n11993, B1 => n11994, B2 => 
                           n13744, ZN => n7976);
   U5491 : OAI22_X1 port map( A1 => n10818, A2 => n11993, B1 => n11995, B2 => 
                           n13743, ZN => n7975);
   U5492 : OAI22_X1 port map( A1 => n10811, A2 => n11993, B1 => n11995, B2 => 
                           n13742, ZN => n7974);
   U5493 : OAI22_X1 port map( A1 => n10804, A2 => n11993, B1 => n11995, B2 => 
                           n13741, ZN => n7973);
   U5494 : OAI22_X1 port map( A1 => n10797, A2 => n11993, B1 => n11995, B2 => 
                           n13740, ZN => n7972);
   U5495 : OAI22_X1 port map( A1 => n10790, A2 => n11992, B1 => n11996, B2 => 
                           n13739, ZN => n7971);
   U5496 : OAI22_X1 port map( A1 => n10783, A2 => n11992, B1 => n11996, B2 => 
                           n13738, ZN => n7970);
   U5497 : OAI22_X1 port map( A1 => n10776, A2 => n11992, B1 => n11996, B2 => 
                           n13737, ZN => n7969);
   U5498 : OAI22_X1 port map( A1 => n10769, A2 => n11992, B1 => n11996, B2 => 
                           n13736, ZN => n7968);
   U5499 : OAI22_X1 port map( A1 => n10762, A2 => n11992, B1 => n11997, B2 => 
                           n13735, ZN => n7967);
   U5500 : OAI22_X1 port map( A1 => n10755, A2 => n11992, B1 => n11997, B2 => 
                           n13734, ZN => n7966);
   U5501 : OAI22_X1 port map( A1 => n10748, A2 => n11992, B1 => n11997, B2 => 
                           n13733, ZN => n7965);
   U5502 : OAI22_X1 port map( A1 => n10741, A2 => n11992, B1 => n11997, B2 => 
                           n13732, ZN => n7964);
   U5503 : OAI22_X1 port map( A1 => n10734, A2 => n11992, B1 => n11998, B2 => 
                           n13731, ZN => n7963);
   U5504 : OAI22_X1 port map( A1 => n10727, A2 => n11992, B1 => n11998, B2 => 
                           n13730, ZN => n7962);
   U5505 : OAI22_X1 port map( A1 => n10720, A2 => n11992, B1 => n11998, B2 => 
                           n13729, ZN => n7961);
   U5506 : OAI22_X1 port map( A1 => n10713, A2 => n11992, B1 => n11998, B2 => 
                           n13728, ZN => n7960);
   U5507 : OAI22_X1 port map( A1 => n10706, A2 => n11991, B1 => n11999, B2 => 
                           n13727, ZN => n7959);
   U5508 : OAI22_X1 port map( A1 => n10699, A2 => n11991, B1 => n11999, B2 => 
                           n13726, ZN => n7958);
   U5509 : OAI22_X1 port map( A1 => n10692, A2 => n11991, B1 => n11999, B2 => 
                           n13725, ZN => n7957);
   U5510 : OAI22_X1 port map( A1 => n10685, A2 => n11991, B1 => n11999, B2 => 
                           n13724, ZN => n7956);
   U5511 : OAI22_X1 port map( A1 => n10678, A2 => n11991, B1 => n12000, B2 => 
                           n13723, ZN => n7955);
   U5512 : OAI22_X1 port map( A1 => n10671, A2 => n11991, B1 => n12000, B2 => 
                           n13722, ZN => n7954);
   U5513 : OAI22_X1 port map( A1 => n10664, A2 => n11991, B1 => n12000, B2 => 
                           n13721, ZN => n7953);
   U5514 : OAI22_X1 port map( A1 => n10657, A2 => n11991, B1 => n12000, B2 => 
                           n13720, ZN => n7952);
   U5515 : OAI22_X1 port map( A1 => n10650, A2 => n11991, B1 => n12001, B2 => 
                           n13719, ZN => n7951);
   U5516 : OAI22_X1 port map( A1 => n10643, A2 => n11991, B1 => n12001, B2 => 
                           n13718, ZN => n7950);
   U5517 : OAI22_X1 port map( A1 => n10636, A2 => n11991, B1 => n12001, B2 => 
                           n13717, ZN => n7949);
   U5518 : OAI22_X1 port map( A1 => n10629, A2 => n11991, B1 => n12001, B2 => 
                           n13716, ZN => n7948);
   U5519 : OAI22_X1 port map( A1 => n10846, A2 => n11981, B1 => n11982, B2 => 
                           n13715, ZN => n7947);
   U5520 : OAI22_X1 port map( A1 => n10839, A2 => n11981, B1 => n11982, B2 => 
                           n13714, ZN => n7946);
   U5521 : OAI22_X1 port map( A1 => n10832, A2 => n11981, B1 => n11982, B2 => 
                           n13713, ZN => n7945);
   U5522 : OAI22_X1 port map( A1 => n10825, A2 => n11981, B1 => n11982, B2 => 
                           n13712, ZN => n7944);
   U5523 : OAI22_X1 port map( A1 => n10818, A2 => n11981, B1 => n11983, B2 => 
                           n13711, ZN => n7943);
   U5524 : OAI22_X1 port map( A1 => n10811, A2 => n11981, B1 => n11983, B2 => 
                           n13710, ZN => n7942);
   U5525 : OAI22_X1 port map( A1 => n10804, A2 => n11981, B1 => n11983, B2 => 
                           n13709, ZN => n7941);
   U5526 : OAI22_X1 port map( A1 => n10797, A2 => n11981, B1 => n11983, B2 => 
                           n13708, ZN => n7940);
   U5527 : OAI22_X1 port map( A1 => n10790, A2 => n11980, B1 => n11984, B2 => 
                           n13707, ZN => n7939);
   U5528 : OAI22_X1 port map( A1 => n10783, A2 => n11980, B1 => n11984, B2 => 
                           n13706, ZN => n7938);
   U5529 : OAI22_X1 port map( A1 => n10776, A2 => n11980, B1 => n11984, B2 => 
                           n13705, ZN => n7937);
   U5530 : OAI22_X1 port map( A1 => n10769, A2 => n11980, B1 => n11984, B2 => 
                           n13704, ZN => n7936);
   U5531 : OAI22_X1 port map( A1 => n10762, A2 => n11980, B1 => n11985, B2 => 
                           n13703, ZN => n7935);
   U5532 : OAI22_X1 port map( A1 => n10755, A2 => n11980, B1 => n11985, B2 => 
                           n13702, ZN => n7934);
   U5533 : OAI22_X1 port map( A1 => n10748, A2 => n11980, B1 => n11985, B2 => 
                           n13701, ZN => n7933);
   U5534 : OAI22_X1 port map( A1 => n10741, A2 => n11980, B1 => n11985, B2 => 
                           n13700, ZN => n7932);
   U5535 : OAI22_X1 port map( A1 => n10734, A2 => n11980, B1 => n11986, B2 => 
                           n13699, ZN => n7931);
   U5536 : OAI22_X1 port map( A1 => n10727, A2 => n11980, B1 => n11986, B2 => 
                           n13698, ZN => n7930);
   U5537 : OAI22_X1 port map( A1 => n10720, A2 => n11980, B1 => n11986, B2 => 
                           n13697, ZN => n7929);
   U5538 : OAI22_X1 port map( A1 => n10713, A2 => n11980, B1 => n11986, B2 => 
                           n13696, ZN => n7928);
   U5539 : OAI22_X1 port map( A1 => n10706, A2 => n11979, B1 => n11987, B2 => 
                           n13695, ZN => n7927);
   U5540 : OAI22_X1 port map( A1 => n10699, A2 => n11979, B1 => n11987, B2 => 
                           n13694, ZN => n7926);
   U5541 : OAI22_X1 port map( A1 => n10692, A2 => n11979, B1 => n11987, B2 => 
                           n13693, ZN => n7925);
   U5542 : OAI22_X1 port map( A1 => n10685, A2 => n11979, B1 => n11987, B2 => 
                           n13692, ZN => n7924);
   U5543 : OAI22_X1 port map( A1 => n10678, A2 => n11979, B1 => n11988, B2 => 
                           n13691, ZN => n7923);
   U5544 : OAI22_X1 port map( A1 => n10671, A2 => n11979, B1 => n11988, B2 => 
                           n13690, ZN => n7922);
   U5545 : OAI22_X1 port map( A1 => n10664, A2 => n11979, B1 => n11988, B2 => 
                           n13689, ZN => n7921);
   U5546 : OAI22_X1 port map( A1 => n10657, A2 => n11979, B1 => n11988, B2 => 
                           n13688, ZN => n7920);
   U5547 : OAI22_X1 port map( A1 => n10650, A2 => n11979, B1 => n11989, B2 => 
                           n13687, ZN => n7919);
   U5548 : OAI22_X1 port map( A1 => n10643, A2 => n11979, B1 => n11989, B2 => 
                           n13686, ZN => n7918);
   U5549 : OAI22_X1 port map( A1 => n10636, A2 => n11979, B1 => n11989, B2 => 
                           n13685, ZN => n7917);
   U5550 : OAI22_X1 port map( A1 => n10629, A2 => n11979, B1 => n11989, B2 => 
                           n13684, ZN => n7916);
   U5551 : OAI22_X1 port map( A1 => n10846, A2 => n11969, B1 => n11970, B2 => 
                           n13683, ZN => n7915);
   U5552 : OAI22_X1 port map( A1 => n10839, A2 => n11969, B1 => n11970, B2 => 
                           n13682, ZN => n7914);
   U5553 : OAI22_X1 port map( A1 => n10832, A2 => n11969, B1 => n11970, B2 => 
                           n13681, ZN => n7913);
   U5554 : OAI22_X1 port map( A1 => n10825, A2 => n11969, B1 => n11970, B2 => 
                           n13680, ZN => n7912);
   U5555 : OAI22_X1 port map( A1 => n10818, A2 => n11969, B1 => n11971, B2 => 
                           n13679, ZN => n7911);
   U5556 : OAI22_X1 port map( A1 => n10811, A2 => n11969, B1 => n11971, B2 => 
                           n13678, ZN => n7910);
   U5557 : OAI22_X1 port map( A1 => n10804, A2 => n11969, B1 => n11971, B2 => 
                           n13677, ZN => n7909);
   U5558 : OAI22_X1 port map( A1 => n10797, A2 => n11969, B1 => n11971, B2 => 
                           n13676, ZN => n7908);
   U5559 : OAI22_X1 port map( A1 => n10790, A2 => n11968, B1 => n11972, B2 => 
                           n13675, ZN => n7907);
   U5560 : OAI22_X1 port map( A1 => n10783, A2 => n11968, B1 => n11972, B2 => 
                           n13674, ZN => n7906);
   U5561 : OAI22_X1 port map( A1 => n10776, A2 => n11968, B1 => n11972, B2 => 
                           n13673, ZN => n7905);
   U5562 : OAI22_X1 port map( A1 => n10769, A2 => n11968, B1 => n11972, B2 => 
                           n13672, ZN => n7904);
   U5563 : OAI22_X1 port map( A1 => n10762, A2 => n11968, B1 => n11973, B2 => 
                           n13671, ZN => n7903);
   U5564 : OAI22_X1 port map( A1 => n10755, A2 => n11968, B1 => n11973, B2 => 
                           n13670, ZN => n7902);
   U5565 : OAI22_X1 port map( A1 => n10748, A2 => n11968, B1 => n11973, B2 => 
                           n13669, ZN => n7901);
   U5566 : OAI22_X1 port map( A1 => n10741, A2 => n11968, B1 => n11973, B2 => 
                           n13668, ZN => n7900);
   U5567 : OAI22_X1 port map( A1 => n10734, A2 => n11968, B1 => n11974, B2 => 
                           n13667, ZN => n7899);
   U5568 : OAI22_X1 port map( A1 => n10727, A2 => n11968, B1 => n11974, B2 => 
                           n13666, ZN => n7898);
   U5569 : OAI22_X1 port map( A1 => n10720, A2 => n11968, B1 => n11974, B2 => 
                           n13665, ZN => n7897);
   U5570 : OAI22_X1 port map( A1 => n10713, A2 => n11968, B1 => n11974, B2 => 
                           n13664, ZN => n7896);
   U5571 : OAI22_X1 port map( A1 => n10706, A2 => n11967, B1 => n11975, B2 => 
                           n13663, ZN => n7895);
   U5572 : OAI22_X1 port map( A1 => n10699, A2 => n11967, B1 => n11975, B2 => 
                           n13662, ZN => n7894);
   U5573 : OAI22_X1 port map( A1 => n10692, A2 => n11967, B1 => n11975, B2 => 
                           n13661, ZN => n7893);
   U5574 : OAI22_X1 port map( A1 => n10685, A2 => n11967, B1 => n11975, B2 => 
                           n13660, ZN => n7892);
   U5575 : OAI22_X1 port map( A1 => n10678, A2 => n11967, B1 => n11976, B2 => 
                           n13659, ZN => n7891);
   U5576 : OAI22_X1 port map( A1 => n10671, A2 => n11967, B1 => n11976, B2 => 
                           n13658, ZN => n7890);
   U5577 : OAI22_X1 port map( A1 => n10664, A2 => n11967, B1 => n11976, B2 => 
                           n13657, ZN => n7889);
   U5578 : OAI22_X1 port map( A1 => n10657, A2 => n11967, B1 => n11976, B2 => 
                           n13656, ZN => n7888);
   U5579 : OAI22_X1 port map( A1 => n10650, A2 => n11967, B1 => n11977, B2 => 
                           n13655, ZN => n7887);
   U5580 : OAI22_X1 port map( A1 => n10643, A2 => n11967, B1 => n11977, B2 => 
                           n13654, ZN => n7886);
   U5581 : OAI22_X1 port map( A1 => n10636, A2 => n11967, B1 => n11977, B2 => 
                           n13653, ZN => n7885);
   U5582 : OAI22_X1 port map( A1 => n10629, A2 => n11967, B1 => n11977, B2 => 
                           n13652, ZN => n7884);
   U5583 : OAI22_X1 port map( A1 => n10847, A2 => n11921, B1 => n11922, B2 => 
                           n13555, ZN => n7787);
   U5584 : OAI22_X1 port map( A1 => n10840, A2 => n11921, B1 => n11922, B2 => 
                           n13554, ZN => n7786);
   U5585 : OAI22_X1 port map( A1 => n10833, A2 => n11921, B1 => n11922, B2 => 
                           n13553, ZN => n7785);
   U5586 : OAI22_X1 port map( A1 => n10826, A2 => n11921, B1 => n11922, B2 => 
                           n13552, ZN => n7784);
   U5587 : OAI22_X1 port map( A1 => n10819, A2 => n11921, B1 => n11923, B2 => 
                           n13551, ZN => n7783);
   U5588 : OAI22_X1 port map( A1 => n10812, A2 => n11921, B1 => n11923, B2 => 
                           n13550, ZN => n7782);
   U5589 : OAI22_X1 port map( A1 => n10805, A2 => n11921, B1 => n11923, B2 => 
                           n13549, ZN => n7781);
   U5590 : OAI22_X1 port map( A1 => n10798, A2 => n11921, B1 => n11923, B2 => 
                           n13548, ZN => n7780);
   U5591 : OAI22_X1 port map( A1 => n10791, A2 => n11920, B1 => n11924, B2 => 
                           n13547, ZN => n7779);
   U5592 : OAI22_X1 port map( A1 => n10784, A2 => n11920, B1 => n11924, B2 => 
                           n13546, ZN => n7778);
   U5593 : OAI22_X1 port map( A1 => n10777, A2 => n11920, B1 => n11924, B2 => 
                           n13545, ZN => n7777);
   U5594 : OAI22_X1 port map( A1 => n10770, A2 => n11920, B1 => n11924, B2 => 
                           n13544, ZN => n7776);
   U5595 : OAI22_X1 port map( A1 => n10763, A2 => n11920, B1 => n11925, B2 => 
                           n13543, ZN => n7775);
   U5596 : OAI22_X1 port map( A1 => n10756, A2 => n11920, B1 => n11925, B2 => 
                           n13542, ZN => n7774);
   U5597 : OAI22_X1 port map( A1 => n10749, A2 => n11920, B1 => n11925, B2 => 
                           n13541, ZN => n7773);
   U5598 : OAI22_X1 port map( A1 => n10742, A2 => n11920, B1 => n11925, B2 => 
                           n13540, ZN => n7772);
   U5599 : OAI22_X1 port map( A1 => n10735, A2 => n11920, B1 => n11926, B2 => 
                           n13539, ZN => n7771);
   U5600 : OAI22_X1 port map( A1 => n10728, A2 => n11920, B1 => n11926, B2 => 
                           n13538, ZN => n7770);
   U5601 : OAI22_X1 port map( A1 => n10721, A2 => n11920, B1 => n11926, B2 => 
                           n13537, ZN => n7769);
   U5602 : OAI22_X1 port map( A1 => n10714, A2 => n11920, B1 => n11926, B2 => 
                           n13536, ZN => n7768);
   U5603 : OAI22_X1 port map( A1 => n10707, A2 => n11919, B1 => n11927, B2 => 
                           n13535, ZN => n7767);
   U5604 : OAI22_X1 port map( A1 => n10700, A2 => n11919, B1 => n11927, B2 => 
                           n13534, ZN => n7766);
   U5605 : OAI22_X1 port map( A1 => n10693, A2 => n11919, B1 => n11927, B2 => 
                           n13533, ZN => n7765);
   U5606 : OAI22_X1 port map( A1 => n10686, A2 => n11919, B1 => n11927, B2 => 
                           n13532, ZN => n7764);
   U5607 : OAI22_X1 port map( A1 => n10679, A2 => n11919, B1 => n11928, B2 => 
                           n13531, ZN => n7763);
   U5608 : OAI22_X1 port map( A1 => n10672, A2 => n11919, B1 => n11928, B2 => 
                           n13530, ZN => n7762);
   U5609 : OAI22_X1 port map( A1 => n10665, A2 => n11919, B1 => n11928, B2 => 
                           n13529, ZN => n7761);
   U5610 : OAI22_X1 port map( A1 => n10658, A2 => n11919, B1 => n11928, B2 => 
                           n13528, ZN => n7760);
   U5611 : OAI22_X1 port map( A1 => n10651, A2 => n11919, B1 => n11929, B2 => 
                           n13527, ZN => n7759);
   U5612 : OAI22_X1 port map( A1 => n10644, A2 => n11919, B1 => n11929, B2 => 
                           n13526, ZN => n7758);
   U5613 : OAI22_X1 port map( A1 => n10637, A2 => n11919, B1 => n11929, B2 => 
                           n13525, ZN => n7757);
   U5614 : OAI22_X1 port map( A1 => n10630, A2 => n11919, B1 => n11929, B2 => 
                           n13524, ZN => n7756);
   U5615 : OAI22_X1 port map( A1 => n10847, A2 => n11909, B1 => n11910, B2 => 
                           n13523, ZN => n7755);
   U5616 : OAI22_X1 port map( A1 => n10840, A2 => n11909, B1 => n11910, B2 => 
                           n13522, ZN => n7754);
   U5617 : OAI22_X1 port map( A1 => n10833, A2 => n11909, B1 => n11910, B2 => 
                           n13521, ZN => n7753);
   U5618 : OAI22_X1 port map( A1 => n10826, A2 => n11909, B1 => n11910, B2 => 
                           n13520, ZN => n7752);
   U5619 : OAI22_X1 port map( A1 => n10819, A2 => n11909, B1 => n11911, B2 => 
                           n13519, ZN => n7751);
   U5620 : OAI22_X1 port map( A1 => n10812, A2 => n11909, B1 => n11911, B2 => 
                           n13518, ZN => n7750);
   U5621 : OAI22_X1 port map( A1 => n10805, A2 => n11909, B1 => n11911, B2 => 
                           n13517, ZN => n7749);
   U5622 : OAI22_X1 port map( A1 => n10798, A2 => n11909, B1 => n11911, B2 => 
                           n13516, ZN => n7748);
   U5623 : OAI22_X1 port map( A1 => n10791, A2 => n11908, B1 => n11912, B2 => 
                           n13515, ZN => n7747);
   U5624 : OAI22_X1 port map( A1 => n10784, A2 => n11908, B1 => n11912, B2 => 
                           n13514, ZN => n7746);
   U5625 : OAI22_X1 port map( A1 => n10777, A2 => n11908, B1 => n11912, B2 => 
                           n13513, ZN => n7745);
   U5626 : OAI22_X1 port map( A1 => n10770, A2 => n11908, B1 => n11912, B2 => 
                           n13512, ZN => n7744);
   U5627 : OAI22_X1 port map( A1 => n10763, A2 => n11908, B1 => n11913, B2 => 
                           n13511, ZN => n7743);
   U5628 : OAI22_X1 port map( A1 => n10756, A2 => n11908, B1 => n11913, B2 => 
                           n13510, ZN => n7742);
   U5629 : OAI22_X1 port map( A1 => n10749, A2 => n11908, B1 => n11913, B2 => 
                           n13509, ZN => n7741);
   U5630 : OAI22_X1 port map( A1 => n10742, A2 => n11908, B1 => n11913, B2 => 
                           n13508, ZN => n7740);
   U5631 : OAI22_X1 port map( A1 => n10735, A2 => n11908, B1 => n11914, B2 => 
                           n13507, ZN => n7739);
   U5632 : OAI22_X1 port map( A1 => n10728, A2 => n11908, B1 => n11914, B2 => 
                           n13506, ZN => n7738);
   U5633 : OAI22_X1 port map( A1 => n10721, A2 => n11908, B1 => n11914, B2 => 
                           n13505, ZN => n7737);
   U5634 : OAI22_X1 port map( A1 => n10714, A2 => n11908, B1 => n11914, B2 => 
                           n13504, ZN => n7736);
   U5635 : OAI22_X1 port map( A1 => n10707, A2 => n11907, B1 => n11915, B2 => 
                           n13503, ZN => n7735);
   U5636 : OAI22_X1 port map( A1 => n10700, A2 => n11907, B1 => n11915, B2 => 
                           n13502, ZN => n7734);
   U5637 : OAI22_X1 port map( A1 => n10693, A2 => n11907, B1 => n11915, B2 => 
                           n13501, ZN => n7733);
   U5638 : OAI22_X1 port map( A1 => n10686, A2 => n11907, B1 => n11915, B2 => 
                           n13500, ZN => n7732);
   U5639 : OAI22_X1 port map( A1 => n10679, A2 => n11907, B1 => n11916, B2 => 
                           n13499, ZN => n7731);
   U5640 : OAI22_X1 port map( A1 => n10672, A2 => n11907, B1 => n11916, B2 => 
                           n13498, ZN => n7730);
   U5641 : OAI22_X1 port map( A1 => n10665, A2 => n11907, B1 => n11916, B2 => 
                           n13497, ZN => n7729);
   U5642 : OAI22_X1 port map( A1 => n10658, A2 => n11907, B1 => n11916, B2 => 
                           n13496, ZN => n7728);
   U5643 : OAI22_X1 port map( A1 => n10651, A2 => n11907, B1 => n11917, B2 => 
                           n13495, ZN => n7727);
   U5644 : OAI22_X1 port map( A1 => n10644, A2 => n11907, B1 => n11917, B2 => 
                           n13494, ZN => n7726);
   U5645 : OAI22_X1 port map( A1 => n10637, A2 => n11907, B1 => n11917, B2 => 
                           n13493, ZN => n7725);
   U5646 : OAI22_X1 port map( A1 => n10630, A2 => n11907, B1 => n11917, B2 => 
                           n13492, ZN => n7724);
   U5647 : OAI22_X1 port map( A1 => n10848, A2 => n11765, B1 => n11766, B2 => 
                           n13395, ZN => n7371);
   U5648 : OAI22_X1 port map( A1 => n10841, A2 => n11765, B1 => n11766, B2 => 
                           n13394, ZN => n7370);
   U5649 : OAI22_X1 port map( A1 => n10834, A2 => n11765, B1 => n11766, B2 => 
                           n13393, ZN => n7369);
   U5650 : OAI22_X1 port map( A1 => n10827, A2 => n11765, B1 => n11766, B2 => 
                           n13392, ZN => n7368);
   U5651 : OAI22_X1 port map( A1 => n10820, A2 => n11765, B1 => n11767, B2 => 
                           n13391, ZN => n7367);
   U5652 : OAI22_X1 port map( A1 => n10813, A2 => n11765, B1 => n11767, B2 => 
                           n13390, ZN => n7366);
   U5653 : OAI22_X1 port map( A1 => n10806, A2 => n11765, B1 => n11767, B2 => 
                           n13389, ZN => n7365);
   U5654 : OAI22_X1 port map( A1 => n10799, A2 => n11765, B1 => n11767, B2 => 
                           n13388, ZN => n7364);
   U5655 : OAI22_X1 port map( A1 => n10792, A2 => n11764, B1 => n11768, B2 => 
                           n13387, ZN => n7363);
   U5656 : OAI22_X1 port map( A1 => n10785, A2 => n11764, B1 => n11768, B2 => 
                           n13386, ZN => n7362);
   U5657 : OAI22_X1 port map( A1 => n10778, A2 => n11764, B1 => n11768, B2 => 
                           n13385, ZN => n7361);
   U5658 : OAI22_X1 port map( A1 => n10771, A2 => n11764, B1 => n11768, B2 => 
                           n13384, ZN => n7360);
   U5659 : OAI22_X1 port map( A1 => n10764, A2 => n11764, B1 => n11769, B2 => 
                           n13383, ZN => n7359);
   U5660 : OAI22_X1 port map( A1 => n10757, A2 => n11764, B1 => n11769, B2 => 
                           n13382, ZN => n7358);
   U5661 : OAI22_X1 port map( A1 => n10750, A2 => n11764, B1 => n11769, B2 => 
                           n13381, ZN => n7357);
   U5662 : OAI22_X1 port map( A1 => n10743, A2 => n11764, B1 => n11769, B2 => 
                           n13380, ZN => n7356);
   U5663 : OAI22_X1 port map( A1 => n10736, A2 => n11764, B1 => n11770, B2 => 
                           n13379, ZN => n7355);
   U5664 : OAI22_X1 port map( A1 => n10729, A2 => n11764, B1 => n11770, B2 => 
                           n13378, ZN => n7354);
   U5665 : OAI22_X1 port map( A1 => n10722, A2 => n11764, B1 => n11770, B2 => 
                           n13377, ZN => n7353);
   U5666 : OAI22_X1 port map( A1 => n10715, A2 => n11764, B1 => n11770, B2 => 
                           n13376, ZN => n7352);
   U5667 : OAI22_X1 port map( A1 => n10708, A2 => n11763, B1 => n11771, B2 => 
                           n13375, ZN => n7351);
   U5668 : OAI22_X1 port map( A1 => n10701, A2 => n11763, B1 => n11771, B2 => 
                           n13374, ZN => n7350);
   U5669 : OAI22_X1 port map( A1 => n10694, A2 => n11763, B1 => n11771, B2 => 
                           n13373, ZN => n7349);
   U5670 : OAI22_X1 port map( A1 => n10687, A2 => n11763, B1 => n11771, B2 => 
                           n13372, ZN => n7348);
   U5671 : OAI22_X1 port map( A1 => n10680, A2 => n11763, B1 => n11772, B2 => 
                           n13371, ZN => n7347);
   U5672 : OAI22_X1 port map( A1 => n10673, A2 => n11763, B1 => n11772, B2 => 
                           n13370, ZN => n7346);
   U5673 : OAI22_X1 port map( A1 => n10666, A2 => n11763, B1 => n11772, B2 => 
                           n13369, ZN => n7345);
   U5674 : OAI22_X1 port map( A1 => n10659, A2 => n11763, B1 => n11772, B2 => 
                           n13368, ZN => n7344);
   U5675 : OAI22_X1 port map( A1 => n10652, A2 => n11763, B1 => n11773, B2 => 
                           n13367, ZN => n7343);
   U5676 : OAI22_X1 port map( A1 => n10645, A2 => n11763, B1 => n11773, B2 => 
                           n13366, ZN => n7342);
   U5677 : OAI22_X1 port map( A1 => n10638, A2 => n11763, B1 => n11773, B2 => 
                           n13365, ZN => n7341);
   U5678 : OAI22_X1 port map( A1 => n10631, A2 => n11763, B1 => n11773, B2 => 
                           n13364, ZN => n7340);
   U5679 : OAI22_X1 port map( A1 => n10806, A2 => n11753, B1 => n11755, B2 => 
                           n13357, ZN => n7333);
   U5680 : OAI22_X1 port map( A1 => n10799, A2 => n11753, B1 => n11755, B2 => 
                           n13356, ZN => n7332);
   U5681 : OAI22_X1 port map( A1 => n10792, A2 => n11752, B1 => n11756, B2 => 
                           n13355, ZN => n7331);
   U5682 : OAI22_X1 port map( A1 => n10785, A2 => n11752, B1 => n11756, B2 => 
                           n13354, ZN => n7330);
   U5683 : OAI22_X1 port map( A1 => n10778, A2 => n11752, B1 => n11756, B2 => 
                           n13353, ZN => n7329);
   U5684 : OAI22_X1 port map( A1 => n10771, A2 => n11752, B1 => n11756, B2 => 
                           n13352, ZN => n7328);
   U5685 : OAI22_X1 port map( A1 => n10764, A2 => n11752, B1 => n11757, B2 => 
                           n13351, ZN => n7327);
   U5686 : OAI22_X1 port map( A1 => n10757, A2 => n11752, B1 => n11757, B2 => 
                           n13350, ZN => n7326);
   U5687 : OAI22_X1 port map( A1 => n10750, A2 => n11752, B1 => n11757, B2 => 
                           n13349, ZN => n7325);
   U5688 : OAI22_X1 port map( A1 => n10743, A2 => n11752, B1 => n11757, B2 => 
                           n13348, ZN => n7324);
   U5689 : OAI22_X1 port map( A1 => n10736, A2 => n11752, B1 => n11758, B2 => 
                           n13347, ZN => n7323);
   U5690 : OAI22_X1 port map( A1 => n10729, A2 => n11752, B1 => n11758, B2 => 
                           n13346, ZN => n7322);
   U5691 : OAI22_X1 port map( A1 => n10722, A2 => n11752, B1 => n11758, B2 => 
                           n13345, ZN => n7321);
   U5692 : OAI22_X1 port map( A1 => n10715, A2 => n11752, B1 => n11758, B2 => 
                           n13344, ZN => n7320);
   U5693 : OAI22_X1 port map( A1 => n10708, A2 => n11751, B1 => n11759, B2 => 
                           n13343, ZN => n7319);
   U5694 : OAI22_X1 port map( A1 => n10701, A2 => n11751, B1 => n11759, B2 => 
                           n13342, ZN => n7318);
   U5695 : OAI22_X1 port map( A1 => n10694, A2 => n11751, B1 => n11759, B2 => 
                           n13341, ZN => n7317);
   U5696 : OAI22_X1 port map( A1 => n10687, A2 => n11751, B1 => n11759, B2 => 
                           n13340, ZN => n7316);
   U5697 : OAI22_X1 port map( A1 => n10680, A2 => n11751, B1 => n11760, B2 => 
                           n13339, ZN => n7315);
   U5698 : OAI22_X1 port map( A1 => n10673, A2 => n11751, B1 => n11760, B2 => 
                           n13338, ZN => n7314);
   U5699 : OAI22_X1 port map( A1 => n10666, A2 => n11751, B1 => n11760, B2 => 
                           n13337, ZN => n7313);
   U5700 : OAI22_X1 port map( A1 => n10659, A2 => n11751, B1 => n11760, B2 => 
                           n13336, ZN => n7312);
   U5701 : OAI22_X1 port map( A1 => n10652, A2 => n11751, B1 => n11761, B2 => 
                           n13335, ZN => n7311);
   U5702 : OAI22_X1 port map( A1 => n10645, A2 => n11751, B1 => n11761, B2 => 
                           n13334, ZN => n7310);
   U5703 : OAI22_X1 port map( A1 => n10638, A2 => n11751, B1 => n11761, B2 => 
                           n13333, ZN => n7309);
   U5704 : OAI22_X1 port map( A1 => n10631, A2 => n11751, B1 => n11761, B2 => 
                           n13332, ZN => n7308);
   U5705 : OAI22_X1 port map( A1 => n10848, A2 => n11741, B1 => n11742, B2 => 
                           n13331, ZN => n7307);
   U5706 : OAI22_X1 port map( A1 => n10841, A2 => n11741, B1 => n11742, B2 => 
                           n13330, ZN => n7306);
   U5707 : OAI22_X1 port map( A1 => n10834, A2 => n11741, B1 => n11742, B2 => 
                           n13329, ZN => n7305);
   U5708 : OAI22_X1 port map( A1 => n10827, A2 => n11741, B1 => n11742, B2 => 
                           n13328, ZN => n7304);
   U5709 : OAI22_X1 port map( A1 => n10820, A2 => n11741, B1 => n11743, B2 => 
                           n13327, ZN => n7303);
   U5710 : OAI22_X1 port map( A1 => n10813, A2 => n11741, B1 => n11743, B2 => 
                           n13326, ZN => n7302);
   U5711 : OAI22_X1 port map( A1 => n10806, A2 => n11741, B1 => n11743, B2 => 
                           n13325, ZN => n7301);
   U5712 : OAI22_X1 port map( A1 => n10799, A2 => n11741, B1 => n11743, B2 => 
                           n13324, ZN => n7300);
   U5713 : OAI22_X1 port map( A1 => n10792, A2 => n11740, B1 => n11744, B2 => 
                           n13323, ZN => n7299);
   U5714 : OAI22_X1 port map( A1 => n10785, A2 => n11740, B1 => n11744, B2 => 
                           n13322, ZN => n7298);
   U5715 : OAI22_X1 port map( A1 => n10778, A2 => n11740, B1 => n11744, B2 => 
                           n13321, ZN => n7297);
   U5716 : OAI22_X1 port map( A1 => n10771, A2 => n11740, B1 => n11744, B2 => 
                           n13320, ZN => n7296);
   U5717 : OAI22_X1 port map( A1 => n10764, A2 => n11740, B1 => n11745, B2 => 
                           n13319, ZN => n7295);
   U5718 : OAI22_X1 port map( A1 => n10757, A2 => n11740, B1 => n11745, B2 => 
                           n13318, ZN => n7294);
   U5719 : OAI22_X1 port map( A1 => n10750, A2 => n11740, B1 => n11745, B2 => 
                           n13317, ZN => n7293);
   U5720 : OAI22_X1 port map( A1 => n10743, A2 => n11740, B1 => n11745, B2 => 
                           n13316, ZN => n7292);
   U5721 : OAI22_X1 port map( A1 => n10736, A2 => n11740, B1 => n11746, B2 => 
                           n13315, ZN => n7291);
   U5722 : OAI22_X1 port map( A1 => n10729, A2 => n11740, B1 => n11746, B2 => 
                           n13314, ZN => n7290);
   U5723 : OAI22_X1 port map( A1 => n10722, A2 => n11740, B1 => n11746, B2 => 
                           n13313, ZN => n7289);
   U5724 : OAI22_X1 port map( A1 => n10715, A2 => n11740, B1 => n11746, B2 => 
                           n13312, ZN => n7288);
   U5725 : OAI22_X1 port map( A1 => n10708, A2 => n11739, B1 => n11747, B2 => 
                           n13311, ZN => n7287);
   U5726 : OAI22_X1 port map( A1 => n10701, A2 => n11739, B1 => n11747, B2 => 
                           n13310, ZN => n7286);
   U5727 : OAI22_X1 port map( A1 => n10694, A2 => n11739, B1 => n11747, B2 => 
                           n13309, ZN => n7285);
   U5728 : OAI22_X1 port map( A1 => n10687, A2 => n11739, B1 => n11747, B2 => 
                           n13308, ZN => n7284);
   U5729 : OAI22_X1 port map( A1 => n10680, A2 => n11739, B1 => n11748, B2 => 
                           n13307, ZN => n7283);
   U5730 : OAI22_X1 port map( A1 => n10673, A2 => n11739, B1 => n11748, B2 => 
                           n13306, ZN => n7282);
   U5731 : OAI22_X1 port map( A1 => n10666, A2 => n11739, B1 => n11748, B2 => 
                           n13305, ZN => n7281);
   U5732 : OAI22_X1 port map( A1 => n10659, A2 => n11739, B1 => n11748, B2 => 
                           n13304, ZN => n7280);
   U5733 : OAI22_X1 port map( A1 => n10652, A2 => n11739, B1 => n11749, B2 => 
                           n13303, ZN => n7279);
   U5734 : OAI22_X1 port map( A1 => n10645, A2 => n11739, B1 => n11749, B2 => 
                           n13302, ZN => n7278);
   U5735 : OAI22_X1 port map( A1 => n10638, A2 => n11739, B1 => n11749, B2 => 
                           n13301, ZN => n7277);
   U5736 : OAI22_X1 port map( A1 => n10631, A2 => n11739, B1 => n11749, B2 => 
                           n13300, ZN => n7276);
   U5737 : OAI22_X1 port map( A1 => n10848, A2 => n11729, B1 => n11730, B2 => 
                           n13299, ZN => n7275);
   U5738 : OAI22_X1 port map( A1 => n10841, A2 => n11729, B1 => n11730, B2 => 
                           n13298, ZN => n7274);
   U5739 : OAI22_X1 port map( A1 => n10834, A2 => n11729, B1 => n11730, B2 => 
                           n13297, ZN => n7273);
   U5740 : OAI22_X1 port map( A1 => n10827, A2 => n11729, B1 => n11730, B2 => 
                           n13296, ZN => n7272);
   U5741 : OAI22_X1 port map( A1 => n10820, A2 => n11729, B1 => n11731, B2 => 
                           n13295, ZN => n7271);
   U5742 : OAI22_X1 port map( A1 => n10813, A2 => n11729, B1 => n11731, B2 => 
                           n13294, ZN => n7270);
   U5743 : OAI22_X1 port map( A1 => n10806, A2 => n11729, B1 => n11731, B2 => 
                           n13293, ZN => n7269);
   U5744 : OAI22_X1 port map( A1 => n10799, A2 => n11729, B1 => n11731, B2 => 
                           n13292, ZN => n7268);
   U5745 : OAI22_X1 port map( A1 => n10792, A2 => n11728, B1 => n11732, B2 => 
                           n13291, ZN => n7267);
   U5746 : OAI22_X1 port map( A1 => n10785, A2 => n11728, B1 => n11732, B2 => 
                           n13290, ZN => n7266);
   U5747 : OAI22_X1 port map( A1 => n10778, A2 => n11728, B1 => n11732, B2 => 
                           n13289, ZN => n7265);
   U5748 : OAI22_X1 port map( A1 => n10771, A2 => n11728, B1 => n11732, B2 => 
                           n13288, ZN => n7264);
   U5749 : OAI22_X1 port map( A1 => n10764, A2 => n11728, B1 => n11733, B2 => 
                           n13287, ZN => n7263);
   U5750 : OAI22_X1 port map( A1 => n10757, A2 => n11728, B1 => n11733, B2 => 
                           n13286, ZN => n7262);
   U5751 : OAI22_X1 port map( A1 => n10750, A2 => n11728, B1 => n11733, B2 => 
                           n13285, ZN => n7261);
   U5752 : OAI22_X1 port map( A1 => n10743, A2 => n11728, B1 => n11733, B2 => 
                           n13284, ZN => n7260);
   U5753 : OAI22_X1 port map( A1 => n10736, A2 => n11728, B1 => n11734, B2 => 
                           n13283, ZN => n7259);
   U5754 : OAI22_X1 port map( A1 => n10729, A2 => n11728, B1 => n11734, B2 => 
                           n13282, ZN => n7258);
   U5755 : OAI22_X1 port map( A1 => n10722, A2 => n11728, B1 => n11734, B2 => 
                           n13281, ZN => n7257);
   U5756 : OAI22_X1 port map( A1 => n10715, A2 => n11728, B1 => n11734, B2 => 
                           n13280, ZN => n7256);
   U5757 : OAI22_X1 port map( A1 => n10708, A2 => n11727, B1 => n11735, B2 => 
                           n13279, ZN => n7255);
   U5758 : OAI22_X1 port map( A1 => n10701, A2 => n11727, B1 => n11735, B2 => 
                           n13278, ZN => n7254);
   U5759 : OAI22_X1 port map( A1 => n10694, A2 => n11727, B1 => n11735, B2 => 
                           n13277, ZN => n7253);
   U5760 : OAI22_X1 port map( A1 => n10687, A2 => n11727, B1 => n11735, B2 => 
                           n13276, ZN => n7252);
   U5761 : OAI22_X1 port map( A1 => n10680, A2 => n11727, B1 => n11736, B2 => 
                           n13275, ZN => n7251);
   U5762 : OAI22_X1 port map( A1 => n10673, A2 => n11727, B1 => n11736, B2 => 
                           n13274, ZN => n7250);
   U5763 : OAI22_X1 port map( A1 => n10666, A2 => n11727, B1 => n11736, B2 => 
                           n13273, ZN => n7249);
   U5764 : OAI22_X1 port map( A1 => n10659, A2 => n11727, B1 => n11736, B2 => 
                           n13272, ZN => n7248);
   U5765 : OAI22_X1 port map( A1 => n10652, A2 => n11727, B1 => n11737, B2 => 
                           n13271, ZN => n7247);
   U5766 : OAI22_X1 port map( A1 => n10645, A2 => n11727, B1 => n11737, B2 => 
                           n13270, ZN => n7246);
   U5767 : OAI22_X1 port map( A1 => n10638, A2 => n11727, B1 => n11737, B2 => 
                           n13269, ZN => n7245);
   U5768 : OAI22_X1 port map( A1 => n10631, A2 => n11727, B1 => n11737, B2 => 
                           n13268, ZN => n7244);
   U5769 : OAI22_X1 port map( A1 => n10848, A2 => n11717, B1 => n11718, B2 => 
                           n13267, ZN => n7243);
   U5770 : OAI22_X1 port map( A1 => n10841, A2 => n11717, B1 => n11718, B2 => 
                           n13266, ZN => n7242);
   U5771 : OAI22_X1 port map( A1 => n10834, A2 => n11717, B1 => n11718, B2 => 
                           n13265, ZN => n7241);
   U5772 : OAI22_X1 port map( A1 => n10827, A2 => n11717, B1 => n11718, B2 => 
                           n13264, ZN => n7240);
   U5773 : OAI22_X1 port map( A1 => n10820, A2 => n11717, B1 => n11719, B2 => 
                           n13263, ZN => n7239);
   U5774 : OAI22_X1 port map( A1 => n10813, A2 => n11717, B1 => n11719, B2 => 
                           n13262, ZN => n7238);
   U5775 : OAI22_X1 port map( A1 => n10806, A2 => n11717, B1 => n11719, B2 => 
                           n13261, ZN => n7237);
   U5776 : OAI22_X1 port map( A1 => n10799, A2 => n11717, B1 => n11719, B2 => 
                           n13260, ZN => n7236);
   U5777 : OAI22_X1 port map( A1 => n10792, A2 => n11716, B1 => n11720, B2 => 
                           n13259, ZN => n7235);
   U5778 : OAI22_X1 port map( A1 => n10785, A2 => n11716, B1 => n11720, B2 => 
                           n13258, ZN => n7234);
   U5779 : OAI22_X1 port map( A1 => n10778, A2 => n11716, B1 => n11720, B2 => 
                           n13257, ZN => n7233);
   U5780 : OAI22_X1 port map( A1 => n10771, A2 => n11716, B1 => n11720, B2 => 
                           n13256, ZN => n7232);
   U5781 : OAI22_X1 port map( A1 => n10764, A2 => n11716, B1 => n11721, B2 => 
                           n13255, ZN => n7231);
   U5782 : OAI22_X1 port map( A1 => n10757, A2 => n11716, B1 => n11721, B2 => 
                           n13254, ZN => n7230);
   U5783 : OAI22_X1 port map( A1 => n10750, A2 => n11716, B1 => n11721, B2 => 
                           n13253, ZN => n7229);
   U5784 : OAI22_X1 port map( A1 => n10743, A2 => n11716, B1 => n11721, B2 => 
                           n13252, ZN => n7228);
   U5785 : OAI22_X1 port map( A1 => n10736, A2 => n11716, B1 => n11722, B2 => 
                           n13251, ZN => n7227);
   U5786 : OAI22_X1 port map( A1 => n10729, A2 => n11716, B1 => n11722, B2 => 
                           n13250, ZN => n7226);
   U5787 : OAI22_X1 port map( A1 => n10722, A2 => n11716, B1 => n11722, B2 => 
                           n13249, ZN => n7225);
   U5788 : OAI22_X1 port map( A1 => n10715, A2 => n11716, B1 => n11722, B2 => 
                           n13248, ZN => n7224);
   U5789 : OAI22_X1 port map( A1 => n10708, A2 => n11715, B1 => n11723, B2 => 
                           n13247, ZN => n7223);
   U5790 : OAI22_X1 port map( A1 => n10701, A2 => n11715, B1 => n11723, B2 => 
                           n13246, ZN => n7222);
   U5791 : OAI22_X1 port map( A1 => n10694, A2 => n11715, B1 => n11723, B2 => 
                           n13245, ZN => n7221);
   U5792 : OAI22_X1 port map( A1 => n10687, A2 => n11715, B1 => n11723, B2 => 
                           n13244, ZN => n7220);
   U5793 : OAI22_X1 port map( A1 => n10680, A2 => n11715, B1 => n11724, B2 => 
                           n13243, ZN => n7219);
   U5794 : OAI22_X1 port map( A1 => n10673, A2 => n11715, B1 => n11724, B2 => 
                           n13242, ZN => n7218);
   U5795 : OAI22_X1 port map( A1 => n10666, A2 => n11715, B1 => n11724, B2 => 
                           n13241, ZN => n7217);
   U5796 : OAI22_X1 port map( A1 => n10659, A2 => n11715, B1 => n11724, B2 => 
                           n13240, ZN => n7216);
   U5797 : OAI22_X1 port map( A1 => n10652, A2 => n11715, B1 => n11725, B2 => 
                           n13239, ZN => n7215);
   U5798 : OAI22_X1 port map( A1 => n10645, A2 => n11715, B1 => n11725, B2 => 
                           n13238, ZN => n7214);
   U5799 : OAI22_X1 port map( A1 => n10638, A2 => n11715, B1 => n11725, B2 => 
                           n13237, ZN => n7213);
   U5800 : OAI22_X1 port map( A1 => n10631, A2 => n11715, B1 => n11725, B2 => 
                           n13236, ZN => n7212);
   U5801 : OAI22_X1 port map( A1 => n10848, A2 => n11705, B1 => n11706, B2 => 
                           n13235, ZN => n7211);
   U5802 : OAI22_X1 port map( A1 => n10841, A2 => n11705, B1 => n11706, B2 => 
                           n13234, ZN => n7210);
   U5803 : OAI22_X1 port map( A1 => n10834, A2 => n11705, B1 => n11706, B2 => 
                           n13233, ZN => n7209);
   U5804 : OAI22_X1 port map( A1 => n10827, A2 => n11705, B1 => n11706, B2 => 
                           n13232, ZN => n7208);
   U5805 : OAI22_X1 port map( A1 => n10820, A2 => n11705, B1 => n11707, B2 => 
                           n13231, ZN => n7207);
   U5806 : OAI22_X1 port map( A1 => n10813, A2 => n11705, B1 => n11707, B2 => 
                           n13230, ZN => n7206);
   U5807 : OAI22_X1 port map( A1 => n10806, A2 => n11705, B1 => n11707, B2 => 
                           n13229, ZN => n7205);
   U5808 : OAI22_X1 port map( A1 => n10799, A2 => n11705, B1 => n11707, B2 => 
                           n13228, ZN => n7204);
   U5809 : OAI22_X1 port map( A1 => n10792, A2 => n11704, B1 => n11708, B2 => 
                           n13227, ZN => n7203);
   U5810 : OAI22_X1 port map( A1 => n10785, A2 => n11704, B1 => n11708, B2 => 
                           n13226, ZN => n7202);
   U5811 : OAI22_X1 port map( A1 => n10778, A2 => n11704, B1 => n11708, B2 => 
                           n13225, ZN => n7201);
   U5812 : OAI22_X1 port map( A1 => n10771, A2 => n11704, B1 => n11708, B2 => 
                           n13224, ZN => n7200);
   U5813 : OAI22_X1 port map( A1 => n10764, A2 => n11704, B1 => n11709, B2 => 
                           n13223, ZN => n7199);
   U5814 : OAI22_X1 port map( A1 => n10757, A2 => n11704, B1 => n11709, B2 => 
                           n13222, ZN => n7198);
   U5815 : OAI22_X1 port map( A1 => n10750, A2 => n11704, B1 => n11709, B2 => 
                           n13221, ZN => n7197);
   U5816 : OAI22_X1 port map( A1 => n10743, A2 => n11704, B1 => n11709, B2 => 
                           n13220, ZN => n7196);
   U5817 : OAI22_X1 port map( A1 => n10736, A2 => n11704, B1 => n11710, B2 => 
                           n13219, ZN => n7195);
   U5818 : OAI22_X1 port map( A1 => n10729, A2 => n11704, B1 => n11710, B2 => 
                           n13218, ZN => n7194);
   U5819 : OAI22_X1 port map( A1 => n10722, A2 => n11704, B1 => n11710, B2 => 
                           n13217, ZN => n7193);
   U5820 : OAI22_X1 port map( A1 => n10715, A2 => n11704, B1 => n11710, B2 => 
                           n13216, ZN => n7192);
   U5821 : OAI22_X1 port map( A1 => n10708, A2 => n11703, B1 => n11711, B2 => 
                           n13215, ZN => n7191);
   U5822 : OAI22_X1 port map( A1 => n10701, A2 => n11703, B1 => n11711, B2 => 
                           n13214, ZN => n7190);
   U5823 : OAI22_X1 port map( A1 => n10694, A2 => n11703, B1 => n11711, B2 => 
                           n13213, ZN => n7189);
   U5824 : OAI22_X1 port map( A1 => n10687, A2 => n11703, B1 => n11711, B2 => 
                           n13212, ZN => n7188);
   U5826 : OAI22_X1 port map( A1 => n10680, A2 => n11703, B1 => n11712, B2 => 
                           n13211, ZN => n7187);
   U5827 : OAI22_X1 port map( A1 => n10673, A2 => n11703, B1 => n11712, B2 => 
                           n13210, ZN => n7186);
   U5828 : OAI22_X1 port map( A1 => n10666, A2 => n11703, B1 => n11712, B2 => 
                           n13209, ZN => n7185);
   U5829 : OAI22_X1 port map( A1 => n10659, A2 => n11703, B1 => n11712, B2 => 
                           n13208, ZN => n7184);
   U5830 : OAI22_X1 port map( A1 => n10652, A2 => n11703, B1 => n11713, B2 => 
                           n13207, ZN => n7183);
   U5831 : OAI22_X1 port map( A1 => n10645, A2 => n11703, B1 => n11713, B2 => 
                           n13206, ZN => n7182);
   U5832 : OAI22_X1 port map( A1 => n10638, A2 => n11703, B1 => n11713, B2 => 
                           n13205, ZN => n7181);
   U5833 : OAI22_X1 port map( A1 => n10631, A2 => n11703, B1 => n11713, B2 => 
                           n13204, ZN => n7180);
   U5834 : OAI22_X1 port map( A1 => n10848, A2 => n11657, B1 => n11658, B2 => 
                           n13107, ZN => n7083);
   U5835 : OAI22_X1 port map( A1 => n10841, A2 => n11657, B1 => n11658, B2 => 
                           n13106, ZN => n7082);
   U5836 : OAI22_X1 port map( A1 => n10834, A2 => n11657, B1 => n11658, B2 => 
                           n13105, ZN => n7081);
   U5837 : OAI22_X1 port map( A1 => n10827, A2 => n11657, B1 => n11658, B2 => 
                           n13104, ZN => n7080);
   U5838 : OAI22_X1 port map( A1 => n10820, A2 => n11657, B1 => n11659, B2 => 
                           n13103, ZN => n7079);
   U5839 : OAI22_X1 port map( A1 => n10813, A2 => n11657, B1 => n11659, B2 => 
                           n13102, ZN => n7078);
   U5840 : OAI22_X1 port map( A1 => n10806, A2 => n11657, B1 => n11659, B2 => 
                           n13101, ZN => n7077);
   U5841 : OAI22_X1 port map( A1 => n10799, A2 => n11657, B1 => n11659, B2 => 
                           n13100, ZN => n7076);
   U5842 : OAI22_X1 port map( A1 => n10792, A2 => n11656, B1 => n11660, B2 => 
                           n13099, ZN => n7075);
   U5843 : OAI22_X1 port map( A1 => n10785, A2 => n11656, B1 => n11660, B2 => 
                           n13098, ZN => n7074);
   U5844 : OAI22_X1 port map( A1 => n10778, A2 => n11656, B1 => n11660, B2 => 
                           n13097, ZN => n7073);
   U5845 : OAI22_X1 port map( A1 => n10771, A2 => n11656, B1 => n11660, B2 => 
                           n13096, ZN => n7072);
   U5846 : OAI22_X1 port map( A1 => n10764, A2 => n11656, B1 => n11661, B2 => 
                           n13095, ZN => n7071);
   U5847 : OAI22_X1 port map( A1 => n10757, A2 => n11656, B1 => n11661, B2 => 
                           n13094, ZN => n7070);
   U5848 : OAI22_X1 port map( A1 => n10750, A2 => n11656, B1 => n11661, B2 => 
                           n13093, ZN => n7069);
   U5849 : OAI22_X1 port map( A1 => n10743, A2 => n11656, B1 => n11661, B2 => 
                           n13092, ZN => n7068);
   U5850 : OAI22_X1 port map( A1 => n10736, A2 => n11656, B1 => n11662, B2 => 
                           n13091, ZN => n7067);
   U5851 : OAI22_X1 port map( A1 => n10729, A2 => n11656, B1 => n11662, B2 => 
                           n13090, ZN => n7066);
   U5852 : OAI22_X1 port map( A1 => n10722, A2 => n11656, B1 => n11662, B2 => 
                           n13089, ZN => n7065);
   U5853 : OAI22_X1 port map( A1 => n10715, A2 => n11656, B1 => n11662, B2 => 
                           n13088, ZN => n7064);
   U5854 : OAI22_X1 port map( A1 => n10708, A2 => n11655, B1 => n11663, B2 => 
                           n13087, ZN => n7063);
   U5855 : OAI22_X1 port map( A1 => n10701, A2 => n11655, B1 => n11663, B2 => 
                           n13086, ZN => n7062);
   U5856 : OAI22_X1 port map( A1 => n10694, A2 => n11655, B1 => n11663, B2 => 
                           n13085, ZN => n7061);
   U5857 : OAI22_X1 port map( A1 => n10687, A2 => n11655, B1 => n11663, B2 => 
                           n13084, ZN => n7060);
   U5858 : OAI22_X1 port map( A1 => n10680, A2 => n11655, B1 => n11664, B2 => 
                           n13083, ZN => n7059);
   U5859 : OAI22_X1 port map( A1 => n10673, A2 => n11655, B1 => n11664, B2 => 
                           n13082, ZN => n7058);
   U5860 : OAI22_X1 port map( A1 => n10666, A2 => n11655, B1 => n11664, B2 => 
                           n13081, ZN => n7057);
   U5861 : OAI22_X1 port map( A1 => n10659, A2 => n11655, B1 => n11664, B2 => 
                           n13080, ZN => n7056);
   U5862 : OAI22_X1 port map( A1 => n10652, A2 => n11655, B1 => n11665, B2 => 
                           n13079, ZN => n7055);
   U5863 : OAI22_X1 port map( A1 => n10645, A2 => n11655, B1 => n11665, B2 => 
                           n13078, ZN => n7054);
   U5864 : OAI22_X1 port map( A1 => n10638, A2 => n11655, B1 => n11665, B2 => 
                           n13077, ZN => n7053);
   U5865 : OAI22_X1 port map( A1 => n10631, A2 => n11655, B1 => n11665, B2 => 
                           n13076, ZN => n7052);
   U5866 : OAI22_X1 port map( A1 => n10849, A2 => n11645, B1 => n11650, B2 => 
                           n13075, ZN => n7051);
   U5867 : OAI22_X1 port map( A1 => n10842, A2 => n11645, B1 => n11653, B2 => 
                           n13074, ZN => n7050);
   U5868 : OAI22_X1 port map( A1 => n10835, A2 => n11645, B1 => n11653, B2 => 
                           n13073, ZN => n7049);
   U5869 : OAI22_X1 port map( A1 => n10828, A2 => n11645, B1 => n11653, B2 => 
                           n13072, ZN => n7048);
   U5870 : OAI22_X1 port map( A1 => n10821, A2 => n11645, B1 => n11652, B2 => 
                           n13071, ZN => n7047);
   U5871 : OAI22_X1 port map( A1 => n10814, A2 => n11645, B1 => n11653, B2 => 
                           n13070, ZN => n7046);
   U5872 : OAI22_X1 port map( A1 => n10807, A2 => n11645, B1 => n11652, B2 => 
                           n13069, ZN => n7045);
   U5873 : OAI22_X1 port map( A1 => n10800, A2 => n11645, B1 => n11652, B2 => 
                           n13068, ZN => n7044);
   U5874 : OAI22_X1 port map( A1 => n10793, A2 => n11644, B1 => n11651, B2 => 
                           n13067, ZN => n7043);
   U5875 : OAI22_X1 port map( A1 => n10786, A2 => n11644, B1 => n11652, B2 => 
                           n13066, ZN => n7042);
   U5876 : OAI22_X1 port map( A1 => n10779, A2 => n11644, B1 => n11651, B2 => 
                           n13065, ZN => n7041);
   U5877 : OAI22_X1 port map( A1 => n10772, A2 => n11644, B1 => n11651, B2 => 
                           n13064, ZN => n7040);
   U5878 : OAI22_X1 port map( A1 => n10765, A2 => n11644, B1 => n11650, B2 => 
                           n13063, ZN => n7039);
   U5879 : OAI22_X1 port map( A1 => n10758, A2 => n11644, B1 => n11651, B2 => 
                           n13062, ZN => n7038);
   U5880 : OAI22_X1 port map( A1 => n10751, A2 => n11644, B1 => n11650, B2 => 
                           n13061, ZN => n7037);
   U5881 : OAI22_X1 port map( A1 => n10744, A2 => n11644, B1 => n11650, B2 => 
                           n13060, ZN => n7036);
   U5882 : AOI21_X1 port map( B1 => n2937, B2 => n2936, A => n14518, ZN => 
                           n2488);
   U5883 : OAI22_X1 port map( A1 => n12419, A2 => n10844, B1 => n2913, B2 => 
                           n12418, ZN => n9131);
   U5884 : OAI22_X1 port map( A1 => n12419, A2 => n10837, B1 => n2912, B2 => 
                           n12418, ZN => n9130);
   U5885 : OAI22_X1 port map( A1 => n12419, A2 => n10830, B1 => n2911, B2 => 
                           n12418, ZN => n9129);
   U5886 : OAI22_X1 port map( A1 => n12419, A2 => n10823, B1 => n2910, B2 => 
                           n12418, ZN => n9128);
   U5887 : OAI22_X1 port map( A1 => n12419, A2 => n10816, B1 => n2909, B2 => 
                           n12418, ZN => n9127);
   U5888 : OAI22_X1 port map( A1 => n12420, A2 => n10809, B1 => n2908, B2 => 
                           n12418, ZN => n9126);
   U5889 : OAI22_X1 port map( A1 => n12420, A2 => n10802, B1 => n2907, B2 => 
                           n12418, ZN => n9125);
   U5890 : OAI22_X1 port map( A1 => n12420, A2 => n10795, B1 => n2906, B2 => 
                           n12418, ZN => n9124);
   U5891 : OAI22_X1 port map( A1 => n12420, A2 => n10788, B1 => n2905, B2 => 
                           n12417, ZN => n9123);
   U5892 : OAI22_X1 port map( A1 => n12420, A2 => n10781, B1 => n2904, B2 => 
                           n12417, ZN => n9122);
   U5893 : OAI22_X1 port map( A1 => n12421, A2 => n10774, B1 => n2903, B2 => 
                           n12417, ZN => n9121);
   U5894 : OAI22_X1 port map( A1 => n12421, A2 => n10767, B1 => n2902, B2 => 
                           n12417, ZN => n9120);
   U5895 : OAI22_X1 port map( A1 => n12421, A2 => n10760, B1 => n2901, B2 => 
                           n12417, ZN => n9119);
   U5896 : OAI22_X1 port map( A1 => n12421, A2 => n10753, B1 => n2900, B2 => 
                           n12417, ZN => n9118);
   U5897 : OAI22_X1 port map( A1 => n12421, A2 => n10746, B1 => n2899, B2 => 
                           n12417, ZN => n9117);
   U5898 : OAI22_X1 port map( A1 => n12422, A2 => n10739, B1 => n2898, B2 => 
                           n12417, ZN => n9116);
   U5899 : OAI22_X1 port map( A1 => n12422, A2 => n10732, B1 => n2897, B2 => 
                           n12417, ZN => n9115);
   U5900 : OAI22_X1 port map( A1 => n12422, A2 => n10725, B1 => n2896, B2 => 
                           n12417, ZN => n9114);
   U5901 : OAI22_X1 port map( A1 => n12422, A2 => n10718, B1 => n2895, B2 => 
                           n12417, ZN => n9113);
   U5902 : OAI22_X1 port map( A1 => n12422, A2 => n10711, B1 => n2894, B2 => 
                           n12417, ZN => n9112);
   U5903 : OAI22_X1 port map( A1 => n12423, A2 => n10704, B1 => n2893, B2 => 
                           n12416, ZN => n9111);
   U5904 : OAI22_X1 port map( A1 => n12423, A2 => n10697, B1 => n2892, B2 => 
                           n12416, ZN => n9110);
   U5905 : OAI22_X1 port map( A1 => n12423, A2 => n10690, B1 => n2891, B2 => 
                           n12416, ZN => n9109);
   U5906 : OAI22_X1 port map( A1 => n12423, A2 => n10683, B1 => n2890, B2 => 
                           n12416, ZN => n9108);
   U5907 : OAI22_X1 port map( A1 => n12423, A2 => n10676, B1 => n2889, B2 => 
                           n12416, ZN => n9107);
   U5908 : OAI22_X1 port map( A1 => n12424, A2 => n10669, B1 => n2888, B2 => 
                           n12416, ZN => n9106);
   U5909 : OAI22_X1 port map( A1 => n12424, A2 => n10662, B1 => n2887, B2 => 
                           n12416, ZN => n9105);
   U5910 : OAI22_X1 port map( A1 => n12424, A2 => n10655, B1 => n2886, B2 => 
                           n12416, ZN => n9104);
   U5911 : OAI22_X1 port map( A1 => n12424, A2 => n10648, B1 => n2885, B2 => 
                           n12416, ZN => n9103);
   U5912 : OAI22_X1 port map( A1 => n12424, A2 => n10641, B1 => n2884, B2 => 
                           n12416, ZN => n9102);
   U5913 : OAI22_X1 port map( A1 => n12425, A2 => n10634, B1 => n2883, B2 => 
                           n12416, ZN => n9101);
   U5914 : OAI22_X1 port map( A1 => n12425, A2 => n10627, B1 => n2882, B2 => 
                           n12416, ZN => n9100);
   U5915 : INV_X1 port map( A => RETRN, ZN => n14518);
   U5916 : NAND2_X1 port map( A1 => U3_U98_Z_5, A2 => r480_carry_5_port, ZN => 
                           r480_n4);
   U5917 : NOR2_X1 port map( A1 => n2935, A2 => r480_A_3_port, ZN => U3_U98_Z_6
                           );
   U5918 : NAND2_X1 port map( A1 => U3_U99_Z_5, A2 => r486_carry_5_port, ZN => 
                           r486_n4);
   U5919 : NOR2_X1 port map( A1 => n2935, A2 => r486_A_3_port, ZN => U3_U99_Z_6
                           );
   U5920 : NOR2_X2 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n5647);
   U5921 : NOR2_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n4214);
   U5922 : NOR2_X2 port map( A1 => n14513, A2 => ADD_RD1(2), ZN => n5649);
   U5923 : NOR2_X2 port map( A1 => n14515, A2 => ADD_RD2(2), ZN => n4216);
   U5924 : NOR3_X1 port map( A1 => n12769, A2 => ADD_RD1(0), A3 => n12771, ZN 
                           => n5705);
   U5925 : NOR3_X1 port map( A1 => n12773, A2 => ADD_RD2(0), A3 => n12775, ZN 
                           => n4272);
   U5926 : AOI222_X1 port map( A1 => n10998, A2 => n9728, B1 => n10995, B2 => 
                           n9664, C1 => n10992, C2 => n13363, ZN => n5667);
   U5927 : AOI222_X1 port map( A1 => n10932, A2 => n9280, B1 => n10929, B2 => 
                           n9216, C1 => n10926, C2 => n13811, ZN => n5680);
   U5928 : AOI222_X1 port map( A1 => n11262, A2 => n9728, B1 => n11259, B2 => 
                           n9664, C1 => n11256, C2 => n13363, ZN => n4234);
   U5929 : AOI222_X1 port map( A1 => n11196, A2 => n9280, B1 => n11193, B2 => 
                           n9216, C1 => n11190, C2 => n13811, ZN => n4247);
   U5930 : AOI222_X1 port map( A1 => n10998, A2 => n9729, B1 => n10995, B2 => 
                           n9665, C1 => n10992, C2 => n13362, ZN => n5607);
   U5931 : AOI222_X1 port map( A1 => n10932, A2 => n9281, B1 => n10929, B2 => 
                           n9217, C1 => n10926, C2 => n13810, ZN => n5616);
   U5932 : AOI222_X1 port map( A1 => n11262, A2 => n9729, B1 => n11259, B2 => 
                           n9665, C1 => n11256, C2 => n13362, ZN => n4174);
   U5933 : AOI222_X1 port map( A1 => n11196, A2 => n9281, B1 => n11193, B2 => 
                           n9217, C1 => n11190, C2 => n13810, ZN => n4183);
   U5934 : AOI222_X1 port map( A1 => n10998, A2 => n9730, B1 => n10995, B2 => 
                           n9666, C1 => n10992, C2 => n13361, ZN => n5566);
   U5935 : AOI222_X1 port map( A1 => n10932, A2 => n9282, B1 => n10929, B2 => 
                           n9218, C1 => n10926, C2 => n13809, ZN => n5575);
   U5936 : AOI222_X1 port map( A1 => n11262, A2 => n9730, B1 => n11259, B2 => 
                           n9666, C1 => n11256, C2 => n13361, ZN => n4133);
   U5937 : AOI222_X1 port map( A1 => n11196, A2 => n9282, B1 => n11193, B2 => 
                           n9218, C1 => n11190, C2 => n13809, ZN => n4142);
   U5938 : AOI222_X1 port map( A1 => n10998, A2 => n9731, B1 => n10995, B2 => 
                           n9667, C1 => n10992, C2 => n13360, ZN => n5525);
   U5939 : AOI222_X1 port map( A1 => n10932, A2 => n9283, B1 => n10929, B2 => 
                           n9219, C1 => n10926, C2 => n13808, ZN => n5534);
   U5940 : AOI222_X1 port map( A1 => n11262, A2 => n9731, B1 => n11259, B2 => 
                           n9667, C1 => n11256, C2 => n13360, ZN => n4092);
   U5941 : AOI222_X1 port map( A1 => n11196, A2 => n9283, B1 => n11193, B2 => 
                           n9219, C1 => n11190, C2 => n13808, ZN => n4101);
   U5942 : AOI222_X1 port map( A1 => n10998, A2 => n9732, B1 => n10995, B2 => 
                           n9668, C1 => n10992, C2 => n13359, ZN => n5484);
   U5943 : AOI222_X1 port map( A1 => n10932, A2 => n9284, B1 => n10929, B2 => 
                           n9220, C1 => n10926, C2 => n13807, ZN => n5493);
   U5944 : AOI222_X1 port map( A1 => n11262, A2 => n9732, B1 => n11259, B2 => 
                           n9668, C1 => n11256, C2 => n13359, ZN => n4051);
   U5945 : AOI222_X1 port map( A1 => n11196, A2 => n9284, B1 => n11193, B2 => 
                           n9220, C1 => n11190, C2 => n13807, ZN => n4060);
   U5946 : AOI222_X1 port map( A1 => n10998, A2 => n9733, B1 => n10995, B2 => 
                           n9669, C1 => n10992, C2 => n13358, ZN => n5443);
   U5947 : AOI222_X1 port map( A1 => n10932, A2 => n9285, B1 => n10929, B2 => 
                           n9221, C1 => n10926, C2 => n13806, ZN => n5452);
   U5948 : AOI222_X1 port map( A1 => n11262, A2 => n9733, B1 => n11259, B2 => 
                           n9669, C1 => n11256, C2 => n13358, ZN => n4010);
   U5949 : AOI222_X1 port map( A1 => n11196, A2 => n9285, B1 => n11193, B2 => 
                           n9221, C1 => n11190, C2 => n13806, ZN => n4019);
   U5950 : AOI222_X1 port map( A1 => n10998, A2 => n9734, B1 => n10995, B2 => 
                           n9670, C1 => n10992, C2 => n9702, ZN => n5402);
   U5951 : AOI222_X1 port map( A1 => n10932, A2 => n9286, B1 => n10929, B2 => 
                           n9222, C1 => n10926, C2 => n13805, ZN => n5411);
   U5952 : AOI222_X1 port map( A1 => n11262, A2 => n9734, B1 => n11259, B2 => 
                           n9670, C1 => n11256, C2 => n9702, ZN => n3969);
   U5953 : AOI222_X1 port map( A1 => n11196, A2 => n9286, B1 => n11193, B2 => 
                           n9222, C1 => n11190, C2 => n13805, ZN => n3978);
   U5954 : AOI222_X1 port map( A1 => n10998, A2 => n9735, B1 => n10995, B2 => 
                           n9671, C1 => n10992, C2 => n9703, ZN => n5361);
   U5955 : AOI222_X1 port map( A1 => n10932, A2 => n9287, B1 => n10929, B2 => 
                           n9223, C1 => n10926, C2 => n13804, ZN => n5370);
   U5956 : AOI222_X1 port map( A1 => n11262, A2 => n9735, B1 => n11259, B2 => 
                           n9671, C1 => n11256, C2 => n9703, ZN => n3928);
   U5957 : AOI222_X1 port map( A1 => n11196, A2 => n9287, B1 => n11193, B2 => 
                           n9223, C1 => n11190, C2 => n13804, ZN => n3937);
   U5958 : AOI222_X1 port map( A1 => n10998, A2 => n9736, B1 => n10995, B2 => 
                           n9672, C1 => n10992, C2 => n9704, ZN => n5320);
   U5959 : AOI222_X1 port map( A1 => n10932, A2 => n9288, B1 => n10929, B2 => 
                           n9224, C1 => n10926, C2 => n13803, ZN => n5329);
   U5960 : AOI222_X1 port map( A1 => n11262, A2 => n9736, B1 => n11259, B2 => 
                           n9672, C1 => n11256, C2 => n9704, ZN => n3887);
   U5961 : AOI222_X1 port map( A1 => n11196, A2 => n9288, B1 => n11193, B2 => 
                           n9224, C1 => n11190, C2 => n13803, ZN => n3896);
   U5962 : AOI222_X1 port map( A1 => n10998, A2 => n9737, B1 => n10995, B2 => 
                           n9673, C1 => n10992, C2 => n9705, ZN => n5279);
   U5963 : AOI222_X1 port map( A1 => n10932, A2 => n9289, B1 => n10929, B2 => 
                           n9225, C1 => n10926, C2 => n13802, ZN => n5288);
   U5964 : AOI222_X1 port map( A1 => n11262, A2 => n9737, B1 => n11259, B2 => 
                           n9673, C1 => n11256, C2 => n9705, ZN => n3846);
   U5965 : AOI222_X1 port map( A1 => n11196, A2 => n9289, B1 => n11193, B2 => 
                           n9225, C1 => n11190, C2 => n13802, ZN => n3855);
   U5966 : AOI222_X1 port map( A1 => n10998, A2 => n9738, B1 => n10995, B2 => 
                           n9674, C1 => n10992, C2 => n9706, ZN => n5238);
   U5967 : AOI222_X1 port map( A1 => n10932, A2 => n9290, B1 => n10929, B2 => 
                           n9226, C1 => n10926, C2 => n13801, ZN => n5247);
   U5968 : AOI222_X1 port map( A1 => n11262, A2 => n9738, B1 => n11259, B2 => 
                           n9674, C1 => n11256, C2 => n9706, ZN => n3805);
   U5969 : AOI222_X1 port map( A1 => n11196, A2 => n9290, B1 => n11193, B2 => 
                           n9226, C1 => n11190, C2 => n13801, ZN => n3814);
   U5970 : AOI222_X1 port map( A1 => n10998, A2 => n9739, B1 => n10995, B2 => 
                           n9675, C1 => n10992, C2 => n9707, ZN => n5197);
   U5971 : AOI222_X1 port map( A1 => n10932, A2 => n9291, B1 => n10929, B2 => 
                           n9227, C1 => n10926, C2 => n13800, ZN => n5206);
   U5972 : AOI222_X1 port map( A1 => n11262, A2 => n9739, B1 => n11259, B2 => 
                           n9675, C1 => n11256, C2 => n9707, ZN => n3764);
   U5973 : AOI222_X1 port map( A1 => n11196, A2 => n9291, B1 => n11193, B2 => 
                           n9227, C1 => n11190, C2 => n13800, ZN => n3773);
   U5974 : AOI222_X1 port map( A1 => n10999, A2 => n9740, B1 => n10996, B2 => 
                           n9676, C1 => n10993, C2 => n9708, ZN => n5156);
   U5975 : AOI222_X1 port map( A1 => n10933, A2 => n9292, B1 => n10930, B2 => 
                           n9228, C1 => n10927, C2 => n13799, ZN => n5165);
   U5976 : AOI222_X1 port map( A1 => n11263, A2 => n9740, B1 => n11260, B2 => 
                           n9676, C1 => n11257, C2 => n9708, ZN => n3723);
   U5977 : AOI222_X1 port map( A1 => n11197, A2 => n9292, B1 => n11194, B2 => 
                           n9228, C1 => n11191, C2 => n13799, ZN => n3732);
   U5978 : AOI222_X1 port map( A1 => n10999, A2 => n9741, B1 => n10996, B2 => 
                           n9677, C1 => n10993, C2 => n9709, ZN => n5115);
   U5979 : AOI222_X1 port map( A1 => n10933, A2 => n9293, B1 => n10930, B2 => 
                           n9229, C1 => n10927, C2 => n13798, ZN => n5124);
   U5980 : AOI222_X1 port map( A1 => n11263, A2 => n9741, B1 => n11260, B2 => 
                           n9677, C1 => n11257, C2 => n9709, ZN => n3682);
   U5981 : AOI222_X1 port map( A1 => n11197, A2 => n9293, B1 => n11194, B2 => 
                           n9229, C1 => n11191, C2 => n13798, ZN => n3691);
   U5982 : AOI222_X1 port map( A1 => n10999, A2 => n9742, B1 => n10996, B2 => 
                           n9678, C1 => n10993, C2 => n9710, ZN => n5074);
   U5983 : AOI222_X1 port map( A1 => n10933, A2 => n9294, B1 => n10930, B2 => 
                           n9230, C1 => n10927, C2 => n13797, ZN => n5083);
   U5984 : AOI222_X1 port map( A1 => n11263, A2 => n9742, B1 => n11260, B2 => 
                           n9678, C1 => n11257, C2 => n9710, ZN => n3641);
   U5985 : AOI222_X1 port map( A1 => n11197, A2 => n9294, B1 => n11194, B2 => 
                           n9230, C1 => n11191, C2 => n13797, ZN => n3650);
   U5986 : AOI222_X1 port map( A1 => n10999, A2 => n9743, B1 => n10996, B2 => 
                           n9679, C1 => n10993, C2 => n9711, ZN => n5033);
   U5987 : AOI222_X1 port map( A1 => n10933, A2 => n9295, B1 => n10930, B2 => 
                           n9231, C1 => n10927, C2 => n13796, ZN => n5042);
   U5988 : AOI222_X1 port map( A1 => n11263, A2 => n9743, B1 => n11260, B2 => 
                           n9679, C1 => n11257, C2 => n9711, ZN => n3600);
   U5989 : AOI222_X1 port map( A1 => n11197, A2 => n9295, B1 => n11194, B2 => 
                           n9231, C1 => n11191, C2 => n13796, ZN => n3609);
   U5990 : AOI222_X1 port map( A1 => n10999, A2 => n9744, B1 => n10996, B2 => 
                           n9680, C1 => n10993, C2 => n9712, ZN => n4992);
   U5991 : AOI222_X1 port map( A1 => n10933, A2 => n9296, B1 => n10930, B2 => 
                           n9232, C1 => n10927, C2 => n13795, ZN => n5001);
   U5992 : AOI222_X1 port map( A1 => n11263, A2 => n9744, B1 => n11260, B2 => 
                           n9680, C1 => n11257, C2 => n9712, ZN => n3559);
   U5993 : AOI222_X1 port map( A1 => n11197, A2 => n9296, B1 => n11194, B2 => 
                           n9232, C1 => n11191, C2 => n13795, ZN => n3568);
   U5994 : AOI222_X1 port map( A1 => n10999, A2 => n9745, B1 => n10996, B2 => 
                           n9681, C1 => n10993, C2 => n9713, ZN => n4951);
   U5995 : AOI222_X1 port map( A1 => n10933, A2 => n9297, B1 => n10930, B2 => 
                           n9233, C1 => n10927, C2 => n9265, ZN => n4960);
   U5996 : AOI222_X1 port map( A1 => n11263, A2 => n9745, B1 => n11260, B2 => 
                           n9681, C1 => n11257, C2 => n9713, ZN => n3518);
   U5997 : AOI222_X1 port map( A1 => n11197, A2 => n9297, B1 => n11194, B2 => 
                           n9233, C1 => n11191, C2 => n9265, ZN => n3527);
   U5998 : AOI222_X1 port map( A1 => n10999, A2 => n9746, B1 => n10996, B2 => 
                           n9682, C1 => n10993, C2 => n9714, ZN => n4910);
   U5999 : AOI222_X1 port map( A1 => n10933, A2 => n9298, B1 => n10930, B2 => 
                           n9234, C1 => n10927, C2 => n9266, ZN => n4919);
   U6000 : AOI222_X1 port map( A1 => n11263, A2 => n9746, B1 => n11260, B2 => 
                           n9682, C1 => n11257, C2 => n9714, ZN => n3477);
   U6001 : AOI222_X1 port map( A1 => n11197, A2 => n9298, B1 => n11194, B2 => 
                           n9234, C1 => n11191, C2 => n9266, ZN => n3486);
   U6002 : AOI222_X1 port map( A1 => n10999, A2 => n9747, B1 => n10996, B2 => 
                           n9683, C1 => n10993, C2 => n9715, ZN => n4869);
   U6003 : AOI222_X1 port map( A1 => n10933, A2 => n9299, B1 => n10930, B2 => 
                           n9235, C1 => n10927, C2 => n9267, ZN => n4878);
   U6004 : AOI222_X1 port map( A1 => n11263, A2 => n9747, B1 => n11260, B2 => 
                           n9683, C1 => n11257, C2 => n9715, ZN => n3436);
   U6005 : AOI222_X1 port map( A1 => n11197, A2 => n9299, B1 => n11194, B2 => 
                           n9235, C1 => n11191, C2 => n9267, ZN => n3445);
   U6006 : AOI222_X1 port map( A1 => n10999, A2 => n9748, B1 => n10996, B2 => 
                           n9684, C1 => n10993, C2 => n9716, ZN => n4828);
   U6007 : AOI222_X1 port map( A1 => n10933, A2 => n9300, B1 => n10930, B2 => 
                           n9236, C1 => n10927, C2 => n9268, ZN => n4837);
   U6008 : AOI222_X1 port map( A1 => n11263, A2 => n9748, B1 => n11260, B2 => 
                           n9684, C1 => n11257, C2 => n9716, ZN => n3395);
   U6009 : AOI222_X1 port map( A1 => n11197, A2 => n9300, B1 => n11194, B2 => 
                           n9236, C1 => n11191, C2 => n9268, ZN => n3404);
   U6010 : AOI222_X1 port map( A1 => n10999, A2 => n9749, B1 => n10996, B2 => 
                           n9685, C1 => n10993, C2 => n9717, ZN => n4787);
   U6011 : AOI222_X1 port map( A1 => n10933, A2 => n9301, B1 => n10930, B2 => 
                           n9237, C1 => n10927, C2 => n9269, ZN => n4796);
   U6012 : AOI222_X1 port map( A1 => n11263, A2 => n9749, B1 => n11260, B2 => 
                           n9685, C1 => n11257, C2 => n9717, ZN => n3354);
   U6013 : AOI222_X1 port map( A1 => n11197, A2 => n9301, B1 => n11194, B2 => 
                           n9237, C1 => n11191, C2 => n9269, ZN => n3363);
   U6014 : AOI222_X1 port map( A1 => n10999, A2 => n9750, B1 => n10996, B2 => 
                           n9686, C1 => n10993, C2 => n9718, ZN => n4746);
   U6015 : AOI222_X1 port map( A1 => n10933, A2 => n9302, B1 => n10930, B2 => 
                           n9238, C1 => n10927, C2 => n9270, ZN => n4755);
   U6016 : AOI222_X1 port map( A1 => n11263, A2 => n9750, B1 => n11260, B2 => 
                           n9686, C1 => n11257, C2 => n9718, ZN => n3313);
   U6017 : AOI222_X1 port map( A1 => n11197, A2 => n9302, B1 => n11194, B2 => 
                           n9238, C1 => n11191, C2 => n9270, ZN => n3322);
   U6018 : AOI222_X1 port map( A1 => n10999, A2 => n9751, B1 => n10996, B2 => 
                           n9687, C1 => n10993, C2 => n9719, ZN => n4705);
   U6019 : AOI222_X1 port map( A1 => n10933, A2 => n9303, B1 => n10930, B2 => 
                           n9239, C1 => n10927, C2 => n9271, ZN => n4714);
   U6020 : AOI222_X1 port map( A1 => n11263, A2 => n9751, B1 => n11260, B2 => 
                           n9687, C1 => n11257, C2 => n9719, ZN => n3272);
   U6021 : AOI222_X1 port map( A1 => n11197, A2 => n9303, B1 => n11194, B2 => 
                           n9239, C1 => n11191, C2 => n9271, ZN => n3281);
   U6022 : AOI222_X1 port map( A1 => n11000, A2 => n9752, B1 => n10997, B2 => 
                           n9688, C1 => n10994, C2 => n9720, ZN => n4664);
   U6023 : AOI222_X1 port map( A1 => n10934, A2 => n9304, B1 => n10931, B2 => 
                           n9240, C1 => n10928, C2 => n9272, ZN => n4673);
   U6024 : AOI222_X1 port map( A1 => n11264, A2 => n9752, B1 => n11261, B2 => 
                           n9688, C1 => n11258, C2 => n9720, ZN => n3231);
   U6025 : AOI222_X1 port map( A1 => n11198, A2 => n9304, B1 => n11195, B2 => 
                           n9240, C1 => n11192, C2 => n9272, ZN => n3240);
   U6026 : AOI222_X1 port map( A1 => n11000, A2 => n9753, B1 => n10997, B2 => 
                           n9689, C1 => n10994, C2 => n9721, ZN => n4623);
   U6027 : AOI222_X1 port map( A1 => n10934, A2 => n9305, B1 => n10931, B2 => 
                           n9241, C1 => n10928, C2 => n9273, ZN => n4632);
   U6028 : AOI222_X1 port map( A1 => n11264, A2 => n9753, B1 => n11261, B2 => 
                           n9689, C1 => n11258, C2 => n9721, ZN => n3190);
   U6029 : AOI222_X1 port map( A1 => n11198, A2 => n9305, B1 => n11195, B2 => 
                           n9241, C1 => n11192, C2 => n9273, ZN => n3199);
   U6030 : AOI222_X1 port map( A1 => n11000, A2 => n9754, B1 => n10997, B2 => 
                           n9690, C1 => n10994, C2 => n9722, ZN => n4582);
   U6031 : AOI222_X1 port map( A1 => n10934, A2 => n9306, B1 => n10931, B2 => 
                           n9242, C1 => n10928, C2 => n9274, ZN => n4591);
   U6032 : AOI222_X1 port map( A1 => n11264, A2 => n9754, B1 => n11261, B2 => 
                           n9690, C1 => n11258, C2 => n9722, ZN => n3149);
   U6033 : AOI222_X1 port map( A1 => n11198, A2 => n9306, B1 => n11195, B2 => 
                           n9242, C1 => n11192, C2 => n9274, ZN => n3158);
   U6034 : AOI222_X1 port map( A1 => n11000, A2 => n9755, B1 => n10997, B2 => 
                           n9691, C1 => n10994, C2 => n9723, ZN => n4541);
   U6035 : AOI222_X1 port map( A1 => n10934, A2 => n9307, B1 => n10931, B2 => 
                           n9243, C1 => n10928, C2 => n9275, ZN => n4550);
   U6036 : AOI222_X1 port map( A1 => n11264, A2 => n9755, B1 => n11261, B2 => 
                           n9691, C1 => n11258, C2 => n9723, ZN => n3108);
   U6037 : AOI222_X1 port map( A1 => n11198, A2 => n9307, B1 => n11195, B2 => 
                           n9243, C1 => n11192, C2 => n9275, ZN => n3117);
   U6038 : AOI222_X1 port map( A1 => n11000, A2 => n9756, B1 => n10997, B2 => 
                           n9692, C1 => n10994, C2 => n9724, ZN => n4500);
   U6039 : AOI222_X1 port map( A1 => n10934, A2 => n9308, B1 => n10931, B2 => 
                           n9244, C1 => n10928, C2 => n9276, ZN => n4509);
   U6040 : AOI222_X1 port map( A1 => n11264, A2 => n9756, B1 => n11261, B2 => 
                           n9692, C1 => n11258, C2 => n9724, ZN => n3067);
   U6041 : AOI222_X1 port map( A1 => n11198, A2 => n9308, B1 => n11195, B2 => 
                           n9244, C1 => n11192, C2 => n9276, ZN => n3076);
   U6042 : AOI222_X1 port map( A1 => n11000, A2 => n9757, B1 => n10997, B2 => 
                           n9693, C1 => n10994, C2 => n9725, ZN => n4459);
   U6043 : AOI222_X1 port map( A1 => n10934, A2 => n9309, B1 => n10931, B2 => 
                           n9245, C1 => n10928, C2 => n9277, ZN => n4468);
   U6044 : AOI222_X1 port map( A1 => n11264, A2 => n9757, B1 => n11261, B2 => 
                           n9693, C1 => n11258, C2 => n9725, ZN => n3026);
   U6045 : AOI222_X1 port map( A1 => n11198, A2 => n9309, B1 => n11195, B2 => 
                           n9245, C1 => n11192, C2 => n9277, ZN => n3035);
   U6046 : AOI222_X1 port map( A1 => n11000, A2 => n9758, B1 => n10997, B2 => 
                           n9694, C1 => n10994, C2 => n9726, ZN => n4418);
   U6047 : AOI222_X1 port map( A1 => n10934, A2 => n9310, B1 => n10931, B2 => 
                           n9246, C1 => n10928, C2 => n9278, ZN => n4427);
   U6048 : AOI222_X1 port map( A1 => n11264, A2 => n9758, B1 => n11261, B2 => 
                           n9694, C1 => n11258, C2 => n9726, ZN => n2985);
   U6049 : AOI222_X1 port map( A1 => n11198, A2 => n9310, B1 => n11195, B2 => 
                           n9246, C1 => n11192, C2 => n9278, ZN => n2994);
   U6050 : AOI222_X1 port map( A1 => n11000, A2 => n9759, B1 => n10997, B2 => 
                           n9695, C1 => n10994, C2 => n9727, ZN => n4311);
   U6051 : AOI222_X1 port map( A1 => n10934, A2 => n13748, B1 => n10931, B2 => 
                           n9247, C1 => n10928, C2 => n9279, ZN => n4342);
   U6052 : AOI222_X1 port map( A1 => n11264, A2 => n9759, B1 => n11261, B2 => 
                           n9695, C1 => n11258, C2 => n9727, ZN => n2811);
   U6053 : AOI222_X1 port map( A1 => n11198, A2 => n13748, B1 => n11195, B2 => 
                           n9247, C1 => n11192, C2 => n9279, ZN => n2874);
   U6054 : OAI222_X1 port map( A1 => n2338, A2 => n11106, B1 => n514, B2 => 
                           n11103, C1 => n1443, C2 => n11100, ZN => n5644);
   U6055 : OAI222_X1 port map( A1 => n10526, A2 => n11040, B1 => n10525, B2 => 
                           n11037, C1 => n10527, C2 => n11034, ZN => n5672);
   U6056 : OAI222_X1 port map( A1 => n10518, A2 => n10974, B1 => n10517, B2 => 
                           n10971, C1 => n10519, C2 => n10968, ZN => n5685);
   U6057 : OAI222_X1 port map( A1 => n2338, A2 => n11370, B1 => n514, B2 => 
                           n11367, C1 => n1443, C2 => n11364, ZN => n4211);
   U6058 : OAI222_X1 port map( A1 => n10526, A2 => n11304, B1 => n10525, B2 => 
                           n11301, C1 => n10527, C2 => n11298, ZN => n4239);
   U6059 : OAI222_X1 port map( A1 => n10518, A2 => n11238, B1 => n10517, B2 => 
                           n11235, C1 => n10519, C2 => n11232, ZN => n4252);
   U6060 : OAI222_X1 port map( A1 => n2326, A2 => n11106, B1 => n502, B2 => 
                           n11103, C1 => n1399, C2 => n11100, ZN => n5603);
   U6061 : OAI222_X1 port map( A1 => n10494, A2 => n11040, B1 => n10493, B2 => 
                           n11037, C1 => n10495, C2 => n11034, ZN => n5612);
   U6062 : OAI222_X1 port map( A1 => n10486, A2 => n10974, B1 => n10485, B2 => 
                           n10971, C1 => n10487, C2 => n10968, ZN => n5621);
   U6063 : OAI222_X1 port map( A1 => n2326, A2 => n11370, B1 => n502, B2 => 
                           n11367, C1 => n1399, C2 => n11364, ZN => n4170);
   U6064 : OAI222_X1 port map( A1 => n10494, A2 => n11304, B1 => n10493, B2 => 
                           n11301, C1 => n10495, C2 => n11298, ZN => n4179);
   U6065 : OAI222_X1 port map( A1 => n10486, A2 => n11238, B1 => n10485, B2 => 
                           n11235, C1 => n10487, C2 => n11232, ZN => n4188);
   U6066 : OAI222_X1 port map( A1 => n2314, A2 => n11106, B1 => n490, B2 => 
                           n11103, C1 => n1387, C2 => n11100, ZN => n5562);
   U6067 : OAI222_X1 port map( A1 => n10462, A2 => n11040, B1 => n10461, B2 => 
                           n11037, C1 => n10463, C2 => n11034, ZN => n5571);
   U6068 : OAI222_X1 port map( A1 => n10454, A2 => n10974, B1 => n10453, B2 => 
                           n10971, C1 => n10455, C2 => n10968, ZN => n5580);
   U6069 : OAI222_X1 port map( A1 => n2314, A2 => n11370, B1 => n490, B2 => 
                           n11367, C1 => n1387, C2 => n11364, ZN => n4129);
   U6070 : OAI222_X1 port map( A1 => n10462, A2 => n11304, B1 => n10461, B2 => 
                           n11301, C1 => n10463, C2 => n11298, ZN => n4138);
   U6071 : OAI222_X1 port map( A1 => n10454, A2 => n11238, B1 => n10453, B2 => 
                           n11235, C1 => n10455, C2 => n11232, ZN => n4147);
   U6072 : OAI222_X1 port map( A1 => n2302, A2 => n11106, B1 => n478, B2 => 
                           n11103, C1 => n1343, C2 => n11100, ZN => n5521);
   U6073 : OAI222_X1 port map( A1 => n10430, A2 => n11040, B1 => n10429, B2 => 
                           n11037, C1 => n10431, C2 => n11034, ZN => n5530);
   U6074 : OAI222_X1 port map( A1 => n10422, A2 => n10974, B1 => n10421, B2 => 
                           n10971, C1 => n10423, C2 => n10968, ZN => n5539);
   U6075 : OAI222_X1 port map( A1 => n2302, A2 => n11370, B1 => n478, B2 => 
                           n11367, C1 => n1343, C2 => n11364, ZN => n4088);
   U6076 : OAI222_X1 port map( A1 => n10430, A2 => n11304, B1 => n10429, B2 => 
                           n11301, C1 => n10431, C2 => n11298, ZN => n4097);
   U6077 : OAI222_X1 port map( A1 => n10422, A2 => n11238, B1 => n10421, B2 => 
                           n11235, C1 => n10423, C2 => n11232, ZN => n4106);
   U6078 : OAI222_X1 port map( A1 => n2290, A2 => n11106, B1 => n466, B2 => 
                           n11103, C1 => n1331, C2 => n11100, ZN => n5480);
   U6079 : OAI222_X1 port map( A1 => n10395, A2 => n11040, B1 => n10394, B2 => 
                           n11037, C1 => n10396, C2 => n11034, ZN => n5489);
   U6080 : OAI222_X1 port map( A1 => n10387, A2 => n10974, B1 => n10386, B2 => 
                           n10971, C1 => n10388, C2 => n10968, ZN => n5498);
   U6081 : OAI222_X1 port map( A1 => n2290, A2 => n11370, B1 => n466, B2 => 
                           n11367, C1 => n1331, C2 => n11364, ZN => n4047);
   U6082 : OAI222_X1 port map( A1 => n10395, A2 => n11304, B1 => n10394, B2 => 
                           n11301, C1 => n10396, C2 => n11298, ZN => n4056);
   U6083 : OAI222_X1 port map( A1 => n10387, A2 => n11238, B1 => n10386, B2 => 
                           n11235, C1 => n10388, C2 => n11232, ZN => n4065);
   U6084 : OAI222_X1 port map( A1 => n2278, A2 => n11106, B1 => n454, B2 => 
                           n11103, C1 => n1319, C2 => n11100, ZN => n5439);
   U6085 : OAI222_X1 port map( A1 => n10363, A2 => n11040, B1 => n10362, B2 => 
                           n11037, C1 => n10364, C2 => n11034, ZN => n5448);
   U6086 : OAI222_X1 port map( A1 => n10355, A2 => n10974, B1 => n10354, B2 => 
                           n10971, C1 => n10356, C2 => n10968, ZN => n5457);
   U6087 : OAI222_X1 port map( A1 => n2278, A2 => n11370, B1 => n454, B2 => 
                           n11367, C1 => n1319, C2 => n11364, ZN => n4006);
   U6088 : OAI222_X1 port map( A1 => n10363, A2 => n11304, B1 => n10362, B2 => 
                           n11301, C1 => n10364, C2 => n11298, ZN => n4015);
   U6089 : OAI222_X1 port map( A1 => n10355, A2 => n11238, B1 => n10354, B2 => 
                           n11235, C1 => n10356, C2 => n11232, ZN => n4024);
   U6090 : OAI222_X1 port map( A1 => n2266, A2 => n11106, B1 => n442, B2 => 
                           n11103, C1 => n1307, C2 => n11100, ZN => n5398);
   U6091 : OAI222_X1 port map( A1 => n10331, A2 => n11040, B1 => n10330, B2 => 
                           n11037, C1 => n10332, C2 => n11034, ZN => n5407);
   U6092 : OAI222_X1 port map( A1 => n10323, A2 => n10974, B1 => n10322, B2 => 
                           n10971, C1 => n10324, C2 => n10968, ZN => n5416);
   U6093 : OAI222_X1 port map( A1 => n2266, A2 => n11370, B1 => n442, B2 => 
                           n11367, C1 => n1307, C2 => n11364, ZN => n3965);
   U6094 : OAI222_X1 port map( A1 => n10331, A2 => n11304, B1 => n10330, B2 => 
                           n11301, C1 => n10332, C2 => n11298, ZN => n3974);
   U6095 : OAI222_X1 port map( A1 => n10323, A2 => n11238, B1 => n10322, B2 => 
                           n11235, C1 => n10324, C2 => n11232, ZN => n3983);
   U6096 : OAI222_X1 port map( A1 => n2254, A2 => n11106, B1 => n430, B2 => 
                           n11103, C1 => n1295, C2 => n11100, ZN => n5357);
   U6097 : OAI222_X1 port map( A1 => n10296, A2 => n11040, B1 => n10295, B2 => 
                           n11037, C1 => n10297, C2 => n11034, ZN => n5366);
   U6098 : OAI222_X1 port map( A1 => n10288, A2 => n10974, B1 => n10287, B2 => 
                           n10971, C1 => n10289, C2 => n10968, ZN => n5375);
   U6099 : OAI222_X1 port map( A1 => n2254, A2 => n11370, B1 => n430, B2 => 
                           n11367, C1 => n1295, C2 => n11364, ZN => n3924);
   U6100 : OAI222_X1 port map( A1 => n10296, A2 => n11304, B1 => n10295, B2 => 
                           n11301, C1 => n10297, C2 => n11298, ZN => n3933);
   U6101 : OAI222_X1 port map( A1 => n10288, A2 => n11238, B1 => n10287, B2 => 
                           n11235, C1 => n10289, C2 => n11232, ZN => n3942);
   U6102 : OAI222_X1 port map( A1 => n2242, A2 => n11106, B1 => n418, B2 => 
                           n11103, C1 => n1283, C2 => n11100, ZN => n5316);
   U6103 : OAI222_X1 port map( A1 => n10264, A2 => n11040, B1 => n10263, B2 => 
                           n11037, C1 => n10265, C2 => n11034, ZN => n5325);
   U6104 : OAI222_X1 port map( A1 => n10256, A2 => n10974, B1 => n10255, B2 => 
                           n10971, C1 => n10257, C2 => n10968, ZN => n5334);
   U6105 : OAI222_X1 port map( A1 => n2242, A2 => n11370, B1 => n418, B2 => 
                           n11367, C1 => n1283, C2 => n11364, ZN => n3883);
   U6106 : OAI222_X1 port map( A1 => n10264, A2 => n11304, B1 => n10263, B2 => 
                           n11301, C1 => n10265, C2 => n11298, ZN => n3892);
   U6107 : OAI222_X1 port map( A1 => n10256, A2 => n11238, B1 => n10255, B2 => 
                           n11235, C1 => n10257, C2 => n11232, ZN => n3901);
   U6108 : OAI222_X1 port map( A1 => n2230, A2 => n11106, B1 => n406, B2 => 
                           n11103, C1 => n1271, C2 => n11100, ZN => n5275);
   U6109 : OAI222_X1 port map( A1 => n10232, A2 => n11040, B1 => n10231, B2 => 
                           n11037, C1 => n10233, C2 => n11034, ZN => n5284);
   U6110 : OAI222_X1 port map( A1 => n10224, A2 => n10974, B1 => n10223, B2 => 
                           n10971, C1 => n10225, C2 => n10968, ZN => n5293);
   U6111 : OAI222_X1 port map( A1 => n2230, A2 => n11370, B1 => n406, B2 => 
                           n11367, C1 => n1271, C2 => n11364, ZN => n3842);
   U6112 : OAI222_X1 port map( A1 => n10232, A2 => n11304, B1 => n10231, B2 => 
                           n11301, C1 => n10233, C2 => n11298, ZN => n3851);
   U6113 : OAI222_X1 port map( A1 => n10224, A2 => n11238, B1 => n10223, B2 => 
                           n11235, C1 => n10225, C2 => n11232, ZN => n3860);
   U6114 : OAI222_X1 port map( A1 => n2218, A2 => n11106, B1 => n394, B2 => 
                           n11103, C1 => n1259, C2 => n11100, ZN => n5234);
   U6115 : OAI222_X1 port map( A1 => n10198, A2 => n11040, B1 => n10197, B2 => 
                           n11037, C1 => n10199, C2 => n11034, ZN => n5243);
   U6116 : OAI222_X1 port map( A1 => n10190, A2 => n10974, B1 => n10189, B2 => 
                           n10971, C1 => n10191, C2 => n10968, ZN => n5252);
   U6117 : OAI222_X1 port map( A1 => n2218, A2 => n11370, B1 => n394, B2 => 
                           n11367, C1 => n1259, C2 => n11364, ZN => n3801);
   U6118 : OAI222_X1 port map( A1 => n10198, A2 => n11304, B1 => n10197, B2 => 
                           n11301, C1 => n10199, C2 => n11298, ZN => n3810);
   U6119 : OAI222_X1 port map( A1 => n10190, A2 => n11238, B1 => n10189, B2 => 
                           n11235, C1 => n10191, C2 => n11232, ZN => n3819);
   U6120 : OAI222_X1 port map( A1 => n2174, A2 => n11106, B1 => n382, B2 => 
                           n11103, C1 => n1247, C2 => n11100, ZN => n5193);
   U6121 : OAI222_X1 port map( A1 => n10166, A2 => n11040, B1 => n10165, B2 => 
                           n11037, C1 => n10167, C2 => n11034, ZN => n5202);
   U6122 : OAI222_X1 port map( A1 => n10158, A2 => n10974, B1 => n10157, B2 => 
                           n10971, C1 => n10159, C2 => n10968, ZN => n5211);
   U6123 : OAI222_X1 port map( A1 => n2174, A2 => n11370, B1 => n382, B2 => 
                           n11367, C1 => n1247, C2 => n11364, ZN => n3760);
   U6124 : OAI222_X1 port map( A1 => n10166, A2 => n11304, B1 => n10165, B2 => 
                           n11301, C1 => n10167, C2 => n11298, ZN => n3769);
   U6125 : OAI222_X1 port map( A1 => n10158, A2 => n11238, B1 => n10157, B2 => 
                           n11235, C1 => n10159, C2 => n11232, ZN => n3778);
   U6126 : OAI222_X1 port map( A1 => n2162, A2 => n11107, B1 => n370, B2 => 
                           n11104, C1 => n1235, C2 => n11101, ZN => n5152);
   U6127 : OAI222_X1 port map( A1 => n10134, A2 => n11041, B1 => n10133, B2 => 
                           n11038, C1 => n10135, C2 => n11035, ZN => n5161);
   U6128 : OAI222_X1 port map( A1 => n10126, A2 => n10975, B1 => n10125, B2 => 
                           n10972, C1 => n10127, C2 => n10969, ZN => n5170);
   U6129 : OAI222_X1 port map( A1 => n2162, A2 => n11371, B1 => n370, B2 => 
                           n11368, C1 => n1235, C2 => n11365, ZN => n3719);
   U6130 : OAI222_X1 port map( A1 => n10134, A2 => n11305, B1 => n10133, B2 => 
                           n11302, C1 => n10135, C2 => n11299, ZN => n3728);
   U6131 : OAI222_X1 port map( A1 => n10126, A2 => n11239, B1 => n10125, B2 => 
                           n11236, C1 => n10127, C2 => n11233, ZN => n3737);
   U6132 : OAI222_X1 port map( A1 => n2150, A2 => n11107, B1 => n358, B2 => 
                           n11104, C1 => n1223, C2 => n11101, ZN => n5111);
   U6133 : OAI222_X1 port map( A1 => n10102, A2 => n11041, B1 => n10101, B2 => 
                           n11038, C1 => n10103, C2 => n11035, ZN => n5120);
   U6134 : OAI222_X1 port map( A1 => n10094, A2 => n10975, B1 => n10093, B2 => 
                           n10972, C1 => n10095, C2 => n10969, ZN => n5129);
   U6135 : OAI222_X1 port map( A1 => n2150, A2 => n11371, B1 => n358, B2 => 
                           n11368, C1 => n1223, C2 => n11365, ZN => n3678);
   U6136 : OAI222_X1 port map( A1 => n10102, A2 => n11305, B1 => n10101, B2 => 
                           n11302, C1 => n10103, C2 => n11299, ZN => n3687);
   U6137 : OAI222_X1 port map( A1 => n10094, A2 => n11239, B1 => n10093, B2 => 
                           n11236, C1 => n10095, C2 => n11233, ZN => n3696);
   U6138 : OAI222_X1 port map( A1 => n2106, A2 => n11107, B1 => n346, B2 => 
                           n11104, C1 => n1211, C2 => n11101, ZN => n5070);
   U6139 : OAI222_X1 port map( A1 => n10070, A2 => n11041, B1 => n10069, B2 => 
                           n11038, C1 => n10071, C2 => n11035, ZN => n5079);
   U6140 : OAI222_X1 port map( A1 => n10062, A2 => n10975, B1 => n10061, B2 => 
                           n10972, C1 => n10063, C2 => n10969, ZN => n5088);
   U6141 : OAI222_X1 port map( A1 => n2106, A2 => n11371, B1 => n346, B2 => 
                           n11368, C1 => n1211, C2 => n11365, ZN => n3637);
   U6142 : OAI222_X1 port map( A1 => n10070, A2 => n11305, B1 => n10069, B2 => 
                           n11302, C1 => n10071, C2 => n11299, ZN => n3646);
   U6143 : OAI222_X1 port map( A1 => n10062, A2 => n11239, B1 => n10061, B2 => 
                           n11236, C1 => n10063, C2 => n11233, ZN => n3655);
   U6144 : OAI222_X1 port map( A1 => n2094, A2 => n11107, B1 => n334, B2 => 
                           n11104, C1 => n1199, C2 => n11101, ZN => n5029);
   U6145 : OAI222_X1 port map( A1 => n10038, A2 => n11041, B1 => n10037, B2 => 
                           n11038, C1 => n10039, C2 => n11035, ZN => n5038);
   U6146 : OAI222_X1 port map( A1 => n10030, A2 => n10975, B1 => n10029, B2 => 
                           n10972, C1 => n10031, C2 => n10969, ZN => n5047);
   U6147 : OAI222_X1 port map( A1 => n2094, A2 => n11371, B1 => n334, B2 => 
                           n11368, C1 => n1199, C2 => n11365, ZN => n3596);
   U6148 : OAI222_X1 port map( A1 => n10038, A2 => n11305, B1 => n10037, B2 => 
                           n11302, C1 => n10039, C2 => n11299, ZN => n3605);
   U6149 : OAI222_X1 port map( A1 => n10030, A2 => n11239, B1 => n10029, B2 => 
                           n11236, C1 => n10031, C2 => n11233, ZN => n3614);
   U6150 : OAI222_X1 port map( A1 => n2082, A2 => n11107, B1 => n322, B2 => 
                           n11104, C1 => n1187, C2 => n11101, ZN => n4988);
   U6151 : OAI222_X1 port map( A1 => n10006, A2 => n11041, B1 => n10005, B2 => 
                           n11038, C1 => n10007, C2 => n11035, ZN => n4997);
   U6152 : OAI222_X1 port map( A1 => n9700, A2 => n10975, B1 => n9699, B2 => 
                           n10972, C1 => n9701, C2 => n10969, ZN => n5006);
   U6153 : OAI222_X1 port map( A1 => n2082, A2 => n11371, B1 => n322, B2 => 
                           n11368, C1 => n1187, C2 => n11365, ZN => n3555);
   U6154 : OAI222_X1 port map( A1 => n10006, A2 => n11305, B1 => n10005, B2 => 
                           n11302, C1 => n10007, C2 => n11299, ZN => n3564);
   U6155 : OAI222_X1 port map( A1 => n9700, A2 => n11239, B1 => n9699, B2 => 
                           n11236, C1 => n9701, C2 => n11233, ZN => n3573);
   U6156 : OAI222_X1 port map( A1 => n2038, A2 => n11107, B1 => n310, B2 => 
                           n11104, C1 => n1175, C2 => n11101, ZN => n4947);
   U6157 : OAI222_X1 port map( A1 => n9644, A2 => n11041, B1 => n9643, B2 => 
                           n11038, C1 => n9645, C2 => n11035, ZN => n4956);
   U6158 : OAI222_X1 port map( A1 => n9636, A2 => n10975, B1 => n9635, B2 => 
                           n10972, C1 => n9637, C2 => n10969, ZN => n4965);
   U6159 : OAI222_X1 port map( A1 => n2038, A2 => n11371, B1 => n310, B2 => 
                           n11368, C1 => n1175, C2 => n11365, ZN => n3514);
   U6160 : OAI222_X1 port map( A1 => n9644, A2 => n11305, B1 => n9643, B2 => 
                           n11302, C1 => n9645, C2 => n11299, ZN => n3523);
   U6161 : OAI222_X1 port map( A1 => n9636, A2 => n11239, B1 => n9635, B2 => 
                           n11236, C1 => n9637, C2 => n11233, ZN => n3532);
   U6162 : OAI222_X1 port map( A1 => n2026, A2 => n11107, B1 => n298, B2 => 
                           n11104, C1 => n1163, C2 => n11101, ZN => n4906);
   U6163 : OAI222_X1 port map( A1 => n9612, A2 => n11041, B1 => n9611, B2 => 
                           n11038, C1 => n9613, C2 => n11035, ZN => n4915);
   U6164 : OAI222_X1 port map( A1 => n9604, A2 => n10975, B1 => n9603, B2 => 
                           n10972, C1 => n9605, C2 => n10969, ZN => n4924);
   U6165 : OAI222_X1 port map( A1 => n2026, A2 => n11371, B1 => n298, B2 => 
                           n11368, C1 => n1163, C2 => n11365, ZN => n3473);
   U6166 : OAI222_X1 port map( A1 => n9612, A2 => n11305, B1 => n9611, B2 => 
                           n11302, C1 => n9613, C2 => n11299, ZN => n3482);
   U6167 : OAI222_X1 port map( A1 => n9604, A2 => n11239, B1 => n9603, B2 => 
                           n11236, C1 => n9605, C2 => n11233, ZN => n3491);
   U6168 : OAI222_X1 port map( A1 => n2014, A2 => n11107, B1 => n286, B2 => 
                           n11104, C1 => n1151, C2 => n11101, ZN => n4865);
   U6169 : OAI222_X1 port map( A1 => n9580, A2 => n11041, B1 => n9579, B2 => 
                           n11038, C1 => n9581, C2 => n11035, ZN => n4874);
   U6170 : OAI222_X1 port map( A1 => n9572, A2 => n10975, B1 => n9571, B2 => 
                           n10972, C1 => n9573, C2 => n10969, ZN => n4883);
   U6171 : OAI222_X1 port map( A1 => n2014, A2 => n11371, B1 => n286, B2 => 
                           n11368, C1 => n1151, C2 => n11365, ZN => n3432);
   U6172 : OAI222_X1 port map( A1 => n9580, A2 => n11305, B1 => n9579, B2 => 
                           n11302, C1 => n9581, C2 => n11299, ZN => n3441);
   U6173 : OAI222_X1 port map( A1 => n9572, A2 => n11239, B1 => n9571, B2 => 
                           n11236, C1 => n9573, C2 => n11233, ZN => n3450);
   U6174 : OAI222_X1 port map( A1 => n2002, A2 => n11107, B1 => n274, B2 => 
                           n11104, C1 => n1139, C2 => n11101, ZN => n4824);
   U6175 : OAI222_X1 port map( A1 => n9214, A2 => n11041, B1 => n9213, B2 => 
                           n11038, C1 => n9215, C2 => n11035, ZN => n4833);
   U6176 : OAI222_X1 port map( A1 => n9206, A2 => n10975, B1 => n9205, B2 => 
                           n10972, C1 => n9207, C2 => n10969, ZN => n4842);
   U6177 : OAI222_X1 port map( A1 => n2002, A2 => n11371, B1 => n274, B2 => 
                           n11368, C1 => n1139, C2 => n11365, ZN => n3391);
   U6178 : OAI222_X1 port map( A1 => n9214, A2 => n11305, B1 => n9213, B2 => 
                           n11302, C1 => n9215, C2 => n11299, ZN => n3400);
   U6179 : OAI222_X1 port map( A1 => n9206, A2 => n11239, B1 => n9205, B2 => 
                           n11236, C1 => n9207, C2 => n11233, ZN => n3409);
   U6180 : OAI222_X1 port map( A1 => n1990, A2 => n11107, B1 => n262, B2 => 
                           n11104, C1 => n1127, C2 => n11101, ZN => n4783);
   U6181 : OAI222_X1 port map( A1 => n9182, A2 => n11041, B1 => n9181, B2 => 
                           n11038, C1 => n9183, C2 => n11035, ZN => n4792);
   U6182 : OAI222_X1 port map( A1 => n9174, A2 => n10975, B1 => n9173, B2 => 
                           n10972, C1 => n9175, C2 => n10969, ZN => n4801);
   U6183 : OAI222_X1 port map( A1 => n1990, A2 => n11371, B1 => n262, B2 => 
                           n11368, C1 => n1127, C2 => n11365, ZN => n3350);
   U6184 : OAI222_X1 port map( A1 => n9182, A2 => n11305, B1 => n9181, B2 => 
                           n11302, C1 => n9183, C2 => n11299, ZN => n3359);
   U6185 : OAI222_X1 port map( A1 => n9174, A2 => n11239, B1 => n9173, B2 => 
                           n11236, C1 => n9175, C2 => n11233, ZN => n3368);
   U6186 : OAI222_X1 port map( A1 => n1978, A2 => n11107, B1 => n250, B2 => 
                           n11104, C1 => n1115, C2 => n11101, ZN => n4742);
   U6187 : OAI222_X1 port map( A1 => n9150, A2 => n11041, B1 => n9149, B2 => 
                           n11038, C1 => n9151, C2 => n11035, ZN => n4751);
   U6188 : OAI222_X1 port map( A1 => n9142, A2 => n10975, B1 => n9141, B2 => 
                           n10972, C1 => n9143, C2 => n10969, ZN => n4760);
   U6189 : OAI222_X1 port map( A1 => n1978, A2 => n11371, B1 => n250, B2 => 
                           n11368, C1 => n1115, C2 => n11365, ZN => n3309);
   U6190 : OAI222_X1 port map( A1 => n9150, A2 => n11305, B1 => n9149, B2 => 
                           n11302, C1 => n9151, C2 => n11299, ZN => n3318);
   U6191 : OAI222_X1 port map( A1 => n9142, A2 => n11239, B1 => n9141, B2 => 
                           n11236, C1 => n9143, C2 => n11233, ZN => n3327);
   U6192 : OAI222_X1 port map( A1 => n1966, A2 => n11107, B1 => n238, B2 => 
                           n11104, C1 => n1103, C2 => n11101, ZN => n4701);
   U6193 : OAI222_X1 port map( A1 => n6236, A2 => n11041, B1 => n6140, B2 => 
                           n11038, C1 => n6301, C2 => n11035, ZN => n4710);
   U6194 : OAI222_X1 port map( A1 => n6007, A2 => n10975, B1 => n6006, B2 => 
                           n10972, C1 => n6008, C2 => n10969, ZN => n4719);
   U6195 : OAI222_X1 port map( A1 => n1966, A2 => n11371, B1 => n238, B2 => 
                           n11368, C1 => n1103, C2 => n11365, ZN => n3268);
   U6196 : OAI222_X1 port map( A1 => n6236, A2 => n11305, B1 => n6140, B2 => 
                           n11302, C1 => n6301, C2 => n11299, ZN => n3277);
   U6197 : OAI222_X1 port map( A1 => n6007, A2 => n11239, B1 => n6006, B2 => 
                           n11236, C1 => n6008, C2 => n11233, ZN => n3286);
   U6198 : OAI222_X1 port map( A1 => n1954, A2 => n11108, B1 => n226, B2 => 
                           n11105, C1 => n1091, C2 => n11102, ZN => n4660);
   U6199 : OAI222_X1 port map( A1 => n5983, A2 => n11042, B1 => n5982, B2 => 
                           n11039, C1 => n5984, C2 => n11036, ZN => n4669);
   U6200 : OAI222_X1 port map( A1 => n5943, A2 => n10976, B1 => n5942, B2 => 
                           n10973, C1 => n5944, C2 => n10970, ZN => n4678);
   U6201 : OAI222_X1 port map( A1 => n1954, A2 => n11372, B1 => n226, B2 => 
                           n11369, C1 => n1091, C2 => n11366, ZN => n3227);
   U6202 : OAI222_X1 port map( A1 => n5983, A2 => n11306, B1 => n5982, B2 => 
                           n11303, C1 => n5984, C2 => n11300, ZN => n3236);
   U6203 : OAI222_X1 port map( A1 => n5943, A2 => n11240, B1 => n5942, B2 => 
                           n11237, C1 => n5944, C2 => n11234, ZN => n3245);
   U6204 : OAI222_X1 port map( A1 => n1942, A2 => n11108, B1 => n214, B2 => 
                           n11105, C1 => n1079, C2 => n11102, ZN => n4619);
   U6205 : OAI222_X1 port map( A1 => n5919, A2 => n11042, B1 => n5918, B2 => 
                           n11039, C1 => n5920, C2 => n11036, ZN => n4628);
   U6206 : OAI222_X1 port map( A1 => n5911, A2 => n10976, B1 => n5910, B2 => 
                           n10973, C1 => n5912, C2 => n10970, ZN => n4637);
   U6207 : OAI222_X1 port map( A1 => n1942, A2 => n11372, B1 => n214, B2 => 
                           n11369, C1 => n1079, C2 => n11366, ZN => n3186);
   U6208 : OAI222_X1 port map( A1 => n5919, A2 => n11306, B1 => n5918, B2 => 
                           n11303, C1 => n5920, C2 => n11300, ZN => n3195);
   U6209 : OAI222_X1 port map( A1 => n5911, A2 => n11240, B1 => n5910, B2 => 
                           n11237, C1 => n5912, C2 => n11234, ZN => n3204);
   U6210 : OAI222_X1 port map( A1 => n1930, A2 => n11108, B1 => n202, B2 => 
                           n11105, C1 => n1067, C2 => n11102, ZN => n4578);
   U6211 : OAI222_X1 port map( A1 => n5887, A2 => n11042, B1 => n5886, B2 => 
                           n11039, C1 => n5888, C2 => n11036, ZN => n4587);
   U6212 : OAI222_X1 port map( A1 => n5879, A2 => n10976, B1 => n5878, B2 => 
                           n10973, C1 => n5880, C2 => n10970, ZN => n4596);
   U6213 : OAI222_X1 port map( A1 => n1930, A2 => n11372, B1 => n202, B2 => 
                           n11369, C1 => n1067, C2 => n11366, ZN => n3145);
   U6214 : OAI222_X1 port map( A1 => n5887, A2 => n11306, B1 => n5886, B2 => 
                           n11303, C1 => n5888, C2 => n11300, ZN => n3154);
   U6215 : OAI222_X1 port map( A1 => n5879, A2 => n11240, B1 => n5878, B2 => 
                           n11237, C1 => n5880, C2 => n11234, ZN => n3163);
   U6216 : OAI222_X1 port map( A1 => n1918, A2 => n11108, B1 => n190, B2 => 
                           n11105, C1 => n1055, C2 => n11102, ZN => n4537);
   U6217 : OAI222_X1 port map( A1 => n5855, A2 => n11042, B1 => n5854, B2 => 
                           n11039, C1 => n5856, C2 => n11036, ZN => n4546);
   U6218 : OAI222_X1 port map( A1 => n5847, A2 => n10976, B1 => n5846, B2 => 
                           n10973, C1 => n5848, C2 => n10970, ZN => n4555);
   U6219 : OAI222_X1 port map( A1 => n1918, A2 => n11372, B1 => n190, B2 => 
                           n11369, C1 => n1055, C2 => n11366, ZN => n3104);
   U6220 : OAI222_X1 port map( A1 => n5855, A2 => n11306, B1 => n5854, B2 => 
                           n11303, C1 => n5856, C2 => n11300, ZN => n3113);
   U6221 : OAI222_X1 port map( A1 => n5847, A2 => n11240, B1 => n5846, B2 => 
                           n11237, C1 => n5848, C2 => n11234, ZN => n3122);
   U6222 : OAI222_X1 port map( A1 => n1906, A2 => n11108, B1 => n178, B2 => 
                           n11105, C1 => n1043, C2 => n11102, ZN => n4496);
   U6223 : OAI222_X1 port map( A1 => n5823, A2 => n11042, B1 => n5822, B2 => 
                           n11039, C1 => n5824, C2 => n11036, ZN => n4505);
   U6224 : OAI222_X1 port map( A1 => n5815, A2 => n10976, B1 => n5814, B2 => 
                           n10973, C1 => n5816, C2 => n10970, ZN => n4514);
   U6225 : OAI222_X1 port map( A1 => n1906, A2 => n11372, B1 => n178, B2 => 
                           n11369, C1 => n1043, C2 => n11366, ZN => n3063);
   U6226 : OAI222_X1 port map( A1 => n5823, A2 => n11306, B1 => n5822, B2 => 
                           n11303, C1 => n5824, C2 => n11300, ZN => n3072);
   U6227 : OAI222_X1 port map( A1 => n5815, A2 => n11240, B1 => n5814, B2 => 
                           n11237, C1 => n5816, C2 => n11234, ZN => n3081);
   U6228 : OAI222_X1 port map( A1 => n5791, A2 => n11042, B1 => n5790, B2 => 
                           n11039, C1 => n5792, C2 => n11036, ZN => n4464);
   U6229 : OAI222_X1 port map( A1 => n5783, A2 => n10976, B1 => n5782, B2 => 
                           n10973, C1 => n5784, C2 => n10970, ZN => n4473);
   U6230 : OAI222_X1 port map( A1 => n5791, A2 => n11306, B1 => n5790, B2 => 
                           n11303, C1 => n5792, C2 => n11300, ZN => n3031);
   U6231 : OAI222_X1 port map( A1 => n5783, A2 => n11240, B1 => n5782, B2 => 
                           n11237, C1 => n5784, C2 => n11234, ZN => n3040);
   U6232 : OAI222_X1 port map( A1 => n5759, A2 => n11042, B1 => n5758, B2 => 
                           n11039, C1 => n5760, C2 => n11036, ZN => n4423);
   U6233 : OAI222_X1 port map( A1 => n5751, A2 => n10976, B1 => n5750, B2 => 
                           n10973, C1 => n5752, C2 => n10970, ZN => n4432);
   U6234 : OAI222_X1 port map( A1 => n5759, A2 => n11306, B1 => n5758, B2 => 
                           n11303, C1 => n5760, C2 => n11300, ZN => n2990);
   U6235 : OAI222_X1 port map( A1 => n5751, A2 => n11240, B1 => n5750, B2 => 
                           n11237, C1 => n5752, C2 => n11234, ZN => n2999);
   U6236 : OAI222_X1 port map( A1 => n5727, A2 => n11042, B1 => n5726, B2 => 
                           n11039, C1 => n5728, C2 => n11036, ZN => n4316);
   U6237 : OAI222_X1 port map( A1 => n5719, A2 => n10976, B1 => n5718, B2 => 
                           n10973, C1 => n5720, C2 => n10970, ZN => n4347);
   U6238 : OAI222_X1 port map( A1 => n14035, A2 => n10910, B1 => n14067, B2 => 
                           n10907, C1 => n998, C2 => n10904, ZN => n4378);
   U6239 : OAI222_X1 port map( A1 => n5727, A2 => n11306, B1 => n5726, B2 => 
                           n11303, C1 => n5728, C2 => n11300, ZN => n2816);
   U6240 : OAI222_X1 port map( A1 => n5719, A2 => n11240, B1 => n5718, B2 => 
                           n11237, C1 => n5720, C2 => n11234, ZN => n2879);
   U6241 : OAI222_X1 port map( A1 => n14035, A2 => n11174, B1 => n14067, B2 => 
                           n11171, C1 => n998, C2 => n11168, ZN => n2945);
   U6242 : OAI222_X1 port map( A1 => n1894, A2 => n11108, B1 => n166, B2 => 
                           n11105, C1 => n12782, C2 => n11102, ZN => n4455);
   U6243 : OAI222_X1 port map( A1 => n1894, A2 => n11372, B1 => n166, B2 => 
                           n11369, C1 => n12782, C2 => n11366, ZN => n3022);
   U6244 : OAI222_X1 port map( A1 => n1882, A2 => n11108, B1 => n154, B2 => 
                           n11105, C1 => n12781, C2 => n11102, ZN => n4414);
   U6245 : OAI222_X1 port map( A1 => n1882, A2 => n11372, B1 => n154, B2 => 
                           n11369, C1 => n12781, C2 => n11366, ZN => n2981);
   U6246 : OAI222_X1 port map( A1 => n1870, A2 => n11108, B1 => n142, B2 => 
                           n11105, C1 => n12780, C2 => n11102, ZN => n4285);
   U6247 : OAI222_X1 port map( A1 => n1870, A2 => n11372, B1 => n142, B2 => 
                           n11369, C1 => n12780, C2 => n11366, ZN => n2753);
   U6248 : OAI222_X1 port map( A1 => n10534, A2 => n11073, B1 => n10533, B2 => 
                           n11070, C1 => n10535, C2 => n11067, ZN => n5658);
   U6249 : OAI222_X1 port map( A1 => n10534, A2 => n11337, B1 => n10533, B2 => 
                           n11334, C1 => n10535, C2 => n11331, ZN => n4225);
   U6250 : OAI222_X1 port map( A1 => n10502, A2 => n11073, B1 => n10501, B2 => 
                           n11070, C1 => n10503, C2 => n11067, ZN => n5605);
   U6251 : OAI222_X1 port map( A1 => n10502, A2 => n11337, B1 => n10501, B2 => 
                           n11334, C1 => n10503, C2 => n11331, ZN => n4172);
   U6252 : OAI222_X1 port map( A1 => n10470, A2 => n11073, B1 => n10469, B2 => 
                           n11070, C1 => n10471, C2 => n11067, ZN => n5564);
   U6253 : OAI222_X1 port map( A1 => n10470, A2 => n11337, B1 => n10469, B2 => 
                           n11334, C1 => n10471, C2 => n11331, ZN => n4131);
   U6254 : OAI222_X1 port map( A1 => n10438, A2 => n11073, B1 => n10437, B2 => 
                           n11070, C1 => n10439, C2 => n11067, ZN => n5523);
   U6255 : OAI222_X1 port map( A1 => n10438, A2 => n11337, B1 => n10437, B2 => 
                           n11334, C1 => n10439, C2 => n11331, ZN => n4090);
   U6256 : OAI222_X1 port map( A1 => n10406, A2 => n11073, B1 => n10405, B2 => 
                           n11070, C1 => n10407, C2 => n11067, ZN => n5482);
   U6257 : OAI222_X1 port map( A1 => n10406, A2 => n11337, B1 => n10405, B2 => 
                           n11334, C1 => n10407, C2 => n11331, ZN => n4049);
   U6258 : OAI222_X1 port map( A1 => n10371, A2 => n11073, B1 => n10370, B2 => 
                           n11070, C1 => n10372, C2 => n11067, ZN => n5441);
   U6259 : OAI222_X1 port map( A1 => n10371, A2 => n11337, B1 => n10370, B2 => 
                           n11334, C1 => n10372, C2 => n11331, ZN => n4008);
   U6260 : OAI222_X1 port map( A1 => n10339, A2 => n11073, B1 => n10338, B2 => 
                           n11070, C1 => n10340, C2 => n11067, ZN => n5400);
   U6261 : OAI222_X1 port map( A1 => n10339, A2 => n11337, B1 => n10338, B2 => 
                           n11334, C1 => n10340, C2 => n11331, ZN => n3967);
   U6262 : OAI222_X1 port map( A1 => n10307, A2 => n11073, B1 => n10306, B2 => 
                           n11070, C1 => n10308, C2 => n11067, ZN => n5359);
   U6263 : OAI222_X1 port map( A1 => n10307, A2 => n11337, B1 => n10306, B2 => 
                           n11334, C1 => n10308, C2 => n11331, ZN => n3926);
   U6264 : OAI222_X1 port map( A1 => n10272, A2 => n11073, B1 => n10271, B2 => 
                           n11070, C1 => n10273, C2 => n11067, ZN => n5318);
   U6265 : OAI222_X1 port map( A1 => n10272, A2 => n11337, B1 => n10271, B2 => 
                           n11334, C1 => n10273, C2 => n11331, ZN => n3885);
   U6266 : OAI222_X1 port map( A1 => n10240, A2 => n11073, B1 => n10239, B2 => 
                           n11070, C1 => n10241, C2 => n11067, ZN => n5277);
   U6267 : OAI222_X1 port map( A1 => n10240, A2 => n11337, B1 => n10239, B2 => 
                           n11334, C1 => n10241, C2 => n11331, ZN => n3844);
   U6268 : OAI222_X1 port map( A1 => n10208, A2 => n11073, B1 => n10205, B2 => 
                           n11070, C1 => n10209, C2 => n11067, ZN => n5236);
   U6269 : OAI222_X1 port map( A1 => n10208, A2 => n11337, B1 => n10205, B2 => 
                           n11334, C1 => n10209, C2 => n11331, ZN => n3803);
   U6270 : OAI222_X1 port map( A1 => n10174, A2 => n11073, B1 => n10173, B2 => 
                           n11070, C1 => n10175, C2 => n11067, ZN => n5195);
   U6271 : OAI222_X1 port map( A1 => n10174, A2 => n11337, B1 => n10173, B2 => 
                           n11334, C1 => n10175, C2 => n11331, ZN => n3762);
   U6272 : OAI222_X1 port map( A1 => n10142, A2 => n11074, B1 => n10141, B2 => 
                           n11071, C1 => n10143, C2 => n11068, ZN => n5154);
   U6273 : OAI222_X1 port map( A1 => n10142, A2 => n11338, B1 => n10141, B2 => 
                           n11335, C1 => n10143, C2 => n11332, ZN => n3721);
   U6274 : OAI222_X1 port map( A1 => n10110, A2 => n11074, B1 => n10109, B2 => 
                           n11071, C1 => n10111, C2 => n11068, ZN => n5113);
   U6275 : OAI222_X1 port map( A1 => n10110, A2 => n11338, B1 => n10109, B2 => 
                           n11335, C1 => n10111, C2 => n11332, ZN => n3680);
   U6276 : OAI222_X1 port map( A1 => n10078, A2 => n11074, B1 => n10077, B2 => 
                           n11071, C1 => n10079, C2 => n11068, ZN => n5072);
   U6277 : OAI222_X1 port map( A1 => n10078, A2 => n11338, B1 => n10077, B2 => 
                           n11335, C1 => n10079, C2 => n11332, ZN => n3639);
   U6278 : OAI222_X1 port map( A1 => n10046, A2 => n11074, B1 => n10045, B2 => 
                           n11071, C1 => n10047, C2 => n11068, ZN => n5031);
   U6279 : OAI222_X1 port map( A1 => n10046, A2 => n11338, B1 => n10045, B2 => 
                           n11335, C1 => n10047, C2 => n11332, ZN => n3598);
   U6280 : OAI222_X1 port map( A1 => n10014, A2 => n11074, B1 => n10013, B2 => 
                           n11071, C1 => n10015, C2 => n11068, ZN => n4990);
   U6281 : OAI222_X1 port map( A1 => n10014, A2 => n11338, B1 => n10013, B2 => 
                           n11335, C1 => n10015, C2 => n11332, ZN => n3557);
   U6282 : OAI222_X1 port map( A1 => n9652, A2 => n11074, B1 => n9651, B2 => 
                           n11071, C1 => n9653, C2 => n11068, ZN => n4949);
   U6283 : OAI222_X1 port map( A1 => n9652, A2 => n11338, B1 => n9651, B2 => 
                           n11335, C1 => n9653, C2 => n11332, ZN => n3516);
   U6284 : OAI222_X1 port map( A1 => n9620, A2 => n11074, B1 => n9619, B2 => 
                           n11071, C1 => n9621, C2 => n11068, ZN => n4908);
   U6285 : OAI222_X1 port map( A1 => n9620, A2 => n11338, B1 => n9619, B2 => 
                           n11335, C1 => n9621, C2 => n11332, ZN => n3475);
   U6286 : OAI222_X1 port map( A1 => n9588, A2 => n11074, B1 => n9587, B2 => 
                           n11071, C1 => n9589, C2 => n11068, ZN => n4867);
   U6287 : OAI222_X1 port map( A1 => n9588, A2 => n11338, B1 => n9587, B2 => 
                           n11335, C1 => n9589, C2 => n11332, ZN => n3434);
   U6288 : OAI222_X1 port map( A1 => n9254, A2 => n11074, B1 => n9253, B2 => 
                           n11071, C1 => n9255, C2 => n11068, ZN => n4826);
   U6289 : OAI222_X1 port map( A1 => n9254, A2 => n11338, B1 => n9253, B2 => 
                           n11335, C1 => n9255, C2 => n11332, ZN => n3393);
   U6290 : OAI222_X1 port map( A1 => n9190, A2 => n11074, B1 => n9189, B2 => 
                           n11071, C1 => n9191, C2 => n11068, ZN => n4785);
   U6291 : OAI222_X1 port map( A1 => n9190, A2 => n11338, B1 => n9189, B2 => 
                           n11335, C1 => n9191, C2 => n11332, ZN => n3352);
   U6292 : OAI222_X1 port map( A1 => n9158, A2 => n11074, B1 => n9157, B2 => 
                           n11071, C1 => n9159, C2 => n11068, ZN => n4744);
   U6293 : OAI222_X1 port map( A1 => n9158, A2 => n11338, B1 => n9157, B2 => 
                           n11335, C1 => n9159, C2 => n11332, ZN => n3311);
   U6294 : OAI222_X1 port map( A1 => n6308, A2 => n11074, B1 => n6307, B2 => 
                           n11071, C1 => n6309, C2 => n11068, ZN => n4703);
   U6295 : OAI222_X1 port map( A1 => n6308, A2 => n11338, B1 => n6307, B2 => 
                           n11335, C1 => n6309, C2 => n11332, ZN => n3270);
   U6296 : OAI222_X1 port map( A1 => n5991, A2 => n11075, B1 => n5990, B2 => 
                           n11072, C1 => n5992, C2 => n11069, ZN => n4662);
   U6297 : OAI222_X1 port map( A1 => n5991, A2 => n11339, B1 => n5990, B2 => 
                           n11336, C1 => n5992, C2 => n11333, ZN => n3229);
   U6298 : OAI222_X1 port map( A1 => n5927, A2 => n11075, B1 => n5926, B2 => 
                           n11072, C1 => n5928, C2 => n11069, ZN => n4621);
   U6299 : OAI222_X1 port map( A1 => n5927, A2 => n11339, B1 => n5926, B2 => 
                           n11336, C1 => n5928, C2 => n11333, ZN => n3188);
   U6300 : OAI222_X1 port map( A1 => n5895, A2 => n11075, B1 => n5894, B2 => 
                           n11072, C1 => n5896, C2 => n11069, ZN => n4580);
   U6301 : OAI222_X1 port map( A1 => n5895, A2 => n11339, B1 => n5894, B2 => 
                           n11336, C1 => n5896, C2 => n11333, ZN => n3147);
   U6302 : OAI222_X1 port map( A1 => n5863, A2 => n11075, B1 => n5862, B2 => 
                           n11072, C1 => n5864, C2 => n11069, ZN => n4539);
   U6303 : OAI222_X1 port map( A1 => n5863, A2 => n11339, B1 => n5862, B2 => 
                           n11336, C1 => n5864, C2 => n11333, ZN => n3106);
   U6304 : OAI222_X1 port map( A1 => n5831, A2 => n11075, B1 => n5830, B2 => 
                           n11072, C1 => n5832, C2 => n11069, ZN => n4498);
   U6305 : OAI222_X1 port map( A1 => n5831, A2 => n11339, B1 => n5830, B2 => 
                           n11336, C1 => n5832, C2 => n11333, ZN => n3065);
   U6306 : OAI222_X1 port map( A1 => n5799, A2 => n11075, B1 => n5798, B2 => 
                           n11072, C1 => n5800, C2 => n11069, ZN => n4457);
   U6307 : OAI222_X1 port map( A1 => n5799, A2 => n11339, B1 => n5798, B2 => 
                           n11336, C1 => n5800, C2 => n11333, ZN => n3024);
   U6308 : OAI222_X1 port map( A1 => n5767, A2 => n11075, B1 => n5766, B2 => 
                           n11072, C1 => n5768, C2 => n11069, ZN => n4416);
   U6309 : OAI222_X1 port map( A1 => n5767, A2 => n11339, B1 => n5766, B2 => 
                           n11336, C1 => n5768, C2 => n11333, ZN => n2983);
   U6310 : OAI222_X1 port map( A1 => n5735, A2 => n11075, B1 => n5734, B2 => 
                           n11072, C1 => n5736, C2 => n11069, ZN => n4300);
   U6311 : OAI222_X1 port map( A1 => n5735, A2 => n11339, B1 => n5734, B2 => 
                           n11336, C1 => n5736, C2 => n11333, ZN => n2800);
   U6312 : OAI222_X1 port map( A1 => n2337, A2 => n11097, B1 => n513, B2 => 
                           n11094, C1 => n1442, C2 => n11091, ZN => n5643);
   U6313 : OAI222_X1 port map( A1 => n10523, A2 => n11031, B1 => n10522, B2 => 
                           n11028, C1 => n10524, C2 => n11025, ZN => n5671);
   U6314 : OAI222_X1 port map( A1 => n2337, A2 => n11361, B1 => n513, B2 => 
                           n11358, C1 => n1442, C2 => n11355, ZN => n4210);
   U6315 : OAI222_X1 port map( A1 => n10523, A2 => n11295, B1 => n10522, B2 => 
                           n11292, C1 => n10524, C2 => n11289, ZN => n4238);
   U6316 : OAI222_X1 port map( A1 => n2325, A2 => n11097, B1 => n501, B2 => 
                           n11094, C1 => n1398, C2 => n11091, ZN => n5602);
   U6317 : OAI222_X1 port map( A1 => n10491, A2 => n11031, B1 => n10490, B2 => 
                           n11028, C1 => n10492, C2 => n11025, ZN => n5611);
   U6318 : OAI222_X1 port map( A1 => n2325, A2 => n11361, B1 => n501, B2 => 
                           n11358, C1 => n1398, C2 => n11355, ZN => n4169);
   U6319 : OAI222_X1 port map( A1 => n10491, A2 => n11295, B1 => n10490, B2 => 
                           n11292, C1 => n10492, C2 => n11289, ZN => n4178);
   U6320 : OAI222_X1 port map( A1 => n2313, A2 => n11097, B1 => n489, B2 => 
                           n11094, C1 => n1386, C2 => n11091, ZN => n5561);
   U6321 : OAI222_X1 port map( A1 => n10459, A2 => n11031, B1 => n10458, B2 => 
                           n11028, C1 => n10460, C2 => n11025, ZN => n5570);
   U6322 : OAI222_X1 port map( A1 => n2313, A2 => n11361, B1 => n489, B2 => 
                           n11358, C1 => n1386, C2 => n11355, ZN => n4128);
   U6323 : OAI222_X1 port map( A1 => n10459, A2 => n11295, B1 => n10458, B2 => 
                           n11292, C1 => n10460, C2 => n11289, ZN => n4137);
   U6324 : OAI222_X1 port map( A1 => n2301, A2 => n11097, B1 => n477, B2 => 
                           n11094, C1 => n1342, C2 => n11091, ZN => n5520);
   U6325 : OAI222_X1 port map( A1 => n10427, A2 => n11031, B1 => n10426, B2 => 
                           n11028, C1 => n10428, C2 => n11025, ZN => n5529);
   U6326 : OAI222_X1 port map( A1 => n2301, A2 => n11361, B1 => n477, B2 => 
                           n11358, C1 => n1342, C2 => n11355, ZN => n4087);
   U6327 : OAI222_X1 port map( A1 => n10427, A2 => n11295, B1 => n10426, B2 => 
                           n11292, C1 => n10428, C2 => n11289, ZN => n4096);
   U6328 : OAI222_X1 port map( A1 => n2289, A2 => n11097, B1 => n465, B2 => 
                           n11094, C1 => n1330, C2 => n11091, ZN => n5479);
   U6329 : OAI222_X1 port map( A1 => n10392, A2 => n11031, B1 => n10391, B2 => 
                           n11028, C1 => n10393, C2 => n11025, ZN => n5488);
   U6330 : OAI222_X1 port map( A1 => n2289, A2 => n11361, B1 => n465, B2 => 
                           n11358, C1 => n1330, C2 => n11355, ZN => n4046);
   U6331 : OAI222_X1 port map( A1 => n10392, A2 => n11295, B1 => n10391, B2 => 
                           n11292, C1 => n10393, C2 => n11289, ZN => n4055);
   U6332 : OAI222_X1 port map( A1 => n2277, A2 => n11097, B1 => n453, B2 => 
                           n11094, C1 => n1318, C2 => n11091, ZN => n5438);
   U6333 : OAI222_X1 port map( A1 => n10360, A2 => n11031, B1 => n10359, B2 => 
                           n11028, C1 => n10361, C2 => n11025, ZN => n5447);
   U6334 : OAI222_X1 port map( A1 => n2277, A2 => n11361, B1 => n453, B2 => 
                           n11358, C1 => n1318, C2 => n11355, ZN => n4005);
   U6335 : OAI222_X1 port map( A1 => n10360, A2 => n11295, B1 => n10359, B2 => 
                           n11292, C1 => n10361, C2 => n11289, ZN => n4014);
   U6336 : OAI222_X1 port map( A1 => n2265, A2 => n11097, B1 => n441, B2 => 
                           n11094, C1 => n1306, C2 => n11091, ZN => n5397);
   U6337 : OAI222_X1 port map( A1 => n10328, A2 => n11031, B1 => n10327, B2 => 
                           n11028, C1 => n10329, C2 => n11025, ZN => n5406);
   U6338 : OAI222_X1 port map( A1 => n2265, A2 => n11361, B1 => n441, B2 => 
                           n11358, C1 => n1306, C2 => n11355, ZN => n3964);
   U6339 : OAI222_X1 port map( A1 => n10328, A2 => n11295, B1 => n10327, B2 => 
                           n11292, C1 => n10329, C2 => n11289, ZN => n3973);
   U6340 : OAI222_X1 port map( A1 => n2253, A2 => n11097, B1 => n429, B2 => 
                           n11094, C1 => n1294, C2 => n11091, ZN => n5356);
   U6341 : OAI222_X1 port map( A1 => n10293, A2 => n11031, B1 => n10292, B2 => 
                           n11028, C1 => n10294, C2 => n11025, ZN => n5365);
   U6342 : OAI222_X1 port map( A1 => n2253, A2 => n11361, B1 => n429, B2 => 
                           n11358, C1 => n1294, C2 => n11355, ZN => n3923);
   U6343 : OAI222_X1 port map( A1 => n10293, A2 => n11295, B1 => n10292, B2 => 
                           n11292, C1 => n10294, C2 => n11289, ZN => n3932);
   U6344 : OAI222_X1 port map( A1 => n2241, A2 => n11097, B1 => n417, B2 => 
                           n11094, C1 => n1282, C2 => n11091, ZN => n5315);
   U6345 : OAI222_X1 port map( A1 => n10261, A2 => n11031, B1 => n10260, B2 => 
                           n11028, C1 => n10262, C2 => n11025, ZN => n5324);
   U6346 : OAI222_X1 port map( A1 => n2241, A2 => n11361, B1 => n417, B2 => 
                           n11358, C1 => n1282, C2 => n11355, ZN => n3882);
   U6347 : OAI222_X1 port map( A1 => n10261, A2 => n11295, B1 => n10260, B2 => 
                           n11292, C1 => n10262, C2 => n11289, ZN => n3891);
   U6348 : OAI222_X1 port map( A1 => n2229, A2 => n11097, B1 => n405, B2 => 
                           n11094, C1 => n1270, C2 => n11091, ZN => n5274);
   U6349 : OAI222_X1 port map( A1 => n10229, A2 => n11031, B1 => n10228, B2 => 
                           n11028, C1 => n10230, C2 => n11025, ZN => n5283);
   U6350 : OAI222_X1 port map( A1 => n2229, A2 => n11361, B1 => n405, B2 => 
                           n11358, C1 => n1270, C2 => n11355, ZN => n3841);
   U6351 : OAI222_X1 port map( A1 => n10229, A2 => n11295, B1 => n10228, B2 => 
                           n11292, C1 => n10230, C2 => n11289, ZN => n3850);
   U6352 : OAI222_X1 port map( A1 => n2217, A2 => n11097, B1 => n393, B2 => 
                           n11094, C1 => n1258, C2 => n11091, ZN => n5233);
   U6353 : OAI222_X1 port map( A1 => n10195, A2 => n11031, B1 => n10194, B2 => 
                           n11028, C1 => n10196, C2 => n11025, ZN => n5242);
   U6354 : OAI222_X1 port map( A1 => n2217, A2 => n11361, B1 => n393, B2 => 
                           n11358, C1 => n1258, C2 => n11355, ZN => n3800);
   U6355 : OAI222_X1 port map( A1 => n10195, A2 => n11295, B1 => n10194, B2 => 
                           n11292, C1 => n10196, C2 => n11289, ZN => n3809);
   U6356 : OAI222_X1 port map( A1 => n2173_port, A2 => n11097, B1 => n381, B2 
                           => n11094, C1 => n1246, C2 => n11091, ZN => n5192);
   U6357 : OAI222_X1 port map( A1 => n10163, A2 => n11031, B1 => n10162, B2 => 
                           n11028, C1 => n10164, C2 => n11025, ZN => n5201);
   U6358 : OAI222_X1 port map( A1 => n2173_port, A2 => n11361, B1 => n381, B2 
                           => n11358, C1 => n1246, C2 => n11355, ZN => n3759);
   U6359 : OAI222_X1 port map( A1 => n10163, A2 => n11295, B1 => n10162, B2 => 
                           n11292, C1 => n10164, C2 => n11289, ZN => n3768);
   U6360 : OAI222_X1 port map( A1 => n2161, A2 => n11098, B1 => n369, B2 => 
                           n11095, C1 => n1234, C2 => n11092, ZN => n5151);
   U6361 : OAI222_X1 port map( A1 => n10131, A2 => n11032, B1 => n10130, B2 => 
                           n11029, C1 => n10132, C2 => n11026, ZN => n5160);
   U6362 : OAI222_X1 port map( A1 => n2161, A2 => n11362, B1 => n369, B2 => 
                           n11359, C1 => n1234, C2 => n11356, ZN => n3718);
   U6363 : OAI222_X1 port map( A1 => n10131, A2 => n11296, B1 => n10130, B2 => 
                           n11293, C1 => n10132, C2 => n11290, ZN => n3727);
   U6364 : OAI222_X1 port map( A1 => n2149, A2 => n11098, B1 => n357, B2 => 
                           n11095, C1 => n1222, C2 => n11092, ZN => n5110);
   U6365 : OAI222_X1 port map( A1 => n10099, A2 => n11032, B1 => n10098, B2 => 
                           n11029, C1 => n10100, C2 => n11026, ZN => n5119);
   U6366 : OAI222_X1 port map( A1 => n2149, A2 => n11362, B1 => n357, B2 => 
                           n11359, C1 => n1222, C2 => n11356, ZN => n3677);
   U6367 : OAI222_X1 port map( A1 => n10099, A2 => n11296, B1 => n10098, B2 => 
                           n11293, C1 => n10100, C2 => n11290, ZN => n3686);
   U6368 : OAI222_X1 port map( A1 => n2105, A2 => n11098, B1 => n345, B2 => 
                           n11095, C1 => n1210, C2 => n11092, ZN => n5069);
   U6369 : OAI222_X1 port map( A1 => n10067, A2 => n11032, B1 => n10066, B2 => 
                           n11029, C1 => n10068, C2 => n11026, ZN => n5078);
   U6370 : OAI222_X1 port map( A1 => n2105, A2 => n11362, B1 => n345, B2 => 
                           n11359, C1 => n1210, C2 => n11356, ZN => n3636);
   U6371 : OAI222_X1 port map( A1 => n10067, A2 => n11296, B1 => n10066, B2 => 
                           n11293, C1 => n10068, C2 => n11290, ZN => n3645);
   U6372 : OAI222_X1 port map( A1 => n2093, A2 => n11098, B1 => n333, B2 => 
                           n11095, C1 => n1198, C2 => n11092, ZN => n5028);
   U6373 : OAI222_X1 port map( A1 => n10035, A2 => n11032, B1 => n10034, B2 => 
                           n11029, C1 => n10036, C2 => n11026, ZN => n5037);
   U6374 : OAI222_X1 port map( A1 => n2093, A2 => n11362, B1 => n333, B2 => 
                           n11359, C1 => n1198, C2 => n11356, ZN => n3595);
   U6375 : OAI222_X1 port map( A1 => n10035, A2 => n11296, B1 => n10034, B2 => 
                           n11293, C1 => n10036, C2 => n11290, ZN => n3604);
   U6376 : OAI222_X1 port map( A1 => n2049, A2 => n11098, B1 => n321, B2 => 
                           n11095, C1 => n1186, C2 => n11092, ZN => n4987);
   U6377 : OAI222_X1 port map( A1 => n10003, A2 => n11032, B1 => n10002, B2 => 
                           n11029, C1 => n10004, C2 => n11026, ZN => n4996);
   U6378 : OAI222_X1 port map( A1 => n2049, A2 => n11362, B1 => n321, B2 => 
                           n11359, C1 => n1186, C2 => n11356, ZN => n3554);
   U6379 : OAI222_X1 port map( A1 => n10003, A2 => n11296, B1 => n10002, B2 => 
                           n11293, C1 => n10004, C2 => n11290, ZN => n3563);
   U6380 : OAI222_X1 port map( A1 => n2037, A2 => n11098, B1 => n309, B2 => 
                           n11095, C1 => n1174, C2 => n11092, ZN => n4946);
   U6381 : OAI222_X1 port map( A1 => n9641, A2 => n11032, B1 => n9640, B2 => 
                           n11029, C1 => n9642, C2 => n11026, ZN => n4955);
   U6382 : OAI222_X1 port map( A1 => n2037, A2 => n11362, B1 => n309, B2 => 
                           n11359, C1 => n1174, C2 => n11356, ZN => n3513);
   U6383 : OAI222_X1 port map( A1 => n9641, A2 => n11296, B1 => n9640, B2 => 
                           n11293, C1 => n9642, C2 => n11290, ZN => n3522);
   U6384 : OAI222_X1 port map( A1 => n2025, A2 => n11098, B1 => n297, B2 => 
                           n11095, C1 => n1162, C2 => n11092, ZN => n4905);
   U6385 : OAI222_X1 port map( A1 => n9609, A2 => n11032, B1 => n9608, B2 => 
                           n11029, C1 => n9610, C2 => n11026, ZN => n4914);
   U6386 : OAI222_X1 port map( A1 => n2025, A2 => n11362, B1 => n297, B2 => 
                           n11359, C1 => n1162, C2 => n11356, ZN => n3472);
   U6387 : OAI222_X1 port map( A1 => n9609, A2 => n11296, B1 => n9608, B2 => 
                           n11293, C1 => n9610, C2 => n11290, ZN => n3481);
   U6388 : OAI222_X1 port map( A1 => n2013, A2 => n11098, B1 => n285, B2 => 
                           n11095, C1 => n1150, C2 => n11092, ZN => n4864);
   U6389 : OAI222_X1 port map( A1 => n9577, A2 => n11032, B1 => n9576, B2 => 
                           n11029, C1 => n9578, C2 => n11026, ZN => n4873);
   U6390 : OAI222_X1 port map( A1 => n2013, A2 => n11362, B1 => n285, B2 => 
                           n11359, C1 => n1150, C2 => n11356, ZN => n3431);
   U6391 : OAI222_X1 port map( A1 => n9577, A2 => n11296, B1 => n9576, B2 => 
                           n11293, C1 => n9578, C2 => n11290, ZN => n3440);
   U6392 : OAI222_X1 port map( A1 => n2001, A2 => n11098, B1 => n273, B2 => 
                           n11095, C1 => n1138, C2 => n11092, ZN => n4823);
   U6393 : OAI222_X1 port map( A1 => n9211, A2 => n11032, B1 => n9210, B2 => 
                           n11029, C1 => n9212, C2 => n11026, ZN => n4832);
   U6394 : OAI222_X1 port map( A1 => n2001, A2 => n11362, B1 => n273, B2 => 
                           n11359, C1 => n1138, C2 => n11356, ZN => n3390);
   U6395 : OAI222_X1 port map( A1 => n9211, A2 => n11296, B1 => n9210, B2 => 
                           n11293, C1 => n9212, C2 => n11290, ZN => n3399);
   U6396 : OAI222_X1 port map( A1 => n1989, A2 => n11098, B1 => n261, B2 => 
                           n11095, C1 => n1126, C2 => n11092, ZN => n4782);
   U6397 : OAI222_X1 port map( A1 => n9179, A2 => n11032, B1 => n9178, B2 => 
                           n11029, C1 => n9180, C2 => n11026, ZN => n4791);
   U6398 : OAI222_X1 port map( A1 => n1989, A2 => n11362, B1 => n261, B2 => 
                           n11359, C1 => n1126, C2 => n11356, ZN => n3349);
   U6399 : OAI222_X1 port map( A1 => n9179, A2 => n11296, B1 => n9178, B2 => 
                           n11293, C1 => n9180, C2 => n11290, ZN => n3358);
   U6400 : OAI222_X1 port map( A1 => n1977, A2 => n11098, B1 => n249, B2 => 
                           n11095, C1 => n1114, C2 => n11092, ZN => n4741);
   U6401 : OAI222_X1 port map( A1 => n9147, A2 => n11032, B1 => n9146, B2 => 
                           n11029, C1 => n9148, C2 => n11026, ZN => n4750);
   U6402 : OAI222_X1 port map( A1 => n1977, A2 => n11362, B1 => n249, B2 => 
                           n11359, C1 => n1114, C2 => n11356, ZN => n3308);
   U6403 : OAI222_X1 port map( A1 => n9147, A2 => n11296, B1 => n9146, B2 => 
                           n11293, C1 => n9148, C2 => n11290, ZN => n3317);
   U6404 : OAI222_X1 port map( A1 => n1965, A2 => n11098, B1 => n237, B2 => 
                           n11095, C1 => n1102, C2 => n11092, ZN => n4700);
   U6405 : OAI222_X1 port map( A1 => n6012, A2 => n11032, B1 => n6011, B2 => 
                           n11029, C1 => n6044, C2 => n11026, ZN => n4709);
   U6406 : OAI222_X1 port map( A1 => n1965, A2 => n11362, B1 => n237, B2 => 
                           n11359, C1 => n1102, C2 => n11356, ZN => n3267);
   U6407 : OAI222_X1 port map( A1 => n6012, A2 => n11296, B1 => n6011, B2 => 
                           n11293, C1 => n6044, C2 => n11290, ZN => n3276);
   U6408 : OAI222_X1 port map( A1 => n1953, A2 => n11099, B1 => n225, B2 => 
                           n11096, C1 => n1090, C2 => n11093, ZN => n4659);
   U6409 : OAI222_X1 port map( A1 => n5948, A2 => n11033, B1 => n5947, B2 => 
                           n11030, C1 => n5981, C2 => n11027, ZN => n4668);
   U6410 : OAI222_X1 port map( A1 => n1953, A2 => n11363, B1 => n225, B2 => 
                           n11360, C1 => n1090, C2 => n11357, ZN => n3226);
   U6411 : OAI222_X1 port map( A1 => n5948, A2 => n11297, B1 => n5947, B2 => 
                           n11294, C1 => n5981, C2 => n11291, ZN => n3235);
   U6412 : OAI222_X1 port map( A1 => n1941, A2 => n11099, B1 => n213, B2 => 
                           n11096, C1 => n1078, C2 => n11093, ZN => n4618);
   U6413 : OAI222_X1 port map( A1 => n5916, A2 => n11033, B1 => n5915, B2 => 
                           n11030, C1 => n5917, C2 => n11027, ZN => n4627);
   U6414 : OAI222_X1 port map( A1 => n1941, A2 => n11363, B1 => n213, B2 => 
                           n11360, C1 => n1078, C2 => n11357, ZN => n3185);
   U6415 : OAI222_X1 port map( A1 => n5916, A2 => n11297, B1 => n5915, B2 => 
                           n11294, C1 => n5917, C2 => n11291, ZN => n3194);
   U6416 : OAI222_X1 port map( A1 => n1929, A2 => n11099, B1 => n201, B2 => 
                           n11096, C1 => n1066, C2 => n11093, ZN => n4577);
   U6417 : OAI222_X1 port map( A1 => n5884, A2 => n11033, B1 => n5883, B2 => 
                           n11030, C1 => n5885, C2 => n11027, ZN => n4586);
   U6418 : OAI222_X1 port map( A1 => n1929, A2 => n11363, B1 => n201, B2 => 
                           n11360, C1 => n1066, C2 => n11357, ZN => n3144);
   U6419 : OAI222_X1 port map( A1 => n5884, A2 => n11297, B1 => n5883, B2 => 
                           n11294, C1 => n5885, C2 => n11291, ZN => n3153);
   U6420 : OAI222_X1 port map( A1 => n1917, A2 => n11099, B1 => n189, B2 => 
                           n11096, C1 => n1054, C2 => n11093, ZN => n4536);
   U6421 : OAI222_X1 port map( A1 => n5852, A2 => n11033, B1 => n5851, B2 => 
                           n11030, C1 => n5853, C2 => n11027, ZN => n4545);
   U6422 : OAI222_X1 port map( A1 => n1917, A2 => n11363, B1 => n189, B2 => 
                           n11360, C1 => n1054, C2 => n11357, ZN => n3103);
   U6423 : OAI222_X1 port map( A1 => n5852, A2 => n11297, B1 => n5851, B2 => 
                           n11294, C1 => n5853, C2 => n11291, ZN => n3112);
   U6424 : OAI222_X1 port map( A1 => n1905, A2 => n11099, B1 => n177, B2 => 
                           n11096, C1 => n1042, C2 => n11093, ZN => n4495);
   U6425 : OAI222_X1 port map( A1 => n5820, A2 => n11033, B1 => n5819, B2 => 
                           n11030, C1 => n5821, C2 => n11027, ZN => n4504);
   U6426 : OAI222_X1 port map( A1 => n1905, A2 => n11363, B1 => n177, B2 => 
                           n11360, C1 => n1042, C2 => n11357, ZN => n3062);
   U6427 : OAI222_X1 port map( A1 => n5820, A2 => n11297, B1 => n5819, B2 => 
                           n11294, C1 => n5821, C2 => n11291, ZN => n3071);
   U6428 : OAI222_X1 port map( A1 => n5788, A2 => n11033, B1 => n5787, B2 => 
                           n11030, C1 => n5789, C2 => n11027, ZN => n4463);
   U6429 : OAI222_X1 port map( A1 => n5788, A2 => n11297, B1 => n5787, B2 => 
                           n11294, C1 => n5789, C2 => n11291, ZN => n3030);
   U6430 : OAI222_X1 port map( A1 => n5756, A2 => n11033, B1 => n5755, B2 => 
                           n11030, C1 => n5757, C2 => n11027, ZN => n4422);
   U6431 : OAI222_X1 port map( A1 => n5756, A2 => n11297, B1 => n5755, B2 => 
                           n11294, C1 => n5757, C2 => n11291, ZN => n2989);
   U6432 : OAI222_X1 port map( A1 => n5724, A2 => n11033, B1 => n5723, B2 => 
                           n11030, C1 => n5725, C2 => n11027, ZN => n4315);
   U6433 : OAI222_X1 port map( A1 => n5724, A2 => n11297, B1 => n5723, B2 => 
                           n11294, C1 => n5725, C2 => n11291, ZN => n2815);
   U6434 : OAI222_X1 port map( A1 => n1893, A2 => n11099, B1 => n165, B2 => 
                           n11096, C1 => n12785, C2 => n11093, ZN => n4454);
   U6435 : OAI222_X1 port map( A1 => n1893, A2 => n11363, B1 => n165, B2 => 
                           n11360, C1 => n12785, C2 => n11357, ZN => n3021);
   U6436 : OAI222_X1 port map( A1 => n1881, A2 => n11099, B1 => n153, B2 => 
                           n11096, C1 => n12784, C2 => n11093, ZN => n4413);
   U6437 : OAI222_X1 port map( A1 => n1881, A2 => n11363, B1 => n153, B2 => 
                           n11360, C1 => n12784, C2 => n11357, ZN => n2980);
   U6438 : OAI222_X1 port map( A1 => n1869, A2 => n11099, B1 => n141, B2 => 
                           n11096, C1 => n12783, C2 => n11093, ZN => n4284);
   U6439 : OAI222_X1 port map( A1 => n1869, A2 => n11363, B1 => n141, B2 => 
                           n11360, C1 => n12783, C2 => n11357, ZN => n2752);
   U6440 : OAI222_X1 port map( A1 => n995, A2 => n11088, B1 => n1859, B2 => 
                           n11085, C1 => n1409, C2 => n11082, ZN => n5642);
   U6441 : OAI222_X1 port map( A1 => n995, A2 => n11352, B1 => n1859, B2 => 
                           n11349, C1 => n1409, C2 => n11346, ZN => n4209);
   U6442 : OAI222_X1 port map( A1 => n991, A2 => n11088, B1 => n1855, B2 => 
                           n11085, C1 => n1397, C2 => n11082, ZN => n5601);
   U6443 : OAI222_X1 port map( A1 => n991, A2 => n11352, B1 => n1855, B2 => 
                           n11349, C1 => n1397, C2 => n11346, ZN => n4168);
   U6444 : OAI222_X1 port map( A1 => n987, A2 => n11088, B1 => n1851, B2 => 
                           n11085, C1 => n1385, C2 => n11082, ZN => n5560);
   U6445 : OAI222_X1 port map( A1 => n987, A2 => n11352, B1 => n1851, B2 => 
                           n11349, C1 => n1385, C2 => n11346, ZN => n4127);
   U6446 : OAI222_X1 port map( A1 => n983, A2 => n11088, B1 => n1847, B2 => 
                           n11085, C1 => n1341, C2 => n11082, ZN => n5519);
   U6447 : OAI222_X1 port map( A1 => n983, A2 => n11352, B1 => n1847, B2 => 
                           n11349, C1 => n1341, C2 => n11346, ZN => n4086);
   U6448 : OAI222_X1 port map( A1 => n979, A2 => n11088, B1 => n1843, B2 => 
                           n11085, C1 => n1329, C2 => n11082, ZN => n5478);
   U6449 : OAI222_X1 port map( A1 => n979, A2 => n11352, B1 => n1843, B2 => 
                           n11349, C1 => n1329, C2 => n11346, ZN => n4045);
   U6450 : OAI222_X1 port map( A1 => n975, A2 => n11088, B1 => n1839, B2 => 
                           n11085, C1 => n1317, C2 => n11082, ZN => n5437);
   U6451 : OAI222_X1 port map( A1 => n975, A2 => n11352, B1 => n1839, B2 => 
                           n11349, C1 => n1317, C2 => n11346, ZN => n4004);
   U6452 : OAI222_X1 port map( A1 => n971, A2 => n11088, B1 => n1835, B2 => 
                           n11085, C1 => n1305, C2 => n11082, ZN => n5396);
   U6453 : OAI222_X1 port map( A1 => n971, A2 => n11352, B1 => n1835, B2 => 
                           n11349, C1 => n1305, C2 => n11346, ZN => n3963);
   U6454 : OAI222_X1 port map( A1 => n967, A2 => n11088, B1 => n1831, B2 => 
                           n11085, C1 => n1293, C2 => n11082, ZN => n5355);
   U6455 : OAI222_X1 port map( A1 => n967, A2 => n11352, B1 => n1831, B2 => 
                           n11349, C1 => n1293, C2 => n11346, ZN => n3922);
   U6456 : OAI222_X1 port map( A1 => n963, A2 => n11088, B1 => n1827, B2 => 
                           n11085, C1 => n1281, C2 => n11082, ZN => n5314);
   U6457 : OAI222_X1 port map( A1 => n963, A2 => n11352, B1 => n1827, B2 => 
                           n11349, C1 => n1281, C2 => n11346, ZN => n3881);
   U6458 : OAI222_X1 port map( A1 => n959, A2 => n11088, B1 => n1823, B2 => 
                           n11085, C1 => n1269, C2 => n11082, ZN => n5273);
   U6459 : OAI222_X1 port map( A1 => n959, A2 => n11352, B1 => n1823, B2 => 
                           n11349, C1 => n1269, C2 => n11346, ZN => n3840);
   U6460 : OAI222_X1 port map( A1 => n955, A2 => n11088, B1 => n1819, B2 => 
                           n11085, C1 => n1257, C2 => n11082, ZN => n5232);
   U6461 : OAI222_X1 port map( A1 => n955, A2 => n11352, B1 => n1819, B2 => 
                           n11349, C1 => n1257, C2 => n11346, ZN => n3799);
   U6462 : OAI222_X1 port map( A1 => n951, A2 => n11088, B1 => n1815, B2 => 
                           n11085, C1 => n1245, C2 => n11082, ZN => n5191);
   U6463 : OAI222_X1 port map( A1 => n951, A2 => n11352, B1 => n1815, B2 => 
                           n11349, C1 => n1245, C2 => n11346, ZN => n3758);
   U6464 : OAI222_X1 port map( A1 => n947, A2 => n11089, B1 => n1811, B2 => 
                           n11086, C1 => n1233, C2 => n11083, ZN => n5150);
   U6465 : OAI222_X1 port map( A1 => n947, A2 => n11353, B1 => n1811, B2 => 
                           n11350, C1 => n1233, C2 => n11347, ZN => n3717);
   U6466 : OAI222_X1 port map( A1 => n943, A2 => n11089, B1 => n1807, B2 => 
                           n11086, C1 => n1221, C2 => n11083, ZN => n5109);
   U6467 : OAI222_X1 port map( A1 => n943, A2 => n11353, B1 => n1807, B2 => 
                           n11350, C1 => n1221, C2 => n11347, ZN => n3676);
   U6468 : OAI222_X1 port map( A1 => n939, A2 => n11089, B1 => n1803, B2 => 
                           n11086, C1 => n1209, C2 => n11083, ZN => n5068);
   U6469 : OAI222_X1 port map( A1 => n939, A2 => n11353, B1 => n1803, B2 => 
                           n11350, C1 => n1209, C2 => n11347, ZN => n3635);
   U6470 : OAI222_X1 port map( A1 => n935, A2 => n11089, B1 => n1799, B2 => 
                           n11086, C1 => n1197, C2 => n11083, ZN => n5027);
   U6471 : OAI222_X1 port map( A1 => n935, A2 => n11353, B1 => n1799, B2 => 
                           n11350, C1 => n1197, C2 => n11347, ZN => n3594);
   U6472 : OAI222_X1 port map( A1 => n931, A2 => n11089, B1 => n1795, B2 => 
                           n11086, C1 => n1185, C2 => n11083, ZN => n4986);
   U6473 : OAI222_X1 port map( A1 => n931, A2 => n11353, B1 => n1795, B2 => 
                           n11350, C1 => n1185, C2 => n11347, ZN => n3553);
   U6474 : OAI222_X1 port map( A1 => n927, A2 => n11089, B1 => n1791, B2 => 
                           n11086, C1 => n1173, C2 => n11083, ZN => n4945);
   U6475 : OAI222_X1 port map( A1 => n927, A2 => n11353, B1 => n1791, B2 => 
                           n11350, C1 => n1173, C2 => n11347, ZN => n3512);
   U6476 : OAI222_X1 port map( A1 => n923, A2 => n11089, B1 => n1787, B2 => 
                           n11086, C1 => n1161, C2 => n11083, ZN => n4904);
   U6477 : OAI222_X1 port map( A1 => n923, A2 => n11353, B1 => n1787, B2 => 
                           n11350, C1 => n1161, C2 => n11347, ZN => n3471);
   U6478 : OAI222_X1 port map( A1 => n919, A2 => n11089, B1 => n1783, B2 => 
                           n11086, C1 => n1149, C2 => n11083, ZN => n4863);
   U6479 : OAI222_X1 port map( A1 => n919, A2 => n11353, B1 => n1783, B2 => 
                           n11350, C1 => n1149, C2 => n11347, ZN => n3430);
   U6480 : OAI222_X1 port map( A1 => n915, A2 => n11089, B1 => n1779, B2 => 
                           n11086, C1 => n1137, C2 => n11083, ZN => n4822);
   U6481 : OAI222_X1 port map( A1 => n915, A2 => n11353, B1 => n1779, B2 => 
                           n11350, C1 => n1137, C2 => n11347, ZN => n3389);
   U6482 : OAI222_X1 port map( A1 => n911, A2 => n11089, B1 => n1775, B2 => 
                           n11086, C1 => n1125, C2 => n11083, ZN => n4781);
   U6483 : OAI222_X1 port map( A1 => n911, A2 => n11353, B1 => n1775, B2 => 
                           n11350, C1 => n1125, C2 => n11347, ZN => n3348);
   U6484 : OAI222_X1 port map( A1 => n907, A2 => n11089, B1 => n1771, B2 => 
                           n11086, C1 => n1113, C2 => n11083, ZN => n4740);
   U6485 : OAI222_X1 port map( A1 => n907, A2 => n11353, B1 => n1771, B2 => 
                           n11350, C1 => n1113, C2 => n11347, ZN => n3307);
   U6486 : OAI222_X1 port map( A1 => n903, A2 => n11089, B1 => n1767, B2 => 
                           n11086, C1 => n1101, C2 => n11083, ZN => n4699);
   U6487 : OAI222_X1 port map( A1 => n903, A2 => n11353, B1 => n1767, B2 => 
                           n11350, C1 => n1101, C2 => n11347, ZN => n3266);
   U6488 : OAI222_X1 port map( A1 => n899, A2 => n11090, B1 => n1763, B2 => 
                           n11087, C1 => n1089, C2 => n11084, ZN => n4658);
   U6489 : OAI222_X1 port map( A1 => n899, A2 => n11354, B1 => n1763, B2 => 
                           n11351, C1 => n1089, C2 => n11348, ZN => n3225);
   U6490 : OAI222_X1 port map( A1 => n895, A2 => n11090, B1 => n1759, B2 => 
                           n11087, C1 => n1077, C2 => n11084, ZN => n4617);
   U6491 : OAI222_X1 port map( A1 => n895, A2 => n11354, B1 => n1759, B2 => 
                           n11351, C1 => n1077, C2 => n11348, ZN => n3184);
   U6492 : OAI222_X1 port map( A1 => n891, A2 => n11090, B1 => n1755, B2 => 
                           n11087, C1 => n1065, C2 => n11084, ZN => n4576);
   U6493 : OAI222_X1 port map( A1 => n891, A2 => n11354, B1 => n1755, B2 => 
                           n11351, C1 => n1065, C2 => n11348, ZN => n3143);
   U6494 : OAI222_X1 port map( A1 => n887, A2 => n11090, B1 => n1751, B2 => 
                           n11087, C1 => n1053, C2 => n11084, ZN => n4535);
   U6495 : OAI222_X1 port map( A1 => n887, A2 => n11354, B1 => n1751, B2 => 
                           n11351, C1 => n1053, C2 => n11348, ZN => n3102);
   U6496 : OAI222_X1 port map( A1 => n883, A2 => n11090, B1 => n1747, B2 => 
                           n11087, C1 => n1041, C2 => n11084, ZN => n4494);
   U6497 : OAI222_X1 port map( A1 => n883, A2 => n11354, B1 => n1747, B2 => 
                           n11351, C1 => n1041, C2 => n11348, ZN => n3061);
   U6498 : OAI222_X1 port map( A1 => n879, A2 => n11090, B1 => n1743, B2 => 
                           n11087, C1 => n1029, C2 => n11084, ZN => n4453);
   U6499 : OAI222_X1 port map( A1 => n879, A2 => n11354, B1 => n1743, B2 => 
                           n11351, C1 => n1029, C2 => n11348, ZN => n3020);
   U6500 : OAI222_X1 port map( A1 => n875, A2 => n11090, B1 => n1739, B2 => 
                           n11087, C1 => n12787, C2 => n11084, ZN => n4412);
   U6501 : OAI222_X1 port map( A1 => n875, A2 => n11354, B1 => n1739, B2 => 
                           n11351, C1 => n12787, C2 => n11348, ZN => n2979);
   U6502 : OAI222_X1 port map( A1 => n871, A2 => n11090, B1 => n1735, B2 => 
                           n11087, C1 => n12786, C2 => n11084, ZN => n4283);
   U6503 : OAI222_X1 port map( A1 => n871, A2 => n11354, B1 => n1735, B2 => 
                           n11351, C1 => n12786, C2 => n11348, ZN => n2751);
   U6504 : AOI222_X1 port map( A1 => n10923, A2 => n9376, B1 => n10920, B2 => 
                           n9312, C1 => n10917, C2 => n9344, ZN => n5679);
   U6505 : AOI222_X1 port map( A1 => n11187, A2 => n9376, B1 => n11184, B2 => 
                           n9312, C1 => n11181, C2 => n9344, ZN => n4246);
   U6506 : AOI222_X1 port map( A1 => n10923, A2 => n9377, B1 => n10920, B2 => 
                           n9313, C1 => n10917, C2 => n9345, ZN => n5615);
   U6507 : AOI222_X1 port map( A1 => n11187, A2 => n9377, B1 => n11184, B2 => 
                           n9313, C1 => n11181, C2 => n9345, ZN => n4182);
   U6508 : AOI222_X1 port map( A1 => n10923, A2 => n9378, B1 => n10920, B2 => 
                           n9314, C1 => n10917, C2 => n9346, ZN => n5574);
   U6509 : AOI222_X1 port map( A1 => n11187, A2 => n9378, B1 => n11184, B2 => 
                           n9314, C1 => n11181, C2 => n9346, ZN => n4141);
   U6510 : AOI222_X1 port map( A1 => n10923, A2 => n9379, B1 => n10920, B2 => 
                           n9315, C1 => n10917, C2 => n9347, ZN => n5533);
   U6511 : AOI222_X1 port map( A1 => n11187, A2 => n9379, B1 => n11184, B2 => 
                           n9315, C1 => n11181, C2 => n9347, ZN => n4100);
   U6512 : AOI222_X1 port map( A1 => n10923, A2 => n9380, B1 => n10920, B2 => 
                           n9316, C1 => n10917, C2 => n9348, ZN => n5492);
   U6513 : AOI222_X1 port map( A1 => n11187, A2 => n9380, B1 => n11184, B2 => 
                           n9316, C1 => n11181, C2 => n9348, ZN => n4059);
   U6514 : AOI222_X1 port map( A1 => n10923, A2 => n9381, B1 => n10920, B2 => 
                           n9317, C1 => n10917, C2 => n9349, ZN => n5451);
   U6515 : AOI222_X1 port map( A1 => n11187, A2 => n9381, B1 => n11184, B2 => 
                           n9317, C1 => n11181, C2 => n9349, ZN => n4018);
   U6516 : AOI222_X1 port map( A1 => n10923, A2 => n9382, B1 => n10920, B2 => 
                           n9318, C1 => n10917, C2 => n9350, ZN => n5410);
   U6517 : AOI222_X1 port map( A1 => n11187, A2 => n9382, B1 => n11184, B2 => 
                           n9318, C1 => n11181, C2 => n9350, ZN => n3977);
   U6518 : AOI222_X1 port map( A1 => n10923, A2 => n9383, B1 => n10920, B2 => 
                           n9319, C1 => n10917, C2 => n9351, ZN => n5369);
   U6519 : AOI222_X1 port map( A1 => n11187, A2 => n9383, B1 => n11184, B2 => 
                           n9319, C1 => n11181, C2 => n9351, ZN => n3936);
   U6520 : AOI222_X1 port map( A1 => n10923, A2 => n9384, B1 => n10920, B2 => 
                           n9320, C1 => n10917, C2 => n9352, ZN => n5328);
   U6521 : AOI222_X1 port map( A1 => n11187, A2 => n9384, B1 => n11184, B2 => 
                           n9320, C1 => n11181, C2 => n9352, ZN => n3895);
   U6522 : AOI222_X1 port map( A1 => n10923, A2 => n9385, B1 => n10920, B2 => 
                           n9321, C1 => n10917, C2 => n9353, ZN => n5287);
   U6523 : AOI222_X1 port map( A1 => n11187, A2 => n9385, B1 => n11184, B2 => 
                           n9321, C1 => n11181, C2 => n9353, ZN => n3854);
   U6524 : AOI222_X1 port map( A1 => n10923, A2 => n9386, B1 => n10920, B2 => 
                           n9322, C1 => n10917, C2 => n9354, ZN => n5246);
   U6525 : AOI222_X1 port map( A1 => n11187, A2 => n9386, B1 => n11184, B2 => 
                           n9322, C1 => n11181, C2 => n9354, ZN => n3813);
   U6526 : AOI222_X1 port map( A1 => n10923, A2 => n9387, B1 => n10920, B2 => 
                           n9323, C1 => n10917, C2 => n9355, ZN => n5205);
   U6527 : AOI222_X1 port map( A1 => n11187, A2 => n9387, B1 => n11184, B2 => 
                           n9323, C1 => n11181, C2 => n9355, ZN => n3772);
   U6528 : AOI222_X1 port map( A1 => n10924, A2 => n9388, B1 => n10921, B2 => 
                           n9324, C1 => n10918, C2 => n9356, ZN => n5164);
   U6529 : AOI222_X1 port map( A1 => n11188, A2 => n9388, B1 => n11185, B2 => 
                           n9324, C1 => n11182, C2 => n9356, ZN => n3731);
   U6530 : AOI222_X1 port map( A1 => n10924, A2 => n9389, B1 => n10921, B2 => 
                           n9325, C1 => n10918, C2 => n9357, ZN => n5123);
   U6531 : AOI222_X1 port map( A1 => n11188, A2 => n9389, B1 => n11185, B2 => 
                           n9325, C1 => n11182, C2 => n9357, ZN => n3690);
   U6532 : AOI222_X1 port map( A1 => n10924, A2 => n9390, B1 => n10921, B2 => 
                           n9326, C1 => n10918, C2 => n9358, ZN => n5082);
   U6533 : AOI222_X1 port map( A1 => n11188, A2 => n9390, B1 => n11185, B2 => 
                           n9326, C1 => n11182, C2 => n9358, ZN => n3649);
   U6534 : AOI222_X1 port map( A1 => n10924, A2 => n9391, B1 => n10921, B2 => 
                           n9327, C1 => n10918, C2 => n9359, ZN => n5041);
   U6535 : AOI222_X1 port map( A1 => n11188, A2 => n9391, B1 => n11185, B2 => 
                           n9327, C1 => n11182, C2 => n9359, ZN => n3608);
   U6536 : AOI222_X1 port map( A1 => n10924, A2 => n9392, B1 => n10921, B2 => 
                           n9328, C1 => n10918, C2 => n9360, ZN => n5000);
   U6537 : AOI222_X1 port map( A1 => n11188, A2 => n9392, B1 => n11185, B2 => 
                           n9328, C1 => n11182, C2 => n9360, ZN => n3567);
   U6538 : AOI222_X1 port map( A1 => n10924, A2 => n9393, B1 => n10921, B2 => 
                           n9329, C1 => n10918, C2 => n9361, ZN => n4959);
   U6539 : AOI222_X1 port map( A1 => n11188, A2 => n9393, B1 => n11185, B2 => 
                           n9329, C1 => n11182, C2 => n9361, ZN => n3526);
   U6540 : AOI222_X1 port map( A1 => n10924, A2 => n9394, B1 => n10921, B2 => 
                           n9330, C1 => n10918, C2 => n9362, ZN => n4918);
   U6541 : AOI222_X1 port map( A1 => n11188, A2 => n9394, B1 => n11185, B2 => 
                           n9330, C1 => n11182, C2 => n9362, ZN => n3485);
   U6542 : AOI222_X1 port map( A1 => n10924, A2 => n9395, B1 => n10921, B2 => 
                           n9331, C1 => n10918, C2 => n9363, ZN => n4877);
   U6543 : AOI222_X1 port map( A1 => n11188, A2 => n9395, B1 => n11185, B2 => 
                           n9331, C1 => n11182, C2 => n9363, ZN => n3444);
   U6544 : AOI222_X1 port map( A1 => n10924, A2 => n9396, B1 => n10921, B2 => 
                           n9332, C1 => n10918, C2 => n9364, ZN => n4836);
   U6545 : AOI222_X1 port map( A1 => n11188, A2 => n9396, B1 => n11185, B2 => 
                           n9332, C1 => n11182, C2 => n9364, ZN => n3403);
   U6546 : AOI222_X1 port map( A1 => n10924, A2 => n9397, B1 => n10921, B2 => 
                           n9333, C1 => n10918, C2 => n9365, ZN => n4795);
   U6547 : AOI222_X1 port map( A1 => n11188, A2 => n9397, B1 => n11185, B2 => 
                           n9333, C1 => n11182, C2 => n9365, ZN => n3362);
   U6548 : AOI222_X1 port map( A1 => n10924, A2 => n9398, B1 => n10921, B2 => 
                           n9334, C1 => n10918, C2 => n9366, ZN => n4754);
   U6549 : AOI222_X1 port map( A1 => n11188, A2 => n9398, B1 => n11185, B2 => 
                           n9334, C1 => n11182, C2 => n9366, ZN => n3321);
   U6550 : AOI222_X1 port map( A1 => n10924, A2 => n9399, B1 => n10921, B2 => 
                           n9335, C1 => n10918, C2 => n9367, ZN => n4713);
   U6551 : AOI222_X1 port map( A1 => n11188, A2 => n9399, B1 => n11185, B2 => 
                           n9335, C1 => n11182, C2 => n9367, ZN => n3280);
   U6552 : AOI222_X1 port map( A1 => n10925, A2 => n9400, B1 => n10922, B2 => 
                           n9336, C1 => n10919, C2 => n9368, ZN => n4672);
   U6553 : AOI222_X1 port map( A1 => n11189, A2 => n9400, B1 => n11186, B2 => 
                           n9336, C1 => n11183, C2 => n9368, ZN => n3239);
   U6554 : AOI222_X1 port map( A1 => n10925, A2 => n9401, B1 => n10922, B2 => 
                           n9337, C1 => n10919, C2 => n9369, ZN => n4631);
   U6555 : AOI222_X1 port map( A1 => n11189, A2 => n9401, B1 => n11186, B2 => 
                           n9337, C1 => n11183, C2 => n9369, ZN => n3198);
   U6556 : AOI222_X1 port map( A1 => n10925, A2 => n9402, B1 => n10922, B2 => 
                           n9338, C1 => n10919, C2 => n9370, ZN => n4590);
   U6557 : AOI222_X1 port map( A1 => n11189, A2 => n9402, B1 => n11186, B2 => 
                           n9338, C1 => n11183, C2 => n9370, ZN => n3157);
   U6558 : AOI222_X1 port map( A1 => n10925, A2 => n9403, B1 => n10922, B2 => 
                           n9339, C1 => n10919, C2 => n9371, ZN => n4549);
   U6559 : AOI222_X1 port map( A1 => n11189, A2 => n9403, B1 => n11186, B2 => 
                           n9339, C1 => n11183, C2 => n9371, ZN => n3116);
   U6560 : AOI222_X1 port map( A1 => n10925, A2 => n9404, B1 => n10922, B2 => 
                           n9340, C1 => n10919, C2 => n9372, ZN => n4508);
   U6561 : AOI222_X1 port map( A1 => n11189, A2 => n9404, B1 => n11186, B2 => 
                           n9340, C1 => n11183, C2 => n9372, ZN => n3075);
   U6562 : AOI222_X1 port map( A1 => n10925, A2 => n9405, B1 => n10922, B2 => 
                           n9341, C1 => n10919, C2 => n9373, ZN => n4467);
   U6563 : AOI222_X1 port map( A1 => n11189, A2 => n9405, B1 => n11186, B2 => 
                           n9341, C1 => n11183, C2 => n9373, ZN => n3034);
   U6564 : AOI222_X1 port map( A1 => n10925, A2 => n9406, B1 => n10922, B2 => 
                           n9342, C1 => n10919, C2 => n9374, ZN => n4426);
   U6565 : AOI222_X1 port map( A1 => n11189, A2 => n9406, B1 => n11186, B2 => 
                           n9342, C1 => n11183, C2 => n9374, ZN => n2993);
   U6566 : AOI222_X1 port map( A1 => n10925, A2 => n9407, B1 => n10922, B2 => 
                           n9343, C1 => n10919, C2 => n9375, ZN => n4341);
   U6567 : AOI222_X1 port map( A1 => n11189, A2 => n9407, B1 => n11186, B2 => 
                           n9343, C1 => n11183, C2 => n9375, ZN => n2873);
   U6568 : NOR4_X1 port map( A1 => n5683, A2 => n5684, A3 => n5685, A4 => n5686
                           , ZN => n5682);
   U6569 : OAI22_X1 port map( A1 => n10521, A2 => n10980, B1 => n10520, B2 => 
                           n10977, ZN => n5686);
   U6570 : OAI222_X1 port map( A1 => n13939, A2 => n10956, B1 => n13875, B2 => 
                           n10953, C1 => n13907, C2 => n10950, ZN => n5683);
   U6571 : OAI222_X1 port map( A1 => n10515, A2 => n10965, B1 => n10514, B2 => 
                           n10962, C1 => n10516, C2 => n10959, ZN => n5684);
   U6572 : NOR4_X1 port map( A1 => n5697, A2 => n5698, A3 => n5699, A4 => n5700
                           , ZN => n5696);
   U6573 : OAI22_X1 port map( A1 => n13971, A2 => n10914, B1 => n14003, B2 => 
                           n10911, ZN => n5700);
   U6574 : OAI222_X1 port map( A1 => n992, A2 => n10890, B1 => n14256, B2 => 
                           n10887, C1 => n14224, C2 => n10884, ZN => n5697);
   U6575 : OAI222_X1 port map( A1 => n14161, A2 => n10899, B1 => n14193, B2 => 
                           n10896, C1 => n14129, C2 => n10893, ZN => n5698);
   U6576 : NOR4_X1 port map( A1 => n4250, A2 => n4251, A3 => n4252, A4 => n4253
                           , ZN => n4249);
   U6577 : OAI22_X1 port map( A1 => n10521, A2 => n11244, B1 => n10520, B2 => 
                           n11241, ZN => n4253);
   U6578 : OAI222_X1 port map( A1 => n13939, A2 => n11220, B1 => n13875, B2 => 
                           n11217, C1 => n13907, C2 => n11214, ZN => n4250);
   U6579 : OAI222_X1 port map( A1 => n10515, A2 => n11229, B1 => n10514, B2 => 
                           n11226, C1 => n10516, C2 => n11223, ZN => n4251);
   U6580 : NOR4_X1 port map( A1 => n4264, A2 => n4265, A3 => n4266, A4 => n4267
                           , ZN => n4263);
   U6581 : OAI22_X1 port map( A1 => n13971, A2 => n11178, B1 => n14003, B2 => 
                           n11175, ZN => n4267);
   U6582 : OAI222_X1 port map( A1 => n992, A2 => n11154, B1 => n14256, B2 => 
                           n11151, C1 => n14224, C2 => n11148, ZN => n4264);
   U6583 : OAI222_X1 port map( A1 => n14161, A2 => n11163, B1 => n14193, B2 => 
                           n11160, C1 => n14129, C2 => n11157, ZN => n4265);
   U6584 : NOR4_X1 port map( A1 => n5619, A2 => n5620, A3 => n5621, A4 => n5622
                           , ZN => n5618);
   U6585 : OAI22_X1 port map( A1 => n10489, A2 => n10980, B1 => n10488, B2 => 
                           n10977, ZN => n5622);
   U6586 : OAI222_X1 port map( A1 => n13938, A2 => n10956, B1 => n13874, B2 => 
                           n10953, C1 => n13906, C2 => n10950, ZN => n5619);
   U6587 : OAI222_X1 port map( A1 => n10483, A2 => n10965, B1 => n10482, B2 => 
                           n10962, C1 => n10484, C2 => n10959, ZN => n5620);
   U6588 : NOR4_X1 port map( A1 => n5628, A2 => n5629, A3 => n5630, A4 => n5631
                           , ZN => n5627);
   U6589 : OAI22_X1 port map( A1 => n13970, A2 => n10914, B1 => n14002, B2 => 
                           n10911, ZN => n5631);
   U6590 : OAI222_X1 port map( A1 => n988, A2 => n10890, B1 => n14255, B2 => 
                           n10887, C1 => n14223, C2 => n10884, ZN => n5628);
   U6591 : OAI222_X1 port map( A1 => n14160, A2 => n10899, B1 => n14192, B2 => 
                           n10896, C1 => n14128, C2 => n10893, ZN => n5629);
   U6592 : NOR4_X1 port map( A1 => n4186, A2 => n4187, A3 => n4188, A4 => n4189
                           , ZN => n4185);
   U6593 : OAI22_X1 port map( A1 => n10489, A2 => n11244, B1 => n10488, B2 => 
                           n11241, ZN => n4189);
   U6594 : OAI222_X1 port map( A1 => n13938, A2 => n11220, B1 => n13874, B2 => 
                           n11217, C1 => n13906, C2 => n11214, ZN => n4186);
   U6595 : OAI222_X1 port map( A1 => n10483, A2 => n11229, B1 => n10482, B2 => 
                           n11226, C1 => n10484, C2 => n11223, ZN => n4187);
   U6596 : NOR4_X1 port map( A1 => n4195, A2 => n4196, A3 => n4197, A4 => n4198
                           , ZN => n4194);
   U6597 : OAI22_X1 port map( A1 => n13970, A2 => n11178, B1 => n14002, B2 => 
                           n11175, ZN => n4198);
   U6598 : OAI222_X1 port map( A1 => n988, A2 => n11154, B1 => n14255, B2 => 
                           n11151, C1 => n14223, C2 => n11148, ZN => n4195);
   U6599 : OAI222_X1 port map( A1 => n14160, A2 => n11163, B1 => n14192, B2 => 
                           n11160, C1 => n14128, C2 => n11157, ZN => n4196);
   U6600 : NOR4_X1 port map( A1 => n5578, A2 => n5579, A3 => n5580, A4 => n5581
                           , ZN => n5577);
   U6601 : OAI22_X1 port map( A1 => n10457, A2 => n10980, B1 => n10456, B2 => 
                           n10977, ZN => n5581);
   U6602 : OAI222_X1 port map( A1 => n13937, A2 => n10956, B1 => n13873, B2 => 
                           n10953, C1 => n13905, C2 => n10950, ZN => n5578);
   U6603 : OAI222_X1 port map( A1 => n10451, A2 => n10965, B1 => n10450, B2 => 
                           n10962, C1 => n10452, C2 => n10959, ZN => n5579);
   U6604 : NOR4_X1 port map( A1 => n5587, A2 => n5588, A3 => n5589, A4 => n5590
                           , ZN => n5586);
   U6605 : OAI22_X1 port map( A1 => n13969, A2 => n10914, B1 => n14001, B2 => 
                           n10911, ZN => n5590);
   U6606 : OAI222_X1 port map( A1 => n984, A2 => n10890, B1 => n14254, B2 => 
                           n10887, C1 => n14222, C2 => n10884, ZN => n5587);
   U6607 : OAI222_X1 port map( A1 => n14159, A2 => n10899, B1 => n14191, B2 => 
                           n10896, C1 => n14127, C2 => n10893, ZN => n5588);
   U6608 : NOR4_X1 port map( A1 => n4145, A2 => n4146, A3 => n4147, A4 => n4148
                           , ZN => n4144);
   U6609 : OAI22_X1 port map( A1 => n10457, A2 => n11244, B1 => n10456, B2 => 
                           n11241, ZN => n4148);
   U6610 : OAI222_X1 port map( A1 => n13937, A2 => n11220, B1 => n13873, B2 => 
                           n11217, C1 => n13905, C2 => n11214, ZN => n4145);
   U6611 : OAI222_X1 port map( A1 => n10451, A2 => n11229, B1 => n10450, B2 => 
                           n11226, C1 => n10452, C2 => n11223, ZN => n4146);
   U6612 : NOR4_X1 port map( A1 => n4154, A2 => n4155, A3 => n4156, A4 => n4157
                           , ZN => n4153);
   U6613 : OAI22_X1 port map( A1 => n13969, A2 => n11178, B1 => n14001, B2 => 
                           n11175, ZN => n4157);
   U6614 : OAI222_X1 port map( A1 => n984, A2 => n11154, B1 => n14254, B2 => 
                           n11151, C1 => n14222, C2 => n11148, ZN => n4154);
   U6615 : OAI222_X1 port map( A1 => n14159, A2 => n11163, B1 => n14191, B2 => 
                           n11160, C1 => n14127, C2 => n11157, ZN => n4155);
   U6616 : NOR4_X1 port map( A1 => n5537, A2 => n5538, A3 => n5539, A4 => n5540
                           , ZN => n5536);
   U6617 : OAI22_X1 port map( A1 => n10425, A2 => n10980, B1 => n10424, B2 => 
                           n10977, ZN => n5540);
   U6618 : OAI222_X1 port map( A1 => n13936, A2 => n10956, B1 => n13872, B2 => 
                           n10953, C1 => n13904, C2 => n10950, ZN => n5537);
   U6619 : OAI222_X1 port map( A1 => n10419, A2 => n10965, B1 => n10418, B2 => 
                           n10962, C1 => n10420, C2 => n10959, ZN => n5538);
   U6620 : NOR4_X1 port map( A1 => n5546, A2 => n5547, A3 => n5548, A4 => n5549
                           , ZN => n5545);
   U6621 : OAI22_X1 port map( A1 => n13968, A2 => n10914, B1 => n14000, B2 => 
                           n10911, ZN => n5549);
   U6622 : OAI222_X1 port map( A1 => n980, A2 => n10890, B1 => n14253, B2 => 
                           n10887, C1 => n14221, C2 => n10884, ZN => n5546);
   U6623 : OAI222_X1 port map( A1 => n14158, A2 => n10899, B1 => n14190, B2 => 
                           n10896, C1 => n14126, C2 => n10893, ZN => n5547);
   U6624 : NOR4_X1 port map( A1 => n4104, A2 => n4105, A3 => n4106, A4 => n4107
                           , ZN => n4103);
   U6625 : OAI22_X1 port map( A1 => n10425, A2 => n11244, B1 => n10424, B2 => 
                           n11241, ZN => n4107);
   U6626 : OAI222_X1 port map( A1 => n13936, A2 => n11220, B1 => n13872, B2 => 
                           n11217, C1 => n13904, C2 => n11214, ZN => n4104);
   U6627 : OAI222_X1 port map( A1 => n10419, A2 => n11229, B1 => n10418, B2 => 
                           n11226, C1 => n10420, C2 => n11223, ZN => n4105);
   U6628 : NOR4_X1 port map( A1 => n4113, A2 => n4114, A3 => n4115, A4 => n4116
                           , ZN => n4112);
   U6629 : OAI22_X1 port map( A1 => n13968, A2 => n11178, B1 => n14000, B2 => 
                           n11175, ZN => n4116);
   U6630 : OAI222_X1 port map( A1 => n980, A2 => n11154, B1 => n14253, B2 => 
                           n11151, C1 => n14221, C2 => n11148, ZN => n4113);
   U6631 : OAI222_X1 port map( A1 => n14158, A2 => n11163, B1 => n14190, B2 => 
                           n11160, C1 => n14126, C2 => n11157, ZN => n4114);
   U6632 : NOR4_X1 port map( A1 => n5496, A2 => n5497, A3 => n5498, A4 => n5499
                           , ZN => n5495);
   U6633 : OAI22_X1 port map( A1 => n10390, A2 => n10980, B1 => n10389, B2 => 
                           n10977, ZN => n5499);
   U6634 : OAI222_X1 port map( A1 => n13935, A2 => n10956, B1 => n13871, B2 => 
                           n10953, C1 => n13903, C2 => n10950, ZN => n5496);
   U6635 : OAI222_X1 port map( A1 => n10384, A2 => n10965, B1 => n10383, B2 => 
                           n10962, C1 => n10385, C2 => n10959, ZN => n5497);
   U6636 : NOR4_X1 port map( A1 => n5505, A2 => n5506, A3 => n5507, A4 => n5508
                           , ZN => n5504);
   U6637 : OAI22_X1 port map( A1 => n13967, A2 => n10914, B1 => n13999, B2 => 
                           n10911, ZN => n5508);
   U6638 : OAI222_X1 port map( A1 => n976, A2 => n10890, B1 => n14252, B2 => 
                           n10887, C1 => n14220, C2 => n10884, ZN => n5505);
   U6639 : OAI222_X1 port map( A1 => n14157, A2 => n10899, B1 => n14189, B2 => 
                           n10896, C1 => n14125, C2 => n10893, ZN => n5506);
   U6640 : NOR4_X1 port map( A1 => n4063, A2 => n4064, A3 => n4065, A4 => n4066
                           , ZN => n4062);
   U6641 : OAI22_X1 port map( A1 => n10390, A2 => n11244, B1 => n10389, B2 => 
                           n11241, ZN => n4066);
   U6642 : OAI222_X1 port map( A1 => n13935, A2 => n11220, B1 => n13871, B2 => 
                           n11217, C1 => n13903, C2 => n11214, ZN => n4063);
   U6643 : OAI222_X1 port map( A1 => n10384, A2 => n11229, B1 => n10383, B2 => 
                           n11226, C1 => n10385, C2 => n11223, ZN => n4064);
   U6644 : NOR4_X1 port map( A1 => n4072, A2 => n4073, A3 => n4074, A4 => n4075
                           , ZN => n4071);
   U6645 : OAI22_X1 port map( A1 => n13967, A2 => n11178, B1 => n13999, B2 => 
                           n11175, ZN => n4075);
   U6646 : OAI222_X1 port map( A1 => n976, A2 => n11154, B1 => n14252, B2 => 
                           n11151, C1 => n14220, C2 => n11148, ZN => n4072);
   U6647 : OAI222_X1 port map( A1 => n14157, A2 => n11163, B1 => n14189, B2 => 
                           n11160, C1 => n14125, C2 => n11157, ZN => n4073);
   U6648 : NOR4_X1 port map( A1 => n5455, A2 => n5456, A3 => n5457, A4 => n5458
                           , ZN => n5454);
   U6649 : OAI22_X1 port map( A1 => n10358, A2 => n10980, B1 => n10357, B2 => 
                           n10977, ZN => n5458);
   U6650 : OAI222_X1 port map( A1 => n13934, A2 => n10956, B1 => n13870, B2 => 
                           n10953, C1 => n13902, C2 => n10950, ZN => n5455);
   U6651 : OAI222_X1 port map( A1 => n10352, A2 => n10965, B1 => n10351, B2 => 
                           n10962, C1 => n10353, C2 => n10959, ZN => n5456);
   U6652 : NOR4_X1 port map( A1 => n5464, A2 => n5465, A3 => n5466, A4 => n5467
                           , ZN => n5463);
   U6653 : OAI22_X1 port map( A1 => n13966, A2 => n10914, B1 => n13998, B2 => 
                           n10911, ZN => n5467);
   U6654 : OAI222_X1 port map( A1 => n972, A2 => n10890, B1 => n14251, B2 => 
                           n10887, C1 => n14219, C2 => n10884, ZN => n5464);
   U6655 : OAI222_X1 port map( A1 => n14156, A2 => n10899, B1 => n14188, B2 => 
                           n10896, C1 => n14124, C2 => n10893, ZN => n5465);
   U6656 : NOR4_X1 port map( A1 => n4022, A2 => n4023, A3 => n4024, A4 => n4025
                           , ZN => n4021);
   U6657 : OAI22_X1 port map( A1 => n10358, A2 => n11244, B1 => n10357, B2 => 
                           n11241, ZN => n4025);
   U6658 : OAI222_X1 port map( A1 => n13934, A2 => n11220, B1 => n13870, B2 => 
                           n11217, C1 => n13902, C2 => n11214, ZN => n4022);
   U6659 : OAI222_X1 port map( A1 => n10352, A2 => n11229, B1 => n10351, B2 => 
                           n11226, C1 => n10353, C2 => n11223, ZN => n4023);
   U6660 : NOR4_X1 port map( A1 => n4031, A2 => n4032, A3 => n4033, A4 => n4034
                           , ZN => n4030);
   U6661 : OAI22_X1 port map( A1 => n13966, A2 => n11178, B1 => n13998, B2 => 
                           n11175, ZN => n4034);
   U6662 : OAI222_X1 port map( A1 => n972, A2 => n11154, B1 => n14251, B2 => 
                           n11151, C1 => n14219, C2 => n11148, ZN => n4031);
   U6663 : OAI222_X1 port map( A1 => n14156, A2 => n11163, B1 => n14188, B2 => 
                           n11160, C1 => n14124, C2 => n11157, ZN => n4032);
   U6664 : NOR4_X1 port map( A1 => n5414, A2 => n5415, A3 => n5416, A4 => n5417
                           , ZN => n5413);
   U6665 : OAI22_X1 port map( A1 => n10326, A2 => n10980, B1 => n10325, B2 => 
                           n10977, ZN => n5417);
   U6666 : OAI222_X1 port map( A1 => n13933, A2 => n10956, B1 => n13869, B2 => 
                           n10953, C1 => n13901, C2 => n10950, ZN => n5414);
   U6667 : OAI222_X1 port map( A1 => n10320, A2 => n10965, B1 => n10319, B2 => 
                           n10962, C1 => n10321, C2 => n10959, ZN => n5415);
   U6668 : NOR4_X1 port map( A1 => n5423, A2 => n5424, A3 => n5425, A4 => n5426
                           , ZN => n5422);
   U6669 : OAI22_X1 port map( A1 => n13965, A2 => n10914, B1 => n13997, B2 => 
                           n10911, ZN => n5426);
   U6670 : OAI222_X1 port map( A1 => n968, A2 => n10890, B1 => n14250, B2 => 
                           n10887, C1 => n14218, C2 => n10884, ZN => n5423);
   U6671 : OAI222_X1 port map( A1 => n14155, A2 => n10899, B1 => n14187, B2 => 
                           n10896, C1 => n14123, C2 => n10893, ZN => n5424);
   U6672 : NOR4_X1 port map( A1 => n3981, A2 => n3982, A3 => n3983, A4 => n3984
                           , ZN => n3980);
   U6673 : OAI22_X1 port map( A1 => n10326, A2 => n11244, B1 => n10325, B2 => 
                           n11241, ZN => n3984);
   U6674 : OAI222_X1 port map( A1 => n13933, A2 => n11220, B1 => n13869, B2 => 
                           n11217, C1 => n13901, C2 => n11214, ZN => n3981);
   U6675 : OAI222_X1 port map( A1 => n10320, A2 => n11229, B1 => n10319, B2 => 
                           n11226, C1 => n10321, C2 => n11223, ZN => n3982);
   U6676 : NOR4_X1 port map( A1 => n3990, A2 => n3991, A3 => n3992, A4 => n3993
                           , ZN => n3989);
   U6677 : OAI22_X1 port map( A1 => n13965, A2 => n11178, B1 => n13997, B2 => 
                           n11175, ZN => n3993);
   U6678 : OAI222_X1 port map( A1 => n968, A2 => n11154, B1 => n14250, B2 => 
                           n11151, C1 => n14218, C2 => n11148, ZN => n3990);
   U6679 : OAI222_X1 port map( A1 => n14155, A2 => n11163, B1 => n14187, B2 => 
                           n11160, C1 => n14123, C2 => n11157, ZN => n3991);
   U6680 : NOR4_X1 port map( A1 => n5373, A2 => n5374, A3 => n5375, A4 => n5376
                           , ZN => n5372);
   U6681 : OAI22_X1 port map( A1 => n10291, A2 => n10980, B1 => n10290, B2 => 
                           n10977, ZN => n5376);
   U6682 : OAI222_X1 port map( A1 => n13932, A2 => n10956, B1 => n13868, B2 => 
                           n10953, C1 => n13900, C2 => n10950, ZN => n5373);
   U6683 : OAI222_X1 port map( A1 => n10285, A2 => n10965, B1 => n10284, B2 => 
                           n10962, C1 => n10286, C2 => n10959, ZN => n5374);
   U6684 : NOR4_X1 port map( A1 => n5382, A2 => n5383, A3 => n5384, A4 => n5385
                           , ZN => n5381);
   U6685 : OAI22_X1 port map( A1 => n13964, A2 => n10914, B1 => n13996, B2 => 
                           n10911, ZN => n5385);
   U6686 : OAI222_X1 port map( A1 => n964, A2 => n10890, B1 => n14249, B2 => 
                           n10887, C1 => n14217, C2 => n10884, ZN => n5382);
   U6687 : OAI222_X1 port map( A1 => n14154, A2 => n10899, B1 => n14186, B2 => 
                           n10896, C1 => n14122, C2 => n10893, ZN => n5383);
   U6688 : NOR4_X1 port map( A1 => n3940, A2 => n3941, A3 => n3942, A4 => n3943
                           , ZN => n3939);
   U6689 : OAI22_X1 port map( A1 => n10291, A2 => n11244, B1 => n10290, B2 => 
                           n11241, ZN => n3943);
   U6690 : OAI222_X1 port map( A1 => n13932, A2 => n11220, B1 => n13868, B2 => 
                           n11217, C1 => n13900, C2 => n11214, ZN => n3940);
   U6691 : OAI222_X1 port map( A1 => n10285, A2 => n11229, B1 => n10284, B2 => 
                           n11226, C1 => n10286, C2 => n11223, ZN => n3941);
   U6692 : NOR4_X1 port map( A1 => n3949, A2 => n3950, A3 => n3951, A4 => n3952
                           , ZN => n3948);
   U6693 : OAI22_X1 port map( A1 => n13964, A2 => n11178, B1 => n13996, B2 => 
                           n11175, ZN => n3952);
   U6694 : OAI222_X1 port map( A1 => n964, A2 => n11154, B1 => n14249, B2 => 
                           n11151, C1 => n14217, C2 => n11148, ZN => n3949);
   U6695 : OAI222_X1 port map( A1 => n14154, A2 => n11163, B1 => n14186, B2 => 
                           n11160, C1 => n14122, C2 => n11157, ZN => n3950);
   U6696 : NOR4_X1 port map( A1 => n5332, A2 => n5333, A3 => n5334, A4 => n5335
                           , ZN => n5331);
   U6697 : OAI22_X1 port map( A1 => n10259, A2 => n10980, B1 => n10258, B2 => 
                           n10977, ZN => n5335);
   U6698 : OAI222_X1 port map( A1 => n13931, A2 => n10956, B1 => n13867, B2 => 
                           n10953, C1 => n13899, C2 => n10950, ZN => n5332);
   U6699 : OAI222_X1 port map( A1 => n10253, A2 => n10965, B1 => n10252, B2 => 
                           n10962, C1 => n10254, C2 => n10959, ZN => n5333);
   U6700 : NOR4_X1 port map( A1 => n5341, A2 => n5342, A3 => n5343, A4 => n5344
                           , ZN => n5340);
   U6701 : OAI22_X1 port map( A1 => n13963, A2 => n10914, B1 => n13995, B2 => 
                           n10911, ZN => n5344);
   U6702 : OAI222_X1 port map( A1 => n960, A2 => n10890, B1 => n14248, B2 => 
                           n10887, C1 => n14216, C2 => n10884, ZN => n5341);
   U6703 : OAI222_X1 port map( A1 => n14153, A2 => n10899, B1 => n14185, B2 => 
                           n10896, C1 => n14121, C2 => n10893, ZN => n5342);
   U6704 : NOR4_X1 port map( A1 => n3899, A2 => n3900, A3 => n3901, A4 => n3902
                           , ZN => n3898);
   U6705 : OAI22_X1 port map( A1 => n10259, A2 => n11244, B1 => n10258, B2 => 
                           n11241, ZN => n3902);
   U6706 : OAI222_X1 port map( A1 => n13931, A2 => n11220, B1 => n13867, B2 => 
                           n11217, C1 => n13899, C2 => n11214, ZN => n3899);
   U6707 : OAI222_X1 port map( A1 => n10253, A2 => n11229, B1 => n10252, B2 => 
                           n11226, C1 => n10254, C2 => n11223, ZN => n3900);
   U6708 : NOR4_X1 port map( A1 => n3908, A2 => n3909, A3 => n3910, A4 => n3911
                           , ZN => n3907);
   U6709 : OAI22_X1 port map( A1 => n13963, A2 => n11178, B1 => n13995, B2 => 
                           n11175, ZN => n3911);
   U6710 : OAI222_X1 port map( A1 => n960, A2 => n11154, B1 => n14248, B2 => 
                           n11151, C1 => n14216, C2 => n11148, ZN => n3908);
   U6711 : OAI222_X1 port map( A1 => n14153, A2 => n11163, B1 => n14185, B2 => 
                           n11160, C1 => n14121, C2 => n11157, ZN => n3909);
   U6712 : NOR4_X1 port map( A1 => n5291, A2 => n5292, A3 => n5293, A4 => n5294
                           , ZN => n5290);
   U6713 : OAI22_X1 port map( A1 => n10227, A2 => n10980, B1 => n10226, B2 => 
                           n10977, ZN => n5294);
   U6714 : OAI222_X1 port map( A1 => n13930, A2 => n10956, B1 => n13866, B2 => 
                           n10953, C1 => n13898, C2 => n10950, ZN => n5291);
   U6715 : OAI222_X1 port map( A1 => n10221, A2 => n10965, B1 => n10220, B2 => 
                           n10962, C1 => n10222, C2 => n10959, ZN => n5292);
   U6716 : NOR4_X1 port map( A1 => n5300, A2 => n5301, A3 => n5302, A4 => n5303
                           , ZN => n5299);
   U6717 : OAI22_X1 port map( A1 => n13962, A2 => n10914, B1 => n13994, B2 => 
                           n10911, ZN => n5303);
   U6718 : OAI222_X1 port map( A1 => n956, A2 => n10890, B1 => n14247, B2 => 
                           n10887, C1 => n14215, C2 => n10884, ZN => n5300);
   U6719 : OAI222_X1 port map( A1 => n14152, A2 => n10899, B1 => n14184, B2 => 
                           n10896, C1 => n14120, C2 => n10893, ZN => n5301);
   U6720 : NOR4_X1 port map( A1 => n3858, A2 => n3859, A3 => n3860, A4 => n3861
                           , ZN => n3857);
   U6721 : OAI22_X1 port map( A1 => n10227, A2 => n11244, B1 => n10226, B2 => 
                           n11241, ZN => n3861);
   U6722 : OAI222_X1 port map( A1 => n13930, A2 => n11220, B1 => n13866, B2 => 
                           n11217, C1 => n13898, C2 => n11214, ZN => n3858);
   U6723 : OAI222_X1 port map( A1 => n10221, A2 => n11229, B1 => n10220, B2 => 
                           n11226, C1 => n10222, C2 => n11223, ZN => n3859);
   U6724 : NOR4_X1 port map( A1 => n3867, A2 => n3868, A3 => n3869, A4 => n3870
                           , ZN => n3866);
   U6725 : OAI22_X1 port map( A1 => n13962, A2 => n11178, B1 => n13994, B2 => 
                           n11175, ZN => n3870);
   U6726 : OAI222_X1 port map( A1 => n956, A2 => n11154, B1 => n14247, B2 => 
                           n11151, C1 => n14215, C2 => n11148, ZN => n3867);
   U6727 : OAI222_X1 port map( A1 => n14152, A2 => n11163, B1 => n14184, B2 => 
                           n11160, C1 => n14120, C2 => n11157, ZN => n3868);
   U6728 : NOR4_X1 port map( A1 => n5250, A2 => n5251, A3 => n5252, A4 => n5253
                           , ZN => n5249);
   U6729 : OAI22_X1 port map( A1 => n10193, A2 => n10980, B1 => n10192, B2 => 
                           n10977, ZN => n5253);
   U6730 : OAI222_X1 port map( A1 => n13929, A2 => n10956, B1 => n13865, B2 => 
                           n10953, C1 => n13897, C2 => n10950, ZN => n5250);
   U6731 : OAI222_X1 port map( A1 => n10187, A2 => n10965, B1 => n10186, B2 => 
                           n10962, C1 => n10188, C2 => n10959, ZN => n5251);
   U6732 : NOR4_X1 port map( A1 => n5259, A2 => n5260, A3 => n5261, A4 => n5262
                           , ZN => n5258);
   U6733 : OAI22_X1 port map( A1 => n13961, A2 => n10914, B1 => n13993, B2 => 
                           n10911, ZN => n5262);
   U6734 : OAI222_X1 port map( A1 => n952, A2 => n10890, B1 => n14246, B2 => 
                           n10887, C1 => n14214, C2 => n10884, ZN => n5259);
   U6735 : OAI222_X1 port map( A1 => n14151, A2 => n10899, B1 => n14183, B2 => 
                           n10896, C1 => n14119, C2 => n10893, ZN => n5260);
   U6736 : NOR4_X1 port map( A1 => n3817, A2 => n3818, A3 => n3819, A4 => n3820
                           , ZN => n3816);
   U6737 : OAI22_X1 port map( A1 => n10193, A2 => n11244, B1 => n10192, B2 => 
                           n11241, ZN => n3820);
   U6738 : OAI222_X1 port map( A1 => n13929, A2 => n11220, B1 => n13865, B2 => 
                           n11217, C1 => n13897, C2 => n11214, ZN => n3817);
   U6739 : OAI222_X1 port map( A1 => n10187, A2 => n11229, B1 => n10186, B2 => 
                           n11226, C1 => n10188, C2 => n11223, ZN => n3818);
   U6740 : NOR4_X1 port map( A1 => n3826, A2 => n3827, A3 => n3828, A4 => n3829
                           , ZN => n3825);
   U6741 : OAI22_X1 port map( A1 => n13961, A2 => n11178, B1 => n13993, B2 => 
                           n11175, ZN => n3829);
   U6742 : OAI222_X1 port map( A1 => n952, A2 => n11154, B1 => n14246, B2 => 
                           n11151, C1 => n14214, C2 => n11148, ZN => n3826);
   U6743 : OAI222_X1 port map( A1 => n14151, A2 => n11163, B1 => n14183, B2 => 
                           n11160, C1 => n14119, C2 => n11157, ZN => n3827);
   U6744 : NOR4_X1 port map( A1 => n5209, A2 => n5210, A3 => n5211, A4 => n5212
                           , ZN => n5208);
   U6745 : OAI22_X1 port map( A1 => n10161, A2 => n10980, B1 => n10160, B2 => 
                           n10977, ZN => n5212);
   U6746 : OAI222_X1 port map( A1 => n13928, A2 => n10956, B1 => n13864, B2 => 
                           n10953, C1 => n13896, C2 => n10950, ZN => n5209);
   U6747 : OAI222_X1 port map( A1 => n10155, A2 => n10965, B1 => n10154, B2 => 
                           n10962, C1 => n10156, C2 => n10959, ZN => n5210);
   U6748 : NOR4_X1 port map( A1 => n5218, A2 => n5219, A3 => n5220, A4 => n5221
                           , ZN => n5217);
   U6749 : OAI22_X1 port map( A1 => n13960, A2 => n10914, B1 => n13992, B2 => 
                           n10911, ZN => n5221);
   U6750 : OAI222_X1 port map( A1 => n948, A2 => n10890, B1 => n14245, B2 => 
                           n10887, C1 => n14213, C2 => n10884, ZN => n5218);
   U6751 : OAI222_X1 port map( A1 => n14150, A2 => n10899, B1 => n14182, B2 => 
                           n10896, C1 => n14118, C2 => n10893, ZN => n5219);
   U6752 : NOR4_X1 port map( A1 => n3776, A2 => n3777, A3 => n3778, A4 => n3779
                           , ZN => n3775);
   U6753 : OAI22_X1 port map( A1 => n10161, A2 => n11244, B1 => n10160, B2 => 
                           n11241, ZN => n3779);
   U6754 : OAI222_X1 port map( A1 => n13928, A2 => n11220, B1 => n13864, B2 => 
                           n11217, C1 => n13896, C2 => n11214, ZN => n3776);
   U6755 : OAI222_X1 port map( A1 => n10155, A2 => n11229, B1 => n10154, B2 => 
                           n11226, C1 => n10156, C2 => n11223, ZN => n3777);
   U6756 : NOR4_X1 port map( A1 => n3785, A2 => n3786, A3 => n3787, A4 => n3788
                           , ZN => n3784);
   U6757 : OAI22_X1 port map( A1 => n13960, A2 => n11178, B1 => n13992, B2 => 
                           n11175, ZN => n3788);
   U6758 : OAI222_X1 port map( A1 => n948, A2 => n11154, B1 => n14245, B2 => 
                           n11151, C1 => n14213, C2 => n11148, ZN => n3785);
   U6759 : OAI222_X1 port map( A1 => n14150, A2 => n11163, B1 => n14182, B2 => 
                           n11160, C1 => n14118, C2 => n11157, ZN => n3786);
   U6760 : NOR4_X1 port map( A1 => n5168, A2 => n5169, A3 => n5170, A4 => n5171
                           , ZN => n5167);
   U6761 : OAI22_X1 port map( A1 => n10129, A2 => n10981, B1 => n10128, B2 => 
                           n10978, ZN => n5171);
   U6762 : OAI222_X1 port map( A1 => n13927, A2 => n10957, B1 => n13863, B2 => 
                           n10954, C1 => n13895, C2 => n10951, ZN => n5168);
   U6763 : OAI222_X1 port map( A1 => n10123, A2 => n10966, B1 => n10122, B2 => 
                           n10963, C1 => n10124, C2 => n10960, ZN => n5169);
   U6764 : NOR4_X1 port map( A1 => n5177, A2 => n5178, A3 => n5179, A4 => n5180
                           , ZN => n5176);
   U6765 : OAI22_X1 port map( A1 => n13959, A2 => n10915, B1 => n13991, B2 => 
                           n10912, ZN => n5180);
   U6766 : OAI222_X1 port map( A1 => n944, A2 => n10891, B1 => n14244, B2 => 
                           n10888, C1 => n14212, C2 => n10885, ZN => n5177);
   U6767 : OAI222_X1 port map( A1 => n14149, A2 => n10900, B1 => n14181, B2 => 
                           n10897, C1 => n14117, C2 => n10894, ZN => n5178);
   U6768 : NOR4_X1 port map( A1 => n3735, A2 => n3736, A3 => n3737, A4 => n3738
                           , ZN => n3734);
   U6769 : OAI22_X1 port map( A1 => n10129, A2 => n11245, B1 => n10128, B2 => 
                           n11242, ZN => n3738);
   U6770 : OAI222_X1 port map( A1 => n13927, A2 => n11221, B1 => n13863, B2 => 
                           n11218, C1 => n13895, C2 => n11215, ZN => n3735);
   U6771 : OAI222_X1 port map( A1 => n10123, A2 => n11230, B1 => n10122, B2 => 
                           n11227, C1 => n10124, C2 => n11224, ZN => n3736);
   U6772 : NOR4_X1 port map( A1 => n3744, A2 => n3745, A3 => n3746, A4 => n3747
                           , ZN => n3743);
   U6773 : OAI22_X1 port map( A1 => n13959, A2 => n11179, B1 => n13991, B2 => 
                           n11176, ZN => n3747);
   U6774 : OAI222_X1 port map( A1 => n944, A2 => n11155, B1 => n14244, B2 => 
                           n11152, C1 => n14212, C2 => n11149, ZN => n3744);
   U6775 : OAI222_X1 port map( A1 => n14149, A2 => n11164, B1 => n14181, B2 => 
                           n11161, C1 => n14117, C2 => n11158, ZN => n3745);
   U6776 : NOR4_X1 port map( A1 => n5127, A2 => n5128, A3 => n5129, A4 => n5130
                           , ZN => n5126);
   U6777 : OAI22_X1 port map( A1 => n10097, A2 => n10981, B1 => n10096, B2 => 
                           n10978, ZN => n5130);
   U6778 : OAI222_X1 port map( A1 => n13926, A2 => n10957, B1 => n13862, B2 => 
                           n10954, C1 => n13894, C2 => n10951, ZN => n5127);
   U6779 : OAI222_X1 port map( A1 => n10091, A2 => n10966, B1 => n10090, B2 => 
                           n10963, C1 => n10092, C2 => n10960, ZN => n5128);
   U6780 : NOR4_X1 port map( A1 => n5136, A2 => n5137, A3 => n5138, A4 => n5139
                           , ZN => n5135);
   U6781 : OAI22_X1 port map( A1 => n13958, A2 => n10915, B1 => n13990, B2 => 
                           n10912, ZN => n5139);
   U6782 : OAI222_X1 port map( A1 => n940, A2 => n10891, B1 => n14243, B2 => 
                           n10888, C1 => n14211, C2 => n10885, ZN => n5136);
   U6783 : OAI222_X1 port map( A1 => n14148, A2 => n10900, B1 => n14180, B2 => 
                           n10897, C1 => n14116, C2 => n10894, ZN => n5137);
   U6784 : NOR4_X1 port map( A1 => n3694, A2 => n3695, A3 => n3696, A4 => n3697
                           , ZN => n3693);
   U6785 : OAI22_X1 port map( A1 => n10097, A2 => n11245, B1 => n10096, B2 => 
                           n11242, ZN => n3697);
   U6786 : OAI222_X1 port map( A1 => n13926, A2 => n11221, B1 => n13862, B2 => 
                           n11218, C1 => n13894, C2 => n11215, ZN => n3694);
   U6787 : OAI222_X1 port map( A1 => n10091, A2 => n11230, B1 => n10090, B2 => 
                           n11227, C1 => n10092, C2 => n11224, ZN => n3695);
   U6788 : NOR4_X1 port map( A1 => n3703, A2 => n3704, A3 => n3705, A4 => n3706
                           , ZN => n3702);
   U6789 : OAI22_X1 port map( A1 => n13958, A2 => n11179, B1 => n13990, B2 => 
                           n11176, ZN => n3706);
   U6790 : OAI222_X1 port map( A1 => n940, A2 => n11155, B1 => n14243, B2 => 
                           n11152, C1 => n14211, C2 => n11149, ZN => n3703);
   U6791 : OAI222_X1 port map( A1 => n14148, A2 => n11164, B1 => n14180, B2 => 
                           n11161, C1 => n14116, C2 => n11158, ZN => n3704);
   U6792 : NOR4_X1 port map( A1 => n5086, A2 => n5087, A3 => n5088, A4 => n5089
                           , ZN => n5085);
   U6793 : OAI22_X1 port map( A1 => n10065, A2 => n10981, B1 => n10064, B2 => 
                           n10978, ZN => n5089);
   U6794 : OAI222_X1 port map( A1 => n13925, A2 => n10957, B1 => n13861, B2 => 
                           n10954, C1 => n13893, C2 => n10951, ZN => n5086);
   U6795 : OAI222_X1 port map( A1 => n10059, A2 => n10966, B1 => n10058, B2 => 
                           n10963, C1 => n10060, C2 => n10960, ZN => n5087);
   U6796 : NOR4_X1 port map( A1 => n5095, A2 => n5096, A3 => n5097, A4 => n5098
                           , ZN => n5094);
   U6797 : OAI22_X1 port map( A1 => n13957, A2 => n10915, B1 => n13989, B2 => 
                           n10912, ZN => n5098);
   U6798 : OAI222_X1 port map( A1 => n936, A2 => n10891, B1 => n14242, B2 => 
                           n10888, C1 => n14210, C2 => n10885, ZN => n5095);
   U6799 : OAI222_X1 port map( A1 => n14147, A2 => n10900, B1 => n14179, B2 => 
                           n10897, C1 => n14115, C2 => n10894, ZN => n5096);
   U6800 : NOR4_X1 port map( A1 => n3653, A2 => n3654, A3 => n3655, A4 => n3656
                           , ZN => n3652);
   U6801 : OAI22_X1 port map( A1 => n10065, A2 => n11245, B1 => n10064, B2 => 
                           n11242, ZN => n3656);
   U6802 : OAI222_X1 port map( A1 => n13925, A2 => n11221, B1 => n13861, B2 => 
                           n11218, C1 => n13893, C2 => n11215, ZN => n3653);
   U6803 : OAI222_X1 port map( A1 => n10059, A2 => n11230, B1 => n10058, B2 => 
                           n11227, C1 => n10060, C2 => n11224, ZN => n3654);
   U6804 : NOR4_X1 port map( A1 => n3662, A2 => n3663, A3 => n3664, A4 => n3665
                           , ZN => n3661);
   U6805 : OAI22_X1 port map( A1 => n13957, A2 => n11179, B1 => n13989, B2 => 
                           n11176, ZN => n3665);
   U6806 : OAI222_X1 port map( A1 => n936, A2 => n11155, B1 => n14242, B2 => 
                           n11152, C1 => n14210, C2 => n11149, ZN => n3662);
   U6807 : OAI222_X1 port map( A1 => n14147, A2 => n11164, B1 => n14179, B2 => 
                           n11161, C1 => n14115, C2 => n11158, ZN => n3663);
   U6808 : NOR4_X1 port map( A1 => n5045, A2 => n5046, A3 => n5047, A4 => n5048
                           , ZN => n5044);
   U6809 : OAI22_X1 port map( A1 => n10033, A2 => n10981, B1 => n10032, B2 => 
                           n10978, ZN => n5048);
   U6810 : OAI222_X1 port map( A1 => n13924, A2 => n10957, B1 => n13860, B2 => 
                           n10954, C1 => n13892, C2 => n10951, ZN => n5045);
   U6811 : OAI222_X1 port map( A1 => n10027, A2 => n10966, B1 => n10026, B2 => 
                           n10963, C1 => n10028, C2 => n10960, ZN => n5046);
   U6812 : NOR4_X1 port map( A1 => n5054, A2 => n5055, A3 => n5056, A4 => n5057
                           , ZN => n5053);
   U6813 : OAI22_X1 port map( A1 => n13956, A2 => n10915, B1 => n13988, B2 => 
                           n10912, ZN => n5057);
   U6814 : OAI222_X1 port map( A1 => n932, A2 => n10891, B1 => n14241, B2 => 
                           n10888, C1 => n14209, C2 => n10885, ZN => n5054);
   U6815 : OAI222_X1 port map( A1 => n14146, A2 => n10900, B1 => n14178, B2 => 
                           n10897, C1 => n14114, C2 => n10894, ZN => n5055);
   U6816 : NOR4_X1 port map( A1 => n3612, A2 => n3613, A3 => n3614, A4 => n3615
                           , ZN => n3611);
   U6817 : OAI22_X1 port map( A1 => n10033, A2 => n11245, B1 => n10032, B2 => 
                           n11242, ZN => n3615);
   U6818 : OAI222_X1 port map( A1 => n13924, A2 => n11221, B1 => n13860, B2 => 
                           n11218, C1 => n13892, C2 => n11215, ZN => n3612);
   U6819 : OAI222_X1 port map( A1 => n10027, A2 => n11230, B1 => n10026, B2 => 
                           n11227, C1 => n10028, C2 => n11224, ZN => n3613);
   U6820 : NOR4_X1 port map( A1 => n3621, A2 => n3622, A3 => n3623, A4 => n3624
                           , ZN => n3620);
   U6821 : OAI22_X1 port map( A1 => n13956, A2 => n11179, B1 => n13988, B2 => 
                           n11176, ZN => n3624);
   U6822 : OAI222_X1 port map( A1 => n932, A2 => n11155, B1 => n14241, B2 => 
                           n11152, C1 => n14209, C2 => n11149, ZN => n3621);
   U6823 : OAI222_X1 port map( A1 => n14146, A2 => n11164, B1 => n14178, B2 => 
                           n11161, C1 => n14114, C2 => n11158, ZN => n3622);
   U6824 : NOR4_X1 port map( A1 => n5004, A2 => n5005, A3 => n5006, A4 => n5007
                           , ZN => n5003);
   U6825 : OAI22_X1 port map( A1 => n10001, A2 => n10981, B1 => n10000, B2 => 
                           n10978, ZN => n5007);
   U6826 : OAI222_X1 port map( A1 => n13923, A2 => n10957, B1 => n13859, B2 => 
                           n10954, C1 => n13891, C2 => n10951, ZN => n5004);
   U6827 : OAI222_X1 port map( A1 => n9697, A2 => n10966, B1 => n9696, B2 => 
                           n10963, C1 => n9698, C2 => n10960, ZN => n5005);
   U6828 : NOR4_X1 port map( A1 => n5013, A2 => n5014, A3 => n5015, A4 => n5016
                           , ZN => n5012);
   U6829 : OAI22_X1 port map( A1 => n13955, A2 => n10915, B1 => n13987, B2 => 
                           n10912, ZN => n5016);
   U6830 : OAI222_X1 port map( A1 => n928, A2 => n10891, B1 => n14240, B2 => 
                           n10888, C1 => n14208, C2 => n10885, ZN => n5013);
   U6831 : OAI222_X1 port map( A1 => n14145, A2 => n10900, B1 => n14177, B2 => 
                           n10897, C1 => n14113, C2 => n10894, ZN => n5014);
   U6832 : NOR4_X1 port map( A1 => n3571, A2 => n3572, A3 => n3573, A4 => n3574
                           , ZN => n3570);
   U6833 : OAI22_X1 port map( A1 => n10001, A2 => n11245, B1 => n10000, B2 => 
                           n11242, ZN => n3574);
   U6834 : OAI222_X1 port map( A1 => n13923, A2 => n11221, B1 => n13859, B2 => 
                           n11218, C1 => n13891, C2 => n11215, ZN => n3571);
   U6835 : OAI222_X1 port map( A1 => n9697, A2 => n11230, B1 => n9696, B2 => 
                           n11227, C1 => n9698, C2 => n11224, ZN => n3572);
   U6836 : NOR4_X1 port map( A1 => n3580, A2 => n3581, A3 => n3582, A4 => n3583
                           , ZN => n3579);
   U6837 : OAI22_X1 port map( A1 => n13955, A2 => n11179, B1 => n13987, B2 => 
                           n11176, ZN => n3583);
   U6838 : OAI222_X1 port map( A1 => n928, A2 => n11155, B1 => n14240, B2 => 
                           n11152, C1 => n14208, C2 => n11149, ZN => n3580);
   U6839 : OAI222_X1 port map( A1 => n14145, A2 => n11164, B1 => n14177, B2 => 
                           n11161, C1 => n14113, C2 => n11158, ZN => n3581);
   U6840 : NOR4_X1 port map( A1 => n4963, A2 => n4964, A3 => n4965, A4 => n4966
                           , ZN => n4962);
   U6841 : OAI22_X1 port map( A1 => n9639, A2 => n10981, B1 => n9638, B2 => 
                           n10978, ZN => n4966);
   U6842 : OAI222_X1 port map( A1 => n13922, A2 => n10957, B1 => n13858, B2 => 
                           n10954, C1 => n13890, C2 => n10951, ZN => n4963);
   U6843 : OAI222_X1 port map( A1 => n9633, A2 => n10966, B1 => n9632, B2 => 
                           n10963, C1 => n9634, C2 => n10960, ZN => n4964);
   U6844 : NOR4_X1 port map( A1 => n4972, A2 => n4973, A3 => n4974, A4 => n4975
                           , ZN => n4971);
   U6845 : OAI22_X1 port map( A1 => n13954, A2 => n10915, B1 => n13986, B2 => 
                           n10912, ZN => n4975);
   U6846 : OAI222_X1 port map( A1 => n924, A2 => n10891, B1 => n14239, B2 => 
                           n10888, C1 => n14207, C2 => n10885, ZN => n4972);
   U6847 : OAI222_X1 port map( A1 => n14144, A2 => n10900, B1 => n14176, B2 => 
                           n10897, C1 => n14112, C2 => n10894, ZN => n4973);
   U6848 : NOR4_X1 port map( A1 => n3530, A2 => n3531, A3 => n3532, A4 => n3533
                           , ZN => n3529);
   U6849 : OAI22_X1 port map( A1 => n9639, A2 => n11245, B1 => n9638, B2 => 
                           n11242, ZN => n3533);
   U6850 : OAI222_X1 port map( A1 => n13922, A2 => n11221, B1 => n13858, B2 => 
                           n11218, C1 => n13890, C2 => n11215, ZN => n3530);
   U6851 : OAI222_X1 port map( A1 => n9633, A2 => n11230, B1 => n9632, B2 => 
                           n11227, C1 => n9634, C2 => n11224, ZN => n3531);
   U6852 : NOR4_X1 port map( A1 => n3539, A2 => n3540, A3 => n3541, A4 => n3542
                           , ZN => n3538);
   U6853 : OAI22_X1 port map( A1 => n13954, A2 => n11179, B1 => n13986, B2 => 
                           n11176, ZN => n3542);
   U6854 : OAI222_X1 port map( A1 => n924, A2 => n11155, B1 => n14239, B2 => 
                           n11152, C1 => n14207, C2 => n11149, ZN => n3539);
   U6855 : OAI222_X1 port map( A1 => n14144, A2 => n11164, B1 => n14176, B2 => 
                           n11161, C1 => n14112, C2 => n11158, ZN => n3540);
   U6856 : NOR4_X1 port map( A1 => n4922, A2 => n4923, A3 => n4924, A4 => n4925
                           , ZN => n4921);
   U6857 : OAI22_X1 port map( A1 => n9607, A2 => n10981, B1 => n9606, B2 => 
                           n10978, ZN => n4925);
   U6858 : OAI222_X1 port map( A1 => n13921, A2 => n10957, B1 => n13857, B2 => 
                           n10954, C1 => n13889, C2 => n10951, ZN => n4922);
   U6859 : OAI222_X1 port map( A1 => n9601, A2 => n10966, B1 => n9600, B2 => 
                           n10963, C1 => n9602, C2 => n10960, ZN => n4923);
   U6860 : NOR4_X1 port map( A1 => n4931, A2 => n4932, A3 => n4933, A4 => n4934
                           , ZN => n4930);
   U6861 : OAI22_X1 port map( A1 => n13953, A2 => n10915, B1 => n13985, B2 => 
                           n10912, ZN => n4934);
   U6862 : OAI222_X1 port map( A1 => n920, A2 => n10891, B1 => n14238, B2 => 
                           n10888, C1 => n14206, C2 => n10885, ZN => n4931);
   U6863 : OAI222_X1 port map( A1 => n14143, A2 => n10900, B1 => n14175, B2 => 
                           n10897, C1 => n14111, C2 => n10894, ZN => n4932);
   U6864 : NOR4_X1 port map( A1 => n3489, A2 => n3490, A3 => n3491, A4 => n3492
                           , ZN => n3488);
   U6865 : OAI22_X1 port map( A1 => n9607, A2 => n11245, B1 => n9606, B2 => 
                           n11242, ZN => n3492);
   U6866 : OAI222_X1 port map( A1 => n13921, A2 => n11221, B1 => n13857, B2 => 
                           n11218, C1 => n13889, C2 => n11215, ZN => n3489);
   U6867 : OAI222_X1 port map( A1 => n9601, A2 => n11230, B1 => n9600, B2 => 
                           n11227, C1 => n9602, C2 => n11224, ZN => n3490);
   U6868 : NOR4_X1 port map( A1 => n3498, A2 => n3499, A3 => n3500, A4 => n3501
                           , ZN => n3497);
   U6869 : OAI22_X1 port map( A1 => n13953, A2 => n11179, B1 => n13985, B2 => 
                           n11176, ZN => n3501);
   U6870 : OAI222_X1 port map( A1 => n920, A2 => n11155, B1 => n14238, B2 => 
                           n11152, C1 => n14206, C2 => n11149, ZN => n3498);
   U6871 : OAI222_X1 port map( A1 => n14143, A2 => n11164, B1 => n14175, B2 => 
                           n11161, C1 => n14111, C2 => n11158, ZN => n3499);
   U6872 : NOR4_X1 port map( A1 => n4881, A2 => n4882, A3 => n4883, A4 => n4884
                           , ZN => n4880);
   U6873 : OAI22_X1 port map( A1 => n9575, A2 => n10981, B1 => n9574, B2 => 
                           n10978, ZN => n4884);
   U6874 : OAI222_X1 port map( A1 => n13920, A2 => n10957, B1 => n13856, B2 => 
                           n10954, C1 => n13888, C2 => n10951, ZN => n4881);
   U6875 : OAI222_X1 port map( A1 => n9569, A2 => n10966, B1 => n9568, B2 => 
                           n10963, C1 => n9570, C2 => n10960, ZN => n4882);
   U6876 : NOR4_X1 port map( A1 => n4890, A2 => n4891, A3 => n4892, A4 => n4893
                           , ZN => n4889);
   U6877 : OAI22_X1 port map( A1 => n13952, A2 => n10915, B1 => n13984, B2 => 
                           n10912, ZN => n4893);
   U6878 : OAI222_X1 port map( A1 => n916, A2 => n10891, B1 => n14237, B2 => 
                           n10888, C1 => n14205, C2 => n10885, ZN => n4890);
   U6879 : OAI222_X1 port map( A1 => n14142, A2 => n10900, B1 => n14174, B2 => 
                           n10897, C1 => n14110, C2 => n10894, ZN => n4891);
   U6880 : NOR4_X1 port map( A1 => n3448, A2 => n3449, A3 => n3450, A4 => n3451
                           , ZN => n3447);
   U6881 : OAI22_X1 port map( A1 => n9575, A2 => n11245, B1 => n9574, B2 => 
                           n11242, ZN => n3451);
   U6882 : OAI222_X1 port map( A1 => n13920, A2 => n11221, B1 => n13856, B2 => 
                           n11218, C1 => n13888, C2 => n11215, ZN => n3448);
   U6883 : OAI222_X1 port map( A1 => n9569, A2 => n11230, B1 => n9568, B2 => 
                           n11227, C1 => n9570, C2 => n11224, ZN => n3449);
   U6884 : NOR4_X1 port map( A1 => n3457, A2 => n3458, A3 => n3459, A4 => n3460
                           , ZN => n3456);
   U6885 : OAI22_X1 port map( A1 => n13952, A2 => n11179, B1 => n13984, B2 => 
                           n11176, ZN => n3460);
   U6886 : OAI222_X1 port map( A1 => n916, A2 => n11155, B1 => n14237, B2 => 
                           n11152, C1 => n14205, C2 => n11149, ZN => n3457);
   U6887 : OAI222_X1 port map( A1 => n14142, A2 => n11164, B1 => n14174, B2 => 
                           n11161, C1 => n14110, C2 => n11158, ZN => n3458);
   U6888 : NOR4_X1 port map( A1 => n4840, A2 => n4841, A3 => n4842, A4 => n4843
                           , ZN => n4839);
   U6889 : OAI22_X1 port map( A1 => n9209, A2 => n10981, B1 => n9208, B2 => 
                           n10978, ZN => n4843);
   U6890 : OAI222_X1 port map( A1 => n13919, A2 => n10957, B1 => n13855, B2 => 
                           n10954, C1 => n13887, C2 => n10951, ZN => n4840);
   U6891 : OAI222_X1 port map( A1 => n9203, A2 => n10966, B1 => n9202, B2 => 
                           n10963, C1 => n9204, C2 => n10960, ZN => n4841);
   U6892 : NOR4_X1 port map( A1 => n4849, A2 => n4850, A3 => n4851, A4 => n4852
                           , ZN => n4848);
   U6893 : OAI22_X1 port map( A1 => n13951, A2 => n10915, B1 => n13983, B2 => 
                           n10912, ZN => n4852);
   U6894 : OAI222_X1 port map( A1 => n912, A2 => n10891, B1 => n14236, B2 => 
                           n10888, C1 => n14204, C2 => n10885, ZN => n4849);
   U6895 : OAI222_X1 port map( A1 => n14141, A2 => n10900, B1 => n14173, B2 => 
                           n10897, C1 => n14109, C2 => n10894, ZN => n4850);
   U6896 : NOR4_X1 port map( A1 => n3407, A2 => n3408, A3 => n3409, A4 => n3410
                           , ZN => n3406);
   U6897 : OAI22_X1 port map( A1 => n9209, A2 => n11245, B1 => n9208, B2 => 
                           n11242, ZN => n3410);
   U6898 : OAI222_X1 port map( A1 => n13919, A2 => n11221, B1 => n13855, B2 => 
                           n11218, C1 => n13887, C2 => n11215, ZN => n3407);
   U6899 : OAI222_X1 port map( A1 => n9203, A2 => n11230, B1 => n9202, B2 => 
                           n11227, C1 => n9204, C2 => n11224, ZN => n3408);
   U6900 : NOR4_X1 port map( A1 => n3416, A2 => n3417, A3 => n3418, A4 => n3419
                           , ZN => n3415);
   U6901 : OAI22_X1 port map( A1 => n13951, A2 => n11179, B1 => n13983, B2 => 
                           n11176, ZN => n3419);
   U6902 : OAI222_X1 port map( A1 => n912, A2 => n11155, B1 => n14236, B2 => 
                           n11152, C1 => n14204, C2 => n11149, ZN => n3416);
   U6903 : OAI222_X1 port map( A1 => n14141, A2 => n11164, B1 => n14173, B2 => 
                           n11161, C1 => n14109, C2 => n11158, ZN => n3417);
   U6904 : NOR4_X1 port map( A1 => n4799, A2 => n4800, A3 => n4801, A4 => n4802
                           , ZN => n4798);
   U6905 : OAI22_X1 port map( A1 => n9177, A2 => n10981, B1 => n9176, B2 => 
                           n10978, ZN => n4802);
   U6906 : OAI222_X1 port map( A1 => n13918, A2 => n10957, B1 => n13854, B2 => 
                           n10954, C1 => n13886, C2 => n10951, ZN => n4799);
   U6907 : OAI222_X1 port map( A1 => n9171, A2 => n10966, B1 => n9170, B2 => 
                           n10963, C1 => n9172, C2 => n10960, ZN => n4800);
   U6908 : NOR4_X1 port map( A1 => n4808, A2 => n4809, A3 => n4810, A4 => n4811
                           , ZN => n4807);
   U6909 : OAI22_X1 port map( A1 => n13950, A2 => n10915, B1 => n13982, B2 => 
                           n10912, ZN => n4811);
   U6910 : OAI222_X1 port map( A1 => n908, A2 => n10891, B1 => n14235, B2 => 
                           n10888, C1 => n14203, C2 => n10885, ZN => n4808);
   U6911 : OAI222_X1 port map( A1 => n14140, A2 => n10900, B1 => n14172, B2 => 
                           n10897, C1 => n14108, C2 => n10894, ZN => n4809);
   U6912 : NOR4_X1 port map( A1 => n3366, A2 => n3367, A3 => n3368, A4 => n3369
                           , ZN => n3365);
   U6913 : OAI22_X1 port map( A1 => n9177, A2 => n11245, B1 => n9176, B2 => 
                           n11242, ZN => n3369);
   U6914 : OAI222_X1 port map( A1 => n13918, A2 => n11221, B1 => n13854, B2 => 
                           n11218, C1 => n13886, C2 => n11215, ZN => n3366);
   U6915 : OAI222_X1 port map( A1 => n9171, A2 => n11230, B1 => n9170, B2 => 
                           n11227, C1 => n9172, C2 => n11224, ZN => n3367);
   U6916 : NOR4_X1 port map( A1 => n3375, A2 => n3376, A3 => n3377, A4 => n3378
                           , ZN => n3374);
   U6917 : OAI22_X1 port map( A1 => n13950, A2 => n11179, B1 => n13982, B2 => 
                           n11176, ZN => n3378);
   U6918 : OAI222_X1 port map( A1 => n908, A2 => n11155, B1 => n14235, B2 => 
                           n11152, C1 => n14203, C2 => n11149, ZN => n3375);
   U6919 : OAI222_X1 port map( A1 => n14140, A2 => n11164, B1 => n14172, B2 => 
                           n11161, C1 => n14108, C2 => n11158, ZN => n3376);
   U6920 : NOR4_X1 port map( A1 => n4758, A2 => n4759, A3 => n4760, A4 => n4761
                           , ZN => n4757);
   U6921 : OAI22_X1 port map( A1 => n9145, A2 => n10981, B1 => n9144, B2 => 
                           n10978, ZN => n4761);
   U6922 : OAI222_X1 port map( A1 => n13917, A2 => n10957, B1 => n13853, B2 => 
                           n10954, C1 => n13885, C2 => n10951, ZN => n4758);
   U6923 : OAI222_X1 port map( A1 => n9139, A2 => n10966, B1 => n9138, B2 => 
                           n10963, C1 => n9140, C2 => n10960, ZN => n4759);
   U6924 : NOR4_X1 port map( A1 => n4767, A2 => n4768, A3 => n4769, A4 => n4770
                           , ZN => n4766);
   U6925 : OAI22_X1 port map( A1 => n13949, A2 => n10915, B1 => n13981, B2 => 
                           n10912, ZN => n4770);
   U6926 : OAI222_X1 port map( A1 => n904, A2 => n10891, B1 => n14234, B2 => 
                           n10888, C1 => n14202, C2 => n10885, ZN => n4767);
   U6927 : OAI222_X1 port map( A1 => n14139, A2 => n10900, B1 => n14171, B2 => 
                           n10897, C1 => n14107, C2 => n10894, ZN => n4768);
   U6928 : NOR4_X1 port map( A1 => n3325, A2 => n3326, A3 => n3327, A4 => n3328
                           , ZN => n3324);
   U6929 : OAI22_X1 port map( A1 => n9145, A2 => n11245, B1 => n9144, B2 => 
                           n11242, ZN => n3328);
   U6930 : OAI222_X1 port map( A1 => n13917, A2 => n11221, B1 => n13853, B2 => 
                           n11218, C1 => n13885, C2 => n11215, ZN => n3325);
   U6931 : OAI222_X1 port map( A1 => n9139, A2 => n11230, B1 => n9138, B2 => 
                           n11227, C1 => n9140, C2 => n11224, ZN => n3326);
   U6932 : NOR4_X1 port map( A1 => n3334, A2 => n3335, A3 => n3336, A4 => n3337
                           , ZN => n3333);
   U6933 : OAI22_X1 port map( A1 => n13949, A2 => n11179, B1 => n13981, B2 => 
                           n11176, ZN => n3337);
   U6934 : OAI222_X1 port map( A1 => n904, A2 => n11155, B1 => n14234, B2 => 
                           n11152, C1 => n14202, C2 => n11149, ZN => n3334);
   U6935 : OAI222_X1 port map( A1 => n14139, A2 => n11164, B1 => n14171, B2 => 
                           n11161, C1 => n14107, C2 => n11158, ZN => n3335);
   U6936 : NOR4_X1 port map( A1 => n4717, A2 => n4718, A3 => n4719, A4 => n4720
                           , ZN => n4716);
   U6937 : OAI22_X1 port map( A1 => n6010, A2 => n10981, B1 => n6009, B2 => 
                           n10978, ZN => n4720);
   U6938 : OAI222_X1 port map( A1 => n13916, A2 => n10957, B1 => n13852, B2 => 
                           n10954, C1 => n13884, C2 => n10951, ZN => n4717);
   U6939 : OAI222_X1 port map( A1 => n6004, A2 => n10966, B1 => n6003, B2 => 
                           n10963, C1 => n6005, C2 => n10960, ZN => n4718);
   U6940 : NOR4_X1 port map( A1 => n4726, A2 => n4727, A3 => n4728, A4 => n4729
                           , ZN => n4725);
   U6941 : OAI22_X1 port map( A1 => n13948, A2 => n10915, B1 => n13980, B2 => 
                           n10912, ZN => n4729);
   U6942 : OAI222_X1 port map( A1 => n900, A2 => n10891, B1 => n14233, B2 => 
                           n10888, C1 => n14201, C2 => n10885, ZN => n4726);
   U6943 : OAI222_X1 port map( A1 => n14138, A2 => n10900, B1 => n14170, B2 => 
                           n10897, C1 => n14106, C2 => n10894, ZN => n4727);
   U6944 : NOR4_X1 port map( A1 => n3284, A2 => n3285, A3 => n3286, A4 => n3287
                           , ZN => n3283);
   U6945 : OAI22_X1 port map( A1 => n6010, A2 => n11245, B1 => n6009, B2 => 
                           n11242, ZN => n3287);
   U6946 : OAI222_X1 port map( A1 => n13916, A2 => n11221, B1 => n13852, B2 => 
                           n11218, C1 => n13884, C2 => n11215, ZN => n3284);
   U6947 : OAI222_X1 port map( A1 => n6004, A2 => n11230, B1 => n6003, B2 => 
                           n11227, C1 => n6005, C2 => n11224, ZN => n3285);
   U6948 : NOR4_X1 port map( A1 => n3293, A2 => n3294, A3 => n3295, A4 => n3296
                           , ZN => n3292);
   U6949 : OAI22_X1 port map( A1 => n13948, A2 => n11179, B1 => n13980, B2 => 
                           n11176, ZN => n3296);
   U6950 : OAI222_X1 port map( A1 => n900, A2 => n11155, B1 => n14233, B2 => 
                           n11152, C1 => n14201, C2 => n11149, ZN => n3293);
   U6951 : OAI222_X1 port map( A1 => n14138, A2 => n11164, B1 => n14170, B2 => 
                           n11161, C1 => n14106, C2 => n11158, ZN => n3294);
   U6952 : NOR4_X1 port map( A1 => n4676, A2 => n4677, A3 => n4678, A4 => n4679
                           , ZN => n4675);
   U6953 : OAI22_X1 port map( A1 => n5946, A2 => n10982, B1 => n5945, B2 => 
                           n10979, ZN => n4679);
   U6954 : OAI222_X1 port map( A1 => n13915, A2 => n10958, B1 => n13851, B2 => 
                           n10955, C1 => n13883, C2 => n10952, ZN => n4676);
   U6955 : OAI222_X1 port map( A1 => n5940, A2 => n10967, B1 => n5939, B2 => 
                           n10964, C1 => n5941, C2 => n10961, ZN => n4677);
   U6956 : NOR4_X1 port map( A1 => n4685, A2 => n4686, A3 => n4687, A4 => n4688
                           , ZN => n4684);
   U6957 : OAI22_X1 port map( A1 => n13947, A2 => n10916, B1 => n13979, B2 => 
                           n10913, ZN => n4688);
   U6958 : OAI222_X1 port map( A1 => n896, A2 => n10892, B1 => n14232, B2 => 
                           n10889, C1 => n14200, C2 => n10886, ZN => n4685);
   U6959 : OAI222_X1 port map( A1 => n14137, A2 => n10901, B1 => n14169, B2 => 
                           n10898, C1 => n14105, C2 => n10895, ZN => n4686);
   U6960 : NOR4_X1 port map( A1 => n3243, A2 => n3244, A3 => n3245, A4 => n3246
                           , ZN => n3242);
   U6961 : OAI22_X1 port map( A1 => n5946, A2 => n11246, B1 => n5945, B2 => 
                           n11243, ZN => n3246);
   U6962 : OAI222_X1 port map( A1 => n13915, A2 => n11222, B1 => n13851, B2 => 
                           n11219, C1 => n13883, C2 => n11216, ZN => n3243);
   U6963 : OAI222_X1 port map( A1 => n5940, A2 => n11231, B1 => n5939, B2 => 
                           n11228, C1 => n5941, C2 => n11225, ZN => n3244);
   U6964 : NOR4_X1 port map( A1 => n3252, A2 => n3253, A3 => n3254, A4 => n3255
                           , ZN => n3251);
   U6965 : OAI22_X1 port map( A1 => n13947, A2 => n11180, B1 => n13979, B2 => 
                           n11177, ZN => n3255);
   U6966 : OAI222_X1 port map( A1 => n896, A2 => n11156, B1 => n14232, B2 => 
                           n11153, C1 => n14200, C2 => n11150, ZN => n3252);
   U6967 : OAI222_X1 port map( A1 => n14137, A2 => n11165, B1 => n14169, B2 => 
                           n11162, C1 => n14105, C2 => n11159, ZN => n3253);
   U6968 : NOR4_X1 port map( A1 => n4635, A2 => n4636, A3 => n4637, A4 => n4638
                           , ZN => n4634);
   U6969 : OAI22_X1 port map( A1 => n5914, A2 => n10982, B1 => n5913, B2 => 
                           n10979, ZN => n4638);
   U6970 : OAI222_X1 port map( A1 => n13914, A2 => n10958, B1 => n13850, B2 => 
                           n10955, C1 => n13882, C2 => n10952, ZN => n4635);
   U6971 : OAI222_X1 port map( A1 => n5908, A2 => n10967, B1 => n5907, B2 => 
                           n10964, C1 => n5909, C2 => n10961, ZN => n4636);
   U6972 : NOR4_X1 port map( A1 => n4644, A2 => n4645, A3 => n4646, A4 => n4647
                           , ZN => n4643);
   U6973 : OAI22_X1 port map( A1 => n13946, A2 => n10916, B1 => n13978, B2 => 
                           n10913, ZN => n4647);
   U6974 : OAI222_X1 port map( A1 => n892, A2 => n10892, B1 => n14231, B2 => 
                           n10889, C1 => n14199, C2 => n10886, ZN => n4644);
   U6975 : OAI222_X1 port map( A1 => n14136, A2 => n10901, B1 => n14168, B2 => 
                           n10898, C1 => n14104, C2 => n10895, ZN => n4645);
   U6976 : NOR4_X1 port map( A1 => n3202, A2 => n3203, A3 => n3204, A4 => n3205
                           , ZN => n3201);
   U6977 : OAI22_X1 port map( A1 => n5914, A2 => n11246, B1 => n5913, B2 => 
                           n11243, ZN => n3205);
   U6978 : OAI222_X1 port map( A1 => n13914, A2 => n11222, B1 => n13850, B2 => 
                           n11219, C1 => n13882, C2 => n11216, ZN => n3202);
   U6979 : OAI222_X1 port map( A1 => n5908, A2 => n11231, B1 => n5907, B2 => 
                           n11228, C1 => n5909, C2 => n11225, ZN => n3203);
   U6980 : NOR4_X1 port map( A1 => n3211, A2 => n3212, A3 => n3213, A4 => n3214
                           , ZN => n3210);
   U6981 : OAI22_X1 port map( A1 => n13946, A2 => n11180, B1 => n13978, B2 => 
                           n11177, ZN => n3214);
   U6982 : OAI222_X1 port map( A1 => n892, A2 => n11156, B1 => n14231, B2 => 
                           n11153, C1 => n14199, C2 => n11150, ZN => n3211);
   U6983 : OAI222_X1 port map( A1 => n14136, A2 => n11165, B1 => n14168, B2 => 
                           n11162, C1 => n14104, C2 => n11159, ZN => n3212);
   U6984 : NOR4_X1 port map( A1 => n4594, A2 => n4595, A3 => n4596, A4 => n4597
                           , ZN => n4593);
   U6985 : OAI22_X1 port map( A1 => n5882, A2 => n10982, B1 => n5881, B2 => 
                           n10979, ZN => n4597);
   U6986 : OAI222_X1 port map( A1 => n13913, A2 => n10958, B1 => n13849, B2 => 
                           n10955, C1 => n13881, C2 => n10952, ZN => n4594);
   U6987 : OAI222_X1 port map( A1 => n5876, A2 => n10967, B1 => n5875, B2 => 
                           n10964, C1 => n5877, C2 => n10961, ZN => n4595);
   U6988 : NOR4_X1 port map( A1 => n4603, A2 => n4604, A3 => n4605, A4 => n4606
                           , ZN => n4602);
   U6989 : OAI22_X1 port map( A1 => n13945, A2 => n10916, B1 => n13977, B2 => 
                           n10913, ZN => n4606);
   U6990 : OAI222_X1 port map( A1 => n888, A2 => n10892, B1 => n14230, B2 => 
                           n10889, C1 => n14198, C2 => n10886, ZN => n4603);
   U6991 : OAI222_X1 port map( A1 => n14135, A2 => n10901, B1 => n14167, B2 => 
                           n10898, C1 => n14103, C2 => n10895, ZN => n4604);
   U6992 : NOR4_X1 port map( A1 => n3161, A2 => n3162, A3 => n3163, A4 => n3164
                           , ZN => n3160);
   U6993 : OAI22_X1 port map( A1 => n5882, A2 => n11246, B1 => n5881, B2 => 
                           n11243, ZN => n3164);
   U6994 : OAI222_X1 port map( A1 => n13913, A2 => n11222, B1 => n13849, B2 => 
                           n11219, C1 => n13881, C2 => n11216, ZN => n3161);
   U6995 : OAI222_X1 port map( A1 => n5876, A2 => n11231, B1 => n5875, B2 => 
                           n11228, C1 => n5877, C2 => n11225, ZN => n3162);
   U6996 : NOR4_X1 port map( A1 => n3170, A2 => n3171, A3 => n3172, A4 => n3173
                           , ZN => n3169);
   U6997 : OAI22_X1 port map( A1 => n13945, A2 => n11180, B1 => n13977, B2 => 
                           n11177, ZN => n3173);
   U6998 : OAI222_X1 port map( A1 => n888, A2 => n11156, B1 => n14230, B2 => 
                           n11153, C1 => n14198, C2 => n11150, ZN => n3170);
   U6999 : OAI222_X1 port map( A1 => n14135, A2 => n11165, B1 => n14167, B2 => 
                           n11162, C1 => n14103, C2 => n11159, ZN => n3171);
   U7000 : NOR4_X1 port map( A1 => n4553, A2 => n4554, A3 => n4555, A4 => n4556
                           , ZN => n4552);
   U7001 : OAI22_X1 port map( A1 => n5850, A2 => n10982, B1 => n5849, B2 => 
                           n10979, ZN => n4556);
   U7002 : OAI222_X1 port map( A1 => n13912, A2 => n10958, B1 => n13848, B2 => 
                           n10955, C1 => n13880, C2 => n10952, ZN => n4553);
   U7003 : OAI222_X1 port map( A1 => n5844, A2 => n10967, B1 => n5843, B2 => 
                           n10964, C1 => n5845, C2 => n10961, ZN => n4554);
   U7004 : NOR4_X1 port map( A1 => n4562, A2 => n4563, A3 => n4564, A4 => n4565
                           , ZN => n4561);
   U7005 : OAI22_X1 port map( A1 => n13944, A2 => n10916, B1 => n13976, B2 => 
                           n10913, ZN => n4565);
   U7006 : OAI222_X1 port map( A1 => n884, A2 => n10892, B1 => n14229, B2 => 
                           n10889, C1 => n14197, C2 => n10886, ZN => n4562);
   U7007 : OAI222_X1 port map( A1 => n14134, A2 => n10901, B1 => n14166, B2 => 
                           n10898, C1 => n14102, C2 => n10895, ZN => n4563);
   U7008 : NOR4_X1 port map( A1 => n3120, A2 => n3121, A3 => n3122, A4 => n3123
                           , ZN => n3119);
   U7009 : OAI22_X1 port map( A1 => n5850, A2 => n11246, B1 => n5849, B2 => 
                           n11243, ZN => n3123);
   U7010 : OAI222_X1 port map( A1 => n13912, A2 => n11222, B1 => n13848, B2 => 
                           n11219, C1 => n13880, C2 => n11216, ZN => n3120);
   U7011 : OAI222_X1 port map( A1 => n5844, A2 => n11231, B1 => n5843, B2 => 
                           n11228, C1 => n5845, C2 => n11225, ZN => n3121);
   U7012 : NOR4_X1 port map( A1 => n3129, A2 => n3130, A3 => n3131, A4 => n3132
                           , ZN => n3128);
   U7013 : OAI22_X1 port map( A1 => n13944, A2 => n11180, B1 => n13976, B2 => 
                           n11177, ZN => n3132);
   U7014 : OAI222_X1 port map( A1 => n884, A2 => n11156, B1 => n14229, B2 => 
                           n11153, C1 => n14197, C2 => n11150, ZN => n3129);
   U7015 : OAI222_X1 port map( A1 => n14134, A2 => n11165, B1 => n14166, B2 => 
                           n11162, C1 => n14102, C2 => n11159, ZN => n3130);
   U7016 : NOR4_X1 port map( A1 => n4512, A2 => n4513, A3 => n4514, A4 => n4515
                           , ZN => n4511);
   U7017 : OAI22_X1 port map( A1 => n5818, A2 => n10982, B1 => n5817, B2 => 
                           n10979, ZN => n4515);
   U7018 : OAI222_X1 port map( A1 => n13911, A2 => n10958, B1 => n13847, B2 => 
                           n10955, C1 => n13879, C2 => n10952, ZN => n4512);
   U7019 : OAI222_X1 port map( A1 => n5812, A2 => n10967, B1 => n5811, B2 => 
                           n10964, C1 => n5813, C2 => n10961, ZN => n4513);
   U7020 : NOR4_X1 port map( A1 => n4521, A2 => n4522, A3 => n4523, A4 => n4524
                           , ZN => n4520);
   U7021 : OAI22_X1 port map( A1 => n13943, A2 => n10916, B1 => n13975, B2 => 
                           n10913, ZN => n4524);
   U7022 : OAI222_X1 port map( A1 => n880, A2 => n10892, B1 => n14228, B2 => 
                           n10889, C1 => n14196, C2 => n10886, ZN => n4521);
   U7023 : OAI222_X1 port map( A1 => n14133, A2 => n10901, B1 => n14165, B2 => 
                           n10898, C1 => n14101, C2 => n10895, ZN => n4522);
   U7024 : NOR4_X1 port map( A1 => n3079, A2 => n3080, A3 => n3081, A4 => n3082
                           , ZN => n3078);
   U7025 : OAI22_X1 port map( A1 => n5818, A2 => n11246, B1 => n5817, B2 => 
                           n11243, ZN => n3082);
   U7026 : OAI222_X1 port map( A1 => n13911, A2 => n11222, B1 => n13847, B2 => 
                           n11219, C1 => n13879, C2 => n11216, ZN => n3079);
   U7027 : OAI222_X1 port map( A1 => n5812, A2 => n11231, B1 => n5811, B2 => 
                           n11228, C1 => n5813, C2 => n11225, ZN => n3080);
   U7028 : NOR4_X1 port map( A1 => n3088, A2 => n3089, A3 => n3090, A4 => n3091
                           , ZN => n3087);
   U7029 : OAI22_X1 port map( A1 => n13943, A2 => n11180, B1 => n13975, B2 => 
                           n11177, ZN => n3091);
   U7030 : OAI222_X1 port map( A1 => n880, A2 => n11156, B1 => n14228, B2 => 
                           n11153, C1 => n14196, C2 => n11150, ZN => n3088);
   U7031 : OAI222_X1 port map( A1 => n14133, A2 => n11165, B1 => n14165, B2 => 
                           n11162, C1 => n14101, C2 => n11159, ZN => n3089);
   U7032 : NOR4_X1 port map( A1 => n4471, A2 => n4472, A3 => n4473, A4 => n4474
                           , ZN => n4470);
   U7033 : OAI22_X1 port map( A1 => n5786, A2 => n10982, B1 => n5785, B2 => 
                           n10979, ZN => n4474);
   U7034 : OAI222_X1 port map( A1 => n13910, A2 => n10958, B1 => n13846, B2 => 
                           n10955, C1 => n13878, C2 => n10952, ZN => n4471);
   U7035 : OAI222_X1 port map( A1 => n5780, A2 => n10967, B1 => n5779, B2 => 
                           n10964, C1 => n5781, C2 => n10961, ZN => n4472);
   U7036 : NOR4_X1 port map( A1 => n4480, A2 => n4481, A3 => n4482, A4 => n4483
                           , ZN => n4479);
   U7037 : OAI22_X1 port map( A1 => n13942, A2 => n10916, B1 => n13974, B2 => 
                           n10913, ZN => n4483);
   U7038 : OAI222_X1 port map( A1 => n876, A2 => n10892, B1 => n14227, B2 => 
                           n10889, C1 => n14195, C2 => n10886, ZN => n4480);
   U7039 : OAI222_X1 port map( A1 => n14132, A2 => n10901, B1 => n14164, B2 => 
                           n10898, C1 => n14100, C2 => n10895, ZN => n4481);
   U7040 : NOR4_X1 port map( A1 => n3038, A2 => n3039, A3 => n3040, A4 => n3041
                           , ZN => n3037);
   U7041 : OAI22_X1 port map( A1 => n5786, A2 => n11246, B1 => n5785, B2 => 
                           n11243, ZN => n3041);
   U7042 : OAI222_X1 port map( A1 => n13910, A2 => n11222, B1 => n13846, B2 => 
                           n11219, C1 => n13878, C2 => n11216, ZN => n3038);
   U7043 : OAI222_X1 port map( A1 => n5780, A2 => n11231, B1 => n5779, B2 => 
                           n11228, C1 => n5781, C2 => n11225, ZN => n3039);
   U7044 : NOR4_X1 port map( A1 => n3047, A2 => n3048, A3 => n3049, A4 => n3050
                           , ZN => n3046);
   U7045 : OAI22_X1 port map( A1 => n13942, A2 => n11180, B1 => n13974, B2 => 
                           n11177, ZN => n3050);
   U7046 : OAI222_X1 port map( A1 => n876, A2 => n11156, B1 => n14227, B2 => 
                           n11153, C1 => n14195, C2 => n11150, ZN => n3047);
   U7047 : OAI222_X1 port map( A1 => n14132, A2 => n11165, B1 => n14164, B2 => 
                           n11162, C1 => n14100, C2 => n11159, ZN => n3048);
   U7048 : NOR4_X1 port map( A1 => n4430, A2 => n4431, A3 => n4432, A4 => n4433
                           , ZN => n4429);
   U7049 : OAI22_X1 port map( A1 => n5754, A2 => n10982, B1 => n5753, B2 => 
                           n10979, ZN => n4433);
   U7050 : OAI222_X1 port map( A1 => n13909, A2 => n10958, B1 => n13845, B2 => 
                           n10955, C1 => n13877, C2 => n10952, ZN => n4430);
   U7051 : OAI222_X1 port map( A1 => n5748, A2 => n10967, B1 => n5747, B2 => 
                           n10964, C1 => n5749, C2 => n10961, ZN => n4431);
   U7052 : NOR4_X1 port map( A1 => n4439, A2 => n4440, A3 => n4441, A4 => n4442
                           , ZN => n4438);
   U7053 : OAI22_X1 port map( A1 => n13941, A2 => n10916, B1 => n13973, B2 => 
                           n10913, ZN => n4442);
   U7054 : OAI222_X1 port map( A1 => n872, A2 => n10892, B1 => n14226, B2 => 
                           n10889, C1 => n14194, C2 => n10886, ZN => n4439);
   U7055 : OAI222_X1 port map( A1 => n14131, A2 => n10901, B1 => n14163, B2 => 
                           n10898, C1 => n14099, C2 => n10895, ZN => n4440);
   U7056 : NOR4_X1 port map( A1 => n2997, A2 => n2998, A3 => n2999, A4 => n3000
                           , ZN => n2996);
   U7057 : OAI22_X1 port map( A1 => n5754, A2 => n11246, B1 => n5753, B2 => 
                           n11243, ZN => n3000);
   U7058 : OAI222_X1 port map( A1 => n13909, A2 => n11222, B1 => n13845, B2 => 
                           n11219, C1 => n13877, C2 => n11216, ZN => n2997);
   U7059 : OAI222_X1 port map( A1 => n5748, A2 => n11231, B1 => n5747, B2 => 
                           n11228, C1 => n5749, C2 => n11225, ZN => n2998);
   U7060 : NOR4_X1 port map( A1 => n3006, A2 => n3007, A3 => n3008, A4 => n3009
                           , ZN => n3005);
   U7061 : OAI22_X1 port map( A1 => n13941, A2 => n11180, B1 => n13973, B2 => 
                           n11177, ZN => n3009);
   U7062 : OAI222_X1 port map( A1 => n872, A2 => n11156, B1 => n14226, B2 => 
                           n11153, C1 => n14194, C2 => n11150, ZN => n3006);
   U7063 : OAI222_X1 port map( A1 => n14131, A2 => n11165, B1 => n14163, B2 => 
                           n11162, C1 => n14099, C2 => n11159, ZN => n3007);
   U7064 : NOR4_X1 port map( A1 => n4345, A2 => n4346, A3 => n4347, A4 => n4348
                           , ZN => n4344);
   U7065 : OAI22_X1 port map( A1 => n5722, A2 => n10982, B1 => n5721, B2 => 
                           n10979, ZN => n4348);
   U7066 : OAI222_X1 port map( A1 => n13908, A2 => n10958, B1 => n13844, B2 => 
                           n10955, C1 => n13876, C2 => n10952, ZN => n4345);
   U7067 : OAI222_X1 port map( A1 => n5716, A2 => n10967, B1 => n5715, B2 => 
                           n10964, C1 => n5717, C2 => n10961, ZN => n4346);
   U7068 : NOR4_X1 port map( A1 => n4376, A2 => n4377, A3 => n4378, A4 => n4379
                           , ZN => n4375);
   U7069 : OAI22_X1 port map( A1 => n13940, A2 => n10916, B1 => n13972, B2 => 
                           n10913, ZN => n4379);
   U7070 : OAI222_X1 port map( A1 => n868, A2 => n10892, B1 => n14225, B2 => 
                           n10889, C1 => n996, C2 => n10886, ZN => n4376);
   U7071 : OAI222_X1 port map( A1 => n14130, A2 => n10901, B1 => n14162, B2 => 
                           n10898, C1 => n997, C2 => n10895, ZN => n4377);
   U7072 : NOR4_X1 port map( A1 => n2877, A2 => n2878, A3 => n2879, A4 => n2880
                           , ZN => n2876);
   U7073 : OAI22_X1 port map( A1 => n5722, A2 => n11246, B1 => n5721, B2 => 
                           n11243, ZN => n2880);
   U7074 : OAI222_X1 port map( A1 => n13908, A2 => n11222, B1 => n13844, B2 => 
                           n11219, C1 => n13876, C2 => n11216, ZN => n2877);
   U7075 : OAI222_X1 port map( A1 => n5716, A2 => n11231, B1 => n5715, B2 => 
                           n11228, C1 => n5717, C2 => n11225, ZN => n2878);
   U7076 : NOR4_X1 port map( A1 => n2943, A2 => n2944, A3 => n2945, A4 => n2946
                           , ZN => n2942);
   U7077 : OAI22_X1 port map( A1 => n13940, A2 => n11180, B1 => n13972, B2 => 
                           n11177, ZN => n2946);
   U7078 : OAI222_X1 port map( A1 => n868, A2 => n11156, B1 => n14225, B2 => 
                           n11153, C1 => n996, C2 => n11150, ZN => n2943);
   U7079 : OAI222_X1 port map( A1 => n14130, A2 => n11165, B1 => n14162, B2 => 
                           n11162, C1 => n997, C2 => n11159, ZN => n2944);
   U7080 : AOI221_X1 port map( B1 => n10947, B2 => n9504, C1 => n10944, C2 => 
                           n9536, A => n5691, ZN => n5681);
   U7081 : OAI222_X1 port map( A1 => n13619, A2 => n10941, B1 => n13651, B2 => 
                           n10938, C1 => n13587, C2 => n10935, ZN => n5691);
   U7082 : AOI221_X1 port map( B1 => n10881, B2 => n14288, C1 => n10878, C2 => 
                           n14480, A => n5704, ZN => n5695);
   U7083 : OAI222_X1 port map( A1 => n10510, A2 => n10875, B1 => n10509, B2 => 
                           n10872, C1 => n10511, C2 => n10869, ZN => n5704);
   U7084 : AOI221_X1 port map( B1 => n11211, B2 => n9504, C1 => n11208, C2 => 
                           n9536, A => n4258, ZN => n4248);
   U7085 : OAI222_X1 port map( A1 => n13619, A2 => n11205, B1 => n13651, B2 => 
                           n11202, C1 => n13587, C2 => n11199, ZN => n4258);
   U7086 : AOI221_X1 port map( B1 => n11145, B2 => n14288, C1 => n11142, C2 => 
                           n14480, A => n4271, ZN => n4262);
   U7087 : OAI222_X1 port map( A1 => n10510, A2 => n11139, B1 => n10509, B2 => 
                           n11136, C1 => n10511, C2 => n11133, ZN => n4271);
   U7088 : AOI221_X1 port map( B1 => n10947, B2 => n9505, C1 => n10944, C2 => 
                           n9537, A => n5623, ZN => n5617);
   U7089 : OAI222_X1 port map( A1 => n13618, A2 => n10941, B1 => n13650, B2 => 
                           n10938, C1 => n13586, C2 => n10935, ZN => n5623);
   U7090 : AOI221_X1 port map( B1 => n10881, B2 => n14287, C1 => n10878, C2 => 
                           n14479, A => n5632, ZN => n5626);
   U7091 : OAI222_X1 port map( A1 => n10478, A2 => n10875, B1 => n10477, B2 => 
                           n10872, C1 => n10479, C2 => n10869, ZN => n5632);
   U7092 : AOI221_X1 port map( B1 => n11211, B2 => n9505, C1 => n11208, C2 => 
                           n9537, A => n4190, ZN => n4184);
   U7093 : OAI222_X1 port map( A1 => n13618, A2 => n11205, B1 => n13650, B2 => 
                           n11202, C1 => n13586, C2 => n11199, ZN => n4190);
   U7094 : AOI221_X1 port map( B1 => n11145, B2 => n14287, C1 => n11142, C2 => 
                           n14479, A => n4199, ZN => n4193);
   U7095 : OAI222_X1 port map( A1 => n10478, A2 => n11139, B1 => n10477, B2 => 
                           n11136, C1 => n10479, C2 => n11133, ZN => n4199);
   U7096 : AOI221_X1 port map( B1 => n10947, B2 => n9506, C1 => n10944, C2 => 
                           n9538, A => n5582, ZN => n5576);
   U7097 : OAI222_X1 port map( A1 => n13617, A2 => n10941, B1 => n13649, B2 => 
                           n10938, C1 => n13585, C2 => n10935, ZN => n5582);
   U7098 : AOI221_X1 port map( B1 => n10881, B2 => n14286, C1 => n10878, C2 => 
                           n14478, A => n5591, ZN => n5585);
   U7099 : OAI222_X1 port map( A1 => n10446, A2 => n10875, B1 => n10445, B2 => 
                           n10872, C1 => n10447, C2 => n10869, ZN => n5591);
   U7100 : AOI221_X1 port map( B1 => n11211, B2 => n9506, C1 => n11208, C2 => 
                           n9538, A => n4149, ZN => n4143);
   U7101 : OAI222_X1 port map( A1 => n13617, A2 => n11205, B1 => n13649, B2 => 
                           n11202, C1 => n13585, C2 => n11199, ZN => n4149);
   U7102 : AOI221_X1 port map( B1 => n11145, B2 => n14286, C1 => n11142, C2 => 
                           n14478, A => n4158, ZN => n4152);
   U7103 : OAI222_X1 port map( A1 => n10446, A2 => n11139, B1 => n10445, B2 => 
                           n11136, C1 => n10447, C2 => n11133, ZN => n4158);
   U7104 : AOI221_X1 port map( B1 => n10947, B2 => n9507, C1 => n10944, C2 => 
                           n9539, A => n5541, ZN => n5535);
   U7105 : OAI222_X1 port map( A1 => n13616, A2 => n10941, B1 => n13648, B2 => 
                           n10938, C1 => n13584, C2 => n10935, ZN => n5541);
   U7106 : AOI221_X1 port map( B1 => n10881, B2 => n14285, C1 => n10878, C2 => 
                           n14477, A => n5550, ZN => n5544);
   U7107 : OAI222_X1 port map( A1 => n10414, A2 => n10875, B1 => n10413, B2 => 
                           n10872, C1 => n10415, C2 => n10869, ZN => n5550);
   U7108 : AOI221_X1 port map( B1 => n11211, B2 => n9507, C1 => n11208, C2 => 
                           n9539, A => n4108, ZN => n4102);
   U7109 : OAI222_X1 port map( A1 => n13616, A2 => n11205, B1 => n13648, B2 => 
                           n11202, C1 => n13584, C2 => n11199, ZN => n4108);
   U7110 : AOI221_X1 port map( B1 => n11145, B2 => n14285, C1 => n11142, C2 => 
                           n14477, A => n4117, ZN => n4111);
   U7111 : OAI222_X1 port map( A1 => n10414, A2 => n11139, B1 => n10413, B2 => 
                           n11136, C1 => n10415, C2 => n11133, ZN => n4117);
   U7112 : AOI221_X1 port map( B1 => n10947, B2 => n9508, C1 => n10944, C2 => 
                           n9540, A => n5500, ZN => n5494);
   U7113 : OAI222_X1 port map( A1 => n13615, A2 => n10941, B1 => n13647, B2 => 
                           n10938, C1 => n13583, C2 => n10935, ZN => n5500);
   U7114 : AOI221_X1 port map( B1 => n10881, B2 => n14284, C1 => n10878, C2 => 
                           n14476, A => n5509, ZN => n5503);
   U7115 : OAI222_X1 port map( A1 => n10379, A2 => n10875, B1 => n10378, B2 => 
                           n10872, C1 => n10380, C2 => n10869, ZN => n5509);
   U7116 : AOI221_X1 port map( B1 => n11211, B2 => n9508, C1 => n11208, C2 => 
                           n9540, A => n4067, ZN => n4061);
   U7117 : OAI222_X1 port map( A1 => n13615, A2 => n11205, B1 => n13647, B2 => 
                           n11202, C1 => n13583, C2 => n11199, ZN => n4067);
   U7118 : AOI221_X1 port map( B1 => n11145, B2 => n14284, C1 => n11142, C2 => 
                           n14476, A => n4076, ZN => n4070);
   U7119 : OAI222_X1 port map( A1 => n10379, A2 => n11139, B1 => n10378, B2 => 
                           n11136, C1 => n10380, C2 => n11133, ZN => n4076);
   U7120 : AOI221_X1 port map( B1 => n10947, B2 => n9509, C1 => n10944, C2 => 
                           n9541, A => n5459, ZN => n5453);
   U7121 : OAI222_X1 port map( A1 => n13614, A2 => n10941, B1 => n13646, B2 => 
                           n10938, C1 => n13582, C2 => n10935, ZN => n5459);
   U7122 : AOI221_X1 port map( B1 => n10881, B2 => n14283, C1 => n10878, C2 => 
                           n14475, A => n5468, ZN => n5462);
   U7123 : OAI222_X1 port map( A1 => n10347, A2 => n10875, B1 => n10346, B2 => 
                           n10872, C1 => n10348, C2 => n10869, ZN => n5468);
   U7124 : AOI221_X1 port map( B1 => n11211, B2 => n9509, C1 => n11208, C2 => 
                           n9541, A => n4026, ZN => n4020);
   U7125 : OAI222_X1 port map( A1 => n13614, A2 => n11205, B1 => n13646, B2 => 
                           n11202, C1 => n13582, C2 => n11199, ZN => n4026);
   U7126 : AOI221_X1 port map( B1 => n11145, B2 => n14283, C1 => n11142, C2 => 
                           n14475, A => n4035, ZN => n4029);
   U7127 : OAI222_X1 port map( A1 => n10347, A2 => n11139, B1 => n10346, B2 => 
                           n11136, C1 => n10348, C2 => n11133, ZN => n4035);
   U7128 : AOI221_X1 port map( B1 => n10947, B2 => n9510, C1 => n10944, C2 => 
                           n9542, A => n5418, ZN => n5412);
   U7129 : OAI222_X1 port map( A1 => n13613, A2 => n10941, B1 => n13645, B2 => 
                           n10938, C1 => n13581, C2 => n10935, ZN => n5418);
   U7130 : AOI221_X1 port map( B1 => n10881, B2 => n14282, C1 => n10878, C2 => 
                           n14474, A => n5427, ZN => n5421);
   U7131 : OAI222_X1 port map( A1 => n10315, A2 => n10875, B1 => n10314, B2 => 
                           n10872, C1 => n10316, C2 => n10869, ZN => n5427);
   U7132 : AOI221_X1 port map( B1 => n11211, B2 => n9510, C1 => n11208, C2 => 
                           n9542, A => n3985, ZN => n3979);
   U7133 : OAI222_X1 port map( A1 => n13613, A2 => n11205, B1 => n13645, B2 => 
                           n11202, C1 => n13581, C2 => n11199, ZN => n3985);
   U7134 : AOI221_X1 port map( B1 => n11145, B2 => n14282, C1 => n11142, C2 => 
                           n14474, A => n3994, ZN => n3988);
   U7135 : OAI222_X1 port map( A1 => n10315, A2 => n11139, B1 => n10314, B2 => 
                           n11136, C1 => n10316, C2 => n11133, ZN => n3994);
   U7136 : AOI221_X1 port map( B1 => n10947, B2 => n9511, C1 => n10944, C2 => 
                           n9543, A => n5377, ZN => n5371);
   U7137 : OAI222_X1 port map( A1 => n13612, A2 => n10941, B1 => n13644, B2 => 
                           n10938, C1 => n13580, C2 => n10935, ZN => n5377);
   U7138 : AOI221_X1 port map( B1 => n10881, B2 => n14281, C1 => n10878, C2 => 
                           n14473, A => n5386, ZN => n5380);
   U7139 : OAI222_X1 port map( A1 => n10280, A2 => n10875, B1 => n10279, B2 => 
                           n10872, C1 => n10281, C2 => n10869, ZN => n5386);
   U7140 : AOI221_X1 port map( B1 => n11211, B2 => n9511, C1 => n11208, C2 => 
                           n9543, A => n3944, ZN => n3938);
   U7141 : OAI222_X1 port map( A1 => n13612, A2 => n11205, B1 => n13644, B2 => 
                           n11202, C1 => n13580, C2 => n11199, ZN => n3944);
   U7142 : AOI221_X1 port map( B1 => n11145, B2 => n14281, C1 => n11142, C2 => 
                           n14473, A => n3953, ZN => n3947);
   U7143 : OAI222_X1 port map( A1 => n10280, A2 => n11139, B1 => n10279, B2 => 
                           n11136, C1 => n10281, C2 => n11133, ZN => n3953);
   U7144 : AOI221_X1 port map( B1 => n10947, B2 => n9512, C1 => n10944, C2 => 
                           n9544, A => n5336, ZN => n5330);
   U7145 : OAI222_X1 port map( A1 => n13611, A2 => n10941, B1 => n13643, B2 => 
                           n10938, C1 => n13579, C2 => n10935, ZN => n5336);
   U7146 : AOI221_X1 port map( B1 => n10881, B2 => n14280, C1 => n10878, C2 => 
                           n14472, A => n5345, ZN => n5339);
   U7147 : OAI222_X1 port map( A1 => n10248, A2 => n10875, B1 => n10247, B2 => 
                           n10872, C1 => n10249, C2 => n10869, ZN => n5345);
   U7148 : AOI221_X1 port map( B1 => n11211, B2 => n9512, C1 => n11208, C2 => 
                           n9544, A => n3903, ZN => n3897);
   U7149 : OAI222_X1 port map( A1 => n13611, A2 => n11205, B1 => n13643, B2 => 
                           n11202, C1 => n13579, C2 => n11199, ZN => n3903);
   U7150 : AOI221_X1 port map( B1 => n11145, B2 => n14280, C1 => n11142, C2 => 
                           n14472, A => n3912, ZN => n3906);
   U7151 : OAI222_X1 port map( A1 => n10248, A2 => n11139, B1 => n10247, B2 => 
                           n11136, C1 => n10249, C2 => n11133, ZN => n3912);
   U7152 : AOI221_X1 port map( B1 => n10947, B2 => n9513, C1 => n10944, C2 => 
                           n9545, A => n5295, ZN => n5289);
   U7153 : OAI222_X1 port map( A1 => n13610, A2 => n10941, B1 => n13642, B2 => 
                           n10938, C1 => n13578, C2 => n10935, ZN => n5295);
   U7154 : AOI221_X1 port map( B1 => n10881, B2 => n14279, C1 => n10878, C2 => 
                           n14471, A => n5304, ZN => n5298);
   U7155 : OAI222_X1 port map( A1 => n10216, A2 => n10875, B1 => n10215, B2 => 
                           n10872, C1 => n10217, C2 => n10869, ZN => n5304);
   U7156 : AOI221_X1 port map( B1 => n11211, B2 => n9513, C1 => n11208, C2 => 
                           n9545, A => n3862, ZN => n3856);
   U7157 : OAI222_X1 port map( A1 => n13610, A2 => n11205, B1 => n13642, B2 => 
                           n11202, C1 => n13578, C2 => n11199, ZN => n3862);
   U7158 : AOI221_X1 port map( B1 => n11145, B2 => n14279, C1 => n11142, C2 => 
                           n14471, A => n3871, ZN => n3865);
   U7159 : OAI222_X1 port map( A1 => n10216, A2 => n11139, B1 => n10215, B2 => 
                           n11136, C1 => n10217, C2 => n11133, ZN => n3871);
   U7160 : AOI221_X1 port map( B1 => n10947, B2 => n9514, C1 => n10944, C2 => 
                           n9546, A => n5254, ZN => n5248);
   U7161 : OAI222_X1 port map( A1 => n13609, A2 => n10941, B1 => n13641, B2 => 
                           n10938, C1 => n13577, C2 => n10935, ZN => n5254);
   U7162 : AOI221_X1 port map( B1 => n10881, B2 => n14278, C1 => n10878, C2 => 
                           n14470, A => n5263, ZN => n5257);
   U7163 : OAI222_X1 port map( A1 => n10182, A2 => n10875, B1 => n10181, B2 => 
                           n10872, C1 => n10183, C2 => n10869, ZN => n5263);
   U7164 : AOI221_X1 port map( B1 => n11211, B2 => n9514, C1 => n11208, C2 => 
                           n9546, A => n3821, ZN => n3815);
   U7165 : OAI222_X1 port map( A1 => n13609, A2 => n11205, B1 => n13641, B2 => 
                           n11202, C1 => n13577, C2 => n11199, ZN => n3821);
   U7166 : AOI221_X1 port map( B1 => n11145, B2 => n14278, C1 => n11142, C2 => 
                           n14470, A => n3830, ZN => n3824);
   U7167 : OAI222_X1 port map( A1 => n10182, A2 => n11139, B1 => n10181, B2 => 
                           n11136, C1 => n10183, C2 => n11133, ZN => n3830);
   U7168 : AOI221_X1 port map( B1 => n10947, B2 => n9515, C1 => n10944, C2 => 
                           n9547, A => n5213, ZN => n5207);
   U7169 : OAI222_X1 port map( A1 => n13608, A2 => n10941, B1 => n13640, B2 => 
                           n10938, C1 => n13576, C2 => n10935, ZN => n5213);
   U7170 : AOI221_X1 port map( B1 => n10881, B2 => n14277, C1 => n10878, C2 => 
                           n14469, A => n5222, ZN => n5216);
   U7171 : OAI222_X1 port map( A1 => n10150, A2 => n10875, B1 => n10149, B2 => 
                           n10872, C1 => n10151, C2 => n10869, ZN => n5222);
   U7172 : AOI221_X1 port map( B1 => n11211, B2 => n9515, C1 => n11208, C2 => 
                           n9547, A => n3780, ZN => n3774);
   U7173 : OAI222_X1 port map( A1 => n13608, A2 => n11205, B1 => n13640, B2 => 
                           n11202, C1 => n13576, C2 => n11199, ZN => n3780);
   U7174 : AOI221_X1 port map( B1 => n11145, B2 => n14277, C1 => n11142, C2 => 
                           n14469, A => n3789, ZN => n3783);
   U7175 : OAI222_X1 port map( A1 => n10150, A2 => n11139, B1 => n10149, B2 => 
                           n11136, C1 => n10151, C2 => n11133, ZN => n3789);
   U7176 : AOI221_X1 port map( B1 => n10948, B2 => n9516, C1 => n10945, C2 => 
                           n9548, A => n5172, ZN => n5166);
   U7177 : OAI222_X1 port map( A1 => n13607, A2 => n10942, B1 => n13639, B2 => 
                           n10939, C1 => n13575, C2 => n10936, ZN => n5172);
   U7178 : AOI221_X1 port map( B1 => n10882, B2 => n14276, C1 => n10879, C2 => 
                           n14468, A => n5181, ZN => n5175);
   U7179 : OAI222_X1 port map( A1 => n10118, A2 => n10876, B1 => n10117, B2 => 
                           n10873, C1 => n10119, C2 => n10870, ZN => n5181);
   U7180 : AOI221_X1 port map( B1 => n11212, B2 => n9516, C1 => n11209, C2 => 
                           n9548, A => n3739, ZN => n3733);
   U7181 : OAI222_X1 port map( A1 => n13607, A2 => n11206, B1 => n13639, B2 => 
                           n11203, C1 => n13575, C2 => n11200, ZN => n3739);
   U7182 : AOI221_X1 port map( B1 => n11146, B2 => n14276, C1 => n11143, C2 => 
                           n14468, A => n3748, ZN => n3742);
   U7183 : OAI222_X1 port map( A1 => n10118, A2 => n11140, B1 => n10117, B2 => 
                           n11137, C1 => n10119, C2 => n11134, ZN => n3748);
   U7184 : AOI221_X1 port map( B1 => n10948, B2 => n9517, C1 => n10945, C2 => 
                           n9549, A => n5131, ZN => n5125);
   U7185 : OAI222_X1 port map( A1 => n13606, A2 => n10942, B1 => n13638, B2 => 
                           n10939, C1 => n13574, C2 => n10936, ZN => n5131);
   U7186 : AOI221_X1 port map( B1 => n10882, B2 => n14275, C1 => n10879, C2 => 
                           n14467, A => n5140, ZN => n5134);
   U7187 : OAI222_X1 port map( A1 => n10086, A2 => n10876, B1 => n10085, B2 => 
                           n10873, C1 => n10087, C2 => n10870, ZN => n5140);
   U7188 : AOI221_X1 port map( B1 => n11212, B2 => n9517, C1 => n11209, C2 => 
                           n9549, A => n3698, ZN => n3692);
   U7189 : OAI222_X1 port map( A1 => n13606, A2 => n11206, B1 => n13638, B2 => 
                           n11203, C1 => n13574, C2 => n11200, ZN => n3698);
   U7190 : AOI221_X1 port map( B1 => n11146, B2 => n14275, C1 => n11143, C2 => 
                           n14467, A => n3707, ZN => n3701);
   U7191 : OAI222_X1 port map( A1 => n10086, A2 => n11140, B1 => n10085, B2 => 
                           n11137, C1 => n10087, C2 => n11134, ZN => n3707);
   U7192 : AOI221_X1 port map( B1 => n10948, B2 => n9518, C1 => n10945, C2 => 
                           n9550, A => n5090, ZN => n5084);
   U7193 : OAI222_X1 port map( A1 => n13605, A2 => n10942, B1 => n13637, B2 => 
                           n10939, C1 => n13573, C2 => n10936, ZN => n5090);
   U7194 : AOI221_X1 port map( B1 => n10882, B2 => n14274, C1 => n10879, C2 => 
                           n14466, A => n5099, ZN => n5093);
   U7195 : OAI222_X1 port map( A1 => n10054, A2 => n10876, B1 => n10053, B2 => 
                           n10873, C1 => n10055, C2 => n10870, ZN => n5099);
   U7196 : AOI221_X1 port map( B1 => n11212, B2 => n9518, C1 => n11209, C2 => 
                           n9550, A => n3657, ZN => n3651);
   U7197 : OAI222_X1 port map( A1 => n13605, A2 => n11206, B1 => n13637, B2 => 
                           n11203, C1 => n13573, C2 => n11200, ZN => n3657);
   U7198 : AOI221_X1 port map( B1 => n11146, B2 => n14274, C1 => n11143, C2 => 
                           n14466, A => n3666, ZN => n3660);
   U7199 : OAI222_X1 port map( A1 => n10054, A2 => n11140, B1 => n10053, B2 => 
                           n11137, C1 => n10055, C2 => n11134, ZN => n3666);
   U7200 : AOI221_X1 port map( B1 => n10948, B2 => n9519, C1 => n10945, C2 => 
                           n9551, A => n5049, ZN => n5043);
   U7201 : OAI222_X1 port map( A1 => n13604, A2 => n10942, B1 => n13636, B2 => 
                           n10939, C1 => n13572, C2 => n10936, ZN => n5049);
   U7202 : AOI221_X1 port map( B1 => n10882, B2 => n14273, C1 => n10879, C2 => 
                           n14465, A => n5058, ZN => n5052);
   U7203 : OAI222_X1 port map( A1 => n10022, A2 => n10876, B1 => n10021, B2 => 
                           n10873, C1 => n10023, C2 => n10870, ZN => n5058);
   U7204 : AOI221_X1 port map( B1 => n11212, B2 => n9519, C1 => n11209, C2 => 
                           n9551, A => n3616, ZN => n3610);
   U7205 : OAI222_X1 port map( A1 => n13604, A2 => n11206, B1 => n13636, B2 => 
                           n11203, C1 => n13572, C2 => n11200, ZN => n3616);
   U7206 : AOI221_X1 port map( B1 => n11146, B2 => n14273, C1 => n11143, C2 => 
                           n14465, A => n3625, ZN => n3619);
   U7207 : OAI222_X1 port map( A1 => n10022, A2 => n11140, B1 => n10021, B2 => 
                           n11137, C1 => n10023, C2 => n11134, ZN => n3625);
   U7208 : AOI221_X1 port map( B1 => n10948, B2 => n9520, C1 => n10945, C2 => 
                           n9552, A => n5008, ZN => n5002);
   U7209 : OAI222_X1 port map( A1 => n13603, A2 => n10942, B1 => n13635, B2 => 
                           n10939, C1 => n13571, C2 => n10936, ZN => n5008);
   U7210 : AOI221_X1 port map( B1 => n10882, B2 => n14272, C1 => n10879, C2 => 
                           n14464, A => n5017, ZN => n5011);
   U7211 : OAI222_X1 port map( A1 => n9660, A2 => n10876, B1 => n9659, B2 => 
                           n10873, C1 => n9661, C2 => n10870, ZN => n5017);
   U7212 : AOI221_X1 port map( B1 => n11212, B2 => n9520, C1 => n11209, C2 => 
                           n9552, A => n3575, ZN => n3569);
   U7213 : OAI222_X1 port map( A1 => n13603, A2 => n11206, B1 => n13635, B2 => 
                           n11203, C1 => n13571, C2 => n11200, ZN => n3575);
   U7214 : AOI221_X1 port map( B1 => n11146, B2 => n14272, C1 => n11143, C2 => 
                           n14464, A => n3584, ZN => n3578);
   U7215 : OAI222_X1 port map( A1 => n9660, A2 => n11140, B1 => n9659, B2 => 
                           n11137, C1 => n9661, C2 => n11134, ZN => n3584);
   U7216 : AOI221_X1 port map( B1 => n10948, B2 => n9521, C1 => n10945, C2 => 
                           n9553, A => n4967, ZN => n4961);
   U7217 : OAI222_X1 port map( A1 => n13602, A2 => n10942, B1 => n13634, B2 => 
                           n10939, C1 => n13570, C2 => n10936, ZN => n4967);
   U7218 : AOI221_X1 port map( B1 => n10882, B2 => n14271, C1 => n10879, C2 => 
                           n14463, A => n4976, ZN => n4970);
   U7219 : OAI222_X1 port map( A1 => n9628, A2 => n10876, B1 => n9627, B2 => 
                           n10873, C1 => n9629, C2 => n10870, ZN => n4976);
   U7220 : AOI221_X1 port map( B1 => n11212, B2 => n9521, C1 => n11209, C2 => 
                           n9553, A => n3534, ZN => n3528);
   U7221 : OAI222_X1 port map( A1 => n13602, A2 => n11206, B1 => n13634, B2 => 
                           n11203, C1 => n13570, C2 => n11200, ZN => n3534);
   U7222 : AOI221_X1 port map( B1 => n11146, B2 => n14271, C1 => n11143, C2 => 
                           n14463, A => n3543, ZN => n3537);
   U7223 : OAI222_X1 port map( A1 => n9628, A2 => n11140, B1 => n9627, B2 => 
                           n11137, C1 => n9629, C2 => n11134, ZN => n3543);
   U7224 : AOI221_X1 port map( B1 => n10948, B2 => n9522, C1 => n10945, C2 => 
                           n9554, A => n4926, ZN => n4920);
   U7225 : OAI222_X1 port map( A1 => n13601, A2 => n10942, B1 => n13633, B2 => 
                           n10939, C1 => n13569, C2 => n10936, ZN => n4926);
   U7226 : AOI221_X1 port map( B1 => n10882, B2 => n14270, C1 => n10879, C2 => 
                           n14462, A => n4935, ZN => n4929);
   U7227 : OAI222_X1 port map( A1 => n9596, A2 => n10876, B1 => n9595, B2 => 
                           n10873, C1 => n9597, C2 => n10870, ZN => n4935);
   U7228 : AOI221_X1 port map( B1 => n11212, B2 => n9522, C1 => n11209, C2 => 
                           n9554, A => n3493, ZN => n3487);
   U7229 : OAI222_X1 port map( A1 => n13601, A2 => n11206, B1 => n13633, B2 => 
                           n11203, C1 => n13569, C2 => n11200, ZN => n3493);
   U7230 : AOI221_X1 port map( B1 => n11146, B2 => n14270, C1 => n11143, C2 => 
                           n14462, A => n3502, ZN => n3496);
   U7231 : OAI222_X1 port map( A1 => n9596, A2 => n11140, B1 => n9595, B2 => 
                           n11137, C1 => n9597, C2 => n11134, ZN => n3502);
   U7232 : AOI221_X1 port map( B1 => n10948, B2 => n9523, C1 => n10945, C2 => 
                           n9555, A => n4885, ZN => n4879);
   U7233 : OAI222_X1 port map( A1 => n13600, A2 => n10942, B1 => n13632, B2 => 
                           n10939, C1 => n13568, C2 => n10936, ZN => n4885);
   U7234 : AOI221_X1 port map( B1 => n10882, B2 => n14269, C1 => n10879, C2 => 
                           n14461, A => n4894, ZN => n4888);
   U7235 : OAI222_X1 port map( A1 => n9262, A2 => n10876, B1 => n9261, B2 => 
                           n10873, C1 => n9263, C2 => n10870, ZN => n4894);
   U7236 : AOI221_X1 port map( B1 => n11212, B2 => n9523, C1 => n11209, C2 => 
                           n9555, A => n3452, ZN => n3446);
   U7237 : OAI222_X1 port map( A1 => n13600, A2 => n11206, B1 => n13632, B2 => 
                           n11203, C1 => n13568, C2 => n11200, ZN => n3452);
   U7238 : AOI221_X1 port map( B1 => n11146, B2 => n14269, C1 => n11143, C2 => 
                           n14461, A => n3461, ZN => n3455);
   U7239 : OAI222_X1 port map( A1 => n9262, A2 => n11140, B1 => n9261, B2 => 
                           n11137, C1 => n9263, C2 => n11134, ZN => n3461);
   U7240 : AOI221_X1 port map( B1 => n10948, B2 => n9524, C1 => n10945, C2 => 
                           n9556, A => n4844, ZN => n4838);
   U7241 : OAI222_X1 port map( A1 => n13599, A2 => n10942, B1 => n13631, B2 => 
                           n10939, C1 => n13567, C2 => n10936, ZN => n4844);
   U7242 : AOI221_X1 port map( B1 => n10882, B2 => n14268, C1 => n10879, C2 => 
                           n14460, A => n4853, ZN => n4847);
   U7243 : OAI222_X1 port map( A1 => n9198, A2 => n10876, B1 => n9197, B2 => 
                           n10873, C1 => n9199, C2 => n10870, ZN => n4853);
   U7244 : AOI221_X1 port map( B1 => n11212, B2 => n9524, C1 => n11209, C2 => 
                           n9556, A => n3411, ZN => n3405);
   U7245 : OAI222_X1 port map( A1 => n13599, A2 => n11206, B1 => n13631, B2 => 
                           n11203, C1 => n13567, C2 => n11200, ZN => n3411);
   U7246 : AOI221_X1 port map( B1 => n11146, B2 => n14268, C1 => n11143, C2 => 
                           n14460, A => n3420, ZN => n3414);
   U7247 : OAI222_X1 port map( A1 => n9198, A2 => n11140, B1 => n9197, B2 => 
                           n11137, C1 => n9199, C2 => n11134, ZN => n3420);
   U7248 : AOI221_X1 port map( B1 => n10948, B2 => n9525, C1 => n10945, C2 => 
                           n9557, A => n4803, ZN => n4797);
   U7249 : OAI222_X1 port map( A1 => n13598, A2 => n10942, B1 => n13630, B2 => 
                           n10939, C1 => n13566, C2 => n10936, ZN => n4803);
   U7250 : AOI221_X1 port map( B1 => n10882, B2 => n14267, C1 => n10879, C2 => 
                           n14459, A => n4812, ZN => n4806);
   U7251 : OAI222_X1 port map( A1 => n9166, A2 => n10876, B1 => n9165, B2 => 
                           n10873, C1 => n9167, C2 => n10870, ZN => n4812);
   U7252 : AOI221_X1 port map( B1 => n11212, B2 => n9525, C1 => n11209, C2 => 
                           n9557, A => n3370, ZN => n3364);
   U7253 : OAI222_X1 port map( A1 => n13598, A2 => n11206, B1 => n13630, B2 => 
                           n11203, C1 => n13566, C2 => n11200, ZN => n3370);
   U7254 : AOI221_X1 port map( B1 => n11146, B2 => n14267, C1 => n11143, C2 => 
                           n14459, A => n3379, ZN => n3373);
   U7255 : OAI222_X1 port map( A1 => n9166, A2 => n11140, B1 => n9165, B2 => 
                           n11137, C1 => n9167, C2 => n11134, ZN => n3379);
   U7256 : AOI221_X1 port map( B1 => n10948, B2 => n9526, C1 => n10945, C2 => 
                           n9558, A => n4762, ZN => n4756);
   U7257 : OAI222_X1 port map( A1 => n13597, A2 => n10942, B1 => n13629, B2 => 
                           n10939, C1 => n13565, C2 => n10936, ZN => n4762);
   U7258 : AOI221_X1 port map( B1 => n10882, B2 => n14266, C1 => n10879, C2 => 
                           n14458, A => n4771, ZN => n4765);
   U7259 : OAI222_X1 port map( A1 => n9134, A2 => n10876, B1 => n6315, B2 => 
                           n10873, C1 => n9135, C2 => n10870, ZN => n4771);
   U7260 : AOI221_X1 port map( B1 => n11212, B2 => n9526, C1 => n11209, C2 => 
                           n9558, A => n3329, ZN => n3323);
   U7261 : OAI222_X1 port map( A1 => n13597, A2 => n11206, B1 => n13629, B2 => 
                           n11203, C1 => n13565, C2 => n11200, ZN => n3329);
   U7262 : AOI221_X1 port map( B1 => n11146, B2 => n14266, C1 => n11143, C2 => 
                           n14458, A => n3338, ZN => n3332);
   U7263 : OAI222_X1 port map( A1 => n9134, A2 => n11140, B1 => n6315, B2 => 
                           n11137, C1 => n9135, C2 => n11134, ZN => n3338);
   U7264 : AOI221_X1 port map( B1 => n10948, B2 => n9527, C1 => n10945, C2 => 
                           n9559, A => n4721, ZN => n4715);
   U7265 : OAI222_X1 port map( A1 => n13596, A2 => n10942, B1 => n13628, B2 => 
                           n10939, C1 => n13564, C2 => n10936, ZN => n4721);
   U7266 : AOI221_X1 port map( B1 => n10882, B2 => n14265, C1 => n10879, C2 => 
                           n14457, A => n4730, ZN => n4724);
   U7267 : OAI222_X1 port map( A1 => n5999, A2 => n10876, B1 => n5998, B2 => 
                           n10873, C1 => n6000, C2 => n10870, ZN => n4730);
   U7268 : AOI221_X1 port map( B1 => n11212, B2 => n9527, C1 => n11209, C2 => 
                           n9559, A => n3288, ZN => n3282);
   U7269 : OAI222_X1 port map( A1 => n13596, A2 => n11206, B1 => n13628, B2 => 
                           n11203, C1 => n13564, C2 => n11200, ZN => n3288);
   U7270 : AOI221_X1 port map( B1 => n11146, B2 => n14265, C1 => n11143, C2 => 
                           n14457, A => n3297, ZN => n3291);
   U7271 : OAI222_X1 port map( A1 => n5999, A2 => n11140, B1 => n5998, B2 => 
                           n11137, C1 => n6000, C2 => n11134, ZN => n3297);
   U7272 : AOI221_X1 port map( B1 => n10949, B2 => n9528, C1 => n10946, C2 => 
                           n9560, A => n4680, ZN => n4674);
   U7273 : OAI222_X1 port map( A1 => n13595, A2 => n10943, B1 => n13627, B2 => 
                           n10940, C1 => n13563, C2 => n10937, ZN => n4680);
   U7274 : AOI221_X1 port map( B1 => n10883, B2 => n14264, C1 => n10880, C2 => 
                           n14456, A => n4689, ZN => n4683);
   U7275 : OAI222_X1 port map( A1 => n5935, A2 => n10877, B1 => n5934, B2 => 
                           n10874, C1 => n5936, C2 => n10871, ZN => n4689);
   U7276 : AOI221_X1 port map( B1 => n11213, B2 => n9528, C1 => n11210, C2 => 
                           n9560, A => n3247, ZN => n3241);
   U7277 : OAI222_X1 port map( A1 => n13595, A2 => n11207, B1 => n13627, B2 => 
                           n11204, C1 => n13563, C2 => n11201, ZN => n3247);
   U7278 : AOI221_X1 port map( B1 => n11147, B2 => n14264, C1 => n11144, C2 => 
                           n14456, A => n3256, ZN => n3250);
   U7279 : OAI222_X1 port map( A1 => n5935, A2 => n11141, B1 => n5934, B2 => 
                           n11138, C1 => n5936, C2 => n11135, ZN => n3256);
   U7280 : AOI221_X1 port map( B1 => n10949, B2 => n9529, C1 => n10946, C2 => 
                           n9561, A => n4639, ZN => n4633);
   U7281 : OAI222_X1 port map( A1 => n13594, A2 => n10943, B1 => n13626, B2 => 
                           n10940, C1 => n13562, C2 => n10937, ZN => n4639);
   U7282 : AOI221_X1 port map( B1 => n10883, B2 => n14263, C1 => n10880, C2 => 
                           n14455, A => n4648, ZN => n4642);
   U7283 : OAI222_X1 port map( A1 => n5903, A2 => n10877, B1 => n5902, B2 => 
                           n10874, C1 => n5904, C2 => n10871, ZN => n4648);
   U7284 : AOI221_X1 port map( B1 => n11213, B2 => n9529, C1 => n11210, C2 => 
                           n9561, A => n3206, ZN => n3200);
   U7285 : OAI222_X1 port map( A1 => n13594, A2 => n11207, B1 => n13626, B2 => 
                           n11204, C1 => n13562, C2 => n11201, ZN => n3206);
   U7286 : AOI221_X1 port map( B1 => n11147, B2 => n14263, C1 => n11144, C2 => 
                           n14455, A => n3215, ZN => n3209);
   U7287 : OAI222_X1 port map( A1 => n5903, A2 => n11141, B1 => n5902, B2 => 
                           n11138, C1 => n5904, C2 => n11135, ZN => n3215);
   U7288 : AOI221_X1 port map( B1 => n10949, B2 => n9530, C1 => n10946, C2 => 
                           n9562, A => n4598, ZN => n4592);
   U7289 : OAI222_X1 port map( A1 => n13593, A2 => n10943, B1 => n13625, B2 => 
                           n10940, C1 => n13561, C2 => n10937, ZN => n4598);
   U7290 : AOI221_X1 port map( B1 => n10883, B2 => n14262, C1 => n10880, C2 => 
                           n14454, A => n4607, ZN => n4601);
   U7291 : OAI222_X1 port map( A1 => n5871, A2 => n10877, B1 => n5870, B2 => 
                           n10874, C1 => n5872, C2 => n10871, ZN => n4607);
   U7292 : AOI221_X1 port map( B1 => n11213, B2 => n9530, C1 => n11210, C2 => 
                           n9562, A => n3165, ZN => n3159);
   U7293 : OAI222_X1 port map( A1 => n13593, A2 => n11207, B1 => n13625, B2 => 
                           n11204, C1 => n13561, C2 => n11201, ZN => n3165);
   U7294 : AOI221_X1 port map( B1 => n11147, B2 => n14262, C1 => n11144, C2 => 
                           n14454, A => n3174, ZN => n3168);
   U7295 : OAI222_X1 port map( A1 => n5871, A2 => n11141, B1 => n5870, B2 => 
                           n11138, C1 => n5872, C2 => n11135, ZN => n3174);
   U7296 : AOI221_X1 port map( B1 => n10949, B2 => n9531, C1 => n10946, C2 => 
                           n9563, A => n4557, ZN => n4551);
   U7297 : OAI222_X1 port map( A1 => n13592, A2 => n10943, B1 => n13624, B2 => 
                           n10940, C1 => n13560, C2 => n10937, ZN => n4557);
   U7298 : AOI221_X1 port map( B1 => n10883, B2 => n14261, C1 => n10880, C2 => 
                           n14453, A => n4566, ZN => n4560);
   U7299 : OAI222_X1 port map( A1 => n5839, A2 => n10877, B1 => n5838, B2 => 
                           n10874, C1 => n5840, C2 => n10871, ZN => n4566);
   U7300 : AOI221_X1 port map( B1 => n11213, B2 => n9531, C1 => n11210, C2 => 
                           n9563, A => n3124, ZN => n3118);
   U7301 : OAI222_X1 port map( A1 => n13592, A2 => n11207, B1 => n13624, B2 => 
                           n11204, C1 => n13560, C2 => n11201, ZN => n3124);
   U7302 : AOI221_X1 port map( B1 => n11147, B2 => n14261, C1 => n11144, C2 => 
                           n14453, A => n3133, ZN => n3127);
   U7303 : OAI222_X1 port map( A1 => n5839, A2 => n11141, B1 => n5838, B2 => 
                           n11138, C1 => n5840, C2 => n11135, ZN => n3133);
   U7304 : AOI221_X1 port map( B1 => n10949, B2 => n9532, C1 => n10946, C2 => 
                           n9564, A => n4516, ZN => n4510);
   U7305 : OAI222_X1 port map( A1 => n13591, A2 => n10943, B1 => n13623, B2 => 
                           n10940, C1 => n13559, C2 => n10937, ZN => n4516);
   U7306 : AOI221_X1 port map( B1 => n10883, B2 => n14260, C1 => n10880, C2 => 
                           n14452, A => n4525, ZN => n4519);
   U7307 : OAI222_X1 port map( A1 => n5807, A2 => n10877, B1 => n5806, B2 => 
                           n10874, C1 => n5808, C2 => n10871, ZN => n4525);
   U7308 : AOI221_X1 port map( B1 => n11213, B2 => n9532, C1 => n11210, C2 => 
                           n9564, A => n3083, ZN => n3077);
   U7309 : OAI222_X1 port map( A1 => n13591, A2 => n11207, B1 => n13623, B2 => 
                           n11204, C1 => n13559, C2 => n11201, ZN => n3083);
   U7310 : AOI221_X1 port map( B1 => n11147, B2 => n14260, C1 => n11144, C2 => 
                           n14452, A => n3092, ZN => n3086);
   U7311 : OAI222_X1 port map( A1 => n5807, A2 => n11141, B1 => n5806, B2 => 
                           n11138, C1 => n5808, C2 => n11135, ZN => n3092);
   U7312 : AOI221_X1 port map( B1 => n10949, B2 => n9533, C1 => n10946, C2 => 
                           n9565, A => n4475, ZN => n4469);
   U7313 : OAI222_X1 port map( A1 => n13590, A2 => n10943, B1 => n13622, B2 => 
                           n10940, C1 => n13558, C2 => n10937, ZN => n4475);
   U7314 : AOI221_X1 port map( B1 => n10883, B2 => n14259, C1 => n10880, C2 => 
                           n14451, A => n4484, ZN => n4478);
   U7315 : OAI222_X1 port map( A1 => n5775, A2 => n10877, B1 => n5774, B2 => 
                           n10874, C1 => n5776, C2 => n10871, ZN => n4484);
   U7316 : AOI221_X1 port map( B1 => n11213, B2 => n9533, C1 => n11210, C2 => 
                           n9565, A => n3042, ZN => n3036);
   U7317 : OAI222_X1 port map( A1 => n13590, A2 => n11207, B1 => n13622, B2 => 
                           n11204, C1 => n13558, C2 => n11201, ZN => n3042);
   U7318 : AOI221_X1 port map( B1 => n11147, B2 => n14259, C1 => n11144, C2 => 
                           n14451, A => n3051, ZN => n3045);
   U7319 : OAI222_X1 port map( A1 => n5775, A2 => n11141, B1 => n5774, B2 => 
                           n11138, C1 => n5776, C2 => n11135, ZN => n3051);
   U7320 : AOI221_X1 port map( B1 => n10949, B2 => n9534, C1 => n10946, C2 => 
                           n9566, A => n4434, ZN => n4428);
   U7321 : OAI222_X1 port map( A1 => n13589, A2 => n10943, B1 => n13621, B2 => 
                           n10940, C1 => n13557, C2 => n10937, ZN => n4434);
   U7322 : AOI221_X1 port map( B1 => n10883, B2 => n14258, C1 => n10880, C2 => 
                           n14450, A => n4443, ZN => n4437);
   U7323 : OAI222_X1 port map( A1 => n5743, A2 => n10877, B1 => n5742, B2 => 
                           n10874, C1 => n5744, C2 => n10871, ZN => n4443);
   U7324 : AOI221_X1 port map( B1 => n11213, B2 => n9534, C1 => n11210, C2 => 
                           n9566, A => n3001, ZN => n2995);
   U7325 : OAI222_X1 port map( A1 => n13589, A2 => n11207, B1 => n13621, B2 => 
                           n11204, C1 => n13557, C2 => n11201, ZN => n3001);
   U7326 : AOI221_X1 port map( B1 => n11147, B2 => n14258, C1 => n11144, C2 => 
                           n14450, A => n3010, ZN => n3004);
   U7327 : OAI222_X1 port map( A1 => n5743, A2 => n11141, B1 => n5742, B2 => 
                           n11138, C1 => n5744, C2 => n11135, ZN => n3010);
   U7328 : AOI221_X1 port map( B1 => n10949, B2 => n9535, C1 => n10946, C2 => 
                           n9567, A => n4362, ZN => n4343);
   U7329 : OAI222_X1 port map( A1 => n13588, A2 => n10943, B1 => n13620, B2 => 
                           n10940, C1 => n13556, C2 => n10937, ZN => n4362);
   U7330 : AOI221_X1 port map( B1 => n10883, B2 => n14257, C1 => n10880, C2 => 
                           n14449, A => n4393, ZN => n4374);
   U7331 : OAI222_X1 port map( A1 => n5711, A2 => n10877, B1 => n5710, B2 => 
                           n10874, C1 => n5712, C2 => n10871, ZN => n4393);
   U7332 : AOI221_X1 port map( B1 => n11213, B2 => n9535, C1 => n11210, C2 => 
                           n9567, A => n2926, ZN => n2875);
   U7333 : OAI222_X1 port map( A1 => n13588, A2 => n11207, B1 => n13620, B2 => 
                           n11204, C1 => n13556, C2 => n11201, ZN => n2926);
   U7334 : AOI221_X1 port map( B1 => n11147, B2 => n14257, C1 => n11144, C2 => 
                           n14449, A => n2960, ZN => n2941);
   U7335 : OAI222_X1 port map( A1 => n5711, A2 => n11141, B1 => n5710, B2 => 
                           n11138, C1 => n5712, C2 => n11135, ZN => n2960);
   U7336 : NOR2_X1 port map( A1 => ADD_RD1(0), A2 => N8434, ZN => n5654);
   U7337 : NOR2_X1 port map( A1 => ADD_RD2(0), A2 => N8578, ZN => n4221);
   U7338 : OAI22_X1 port map( A1 => n1955, A2 => n11114, B1 => n227, B2 => 
                           n11111, ZN => n4661);
   U7339 : OAI22_X1 port map( A1 => n5986, A2 => n11048, B1 => n5985, B2 => 
                           n11045, ZN => n4670);
   U7340 : OAI22_X1 port map( A1 => n1955, A2 => n11378, B1 => n227, B2 => 
                           n11375, ZN => n3228);
   U7341 : OAI22_X1 port map( A1 => n5986, A2 => n11312, B1 => n5985, B2 => 
                           n11309, ZN => n3237);
   U7342 : OAI22_X1 port map( A1 => n1943, A2 => n11114, B1 => n215, B2 => 
                           n11111, ZN => n4620);
   U7343 : OAI22_X1 port map( A1 => n5922, A2 => n11048, B1 => n5921, B2 => 
                           n11045, ZN => n4629);
   U7344 : OAI22_X1 port map( A1 => n1943, A2 => n11378, B1 => n215, B2 => 
                           n11375, ZN => n3187);
   U7345 : OAI22_X1 port map( A1 => n5922, A2 => n11312, B1 => n5921, B2 => 
                           n11309, ZN => n3196);
   U7346 : OAI22_X1 port map( A1 => n1931, A2 => n11114, B1 => n203, B2 => 
                           n11111, ZN => n4579);
   U7347 : OAI22_X1 port map( A1 => n5890, A2 => n11048, B1 => n5889, B2 => 
                           n11045, ZN => n4588);
   U7348 : OAI22_X1 port map( A1 => n1931, A2 => n11378, B1 => n203, B2 => 
                           n11375, ZN => n3146);
   U7349 : OAI22_X1 port map( A1 => n5890, A2 => n11312, B1 => n5889, B2 => 
                           n11309, ZN => n3155);
   U7350 : OAI22_X1 port map( A1 => n1919, A2 => n11114, B1 => n191, B2 => 
                           n11111, ZN => n4538);
   U7351 : OAI22_X1 port map( A1 => n5858, A2 => n11048, B1 => n5857, B2 => 
                           n11045, ZN => n4547);
   U7352 : OAI22_X1 port map( A1 => n1919, A2 => n11378, B1 => n191, B2 => 
                           n11375, ZN => n3105);
   U7353 : OAI22_X1 port map( A1 => n5858, A2 => n11312, B1 => n5857, B2 => 
                           n11309, ZN => n3114);
   U7354 : OAI22_X1 port map( A1 => n1907, A2 => n11114, B1 => n179, B2 => 
                           n11111, ZN => n4497);
   U7355 : OAI22_X1 port map( A1 => n5826, A2 => n11048, B1 => n5825, B2 => 
                           n11045, ZN => n4506);
   U7356 : OAI22_X1 port map( A1 => n1907, A2 => n11378, B1 => n179, B2 => 
                           n11375, ZN => n3064);
   U7357 : OAI22_X1 port map( A1 => n5826, A2 => n11312, B1 => n5825, B2 => 
                           n11309, ZN => n3073);
   U7358 : OAI22_X1 port map( A1 => n1895, A2 => n11114, B1 => n167, B2 => 
                           n11111, ZN => n4456);
   U7359 : OAI22_X1 port map( A1 => n5794, A2 => n11048, B1 => n5793, B2 => 
                           n11045, ZN => n4465);
   U7360 : OAI22_X1 port map( A1 => n1895, A2 => n11378, B1 => n167, B2 => 
                           n11375, ZN => n3023);
   U7361 : OAI22_X1 port map( A1 => n5794, A2 => n11312, B1 => n5793, B2 => 
                           n11309, ZN => n3032);
   U7362 : OAI22_X1 port map( A1 => n1883, A2 => n11114, B1 => n155, B2 => 
                           n11111, ZN => n4415);
   U7363 : OAI22_X1 port map( A1 => n5762, A2 => n11048, B1 => n5761, B2 => 
                           n11045, ZN => n4424);
   U7364 : OAI22_X1 port map( A1 => n1883, A2 => n11378, B1 => n155, B2 => 
                           n11375, ZN => n2982);
   U7365 : OAI22_X1 port map( A1 => n5762, A2 => n11312, B1 => n5761, B2 => 
                           n11309, ZN => n2991);
   U7366 : OAI22_X1 port map( A1 => n1871, A2 => n11114, B1 => n143, B2 => 
                           n11111, ZN => n4286);
   U7367 : OAI22_X1 port map( A1 => n5730, A2 => n11048, B1 => n5729, B2 => 
                           n11045, ZN => n4317);
   U7368 : OAI22_X1 port map( A1 => n1871, A2 => n11378, B1 => n143, B2 => 
                           n11375, ZN => n2786);
   U7369 : OAI22_X1 port map( A1 => n5730, A2 => n11312, B1 => n5729, B2 => 
                           n11309, ZN => n2817);
   U7370 : OAI22_X1 port map( A1 => n2339, A2 => n11112, B1 => n515, B2 => 
                           n11109, ZN => n5645);
   U7371 : OAI22_X1 port map( A1 => n10529, A2 => n11046, B1 => n10528, B2 => 
                           n11043, ZN => n5673);
   U7372 : OAI22_X1 port map( A1 => n2339, A2 => n11376, B1 => n515, B2 => 
                           n11373, ZN => n4212);
   U7373 : OAI22_X1 port map( A1 => n10529, A2 => n11310, B1 => n10528, B2 => 
                           n11307, ZN => n4240);
   U7374 : OAI22_X1 port map( A1 => n2327, A2 => n11112, B1 => n503, B2 => 
                           n11109, ZN => n5604);
   U7375 : OAI22_X1 port map( A1 => n10497, A2 => n11046, B1 => n10496, B2 => 
                           n11043, ZN => n5613);
   U7376 : OAI22_X1 port map( A1 => n2327, A2 => n11376, B1 => n503, B2 => 
                           n11373, ZN => n4171);
   U7377 : OAI22_X1 port map( A1 => n10497, A2 => n11310, B1 => n10496, B2 => 
                           n11307, ZN => n4180);
   U7378 : OAI22_X1 port map( A1 => n2315, A2 => n11112, B1 => n491, B2 => 
                           n11109, ZN => n5563);
   U7379 : OAI22_X1 port map( A1 => n10465, A2 => n11046, B1 => n10464, B2 => 
                           n11043, ZN => n5572);
   U7380 : OAI22_X1 port map( A1 => n2315, A2 => n11376, B1 => n491, B2 => 
                           n11373, ZN => n4130);
   U7381 : OAI22_X1 port map( A1 => n10465, A2 => n11310, B1 => n10464, B2 => 
                           n11307, ZN => n4139);
   U7382 : OAI22_X1 port map( A1 => n2303, A2 => n11112, B1 => n479, B2 => 
                           n11109, ZN => n5522);
   U7383 : OAI22_X1 port map( A1 => n10433, A2 => n11046, B1 => n10432, B2 => 
                           n11043, ZN => n5531);
   U7384 : OAI22_X1 port map( A1 => n2303, A2 => n11376, B1 => n479, B2 => 
                           n11373, ZN => n4089);
   U7385 : OAI22_X1 port map( A1 => n10433, A2 => n11310, B1 => n10432, B2 => 
                           n11307, ZN => n4098);
   U7386 : OAI22_X1 port map( A1 => n2291, A2 => n11112, B1 => n467, B2 => 
                           n11109, ZN => n5481);
   U7387 : OAI22_X1 port map( A1 => n10401, A2 => n11046, B1 => n10400, B2 => 
                           n11043, ZN => n5490);
   U7388 : OAI22_X1 port map( A1 => n2291, A2 => n11376, B1 => n467, B2 => 
                           n11373, ZN => n4048);
   U7389 : OAI22_X1 port map( A1 => n10401, A2 => n11310, B1 => n10400, B2 => 
                           n11307, ZN => n4057);
   U7390 : OAI22_X1 port map( A1 => n2279, A2 => n11112, B1 => n455, B2 => 
                           n11109, ZN => n5440);
   U7391 : OAI22_X1 port map( A1 => n10366, A2 => n11046, B1 => n10365, B2 => 
                           n11043, ZN => n5449);
   U7392 : OAI22_X1 port map( A1 => n2279, A2 => n11376, B1 => n455, B2 => 
                           n11373, ZN => n4007);
   U7393 : OAI22_X1 port map( A1 => n10366, A2 => n11310, B1 => n10365, B2 => 
                           n11307, ZN => n4016);
   U7394 : OAI22_X1 port map( A1 => n2267, A2 => n11112, B1 => n443, B2 => 
                           n11109, ZN => n5399);
   U7395 : OAI22_X1 port map( A1 => n10334, A2 => n11046, B1 => n10333, B2 => 
                           n11043, ZN => n5408);
   U7396 : OAI22_X1 port map( A1 => n2267, A2 => n11376, B1 => n443, B2 => 
                           n11373, ZN => n3966);
   U7397 : OAI22_X1 port map( A1 => n10334, A2 => n11310, B1 => n10333, B2 => 
                           n11307, ZN => n3975);
   U7398 : OAI22_X1 port map( A1 => n2255, A2 => n11112, B1 => n431, B2 => 
                           n11109, ZN => n5358);
   U7399 : OAI22_X1 port map( A1 => n10299, A2 => n11046, B1 => n10298, B2 => 
                           n11043, ZN => n5367);
   U7400 : OAI22_X1 port map( A1 => n2255, A2 => n11376, B1 => n431, B2 => 
                           n11373, ZN => n3925);
   U7401 : OAI22_X1 port map( A1 => n10299, A2 => n11310, B1 => n10298, B2 => 
                           n11307, ZN => n3934);
   U7402 : OAI22_X1 port map( A1 => n2243, A2 => n11112, B1 => n419, B2 => 
                           n11109, ZN => n5317);
   U7403 : OAI22_X1 port map( A1 => n10267, A2 => n11046, B1 => n10266, B2 => 
                           n11043, ZN => n5326);
   U7404 : OAI22_X1 port map( A1 => n2243, A2 => n11376, B1 => n419, B2 => 
                           n11373, ZN => n3884);
   U7405 : OAI22_X1 port map( A1 => n10267, A2 => n11310, B1 => n10266, B2 => 
                           n11307, ZN => n3893);
   U7406 : OAI22_X1 port map( A1 => n2231, A2 => n11112, B1 => n407, B2 => 
                           n11109, ZN => n5276);
   U7407 : OAI22_X1 port map( A1 => n10235, A2 => n11046, B1 => n10234, B2 => 
                           n11043, ZN => n5285);
   U7408 : OAI22_X1 port map( A1 => n2231, A2 => n11376, B1 => n407, B2 => 
                           n11373, ZN => n3843);
   U7409 : OAI22_X1 port map( A1 => n10235, A2 => n11310, B1 => n10234, B2 => 
                           n11307, ZN => n3852);
   U7410 : OAI22_X1 port map( A1 => n2219, A2 => n11112, B1 => n395, B2 => 
                           n11109, ZN => n5235);
   U7411 : OAI22_X1 port map( A1 => n10201, A2 => n11046, B1 => n10200, B2 => 
                           n11043, ZN => n5244);
   U7412 : OAI22_X1 port map( A1 => n2219, A2 => n11376, B1 => n395, B2 => 
                           n11373, ZN => n3802);
   U7413 : OAI22_X1 port map( A1 => n10201, A2 => n11310, B1 => n10200, B2 => 
                           n11307, ZN => n3811);
   U7414 : OAI22_X1 port map( A1 => n2175, A2 => n11112, B1 => n383, B2 => 
                           n11109, ZN => n5194);
   U7415 : OAI22_X1 port map( A1 => n10169, A2 => n11046, B1 => n10168, B2 => 
                           n11043, ZN => n5203);
   U7416 : OAI22_X1 port map( A1 => n2175, A2 => n11376, B1 => n383, B2 => 
                           n11373, ZN => n3761);
   U7417 : OAI22_X1 port map( A1 => n10169, A2 => n11310, B1 => n10168, B2 => 
                           n11307, ZN => n3770);
   U7418 : OAI22_X1 port map( A1 => n2163, A2 => n11113, B1 => n371, B2 => 
                           n11110, ZN => n5153);
   U7419 : OAI22_X1 port map( A1 => n10137, A2 => n11047, B1 => n10136, B2 => 
                           n11044, ZN => n5162);
   U7420 : OAI22_X1 port map( A1 => n2163, A2 => n11377, B1 => n371, B2 => 
                           n11374, ZN => n3720);
   U7421 : OAI22_X1 port map( A1 => n10137, A2 => n11311, B1 => n10136, B2 => 
                           n11308, ZN => n3729);
   U7422 : OAI22_X1 port map( A1 => n2151, A2 => n11113, B1 => n359, B2 => 
                           n11110, ZN => n5112);
   U7423 : OAI22_X1 port map( A1 => n10105, A2 => n11047, B1 => n10104, B2 => 
                           n11044, ZN => n5121);
   U7424 : OAI22_X1 port map( A1 => n2151, A2 => n11377, B1 => n359, B2 => 
                           n11374, ZN => n3679);
   U7425 : OAI22_X1 port map( A1 => n10105, A2 => n11311, B1 => n10104, B2 => 
                           n11308, ZN => n3688);
   U7426 : OAI22_X1 port map( A1 => n2107, A2 => n11113, B1 => n347, B2 => 
                           n11110, ZN => n5071);
   U7427 : OAI22_X1 port map( A1 => n10073, A2 => n11047, B1 => n10072, B2 => 
                           n11044, ZN => n5080);
   U7428 : OAI22_X1 port map( A1 => n2107, A2 => n11377, B1 => n347, B2 => 
                           n11374, ZN => n3638);
   U7429 : OAI22_X1 port map( A1 => n10073, A2 => n11311, B1 => n10072, B2 => 
                           n11308, ZN => n3647);
   U7430 : OAI22_X1 port map( A1 => n2095, A2 => n11113, B1 => n335, B2 => 
                           n11110, ZN => n5030);
   U7431 : OAI22_X1 port map( A1 => n10041, A2 => n11047, B1 => n10040, B2 => 
                           n11044, ZN => n5039);
   U7432 : OAI22_X1 port map( A1 => n2095, A2 => n11377, B1 => n335, B2 => 
                           n11374, ZN => n3597);
   U7433 : OAI22_X1 port map( A1 => n10041, A2 => n11311, B1 => n10040, B2 => 
                           n11308, ZN => n3606);
   U7434 : OAI22_X1 port map( A1 => n2083, A2 => n11113, B1 => n323, B2 => 
                           n11110, ZN => n4989);
   U7435 : OAI22_X1 port map( A1 => n10009, A2 => n11047, B1 => n10008, B2 => 
                           n11044, ZN => n4998);
   U7436 : OAI22_X1 port map( A1 => n2083, A2 => n11377, B1 => n323, B2 => 
                           n11374, ZN => n3556);
   U7437 : OAI22_X1 port map( A1 => n10009, A2 => n11311, B1 => n10008, B2 => 
                           n11308, ZN => n3565);
   U7438 : OAI22_X1 port map( A1 => n2039, A2 => n11113, B1 => n311, B2 => 
                           n11110, ZN => n4948);
   U7439 : OAI22_X1 port map( A1 => n9647, A2 => n11047, B1 => n9646, B2 => 
                           n11044, ZN => n4957);
   U7440 : OAI22_X1 port map( A1 => n2039, A2 => n11377, B1 => n311, B2 => 
                           n11374, ZN => n3515);
   U7441 : OAI22_X1 port map( A1 => n9647, A2 => n11311, B1 => n9646, B2 => 
                           n11308, ZN => n3524);
   U7442 : OAI22_X1 port map( A1 => n2027, A2 => n11113, B1 => n299, B2 => 
                           n11110, ZN => n4907);
   U7443 : OAI22_X1 port map( A1 => n9615, A2 => n11047, B1 => n9614, B2 => 
                           n11044, ZN => n4916);
   U7444 : OAI22_X1 port map( A1 => n2027, A2 => n11377, B1 => n299, B2 => 
                           n11374, ZN => n3474);
   U7445 : OAI22_X1 port map( A1 => n9615, A2 => n11311, B1 => n9614, B2 => 
                           n11308, ZN => n3483);
   U7446 : OAI22_X1 port map( A1 => n2015, A2 => n11113, B1 => n287, B2 => 
                           n11110, ZN => n4866);
   U7447 : OAI22_X1 port map( A1 => n9583, A2 => n11047, B1 => n9582, B2 => 
                           n11044, ZN => n4875);
   U7448 : OAI22_X1 port map( A1 => n2015, A2 => n11377, B1 => n287, B2 => 
                           n11374, ZN => n3433);
   U7449 : OAI22_X1 port map( A1 => n9583, A2 => n11311, B1 => n9582, B2 => 
                           n11308, ZN => n3442);
   U7450 : OAI22_X1 port map( A1 => n2003, A2 => n11113, B1 => n275, B2 => 
                           n11110, ZN => n4825);
   U7451 : OAI22_X1 port map( A1 => n9249, A2 => n11047, B1 => n9248, B2 => 
                           n11044, ZN => n4834);
   U7452 : OAI22_X1 port map( A1 => n2003, A2 => n11377, B1 => n275, B2 => 
                           n11374, ZN => n3392);
   U7453 : OAI22_X1 port map( A1 => n9249, A2 => n11311, B1 => n9248, B2 => 
                           n11308, ZN => n3401);
   U7454 : OAI22_X1 port map( A1 => n1991, A2 => n11113, B1 => n263, B2 => 
                           n11110, ZN => n4784);
   U7455 : OAI22_X1 port map( A1 => n9185, A2 => n11047, B1 => n9184, B2 => 
                           n11044, ZN => n4793);
   U7456 : OAI22_X1 port map( A1 => n1991, A2 => n11377, B1 => n263, B2 => 
                           n11374, ZN => n3351);
   U7457 : OAI22_X1 port map( A1 => n9185, A2 => n11311, B1 => n9184, B2 => 
                           n11308, ZN => n3360);
   U7458 : OAI22_X1 port map( A1 => n1979, A2 => n11113, B1 => n251, B2 => 
                           n11110, ZN => n4743);
   U7459 : OAI22_X1 port map( A1 => n9153, A2 => n11047, B1 => n9152, B2 => 
                           n11044, ZN => n4752);
   U7460 : OAI22_X1 port map( A1 => n1979, A2 => n11377, B1 => n251, B2 => 
                           n11374, ZN => n3310);
   U7461 : OAI22_X1 port map( A1 => n9153, A2 => n11311, B1 => n9152, B2 => 
                           n11308, ZN => n3319);
   U7462 : OAI22_X1 port map( A1 => n1967, A2 => n11113, B1 => n239, B2 => 
                           n11110, ZN => n4702);
   U7463 : OAI22_X1 port map( A1 => n6303, A2 => n11047, B1 => n6302, B2 => 
                           n11044, ZN => n4711);
   U7464 : OAI22_X1 port map( A1 => n1967, A2 => n11377, B1 => n239, B2 => 
                           n11374, ZN => n3269);
   U7465 : OAI22_X1 port map( A1 => n6303, A2 => n11311, B1 => n6302, B2 => 
                           n11308, ZN => n3278);
   U7466 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n5651);
   U7467 : AND2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n4218);
   U7468 : AND2_X1 port map( A1 => ADD_RD1(2), A2 => n14513, ZN => n5650);
   U7469 : AND2_X1 port map( A1 => ADD_RD2(2), A2 => n14515, ZN => n4217);
   U7470 : NOR2_X1 port map( A1 => n12772, A2 => ADD_RD1(0), ZN => n5703);
   U7471 : NOR2_X1 port map( A1 => n12776, A2 => ADD_RD2(0), ZN => n4270);
   U7472 : XNOR2_X1 port map( A => U3_U97_Z_6, B => r472_n4, ZN => N2173);
   U7473 : NAND2_X1 port map( A1 => U3_U97_Z_5, A2 => r472_carry_5_port, ZN => 
                           r472_n4);
   U7474 : NOR2_X1 port map( A1 => n2935, A2 => r472_B_3_port, ZN => U3_U97_Z_6
                           );
   U7475 : NOR2_X1 port map( A1 => n12735, A2 => ADD_WR(0), ZN => n2719);
   U7476 : NOR2_X1 port map( A1 => n12736, A2 => ADD_WR(1), ZN => n2721);
   U7477 : NOR2_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), ZN => n2723);
   U7478 : NOR2_X1 port map( A1 => ADD_WR(2), A2 => N2170, ZN => n2735);
   U7479 : NAND4_X1 port map( A1 => n5666, A2 => n5667, A3 => n5668, A4 => 
                           n5669, ZN => n5636);
   U7480 : AOI221_X1 port map( B1 => n11013, B2 => n9952, C1 => n11010, C2 => 
                           n9984, A => n5677, ZN => n5668);
   U7481 : NOR4_X1 port map( A1 => n5670, A2 => n5671, A3 => n5672, A4 => n5673
                           , ZN => n5669);
   U7482 : AOI222_X1 port map( A1 => n10989, A2 => n9824, B1 => n10986, B2 => 
                           n9760, C1 => n10983, C2 => n9792, ZN => n5666);
   U7483 : NAND4_X1 port map( A1 => n4233, A2 => n4234, A3 => n4235, A4 => 
                           n4236, ZN => n4203);
   U7484 : AOI221_X1 port map( B1 => n11277, B2 => n9952, C1 => n11274, C2 => 
                           n9984, A => n4244, ZN => n4235);
   U7485 : NOR4_X1 port map( A1 => n4237, A2 => n4238, A3 => n4239, A4 => n4240
                           , ZN => n4236);
   U7486 : AOI222_X1 port map( A1 => n11253, A2 => n9824, B1 => n11250, B2 => 
                           n9760, C1 => n11247, C2 => n9792, ZN => n4233);
   U7487 : NAND4_X1 port map( A1 => n5606, A2 => n5607, A3 => n5608, A4 => 
                           n5609, ZN => n5595);
   U7488 : AOI221_X1 port map( B1 => n11013, B2 => n9953, C1 => n11010, C2 => 
                           n9985, A => n5614, ZN => n5608);
   U7489 : NOR4_X1 port map( A1 => n5610, A2 => n5611, A3 => n5612, A4 => n5613
                           , ZN => n5609);
   U7490 : AOI222_X1 port map( A1 => n10989, A2 => n9825, B1 => n10986, B2 => 
                           n9761, C1 => n10983, C2 => n9793, ZN => n5606);
   U7491 : NAND4_X1 port map( A1 => n4173, A2 => n4174, A3 => n4175, A4 => 
                           n4176, ZN => n4162);
   U7492 : AOI221_X1 port map( B1 => n11277, B2 => n9953, C1 => n11274, C2 => 
                           n9985, A => n4181, ZN => n4175);
   U7493 : NOR4_X1 port map( A1 => n4177, A2 => n4178, A3 => n4179, A4 => n4180
                           , ZN => n4176);
   U7494 : AOI222_X1 port map( A1 => n11253, A2 => n9825, B1 => n11250, B2 => 
                           n9761, C1 => n11247, C2 => n9793, ZN => n4173);
   U7495 : NAND4_X1 port map( A1 => n5565, A2 => n5566, A3 => n5567, A4 => 
                           n5568, ZN => n5554);
   U7496 : AOI221_X1 port map( B1 => n11013, B2 => n9954, C1 => n11010, C2 => 
                           n9986, A => n5573, ZN => n5567);
   U7497 : NOR4_X1 port map( A1 => n5569, A2 => n5570, A3 => n5571, A4 => n5572
                           , ZN => n5568);
   U7498 : AOI222_X1 port map( A1 => n10989, A2 => n9826, B1 => n10986, B2 => 
                           n9762, C1 => n10983, C2 => n9794, ZN => n5565);
   U7499 : NAND4_X1 port map( A1 => n4132, A2 => n4133, A3 => n4134, A4 => 
                           n4135, ZN => n4121);
   U7500 : AOI221_X1 port map( B1 => n11277, B2 => n9954, C1 => n11274, C2 => 
                           n9986, A => n4140, ZN => n4134);
   U7501 : NOR4_X1 port map( A1 => n4136, A2 => n4137, A3 => n4138, A4 => n4139
                           , ZN => n4135);
   U7502 : AOI222_X1 port map( A1 => n11253, A2 => n9826, B1 => n11250, B2 => 
                           n9762, C1 => n11247, C2 => n9794, ZN => n4132);
   U7503 : NAND4_X1 port map( A1 => n5524, A2 => n5525, A3 => n5526, A4 => 
                           n5527, ZN => n5513);
   U7504 : AOI221_X1 port map( B1 => n11013, B2 => n9955, C1 => n11010, C2 => 
                           n9987, A => n5532, ZN => n5526);
   U7505 : NOR4_X1 port map( A1 => n5528, A2 => n5529, A3 => n5530, A4 => n5531
                           , ZN => n5527);
   U7506 : AOI222_X1 port map( A1 => n10989, A2 => n9827, B1 => n10986, B2 => 
                           n9763, C1 => n10983, C2 => n9795, ZN => n5524);
   U7507 : NAND4_X1 port map( A1 => n4091, A2 => n4092, A3 => n4093, A4 => 
                           n4094, ZN => n4080);
   U7508 : AOI221_X1 port map( B1 => n11277, B2 => n9955, C1 => n11274, C2 => 
                           n9987, A => n4099, ZN => n4093);
   U7509 : NOR4_X1 port map( A1 => n4095, A2 => n4096, A3 => n4097, A4 => n4098
                           , ZN => n4094);
   U7510 : AOI222_X1 port map( A1 => n11253, A2 => n9827, B1 => n11250, B2 => 
                           n9763, C1 => n11247, C2 => n9795, ZN => n4091);
   U7511 : NAND4_X1 port map( A1 => n5483, A2 => n5484, A3 => n5485, A4 => 
                           n5486, ZN => n5472);
   U7512 : AOI221_X1 port map( B1 => n11013, B2 => n9956, C1 => n11010, C2 => 
                           n9988, A => n5491, ZN => n5485);
   U7513 : NOR4_X1 port map( A1 => n5487, A2 => n5488, A3 => n5489, A4 => n5490
                           , ZN => n5486);
   U7514 : AOI222_X1 port map( A1 => n10989, A2 => n9828, B1 => n10986, B2 => 
                           n9764, C1 => n10983, C2 => n9796, ZN => n5483);
   U7515 : NAND4_X1 port map( A1 => n4050, A2 => n4051, A3 => n4052, A4 => 
                           n4053, ZN => n4039);
   U7516 : AOI221_X1 port map( B1 => n11277, B2 => n9956, C1 => n11274, C2 => 
                           n9988, A => n4058, ZN => n4052);
   U7517 : NOR4_X1 port map( A1 => n4054, A2 => n4055, A3 => n4056, A4 => n4057
                           , ZN => n4053);
   U7518 : AOI222_X1 port map( A1 => n11253, A2 => n9828, B1 => n11250, B2 => 
                           n9764, C1 => n11247, C2 => n9796, ZN => n4050);
   U7519 : NAND4_X1 port map( A1 => n5442, A2 => n5443, A3 => n5444, A4 => 
                           n5445, ZN => n5431);
   U7520 : AOI221_X1 port map( B1 => n11013, B2 => n9957, C1 => n11010, C2 => 
                           n9989, A => n5450, ZN => n5444);
   U7521 : NOR4_X1 port map( A1 => n5446, A2 => n5447, A3 => n5448, A4 => n5449
                           , ZN => n5445);
   U7522 : AOI222_X1 port map( A1 => n10989, A2 => n9829, B1 => n10986, B2 => 
                           n9765, C1 => n10983, C2 => n9797, ZN => n5442);
   U7523 : NAND4_X1 port map( A1 => n4009, A2 => n4010, A3 => n4011, A4 => 
                           n4012, ZN => n3998);
   U7524 : AOI221_X1 port map( B1 => n11277, B2 => n9957, C1 => n11274, C2 => 
                           n9989, A => n4017, ZN => n4011);
   U7525 : NOR4_X1 port map( A1 => n4013, A2 => n4014, A3 => n4015, A4 => n4016
                           , ZN => n4012);
   U7526 : AOI222_X1 port map( A1 => n11253, A2 => n9829, B1 => n11250, B2 => 
                           n9765, C1 => n11247, C2 => n9797, ZN => n4009);
   U7527 : NAND4_X1 port map( A1 => n5401, A2 => n5402, A3 => n5403, A4 => 
                           n5404, ZN => n5390);
   U7528 : AOI221_X1 port map( B1 => n11013, B2 => n9958, C1 => n11010, C2 => 
                           n9990, A => n5409, ZN => n5403);
   U7529 : NOR4_X1 port map( A1 => n5405, A2 => n5406, A3 => n5407, A4 => n5408
                           , ZN => n5404);
   U7530 : AOI222_X1 port map( A1 => n10989, A2 => n9830, B1 => n10986, B2 => 
                           n9766, C1 => n10983, C2 => n9798, ZN => n5401);
   U7531 : NAND4_X1 port map( A1 => n3968, A2 => n3969, A3 => n3970, A4 => 
                           n3971, ZN => n3957);
   U7532 : AOI221_X1 port map( B1 => n11277, B2 => n9958, C1 => n11274, C2 => 
                           n9990, A => n3976, ZN => n3970);
   U7533 : NOR4_X1 port map( A1 => n3972, A2 => n3973, A3 => n3974, A4 => n3975
                           , ZN => n3971);
   U7534 : AOI222_X1 port map( A1 => n11253, A2 => n9830, B1 => n11250, B2 => 
                           n9766, C1 => n11247, C2 => n9798, ZN => n3968);
   U7535 : NAND4_X1 port map( A1 => n5360, A2 => n5361, A3 => n5362, A4 => 
                           n5363, ZN => n5349);
   U7536 : AOI221_X1 port map( B1 => n11013, B2 => n9959, C1 => n11010, C2 => 
                           n9991, A => n5368, ZN => n5362);
   U7537 : NOR4_X1 port map( A1 => n5364, A2 => n5365, A3 => n5366, A4 => n5367
                           , ZN => n5363);
   U7538 : AOI222_X1 port map( A1 => n10989, A2 => n9831, B1 => n10986, B2 => 
                           n9767, C1 => n10983, C2 => n9799, ZN => n5360);
   U7539 : NAND4_X1 port map( A1 => n3927, A2 => n3928, A3 => n3929, A4 => 
                           n3930, ZN => n3916);
   U7540 : AOI221_X1 port map( B1 => n11277, B2 => n9959, C1 => n11274, C2 => 
                           n9991, A => n3935, ZN => n3929);
   U7541 : NOR4_X1 port map( A1 => n3931, A2 => n3932, A3 => n3933, A4 => n3934
                           , ZN => n3930);
   U7542 : AOI222_X1 port map( A1 => n11253, A2 => n9831, B1 => n11250, B2 => 
                           n9767, C1 => n11247, C2 => n9799, ZN => n3927);
   U7543 : NAND4_X1 port map( A1 => n5319, A2 => n5320, A3 => n5321, A4 => 
                           n5322, ZN => n5308);
   U7544 : AOI221_X1 port map( B1 => n11013, B2 => n9960, C1 => n11010, C2 => 
                           n9992, A => n5327, ZN => n5321);
   U7545 : NOR4_X1 port map( A1 => n5323, A2 => n5324, A3 => n5325, A4 => n5326
                           , ZN => n5322);
   U7546 : AOI222_X1 port map( A1 => n10989, A2 => n9832, B1 => n10986, B2 => 
                           n9768, C1 => n10983, C2 => n9800, ZN => n5319);
   U7547 : NAND4_X1 port map( A1 => n3886, A2 => n3887, A3 => n3888, A4 => 
                           n3889, ZN => n3875);
   U7548 : AOI221_X1 port map( B1 => n11277, B2 => n9960, C1 => n11274, C2 => 
                           n9992, A => n3894, ZN => n3888);
   U7549 : NOR4_X1 port map( A1 => n3890, A2 => n3891, A3 => n3892, A4 => n3893
                           , ZN => n3889);
   U7550 : AOI222_X1 port map( A1 => n11253, A2 => n9832, B1 => n11250, B2 => 
                           n9768, C1 => n11247, C2 => n9800, ZN => n3886);
   U7551 : NAND4_X1 port map( A1 => n5278, A2 => n5279, A3 => n5280, A4 => 
                           n5281, ZN => n5267);
   U7552 : AOI221_X1 port map( B1 => n11013, B2 => n9961, C1 => n11010, C2 => 
                           n9993, A => n5286, ZN => n5280);
   U7553 : NOR4_X1 port map( A1 => n5282, A2 => n5283, A3 => n5284, A4 => n5285
                           , ZN => n5281);
   U7554 : AOI222_X1 port map( A1 => n10989, A2 => n9833, B1 => n10986, B2 => 
                           n9769, C1 => n10983, C2 => n9801, ZN => n5278);
   U7555 : NAND4_X1 port map( A1 => n3845, A2 => n3846, A3 => n3847, A4 => 
                           n3848, ZN => n3834);
   U7556 : AOI221_X1 port map( B1 => n11277, B2 => n9961, C1 => n11274, C2 => 
                           n9993, A => n3853, ZN => n3847);
   U7557 : NOR4_X1 port map( A1 => n3849, A2 => n3850, A3 => n3851, A4 => n3852
                           , ZN => n3848);
   U7558 : AOI222_X1 port map( A1 => n11253, A2 => n9833, B1 => n11250, B2 => 
                           n9769, C1 => n11247, C2 => n9801, ZN => n3845);
   U7559 : NAND4_X1 port map( A1 => n5237, A2 => n5238, A3 => n5239, A4 => 
                           n5240, ZN => n5226);
   U7560 : AOI221_X1 port map( B1 => n11013, B2 => n9962, C1 => n11010, C2 => 
                           n9994, A => n5245, ZN => n5239);
   U7561 : NOR4_X1 port map( A1 => n5241, A2 => n5242, A3 => n5243, A4 => n5244
                           , ZN => n5240);
   U7562 : AOI222_X1 port map( A1 => n10989, A2 => n9834, B1 => n10986, B2 => 
                           n9770, C1 => n10983, C2 => n9802, ZN => n5237);
   U7563 : NAND4_X1 port map( A1 => n3804, A2 => n3805, A3 => n3806, A4 => 
                           n3807, ZN => n3793);
   U7564 : AOI221_X1 port map( B1 => n11277, B2 => n9962, C1 => n11274, C2 => 
                           n9994, A => n3812, ZN => n3806);
   U7565 : NOR4_X1 port map( A1 => n3808, A2 => n3809, A3 => n3810, A4 => n3811
                           , ZN => n3807);
   U7566 : AOI222_X1 port map( A1 => n11253, A2 => n9834, B1 => n11250, B2 => 
                           n9770, C1 => n11247, C2 => n9802, ZN => n3804);
   U7567 : NAND4_X1 port map( A1 => n5196, A2 => n5197, A3 => n5198, A4 => 
                           n5199, ZN => n5185);
   U7568 : AOI221_X1 port map( B1 => n11013, B2 => n9963, C1 => n11010, C2 => 
                           n9995, A => n5204, ZN => n5198);
   U7569 : NOR4_X1 port map( A1 => n5200, A2 => n5201, A3 => n5202, A4 => n5203
                           , ZN => n5199);
   U7570 : AOI222_X1 port map( A1 => n10989, A2 => n9835, B1 => n10986, B2 => 
                           n9771, C1 => n10983, C2 => n9803, ZN => n5196);
   U7571 : NAND4_X1 port map( A1 => n3763, A2 => n3764, A3 => n3765, A4 => 
                           n3766, ZN => n3752);
   U7572 : AOI221_X1 port map( B1 => n11277, B2 => n9963, C1 => n11274, C2 => 
                           n9995, A => n3771, ZN => n3765);
   U7573 : NOR4_X1 port map( A1 => n3767, A2 => n3768, A3 => n3769, A4 => n3770
                           , ZN => n3766);
   U7574 : AOI222_X1 port map( A1 => n11253, A2 => n9835, B1 => n11250, B2 => 
                           n9771, C1 => n11247, C2 => n9803, ZN => n3763);
   U7575 : NAND4_X1 port map( A1 => n5155, A2 => n5156, A3 => n5157, A4 => 
                           n5158, ZN => n5144);
   U7576 : AOI221_X1 port map( B1 => n11014, B2 => n9964, C1 => n11011, C2 => 
                           n9996, A => n5163, ZN => n5157);
   U7577 : NOR4_X1 port map( A1 => n5159, A2 => n5160, A3 => n5161, A4 => n5162
                           , ZN => n5158);
   U7578 : AOI222_X1 port map( A1 => n10990, A2 => n9836, B1 => n10987, B2 => 
                           n9772, C1 => n10984, C2 => n9804, ZN => n5155);
   U7579 : NAND4_X1 port map( A1 => n3722, A2 => n3723, A3 => n3724, A4 => 
                           n3725, ZN => n3711);
   U7580 : AOI221_X1 port map( B1 => n11278, B2 => n9964, C1 => n11275, C2 => 
                           n9996, A => n3730, ZN => n3724);
   U7581 : NOR4_X1 port map( A1 => n3726, A2 => n3727, A3 => n3728, A4 => n3729
                           , ZN => n3725);
   U7582 : AOI222_X1 port map( A1 => n11254, A2 => n9836, B1 => n11251, B2 => 
                           n9772, C1 => n11248, C2 => n9804, ZN => n3722);
   U7583 : NAND4_X1 port map( A1 => n5114, A2 => n5115, A3 => n5116, A4 => 
                           n5117, ZN => n5103);
   U7584 : AOI221_X1 port map( B1 => n11014, B2 => n9965, C1 => n11011, C2 => 
                           n9997, A => n5122, ZN => n5116);
   U7585 : NOR4_X1 port map( A1 => n5118, A2 => n5119, A3 => n5120, A4 => n5121
                           , ZN => n5117);
   U7586 : AOI222_X1 port map( A1 => n10990, A2 => n9837, B1 => n10987, B2 => 
                           n9773, C1 => n10984, C2 => n9805, ZN => n5114);
   U7587 : NAND4_X1 port map( A1 => n3681, A2 => n3682, A3 => n3683, A4 => 
                           n3684, ZN => n3670);
   U7588 : AOI221_X1 port map( B1 => n11278, B2 => n9965, C1 => n11275, C2 => 
                           n9997, A => n3689, ZN => n3683);
   U7589 : NOR4_X1 port map( A1 => n3685, A2 => n3686, A3 => n3687, A4 => n3688
                           , ZN => n3684);
   U7590 : AOI222_X1 port map( A1 => n11254, A2 => n9837, B1 => n11251, B2 => 
                           n9773, C1 => n11248, C2 => n9805, ZN => n3681);
   U7591 : NAND4_X1 port map( A1 => n5073, A2 => n5074, A3 => n5075, A4 => 
                           n5076, ZN => n5062);
   U7592 : AOI221_X1 port map( B1 => n11014, B2 => n9966, C1 => n11011, C2 => 
                           n9998, A => n5081, ZN => n5075);
   U7593 : NOR4_X1 port map( A1 => n5077, A2 => n5078, A3 => n5079, A4 => n5080
                           , ZN => n5076);
   U7594 : AOI222_X1 port map( A1 => n10990, A2 => n9838, B1 => n10987, B2 => 
                           n9774, C1 => n10984, C2 => n9806, ZN => n5073);
   U7595 : NAND4_X1 port map( A1 => n3640, A2 => n3641, A3 => n3642, A4 => 
                           n3643, ZN => n3629);
   U7596 : AOI221_X1 port map( B1 => n11278, B2 => n9966, C1 => n11275, C2 => 
                           n9998, A => n3648, ZN => n3642);
   U7597 : NOR4_X1 port map( A1 => n3644, A2 => n3645, A3 => n3646, A4 => n3647
                           , ZN => n3643);
   U7598 : AOI222_X1 port map( A1 => n11254, A2 => n9838, B1 => n11251, B2 => 
                           n9774, C1 => n11248, C2 => n9806, ZN => n3640);
   U7599 : NAND4_X1 port map( A1 => n5032, A2 => n5033, A3 => n5034, A4 => 
                           n5035, ZN => n5021);
   U7600 : AOI221_X1 port map( B1 => n11014, B2 => n9967, C1 => n11011, C2 => 
                           n9999, A => n5040, ZN => n5034);
   U7601 : NOR4_X1 port map( A1 => n5036, A2 => n5037, A3 => n5038, A4 => n5039
                           , ZN => n5035);
   U7602 : AOI222_X1 port map( A1 => n10990, A2 => n9839, B1 => n10987, B2 => 
                           n9775, C1 => n10984, C2 => n9807, ZN => n5032);
   U7603 : NAND4_X1 port map( A1 => n3599, A2 => n3600, A3 => n3601, A4 => 
                           n3602, ZN => n3588);
   U7604 : AOI221_X1 port map( B1 => n11278, B2 => n9967, C1 => n11275, C2 => 
                           n9999, A => n3607, ZN => n3601);
   U7605 : NOR4_X1 port map( A1 => n3603, A2 => n3604, A3 => n3605, A4 => n3606
                           , ZN => n3602);
   U7606 : AOI222_X1 port map( A1 => n11254, A2 => n9839, B1 => n11251, B2 => 
                           n9775, C1 => n11248, C2 => n9807, ZN => n3599);
   U7607 : NAND4_X1 port map( A1 => n4991, A2 => n4992, A3 => n4993, A4 => 
                           n4994, ZN => n4980);
   U7608 : AOI221_X1 port map( B1 => n11014, B2 => n9968, C1 => n11011, C2 => 
                           n13059, A => n4999, ZN => n4993);
   U7609 : NOR4_X1 port map( A1 => n4995, A2 => n4996, A3 => n4997, A4 => n4998
                           , ZN => n4994);
   U7610 : AOI222_X1 port map( A1 => n10990, A2 => n9840, B1 => n10987, B2 => 
                           n9776, C1 => n10984, C2 => n9808, ZN => n4991);
   U7611 : NAND4_X1 port map( A1 => n3558, A2 => n3559, A3 => n3560, A4 => 
                           n3561, ZN => n3547);
   U7612 : AOI221_X1 port map( B1 => n11278, B2 => n9968, C1 => n11275, C2 => 
                           n13059, A => n3566, ZN => n3560);
   U7613 : NOR4_X1 port map( A1 => n3562, A2 => n3563, A3 => n3564, A4 => n3565
                           , ZN => n3561);
   U7614 : AOI222_X1 port map( A1 => n11254, A2 => n9840, B1 => n11251, B2 => 
                           n9776, C1 => n11248, C2 => n9808, ZN => n3558);
   U7615 : NAND4_X1 port map( A1 => n4950, A2 => n4951, A3 => n4952, A4 => 
                           n4953, ZN => n4939);
   U7616 : AOI221_X1 port map( B1 => n11014, B2 => n9969, C1 => n11011, C2 => 
                           n13058, A => n4958, ZN => n4952);
   U7617 : NOR4_X1 port map( A1 => n4954, A2 => n4955, A3 => n4956, A4 => n4957
                           , ZN => n4953);
   U7618 : AOI222_X1 port map( A1 => n10990, A2 => n9841, B1 => n10987, B2 => 
                           n9777, C1 => n10984, C2 => n9809, ZN => n4950);
   U7619 : NAND4_X1 port map( A1 => n3517, A2 => n3518, A3 => n3519, A4 => 
                           n3520, ZN => n3506);
   U7620 : AOI221_X1 port map( B1 => n11278, B2 => n9969, C1 => n11275, C2 => 
                           n13058, A => n3525, ZN => n3519);
   U7621 : NOR4_X1 port map( A1 => n3521, A2 => n3522, A3 => n3523, A4 => n3524
                           , ZN => n3520);
   U7622 : AOI222_X1 port map( A1 => n11254, A2 => n9841, B1 => n11251, B2 => 
                           n9777, C1 => n11248, C2 => n9809, ZN => n3517);
   U7623 : NAND4_X1 port map( A1 => n4909, A2 => n4910, A3 => n4911, A4 => 
                           n4912, ZN => n4898);
   U7624 : AOI221_X1 port map( B1 => n11014, B2 => n9970, C1 => n11011, C2 => 
                           n13057, A => n4917, ZN => n4911);
   U7625 : NOR4_X1 port map( A1 => n4913, A2 => n4914, A3 => n4915, A4 => n4916
                           , ZN => n4912);
   U7626 : AOI222_X1 port map( A1 => n10990, A2 => n9842, B1 => n10987, B2 => 
                           n9778, C1 => n10984, C2 => n9810, ZN => n4909);
   U7627 : NAND4_X1 port map( A1 => n3476, A2 => n3477, A3 => n3478, A4 => 
                           n3479, ZN => n3465);
   U7628 : AOI221_X1 port map( B1 => n11278, B2 => n9970, C1 => n11275, C2 => 
                           n13057, A => n3484, ZN => n3478);
   U7629 : NOR4_X1 port map( A1 => n3480, A2 => n3481, A3 => n3482, A4 => n3483
                           , ZN => n3479);
   U7630 : AOI222_X1 port map( A1 => n11254, A2 => n9842, B1 => n11251, B2 => 
                           n9778, C1 => n11248, C2 => n9810, ZN => n3476);
   U7631 : NAND4_X1 port map( A1 => n4868, A2 => n4869, A3 => n4870, A4 => 
                           n4871, ZN => n4857);
   U7632 : AOI221_X1 port map( B1 => n11014, B2 => n9971, C1 => n11011, C2 => 
                           n13056, A => n4876, ZN => n4870);
   U7633 : NOR4_X1 port map( A1 => n4872, A2 => n4873, A3 => n4874, A4 => n4875
                           , ZN => n4871);
   U7634 : AOI222_X1 port map( A1 => n10990, A2 => n9843, B1 => n10987, B2 => 
                           n9779, C1 => n10984, C2 => n9811, ZN => n4868);
   U7635 : NAND4_X1 port map( A1 => n3435, A2 => n3436, A3 => n3437, A4 => 
                           n3438, ZN => n3424);
   U7636 : AOI221_X1 port map( B1 => n11278, B2 => n9971, C1 => n11275, C2 => 
                           n13056, A => n3443, ZN => n3437);
   U7637 : NOR4_X1 port map( A1 => n3439, A2 => n3440, A3 => n3441, A4 => n3442
                           , ZN => n3438);
   U7638 : AOI222_X1 port map( A1 => n11254, A2 => n9843, B1 => n11251, B2 => 
                           n9779, C1 => n11248, C2 => n9811, ZN => n3435);
   U7639 : NAND4_X1 port map( A1 => n4827, A2 => n4828, A3 => n4829, A4 => 
                           n4830, ZN => n4816);
   U7640 : AOI221_X1 port map( B1 => n11014, B2 => n9972, C1 => n11011, C2 => 
                           n13055, A => n4835, ZN => n4829);
   U7641 : NOR4_X1 port map( A1 => n4831, A2 => n4832, A3 => n4833, A4 => n4834
                           , ZN => n4830);
   U7642 : AOI222_X1 port map( A1 => n10990, A2 => n9844, B1 => n10987, B2 => 
                           n9780, C1 => n10984, C2 => n9812, ZN => n4827);
   U7643 : NAND4_X1 port map( A1 => n3394, A2 => n3395, A3 => n3396, A4 => 
                           n3397, ZN => n3383);
   U7644 : AOI221_X1 port map( B1 => n11278, B2 => n9972, C1 => n11275, C2 => 
                           n13055, A => n3402, ZN => n3396);
   U7645 : NOR4_X1 port map( A1 => n3398, A2 => n3399, A3 => n3400, A4 => n3401
                           , ZN => n3397);
   U7646 : AOI222_X1 port map( A1 => n11254, A2 => n9844, B1 => n11251, B2 => 
                           n9780, C1 => n11248, C2 => n9812, ZN => n3394);
   U7647 : NAND4_X1 port map( A1 => n4786, A2 => n4787, A3 => n4788, A4 => 
                           n4789, ZN => n4775);
   U7648 : AOI221_X1 port map( B1 => n11014, B2 => n9973, C1 => n11011, C2 => 
                           n13054, A => n4794, ZN => n4788);
   U7649 : NOR4_X1 port map( A1 => n4790, A2 => n4791, A3 => n4792, A4 => n4793
                           , ZN => n4789);
   U7650 : AOI222_X1 port map( A1 => n10990, A2 => n9845, B1 => n10987, B2 => 
                           n9781, C1 => n10984, C2 => n9813, ZN => n4786);
   U7651 : NAND4_X1 port map( A1 => n3353, A2 => n3354, A3 => n3355, A4 => 
                           n3356, ZN => n3342);
   U7652 : AOI221_X1 port map( B1 => n11278, B2 => n9973, C1 => n11275, C2 => 
                           n13054, A => n3361, ZN => n3355);
   U7653 : NOR4_X1 port map( A1 => n3357, A2 => n3358, A3 => n3359, A4 => n3360
                           , ZN => n3356);
   U7654 : AOI222_X1 port map( A1 => n11254, A2 => n9845, B1 => n11251, B2 => 
                           n9781, C1 => n11248, C2 => n9813, ZN => n3353);
   U7655 : NAND4_X1 port map( A1 => n4745, A2 => n4746, A3 => n4747, A4 => 
                           n4748, ZN => n4734);
   U7656 : AOI221_X1 port map( B1 => n11014, B2 => n9974, C1 => n11011, C2 => 
                           n13053, A => n4753, ZN => n4747);
   U7657 : NOR4_X1 port map( A1 => n4749, A2 => n4750, A3 => n4751, A4 => n4752
                           , ZN => n4748);
   U7658 : AOI222_X1 port map( A1 => n10990, A2 => n9846, B1 => n10987, B2 => 
                           n9782, C1 => n10984, C2 => n9814, ZN => n4745);
   U7659 : NAND4_X1 port map( A1 => n3312, A2 => n3313, A3 => n3314, A4 => 
                           n3315, ZN => n3301);
   U7660 : AOI221_X1 port map( B1 => n11278, B2 => n9974, C1 => n11275, C2 => 
                           n13053, A => n3320, ZN => n3314);
   U7661 : NOR4_X1 port map( A1 => n3316, A2 => n3317, A3 => n3318, A4 => n3319
                           , ZN => n3315);
   U7662 : AOI222_X1 port map( A1 => n11254, A2 => n9846, B1 => n11251, B2 => 
                           n9782, C1 => n11248, C2 => n9814, ZN => n3312);
   U7663 : NAND4_X1 port map( A1 => n4704, A2 => n4705, A3 => n4706, A4 => 
                           n4707, ZN => n4693);
   U7664 : AOI221_X1 port map( B1 => n11014, B2 => n9975, C1 => n11011, C2 => 
                           n13052, A => n4712, ZN => n4706);
   U7665 : NOR4_X1 port map( A1 => n4708, A2 => n4709, A3 => n4710, A4 => n4711
                           , ZN => n4707);
   U7666 : AOI222_X1 port map( A1 => n10990, A2 => n9847, B1 => n10987, B2 => 
                           n9783, C1 => n10984, C2 => n9815, ZN => n4704);
   U7667 : NAND4_X1 port map( A1 => n3271, A2 => n3272, A3 => n3273, A4 => 
                           n3274, ZN => n3260);
   U7668 : AOI221_X1 port map( B1 => n11278, B2 => n9975, C1 => n11275, C2 => 
                           n13052, A => n3279, ZN => n3273);
   U7669 : NOR4_X1 port map( A1 => n3275, A2 => n3276, A3 => n3277, A4 => n3278
                           , ZN => n3274);
   U7670 : AOI222_X1 port map( A1 => n11254, A2 => n9847, B1 => n11251, B2 => 
                           n9783, C1 => n11248, C2 => n9815, ZN => n3271);
   U7671 : NAND4_X1 port map( A1 => n4663, A2 => n4664, A3 => n4665, A4 => 
                           n4666, ZN => n4652);
   U7672 : AOI221_X1 port map( B1 => n11015, B2 => n9976, C1 => n11012, C2 => 
                           n13051, A => n4671, ZN => n4665);
   U7673 : NOR4_X1 port map( A1 => n4667, A2 => n4668, A3 => n4669, A4 => n4670
                           , ZN => n4666);
   U7674 : AOI222_X1 port map( A1 => n10991, A2 => n9848, B1 => n10988, B2 => 
                           n9784, C1 => n10985, C2 => n9816, ZN => n4663);
   U7675 : NAND4_X1 port map( A1 => n3230, A2 => n3231, A3 => n3232, A4 => 
                           n3233, ZN => n3219);
   U7676 : AOI221_X1 port map( B1 => n11279, B2 => n9976, C1 => n11276, C2 => 
                           n13051, A => n3238, ZN => n3232);
   U7677 : NOR4_X1 port map( A1 => n3234, A2 => n3235, A3 => n3236, A4 => n3237
                           , ZN => n3233);
   U7678 : AOI222_X1 port map( A1 => n11255, A2 => n9848, B1 => n11252, B2 => 
                           n9784, C1 => n11249, C2 => n9816, ZN => n3230);
   U7679 : NAND4_X1 port map( A1 => n4622, A2 => n4623, A3 => n4624, A4 => 
                           n4625, ZN => n4611);
   U7680 : AOI221_X1 port map( B1 => n11015, B2 => n9977, C1 => n11012, C2 => 
                           n13050, A => n4630, ZN => n4624);
   U7681 : NOR4_X1 port map( A1 => n4626, A2 => n4627, A3 => n4628, A4 => n4629
                           , ZN => n4625);
   U7682 : AOI222_X1 port map( A1 => n10991, A2 => n9849, B1 => n10988, B2 => 
                           n9785, C1 => n10985, C2 => n9817, ZN => n4622);
   U7683 : NAND4_X1 port map( A1 => n3189, A2 => n3190, A3 => n3191, A4 => 
                           n3192, ZN => n3178);
   U7684 : AOI221_X1 port map( B1 => n11279, B2 => n9977, C1 => n11276, C2 => 
                           n13050, A => n3197, ZN => n3191);
   U7685 : NOR4_X1 port map( A1 => n3193, A2 => n3194, A3 => n3195, A4 => n3196
                           , ZN => n3192);
   U7686 : AOI222_X1 port map( A1 => n11255, A2 => n9849, B1 => n11252, B2 => 
                           n9785, C1 => n11249, C2 => n9817, ZN => n3189);
   U7687 : NAND4_X1 port map( A1 => n4581, A2 => n4582, A3 => n4583, A4 => 
                           n4584, ZN => n4570);
   U7688 : AOI221_X1 port map( B1 => n11015, B2 => n9978, C1 => n11012, C2 => 
                           n13049, A => n4589, ZN => n4583);
   U7689 : NOR4_X1 port map( A1 => n4585, A2 => n4586, A3 => n4587, A4 => n4588
                           , ZN => n4584);
   U7690 : AOI222_X1 port map( A1 => n10991, A2 => n9850, B1 => n10988, B2 => 
                           n9786, C1 => n10985, C2 => n9818, ZN => n4581);
   U7691 : NAND4_X1 port map( A1 => n3148, A2 => n3149, A3 => n3150, A4 => 
                           n3151, ZN => n3137);
   U7692 : AOI221_X1 port map( B1 => n11279, B2 => n9978, C1 => n11276, C2 => 
                           n13049, A => n3156, ZN => n3150);
   U7693 : NOR4_X1 port map( A1 => n3152, A2 => n3153, A3 => n3154, A4 => n3155
                           , ZN => n3151);
   U7694 : AOI222_X1 port map( A1 => n11255, A2 => n9850, B1 => n11252, B2 => 
                           n9786, C1 => n11249, C2 => n9818, ZN => n3148);
   U7695 : NAND4_X1 port map( A1 => n4540, A2 => n4541, A3 => n4542, A4 => 
                           n4543, ZN => n4529);
   U7696 : AOI221_X1 port map( B1 => n11015, B2 => n9979, C1 => n11012, C2 => 
                           n13048, A => n4548, ZN => n4542);
   U7697 : NOR4_X1 port map( A1 => n4544, A2 => n4545, A3 => n4546, A4 => n4547
                           , ZN => n4543);
   U7698 : AOI222_X1 port map( A1 => n10991, A2 => n9851, B1 => n10988, B2 => 
                           n9787, C1 => n10985, C2 => n9819, ZN => n4540);
   U7699 : NAND4_X1 port map( A1 => n3107, A2 => n3108, A3 => n3109, A4 => 
                           n3110, ZN => n3096);
   U7700 : AOI221_X1 port map( B1 => n11279, B2 => n9979, C1 => n11276, C2 => 
                           n13048, A => n3115, ZN => n3109);
   U7701 : NOR4_X1 port map( A1 => n3111, A2 => n3112, A3 => n3113, A4 => n3114
                           , ZN => n3110);
   U7702 : AOI222_X1 port map( A1 => n11255, A2 => n9851, B1 => n11252, B2 => 
                           n9787, C1 => n11249, C2 => n9819, ZN => n3107);
   U7703 : NAND4_X1 port map( A1 => n4499, A2 => n4500, A3 => n4501, A4 => 
                           n4502, ZN => n4488);
   U7704 : AOI221_X1 port map( B1 => n11015, B2 => n9980, C1 => n11012, C2 => 
                           n13047, A => n4507, ZN => n4501);
   U7705 : NOR4_X1 port map( A1 => n4503, A2 => n4504, A3 => n4505, A4 => n4506
                           , ZN => n4502);
   U7706 : AOI222_X1 port map( A1 => n10991, A2 => n9852, B1 => n10988, B2 => 
                           n9788, C1 => n10985, C2 => n9820, ZN => n4499);
   U7707 : NAND4_X1 port map( A1 => n3066, A2 => n3067, A3 => n3068, A4 => 
                           n3069, ZN => n3055);
   U7708 : AOI221_X1 port map( B1 => n11279, B2 => n9980, C1 => n11276, C2 => 
                           n13047, A => n3074, ZN => n3068);
   U7709 : NOR4_X1 port map( A1 => n3070, A2 => n3071, A3 => n3072, A4 => n3073
                           , ZN => n3069);
   U7710 : AOI222_X1 port map( A1 => n11255, A2 => n9852, B1 => n11252, B2 => 
                           n9788, C1 => n11249, C2 => n9820, ZN => n3066);
   U7711 : NAND4_X1 port map( A1 => n4458, A2 => n4459, A3 => n4460, A4 => 
                           n4461, ZN => n4447);
   U7712 : AOI221_X1 port map( B1 => n11015, B2 => n9981, C1 => n11012, C2 => 
                           n13046, A => n4466, ZN => n4460);
   U7713 : NOR4_X1 port map( A1 => n4462, A2 => n4463, A3 => n4464, A4 => n4465
                           , ZN => n4461);
   U7714 : AOI222_X1 port map( A1 => n10991, A2 => n9853, B1 => n10988, B2 => 
                           n9789, C1 => n10985, C2 => n9821, ZN => n4458);
   U7715 : NAND4_X1 port map( A1 => n3025, A2 => n3026, A3 => n3027, A4 => 
                           n3028, ZN => n3014);
   U7716 : AOI221_X1 port map( B1 => n11279, B2 => n9981, C1 => n11276, C2 => 
                           n13046, A => n3033, ZN => n3027);
   U7717 : NOR4_X1 port map( A1 => n3029, A2 => n3030, A3 => n3031, A4 => n3032
                           , ZN => n3028);
   U7718 : AOI222_X1 port map( A1 => n11255, A2 => n9853, B1 => n11252, B2 => 
                           n9789, C1 => n11249, C2 => n9821, ZN => n3025);
   U7719 : NAND4_X1 port map( A1 => n4417, A2 => n4418, A3 => n4419, A4 => 
                           n4420, ZN => n4406);
   U7720 : AOI221_X1 port map( B1 => n11015, B2 => n9982, C1 => n11012, C2 => 
                           n13045, A => n4425, ZN => n4419);
   U7721 : NOR4_X1 port map( A1 => n4421, A2 => n4422, A3 => n4423, A4 => n4424
                           , ZN => n4420);
   U7722 : AOI222_X1 port map( A1 => n10991, A2 => n9854, B1 => n10988, B2 => 
                           n9790, C1 => n10985, C2 => n9822, ZN => n4417);
   U7723 : NAND4_X1 port map( A1 => n2984, A2 => n2985, A3 => n2986, A4 => 
                           n2987, ZN => n2973);
   U7724 : AOI221_X1 port map( B1 => n11279, B2 => n9982, C1 => n11276, C2 => 
                           n13045, A => n2992, ZN => n2986);
   U7725 : NOR4_X1 port map( A1 => n2988, A2 => n2989, A3 => n2990, A4 => n2991
                           , ZN => n2987);
   U7726 : AOI222_X1 port map( A1 => n11255, A2 => n9854, B1 => n11252, B2 => 
                           n9790, C1 => n11249, C2 => n9822, ZN => n2984);
   U7727 : NAND4_X1 port map( A1 => n4310, A2 => n4311, A3 => n4312, A4 => 
                           n4313, ZN => n4277);
   U7728 : AOI221_X1 port map( B1 => n11015, B2 => n9983, C1 => n11012, C2 => 
                           n13044, A => n4331, ZN => n4312);
   U7729 : NOR4_X1 port map( A1 => n4314, A2 => n4315, A3 => n4316, A4 => n4317
                           , ZN => n4313);
   U7730 : AOI222_X1 port map( A1 => n10991, A2 => n9855, B1 => n10988, B2 => 
                           n9791, C1 => n10985, C2 => n9823, ZN => n4310);
   U7731 : NAND4_X1 port map( A1 => n2810, A2 => n2811, A3 => n2812, A4 => 
                           n2813, ZN => n2745);
   U7732 : AOI221_X1 port map( B1 => n11279, B2 => n9983, C1 => n11276, C2 => 
                           n13044, A => n2863, ZN => n2812);
   U7733 : NOR4_X1 port map( A1 => n2814, A2 => n2815, A3 => n2816, A4 => n2817
                           , ZN => n2813);
   U7734 : AOI222_X1 port map( A1 => n11255, A2 => n9855, B1 => n11252, B2 => 
                           n9791, C1 => n11249, C2 => n9823, ZN => n2810);
   U7735 : NAND2_X1 port map( A1 => n2937, A2 => n2740, ZN => U3_U98_Z_4);
   U7736 : NAND2_X1 port map( A1 => n2937, A2 => n2739, ZN => U3_U99_Z_4);
   U7737 : NAND2_X1 port map( A1 => n2937, A2 => n2741, ZN => U3_U97_Z_4);
   U7738 : NAND2_X1 port map( A1 => n2936, A2 => n2740, ZN => U3_U98_Z_5);
   U7739 : NAND2_X1 port map( A1 => n2936, A2 => n2739, ZN => U3_U99_Z_5);
   U7740 : NAND2_X1 port map( A1 => n2936, A2 => n2741, ZN => U3_U97_Z_5);
   U7741 : INV_X1 port map( A => DATAIN(0), ZN => n12768);
   U7742 : INV_X1 port map( A => DATAIN(1), ZN => n12767);
   U7743 : INV_X1 port map( A => DATAIN(2), ZN => n12766);
   U7744 : INV_X1 port map( A => DATAIN(3), ZN => n12765);
   U7745 : INV_X1 port map( A => DATAIN(4), ZN => n12764);
   U7746 : INV_X1 port map( A => DATAIN(5), ZN => n12763);
   U7747 : INV_X1 port map( A => DATAIN(6), ZN => n12762);
   U7748 : INV_X1 port map( A => DATAIN(7), ZN => n12761);
   U7749 : INV_X1 port map( A => DATAIN(8), ZN => n12760);
   U7750 : INV_X1 port map( A => DATAIN(9), ZN => n12759);
   U7751 : INV_X1 port map( A => DATAIN(10), ZN => n12758);
   U7752 : INV_X1 port map( A => DATAIN(11), ZN => n12757);
   U7753 : INV_X1 port map( A => DATAIN(12), ZN => n12756);
   U7754 : INV_X1 port map( A => DATAIN(13), ZN => n12755);
   U7755 : INV_X1 port map( A => DATAIN(14), ZN => n12754);
   U7756 : INV_X1 port map( A => DATAIN(15), ZN => n12753);
   U7757 : INV_X1 port map( A => DATAIN(16), ZN => n12752);
   U7758 : INV_X1 port map( A => DATAIN(17), ZN => n12751);
   U7759 : INV_X1 port map( A => DATAIN(18), ZN => n12750);
   U7760 : INV_X1 port map( A => DATAIN(19), ZN => n12749);
   U7761 : INV_X1 port map( A => DATAIN(20), ZN => n12748);
   U7762 : INV_X1 port map( A => DATAIN(21), ZN => n12747);
   U7763 : INV_X1 port map( A => DATAIN(22), ZN => n12746);
   U7764 : INV_X1 port map( A => DATAIN(23), ZN => n12745);
   U7765 : INV_X1 port map( A => DATAIN(24), ZN => n12744);
   U7766 : INV_X1 port map( A => DATAIN(25), ZN => n12743);
   U7767 : INV_X1 port map( A => DATAIN(26), ZN => n12742);
   U7768 : INV_X1 port map( A => DATAIN(27), ZN => n12741);
   U7769 : INV_X1 port map( A => DATAIN(28), ZN => n12740);
   U7770 : INV_X1 port map( A => DATAIN(29), ZN => n12739);
   U7771 : INV_X1 port map( A => DATAIN(30), ZN => n12738);
   U7772 : INV_X1 port map( A => DATAIN(31), ZN => n12737);
   U7773 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n2740);
   U7774 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n2739);
   U7775 : NAND2_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), ZN => n2741);
   U7776 : INV_X1 port map( A => ADD_RD1(0), ZN => n14514);
   U7777 : INV_X1 port map( A => ADD_RD2(0), ZN => n14516);
   U7778 : INV_X1 port map( A => ADD_RD1(1), ZN => n14513);
   U7779 : INV_X1 port map( A => ADD_RD2(1), ZN => n14515);
   U7780 : AND2_X1 port map( A1 => N2170, A2 => ADD_WR(2), ZN => n2716);
   U7781 : INV_X1 port map( A => ADD_WR(0), ZN => n12736);
   U7782 : INV_X1 port map( A => ADD_WR(1), ZN => n12735);
   U7783 : INV_X1 port map( A => ADD_WR(2), ZN => n12734);
   U7784 : OR2_X1 port map( A1 => RD1, A2 => n12712, ZN => N8702);
   U7785 : OR2_X1 port map( A1 => RD2, A2 => n12712, ZN => N8735);
   U7786 : INV_X1 port map( A => n11390, ZN => n11381);
   U7787 : INV_X1 port map( A => n11402, ZN => n11393);
   U7788 : INV_X1 port map( A => n11414, ZN => n11405);
   U7789 : INV_X1 port map( A => n11426, ZN => n11417);
   U7790 : INV_X1 port map( A => n11438, ZN => n11429);
   U7791 : INV_X1 port map( A => n11450, ZN => n11441);
   U7792 : INV_X1 port map( A => n11462, ZN => n11453);
   U7793 : INV_X1 port map( A => n11474, ZN => n11465);
   U7794 : INV_X1 port map( A => n11486, ZN => n11477);
   U7795 : INV_X1 port map( A => n11498, ZN => n11489);
   U7796 : INV_X1 port map( A => n11510, ZN => n11501);
   U7797 : INV_X1 port map( A => n11522, ZN => n11513);
   U7798 : INV_X1 port map( A => n11534, ZN => n11525);
   U7799 : INV_X1 port map( A => n11546, ZN => n11537);
   U7800 : INV_X1 port map( A => n11558, ZN => n11549);
   U7801 : INV_X1 port map( A => n11570, ZN => n11561);
   U7802 : INV_X1 port map( A => n11582, ZN => n11573);
   U7803 : INV_X1 port map( A => n11594, ZN => n11585);
   U7804 : INV_X1 port map( A => n11606, ZN => n11597);
   U7805 : INV_X1 port map( A => n11618, ZN => n11609);
   U7806 : INV_X1 port map( A => n11630, ZN => n11621);
   U7807 : INV_X1 port map( A => n11642, ZN => n11633);
   U7808 : INV_X1 port map( A => n11654, ZN => n11645);
   U7809 : INV_X1 port map( A => n11666, ZN => n11657);
   U7810 : INV_X1 port map( A => n11678, ZN => n11669);
   U7811 : INV_X1 port map( A => n11690, ZN => n11681);
   U7812 : INV_X1 port map( A => n11702, ZN => n11693);
   U7813 : INV_X1 port map( A => n11714, ZN => n11705);
   U7814 : INV_X1 port map( A => n11726, ZN => n11717);
   U7815 : INV_X1 port map( A => n11738, ZN => n11729);
   U7816 : INV_X1 port map( A => n11750, ZN => n11741);
   U7817 : INV_X1 port map( A => n11762, ZN => n11753);
   U7818 : INV_X1 port map( A => n11774, ZN => n11765);
   U7819 : INV_X1 port map( A => n11786, ZN => n11777);
   U7820 : INV_X1 port map( A => n11798, ZN => n11789);
   U7821 : INV_X1 port map( A => n11810, ZN => n11801);
   U7822 : INV_X1 port map( A => n11822, ZN => n11813);
   U7823 : INV_X1 port map( A => n11834, ZN => n11825);
   U7824 : INV_X1 port map( A => n11846, ZN => n11837);
   U7825 : INV_X1 port map( A => n11858, ZN => n11849);
   U7826 : INV_X1 port map( A => n11870, ZN => n11861);
   U7827 : INV_X1 port map( A => n11882, ZN => n11873);
   U7828 : INV_X1 port map( A => n11894, ZN => n11885);
   U7829 : INV_X1 port map( A => n11906, ZN => n11897);
   U7830 : INV_X1 port map( A => n11918, ZN => n11909);
   U7831 : INV_X1 port map( A => n11930, ZN => n11921);
   U7832 : INV_X1 port map( A => n11942, ZN => n11933);
   U7833 : INV_X1 port map( A => n11954, ZN => n11945);
   U7834 : INV_X1 port map( A => n11966, ZN => n11957);
   U7839 : INV_X1 port map( A => n11978, ZN => n11969);
   U7840 : INV_X1 port map( A => n11990, ZN => n11981);
   U7841 : INV_X1 port map( A => n12002, ZN => n11993);
   U7842 : INV_X1 port map( A => n12014, ZN => n12005);
   U7843 : INV_X1 port map( A => n12026, ZN => n12017);
   U7844 : INV_X1 port map( A => n12038, ZN => n12029);
   U7845 : INV_X1 port map( A => n12050, ZN => n12041);
   U7846 : INV_X1 port map( A => n12062, ZN => n12053);
   U7847 : INV_X1 port map( A => n12074, ZN => n12065);
   U7848 : INV_X1 port map( A => n12086, ZN => n12077);
   U7849 : INV_X1 port map( A => n12098, ZN => n12089);
   U7850 : INV_X1 port map( A => n12110, ZN => n12101);
   U7851 : INV_X1 port map( A => n12122, ZN => n12113);
   U7852 : INV_X1 port map( A => n12134, ZN => n12125);
   U7853 : INV_X1 port map( A => n12146, ZN => n12137);
   U7854 : INV_X1 port map( A => n12158, ZN => n12149);
   U7855 : INV_X1 port map( A => n12170, ZN => n12161);
   U7856 : INV_X1 port map( A => n12182, ZN => n12173);
   U7857 : INV_X1 port map( A => n12194, ZN => n12185);
   U7858 : INV_X1 port map( A => n12206, ZN => n12197);
   U7859 : INV_X1 port map( A => n12218, ZN => n12209);
   U7860 : INV_X1 port map( A => n12230, ZN => n12221);
   U7861 : INV_X1 port map( A => n12242, ZN => n12233);
   U7862 : INV_X1 port map( A => n12254, ZN => n12245);
   U7863 : INV_X1 port map( A => n12266, ZN => n12257);
   U7864 : INV_X1 port map( A => n12278, ZN => n12269);
   U7865 : INV_X1 port map( A => n12290, ZN => n12281);
   U7866 : INV_X1 port map( A => n12302, ZN => n12293);
   U7867 : INV_X1 port map( A => n12314, ZN => n12305);
   U7868 : INV_X1 port map( A => n12326, ZN => n12317);
   U7869 : INV_X1 port map( A => n12338, ZN => n12329);
   U7870 : INV_X1 port map( A => n12425, ZN => n12418);
   U7871 : INV_X1 port map( A => n12691, ZN => n12433);
   U7872 : INV_X1 port map( A => n12691, ZN => n12434);
   U7873 : INV_X1 port map( A => n12690, ZN => n12435);
   U7874 : INV_X1 port map( A => n12690, ZN => n12436);
   U7875 : INV_X1 port map( A => n12690, ZN => n12437);
   U7876 : INV_X1 port map( A => n12690, ZN => n12438);
   U7877 : INV_X1 port map( A => n12690, ZN => n12439);
   U7878 : INV_X1 port map( A => n12690, ZN => n12440);
   U7879 : INV_X1 port map( A => n12690, ZN => n12441);
   U7880 : INV_X1 port map( A => n12689, ZN => n12442);
   U7881 : INV_X1 port map( A => n12689, ZN => n12443);
   U7882 : INV_X1 port map( A => n12689, ZN => n12444);
   U7883 : INV_X1 port map( A => n12689, ZN => n12445);
   U7884 : INV_X1 port map( A => n12689, ZN => n12446);
   U7885 : INV_X1 port map( A => n12689, ZN => n12447);
   U7886 : INV_X1 port map( A => n12689, ZN => n12448);
   U7887 : INV_X1 port map( A => n12688, ZN => n12449);
   U7888 : INV_X1 port map( A => n12688, ZN => n12450);
   U7889 : INV_X1 port map( A => n12688, ZN => n12451);
   U7890 : INV_X1 port map( A => n12688, ZN => n12452);
   U7891 : INV_X1 port map( A => n12688, ZN => n12453);
   U7892 : INV_X1 port map( A => n12688, ZN => n12454);
   U7893 : INV_X1 port map( A => n12687, ZN => n12455);
   U7894 : INV_X1 port map( A => n12687, ZN => n12456);
   U7895 : INV_X1 port map( A => n12687, ZN => n12457);
   U7896 : INV_X1 port map( A => n12687, ZN => n12458);
   U7897 : INV_X1 port map( A => n12687, ZN => n12459);
   U7898 : INV_X1 port map( A => n12687, ZN => n12460);
   U7899 : INV_X1 port map( A => n12687, ZN => n12461);
   U7900 : INV_X1 port map( A => n12686, ZN => n12462);
   U7901 : INV_X1 port map( A => n12686, ZN => n12463);
   U7902 : INV_X1 port map( A => n12686, ZN => n12464);
   U7903 : INV_X1 port map( A => n12686, ZN => n12465);
   U7904 : INV_X1 port map( A => n12686, ZN => n12466);
   U7905 : INV_X1 port map( A => n12686, ZN => n12467);
   U7906 : INV_X1 port map( A => n12686, ZN => n12468);
   U7907 : INV_X1 port map( A => n12685, ZN => n12469);
   U7908 : INV_X1 port map( A => n12685, ZN => n12470);
   U7909 : INV_X1 port map( A => n12685, ZN => n12471);
   U7910 : INV_X1 port map( A => n12685, ZN => n12472);
   U7911 : INV_X1 port map( A => n12685, ZN => n12473);
   U7912 : INV_X1 port map( A => n12685, ZN => n12474);
   U7913 : INV_X1 port map( A => n12684, ZN => n12475);
   U7914 : INV_X1 port map( A => n12684, ZN => n12476);
   U7915 : INV_X1 port map( A => n12684, ZN => n12477);
   U7916 : INV_X1 port map( A => n12684, ZN => n12478);
   U7917 : INV_X1 port map( A => n12684, ZN => n12479);
   U7918 : INV_X1 port map( A => n12684, ZN => n12480);
   U7919 : INV_X1 port map( A => n12684, ZN => n12481);
   U7920 : INV_X1 port map( A => n12683, ZN => n12482);
   U7921 : INV_X1 port map( A => n12683, ZN => n12483);
   U7922 : INV_X1 port map( A => n12683, ZN => n12484);
   U7923 : INV_X1 port map( A => n12683, ZN => n12485);
   U7924 : INV_X1 port map( A => n12683, ZN => n12486);
   U7925 : INV_X1 port map( A => n12683, ZN => n12487);
   U7926 : INV_X1 port map( A => n12683, ZN => n12488);
   U7927 : INV_X1 port map( A => n12682, ZN => n12489);
   U7928 : INV_X1 port map( A => n12682, ZN => n12490);
   U7929 : INV_X1 port map( A => n12682, ZN => n12491);
   U7930 : INV_X1 port map( A => n12682, ZN => n12492);
   U7931 : INV_X1 port map( A => n12682, ZN => n12493);
   U7932 : INV_X1 port map( A => n12682, ZN => n12494);
   U7933 : INV_X1 port map( A => n12682, ZN => n12495);
   U7934 : INV_X1 port map( A => n12681, ZN => n12496);
   U7935 : INV_X1 port map( A => n12681, ZN => n12497);
   U7936 : INV_X1 port map( A => n12681, ZN => n12498);
   U7937 : INV_X1 port map( A => n12681, ZN => n12499);
   U7938 : INV_X1 port map( A => n12681, ZN => n12500);
   U7939 : INV_X1 port map( A => n12681, ZN => n12501);
   U7940 : INV_X1 port map( A => n12681, ZN => n12502);
   U7941 : INV_X1 port map( A => n12680, ZN => n12503);
   U7942 : INV_X1 port map( A => n12680, ZN => n12504);
   U7943 : INV_X1 port map( A => n12680, ZN => n12505);
   U7944 : INV_X1 port map( A => n12680, ZN => n12506);
   U7945 : INV_X1 port map( A => n12680, ZN => n12507);
   U7946 : INV_X1 port map( A => n12680, ZN => n12508);
   U7947 : INV_X1 port map( A => n12680, ZN => n12509);
   U7948 : INV_X1 port map( A => n12679, ZN => n12510);
   U7949 : INV_X1 port map( A => n12679, ZN => n12511);
   U7950 : INV_X1 port map( A => n12679, ZN => n12512);
   U7951 : INV_X1 port map( A => n12679, ZN => n12513);
   U7952 : INV_X1 port map( A => n12679, ZN => n12514);
   U7953 : INV_X1 port map( A => n12679, ZN => n12515);
   U7954 : INV_X1 port map( A => n12685, ZN => n12516);
   U7955 : INV_X1 port map( A => n12711, ZN => n12517);
   U7956 : INV_X1 port map( A => n12711, ZN => n12518);
   U7957 : INV_X1 port map( A => n12711, ZN => n12519);
   U7958 : INV_X1 port map( A => n12711, ZN => n12520);
   U7959 : INV_X1 port map( A => n12711, ZN => n12521);
   U7960 : INV_X1 port map( A => n12711, ZN => n12522);
   U7961 : INV_X1 port map( A => n12710, ZN => n12523);
   U7962 : INV_X1 port map( A => n12711, ZN => n12524);
   U7963 : INV_X1 port map( A => n12710, ZN => n12525);
   U7964 : INV_X1 port map( A => n12710, ZN => n12526);
   U7965 : INV_X1 port map( A => n12710, ZN => n12527);
   U7966 : INV_X1 port map( A => n12710, ZN => n12528);
   U7967 : INV_X1 port map( A => n12710, ZN => n12529);
   U7968 : INV_X1 port map( A => n12710, ZN => n12530);
   U7969 : INV_X1 port map( A => n12709, ZN => n12531);
   U7970 : INV_X1 port map( A => n12709, ZN => n12532);
   U7971 : INV_X1 port map( A => n12709, ZN => n12533);
   U7972 : INV_X1 port map( A => n12709, ZN => n12534);
   U7973 : INV_X1 port map( A => n12709, ZN => n12535);
   U7974 : INV_X1 port map( A => n12709, ZN => n12536);
   U7975 : INV_X1 port map( A => n12708, ZN => n12537);
   U7976 : INV_X1 port map( A => n12709, ZN => n12538);
   U7977 : INV_X1 port map( A => n12708, ZN => n12539);
   U7978 : INV_X1 port map( A => n12708, ZN => n12540);
   U7979 : INV_X1 port map( A => n12708, ZN => n12541);
   U7980 : INV_X1 port map( A => n12708, ZN => n12542);
   U7981 : INV_X1 port map( A => n12708, ZN => n12543);
   U7982 : INV_X1 port map( A => n12708, ZN => n12544);
   U7983 : INV_X1 port map( A => n12707, ZN => n12545);
   U7984 : INV_X1 port map( A => n12707, ZN => n12546);
   U7985 : INV_X1 port map( A => n12707, ZN => n12547);
   U7986 : INV_X1 port map( A => n12707, ZN => n12548);
   U7987 : INV_X1 port map( A => n12707, ZN => n12549);
   U7988 : INV_X1 port map( A => n12707, ZN => n12550);
   U7989 : INV_X1 port map( A => n12707, ZN => n12551);
   U7990 : INV_X1 port map( A => n12706, ZN => n12552);
   U7991 : INV_X1 port map( A => n12706, ZN => n12553);
   U7992 : INV_X1 port map( A => n12706, ZN => n12554);
   U7993 : INV_X1 port map( A => n12706, ZN => n12555);
   U7994 : INV_X1 port map( A => n12706, ZN => n12556);
   U7995 : INV_X1 port map( A => n12706, ZN => n12557);
   U7996 : INV_X1 port map( A => n12706, ZN => n12558);
   U7997 : INV_X1 port map( A => n12705, ZN => n12559);
   U7998 : INV_X1 port map( A => n12705, ZN => n12560);
   U7999 : INV_X1 port map( A => n12705, ZN => n12561);
   U8000 : INV_X1 port map( A => n12705, ZN => n12562);
   U8001 : INV_X1 port map( A => n12705, ZN => n12563);
   U8002 : INV_X1 port map( A => n12705, ZN => n12564);
   U8003 : INV_X1 port map( A => n12705, ZN => n12565);
   U8004 : INV_X1 port map( A => n12704, ZN => n12566);
   U8005 : INV_X1 port map( A => n12704, ZN => n12567);
   U8006 : INV_X1 port map( A => n12704, ZN => n12568);
   U8007 : INV_X1 port map( A => n12704, ZN => n12569);
   U8008 : INV_X1 port map( A => n12704, ZN => n12570);
   U8009 : INV_X1 port map( A => n12704, ZN => n12571);
   U8010 : INV_X1 port map( A => n12704, ZN => n12572);
   U8011 : INV_X1 port map( A => n12703, ZN => n12573);
   U8012 : INV_X1 port map( A => n12703, ZN => n12574);
   U8013 : INV_X1 port map( A => n12703, ZN => n12575);
   U8014 : INV_X1 port map( A => n12703, ZN => n12576);
   U8015 : INV_X1 port map( A => n12703, ZN => n12577);
   U8016 : INV_X1 port map( A => n12703, ZN => n12578);
   U8017 : INV_X1 port map( A => n12703, ZN => n12579);
   U8018 : INV_X1 port map( A => n12702, ZN => n12580);
   U8019 : INV_X1 port map( A => n12702, ZN => n12581);
   U8020 : INV_X1 port map( A => n12702, ZN => n12582);
   U8021 : INV_X1 port map( A => n12702, ZN => n12583);
   U8022 : INV_X1 port map( A => n12702, ZN => n12584);
   U8023 : INV_X1 port map( A => n12702, ZN => n12585);
   U8024 : INV_X1 port map( A => n12702, ZN => n12586);
   U8025 : INV_X1 port map( A => n12701, ZN => n12587);
   U8026 : INV_X1 port map( A => n12701, ZN => n12588);
   U8027 : INV_X1 port map( A => n12701, ZN => n12589);
   U8028 : INV_X1 port map( A => n12701, ZN => n12590);
   U8029 : INV_X1 port map( A => n12701, ZN => n12591);
   U8030 : INV_X1 port map( A => n12701, ZN => n12592);
   U8031 : INV_X1 port map( A => n12700, ZN => n12593);
   U8032 : INV_X1 port map( A => n12700, ZN => n12594);
   U8033 : INV_X1 port map( A => n12700, ZN => n12595);
   U8034 : INV_X1 port map( A => n12700, ZN => n12596);
   U8035 : INV_X1 port map( A => n12700, ZN => n12597);
   U8036 : INV_X1 port map( A => n12700, ZN => n12598);
   U8037 : INV_X1 port map( A => n12700, ZN => n12599);
   U8038 : INV_X1 port map( A => n12699, ZN => n12600);
   U8039 : INV_X1 port map( A => n12699, ZN => n12601);
   U8040 : INV_X1 port map( A => n12699, ZN => n12602);
   U8041 : INV_X1 port map( A => n12699, ZN => n12603);
   U8042 : INV_X1 port map( A => n12699, ZN => n12604);
   U8043 : INV_X1 port map( A => n12699, ZN => n12605);
   U8044 : INV_X1 port map( A => n12699, ZN => n12606);
   U8045 : INV_X1 port map( A => n12698, ZN => n12607);
   U8046 : INV_X1 port map( A => n12698, ZN => n12608);
   U8047 : INV_X1 port map( A => n12698, ZN => n12609);
   U8048 : INV_X1 port map( A => n12698, ZN => n12610);
   U8049 : INV_X1 port map( A => n12698, ZN => n12611);
   U8050 : INV_X1 port map( A => n12698, ZN => n12612);
   U8051 : INV_X1 port map( A => n12698, ZN => n12613);
   U8052 : INV_X1 port map( A => n12697, ZN => n12614);
   U8053 : INV_X1 port map( A => n12697, ZN => n12615);
   U8054 : INV_X1 port map( A => n12697, ZN => n12616);
   U8055 : INV_X1 port map( A => n12697, ZN => n12617);
   U8056 : INV_X1 port map( A => n12697, ZN => n12618);
   U8057 : INV_X1 port map( A => n12697, ZN => n12619);
   U8058 : INV_X1 port map( A => n12697, ZN => n12620);
   U8059 : INV_X1 port map( A => n12696, ZN => n12621);
   U8060 : INV_X1 port map( A => n12696, ZN => n12622);
   U8061 : INV_X1 port map( A => n12696, ZN => n12623);
   U8062 : INV_X1 port map( A => n12696, ZN => n12624);
   U8063 : INV_X1 port map( A => n12696, ZN => n12625);
   U8064 : INV_X1 port map( A => n12696, ZN => n12626);
   U8065 : INV_X1 port map( A => n12696, ZN => n12627);
   U8066 : INV_X1 port map( A => n12695, ZN => n12628);
   U8067 : INV_X1 port map( A => n12695, ZN => n12629);
   U8068 : INV_X1 port map( A => n12695, ZN => n12630);
   U8069 : INV_X1 port map( A => n12695, ZN => n12631);
   U8070 : INV_X1 port map( A => n12695, ZN => n12632);
   U8071 : INV_X1 port map( A => n12695, ZN => n12633);
   U8072 : INV_X1 port map( A => n12695, ZN => n12634);
   U8073 : INV_X1 port map( A => n12694, ZN => n12635);
   U8074 : INV_X1 port map( A => n12694, ZN => n12636);
   U8075 : INV_X1 port map( A => n12694, ZN => n12637);
   U8076 : INV_X1 port map( A => n12694, ZN => n12638);
   U8077 : INV_X1 port map( A => n12694, ZN => n12639);
   U8078 : INV_X1 port map( A => n12694, ZN => n12640);
   U8079 : INV_X1 port map( A => n12694, ZN => n12641);
   U8080 : INV_X1 port map( A => n12693, ZN => n12642);
   U8081 : INV_X1 port map( A => n12693, ZN => n12643);
   U8082 : INV_X1 port map( A => n12693, ZN => n12644);
   U8083 : INV_X1 port map( A => n12693, ZN => n12645);
   U8084 : INV_X1 port map( A => n12693, ZN => n12646);
   U8085 : INV_X1 port map( A => n12693, ZN => n12647);
   U8086 : INV_X1 port map( A => n12693, ZN => n12648);
   U8087 : INV_X1 port map( A => n12692, ZN => n12649);
   U8088 : INV_X1 port map( A => n12692, ZN => n12650);
   U8089 : INV_X1 port map( A => n12692, ZN => n12651);
   U8090 : INV_X1 port map( A => n12692, ZN => n12652);
   U8091 : INV_X1 port map( A => n12692, ZN => n12653);
   U8092 : INV_X1 port map( A => n12692, ZN => n12654);
   U8093 : INV_X1 port map( A => n12692, ZN => n12655);
   U8094 : INV_X1 port map( A => n12691, ZN => n12656);
   U8095 : INV_X1 port map( A => n12691, ZN => n12657);
   U8096 : INV_X1 port map( A => n12691, ZN => n12658);
   U8097 : INV_X1 port map( A => n12691, ZN => n12659);
   U8098 : INV_X1 port map( A => n12701, ZN => n12660);
   U8099 : INV_X1 port map( A => n12679, ZN => n12661);
   U8100 : INV_X1 port map( A => n12691, ZN => n12662);
   U8101 : AND2_X1 port map( A1 => r480_A_3_port, A2 => ADD_RD1(3), ZN => 
                           r480_carry_4_port);
   U8102 : XOR2_X1 port map( A => ADD_RD1(3), B => r480_A_3_port, Z => N8434);
   U8103 : AND2_X1 port map( A1 => r486_A_3_port, A2 => ADD_RD2(3), ZN => 
                           r486_carry_4_port);
   U8104 : XOR2_X1 port map( A => ADD_RD2(3), B => r486_A_3_port, Z => N8578);
   U8105 : AND2_X1 port map( A1 => ADD_WR(3), A2 => r472_B_3_port, ZN => 
                           r472_carry_4_port);
   U8106 : XOR2_X1 port map( A => r472_B_3_port, B => ADD_WR(3), Z => N2170);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IR_DECODE_NBIT32_opBIT6_regBIT5 is

   port( CLK : in std_logic;  IR_26 : in std_logic_vector (25 downto 0);  
         OPCODE : in std_logic_vector (5 downto 0);  is_signed : in std_logic; 
         RS1, RS2, RD : out std_logic_vector (4 downto 0);  IMMEDIATE : out 
         std_logic_vector (31 downto 0));

end IR_DECODE_NBIT32_opBIT6_regBIT5;

architecture SYN_BEHAV of IR_DECODE_NBIT32_opBIT6_regBIT5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component sign_eval_N_in26_N_out32
      port( IR_out : in std_logic_vector (25 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_eval_N_in16_N_out32
      port( IR_out : in std_logic_vector (15 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_eval_N_in5_N_out32
      port( IR_out : in std_logic_vector (4 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic0_port, IMMEDIATE_16_31_port, IMMEDIATE_16_15_port, 
      IMMEDIATE_16_14_port, IMMEDIATE_16_13_port, IMMEDIATE_16_12_port, 
      IMMEDIATE_16_11_port, IMMEDIATE_16_10_port, IMMEDIATE_16_9_port, 
      IMMEDIATE_16_8_port, IMMEDIATE_16_7_port, IMMEDIATE_16_6_port, 
      IMMEDIATE_16_5_port, IMMEDIATE_16_4_port, IMMEDIATE_16_3_port, 
      IMMEDIATE_16_2_port, IMMEDIATE_16_1_port, IMMEDIATE_16_0_port, n3, n4, n5
      , n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, 
      n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, 
      n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, 
      n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, 
      n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, 
      n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, 
      n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, 
      n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, 
      n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   RD_reg_4_inst : DLH_X1 port map( G => CLK, D => n34, Q => RD(4));
   RD_reg_3_inst : DLH_X1 port map( G => CLK, D => n35, Q => RD(3));
   RD_reg_2_inst : DLH_X1 port map( G => CLK, D => n36, Q => RD(2));
   RD_reg_1_inst : DLH_X1 port map( G => CLK, D => n37, Q => RD(1));
   RD_reg_0_inst : DLH_X1 port map( G => CLK, D => n38, Q => RD(0));
   IMMEDIATE_reg_31_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(31));
   IMMEDIATE_reg_30_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(30));
   IMMEDIATE_reg_29_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(29));
   IMMEDIATE_reg_28_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(28));
   IMMEDIATE_reg_27_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(27));
   IMMEDIATE_reg_26_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(26));
   IMMEDIATE_reg_25_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(25));
   IMMEDIATE_reg_24_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(24));
   IMMEDIATE_reg_23_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(23));
   IMMEDIATE_reg_22_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(22));
   IMMEDIATE_reg_21_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(21));
   IMMEDIATE_reg_20_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(20));
   IMMEDIATE_reg_19_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(19));
   IMMEDIATE_reg_18_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(18));
   IMMEDIATE_reg_17_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(17));
   IMMEDIATE_reg_16_inst : DLH_X1 port map( G => CLK, D => n33, Q => 
                           IMMEDIATE(16));
   IMMEDIATE_reg_15_inst : DLH_X1 port map( G => CLK, D => n18, Q => 
                           IMMEDIATE(15));
   IMMEDIATE_reg_14_inst : DLH_X1 port map( G => CLK, D => n17, Q => 
                           IMMEDIATE(14));
   IMMEDIATE_reg_13_inst : DLH_X1 port map( G => CLK, D => n16, Q => 
                           IMMEDIATE(13));
   IMMEDIATE_reg_12_inst : DLH_X1 port map( G => CLK, D => n15, Q => 
                           IMMEDIATE(12));
   IMMEDIATE_reg_11_inst : DLH_X1 port map( G => CLK, D => n14, Q => 
                           IMMEDIATE(11));
   IMMEDIATE_reg_10_inst : DLH_X1 port map( G => CLK, D => n13, Q => 
                           IMMEDIATE(10));
   IMMEDIATE_reg_9_inst : DLH_X1 port map( G => CLK, D => n12, Q => 
                           IMMEDIATE(9));
   IMMEDIATE_reg_8_inst : DLH_X1 port map( G => CLK, D => n11, Q => 
                           IMMEDIATE(8));
   IMMEDIATE_reg_7_inst : DLH_X1 port map( G => CLK, D => n10, Q => 
                           IMMEDIATE(7));
   IMMEDIATE_reg_6_inst : DLH_X1 port map( G => CLK, D => n9, Q => IMMEDIATE(6)
                           );
   IMMEDIATE_reg_5_inst : DLH_X1 port map( G => CLK, D => n8, Q => IMMEDIATE(5)
                           );
   IMMEDIATE_reg_4_inst : DLH_X1 port map( G => CLK, D => n7, Q => IMMEDIATE(4)
                           );
   IMMEDIATE_reg_3_inst : DLH_X1 port map( G => CLK, D => n6, Q => IMMEDIATE(3)
                           );
   IMMEDIATE_reg_2_inst : DLH_X1 port map( G => CLK, D => n5, Q => IMMEDIATE(2)
                           );
   IMMEDIATE_reg_1_inst : DLH_X1 port map( G => CLK, D => n4, Q => IMMEDIATE(1)
                           );
   IMMEDIATE_reg_0_inst : DLH_X1 port map( G => CLK, D => n3, Q => IMMEDIATE(0)
                           );
   RS1_reg_4_inst : DLH_X1 port map( G => CLK, D => IR_26(25), Q => RS1(4));
   RS1_reg_3_inst : DLH_X1 port map( G => CLK, D => IR_26(24), Q => RS1(3));
   RS1_reg_2_inst : DLH_X1 port map( G => CLK, D => IR_26(23), Q => RS1(2));
   RS1_reg_1_inst : DLH_X1 port map( G => CLK, D => IR_26(22), Q => RS1(1));
   RS1_reg_0_inst : DLH_X1 port map( G => CLK, D => IR_26(21), Q => RS1(0));
   RS2_reg_4_inst : DLH_X1 port map( G => CLK, D => IR_26(20), Q => RS2(4));
   RS2_reg_3_inst : DLH_X1 port map( G => CLK, D => IR_26(19), Q => RS2(3));
   RS2_reg_2_inst : DLH_X1 port map( G => CLK, D => IR_26(18), Q => RS2(2));
   RS2_reg_1_inst : DLH_X1 port map( G => CLK, D => IR_26(17), Q => RS2(1));
   RS2_reg_0_inst : DLH_X1 port map( G => CLK, D => IR_26(16), Q => RS2(0));
   SIGN_EXTENSION_imm5 : sign_eval_N_in5_N_out32 port map( IR_out(4) => 
                           IR_26(15), IR_out(3) => IR_26(14), IR_out(2) => 
                           IR_26(13), IR_out(1) => IR_26(12), IR_out(0) => 
                           IR_26(11), signed_val => is_signed, Immediate(31) =>
                           n_2966, Immediate(30) => n_2967, Immediate(29) => 
                           n_2968, Immediate(28) => n_2969, Immediate(27) => 
                           n_2970, Immediate(26) => n_2971, Immediate(25) => 
                           n_2972, Immediate(24) => n_2973, Immediate(23) => 
                           n_2974, Immediate(22) => n_2975, Immediate(21) => 
                           n_2976, Immediate(20) => n_2977, Immediate(19) => 
                           n_2978, Immediate(18) => n_2979, Immediate(17) => 
                           n_2980, Immediate(16) => n_2981, Immediate(15) => 
                           n_2982, Immediate(14) => n_2983, Immediate(13) => 
                           n_2984, Immediate(12) => n_2985, Immediate(11) => 
                           n_2986, Immediate(10) => n_2987, Immediate(9) => 
                           n_2988, Immediate(8) => n_2989, Immediate(7) => 
                           n_2990, Immediate(6) => n_2991, Immediate(5) => 
                           n_2992, Immediate(4) => n_2993, Immediate(3) => 
                           n_2994, Immediate(2) => n_2995, Immediate(1) => 
                           n_2996, Immediate(0) => n_2997);
   SIGN_EXTENSION_imm16 : sign_eval_N_in16_N_out32 port map( IR_out(15) => 
                           IR_26(15), IR_out(14) => IR_26(14), IR_out(13) => 
                           IR_26(13), IR_out(12) => IR_26(12), IR_out(11) => 
                           IR_26(11), IR_out(10) => IR_26(10), IR_out(9) => 
                           IR_26(9), IR_out(8) => IR_26(8), IR_out(7) => 
                           IR_26(7), IR_out(6) => IR_26(6), IR_out(5) => 
                           IR_26(5), IR_out(4) => IR_26(4), IR_out(3) => 
                           IR_26(3), IR_out(2) => IR_26(2), IR_out(1) => 
                           IR_26(1), IR_out(0) => IR_26(0), signed_val => 
                           is_signed, Immediate(31) => IMMEDIATE_16_31_port, 
                           Immediate(30) => n_2998, Immediate(29) => n_2999, 
                           Immediate(28) => n_3000, Immediate(27) => n_3001, 
                           Immediate(26) => n_3002, Immediate(25) => n_3003, 
                           Immediate(24) => n_3004, Immediate(23) => n_3005, 
                           Immediate(22) => n_3006, Immediate(21) => n_3007, 
                           Immediate(20) => n_3008, Immediate(19) => n_3009, 
                           Immediate(18) => n_3010, Immediate(17) => n_3011, 
                           Immediate(16) => n_3012, Immediate(15) => 
                           IMMEDIATE_16_15_port, Immediate(14) => 
                           IMMEDIATE_16_14_port, Immediate(13) => 
                           IMMEDIATE_16_13_port, Immediate(12) => 
                           IMMEDIATE_16_12_port, Immediate(11) => 
                           IMMEDIATE_16_11_port, Immediate(10) => 
                           IMMEDIATE_16_10_port, Immediate(9) => 
                           IMMEDIATE_16_9_port, Immediate(8) => 
                           IMMEDIATE_16_8_port, Immediate(7) => 
                           IMMEDIATE_16_7_port, Immediate(6) => 
                           IMMEDIATE_16_6_port, Immediate(5) => 
                           IMMEDIATE_16_5_port, Immediate(4) => 
                           IMMEDIATE_16_4_port, Immediate(3) => 
                           IMMEDIATE_16_3_port, Immediate(2) => 
                           IMMEDIATE_16_2_port, Immediate(1) => 
                           IMMEDIATE_16_1_port, Immediate(0) => 
                           IMMEDIATE_16_0_port);
   SIGN_EXTENSION_imm26 : sign_eval_N_in26_N_out32 port map( IR_out(25) => 
                           IR_26(25), IR_out(24) => IR_26(24), IR_out(23) => 
                           IR_26(23), IR_out(22) => IR_26(22), IR_out(21) => 
                           IR_26(21), IR_out(20) => IR_26(20), IR_out(19) => 
                           IR_26(19), IR_out(18) => IR_26(18), IR_out(17) => 
                           IR_26(17), IR_out(16) => IR_26(16), IR_out(15) => 
                           IR_26(15), IR_out(14) => IR_26(14), IR_out(13) => 
                           IR_26(13), IR_out(12) => IR_26(12), IR_out(11) => 
                           IR_26(11), IR_out(10) => IR_26(10), IR_out(9) => 
                           IR_26(9), IR_out(8) => IR_26(8), IR_out(7) => 
                           IR_26(7), IR_out(6) => IR_26(6), IR_out(5) => 
                           IR_26(5), IR_out(4) => IR_26(4), IR_out(3) => 
                           IR_26(3), IR_out(2) => IR_26(2), IR_out(1) => 
                           IR_26(1), IR_out(0) => IR_26(0), signed_val => 
                           X_Logic0_port, Immediate(31) => n_3013, 
                           Immediate(30) => n_3014, Immediate(29) => n_3015, 
                           Immediate(28) => n_3016, Immediate(27) => n_3017, 
                           Immediate(26) => n_3018, Immediate(25) => n_3019, 
                           Immediate(24) => n_3020, Immediate(23) => n_3021, 
                           Immediate(22) => n_3022, Immediate(21) => n_3023, 
                           Immediate(20) => n_3024, Immediate(19) => n_3025, 
                           Immediate(18) => n_3026, Immediate(17) => n_3027, 
                           Immediate(16) => n_3028, Immediate(15) => n_3029, 
                           Immediate(14) => n_3030, Immediate(13) => n_3031, 
                           Immediate(12) => n_3032, Immediate(11) => n_3033, 
                           Immediate(10) => n_3034, Immediate(9) => n_3035, 
                           Immediate(8) => n_3036, Immediate(7) => n_3037, 
                           Immediate(6) => n_3038, Immediate(5) => n_3039, 
                           Immediate(4) => n_3040, Immediate(3) => n_3041, 
                           Immediate(2) => n_3042, Immediate(1) => n_3043, 
                           Immediate(0) => n_3044);
   U3 : INV_X1 port map( A => n31, ZN => n20);
   U4 : INV_X1 port map( A => n31, ZN => n21);
   U5 : OR2_X2 port map( A1 => n29, A2 => n28, ZN => n31);
   U6 : OR2_X2 port map( A1 => n29, A2 => n28, ZN => n22);
   U7 : INV_X1 port map( A => n30, ZN => n33);
   U8 : NOR2_X1 port map( A1 => OPCODE(5), A2 => OPCODE(3), ZN => n25);
   U9 : NAND2_X1 port map( A1 => n27, A2 => n26, ZN => n28);
   U10 : INV_X1 port map( A => OPCODE(1), ZN => n26);
   U11 : INV_X1 port map( A => OPCODE(0), ZN => n27);
   U12 : INV_X1 port map( A => OPCODE(2), ZN => n23);
   U13 : INV_X1 port map( A => OPCODE(4), ZN => n24);
   U14 : NAND3_X1 port map( A1 => n25, A2 => n24, A3 => n23, ZN => n29);
   U15 : AND2_X1 port map( A1 => IMMEDIATE_16_0_port, A2 => n22, ZN => n3);
   U16 : AND2_X1 port map( A1 => IMMEDIATE_16_1_port, A2 => n22, ZN => n4);
   U17 : AND2_X1 port map( A1 => IMMEDIATE_16_2_port, A2 => n22, ZN => n5);
   U18 : AND2_X1 port map( A1 => IMMEDIATE_16_3_port, A2 => n22, ZN => n6);
   U19 : AND2_X1 port map( A1 => IMMEDIATE_16_4_port, A2 => n22, ZN => n7);
   U20 : AND2_X1 port map( A1 => IMMEDIATE_16_5_port, A2 => n22, ZN => n8);
   U21 : AND2_X1 port map( A1 => IMMEDIATE_16_6_port, A2 => n22, ZN => n9);
   U22 : AND2_X1 port map( A1 => IMMEDIATE_16_7_port, A2 => n22, ZN => n10);
   U23 : AND2_X1 port map( A1 => IMMEDIATE_16_8_port, A2 => n22, ZN => n11);
   U24 : AND2_X1 port map( A1 => IMMEDIATE_16_9_port, A2 => n22, ZN => n12);
   U25 : AND2_X1 port map( A1 => IMMEDIATE_16_10_port, A2 => n22, ZN => n13);
   U26 : AND2_X1 port map( A1 => IMMEDIATE_16_11_port, A2 => n22, ZN => n14);
   U27 : AND2_X1 port map( A1 => IMMEDIATE_16_12_port, A2 => n22, ZN => n15);
   U28 : AND2_X1 port map( A1 => IMMEDIATE_16_13_port, A2 => n22, ZN => n16);
   U29 : AND2_X1 port map( A1 => IMMEDIATE_16_14_port, A2 => n22, ZN => n17);
   U30 : AND2_X1 port map( A1 => IMMEDIATE_16_15_port, A2 => n22, ZN => n18);
   U31 : NAND2_X1 port map( A1 => n31, A2 => IMMEDIATE_16_31_port, ZN => n30);
   U32 : INV_X1 port map( A => n31, ZN => n32);
   U33 : MUX2_X1 port map( A => IR_26(16), B => IR_26(11), S => n32, Z => n38);
   U34 : MUX2_X1 port map( A => IR_26(17), B => IR_26(12), S => n32, Z => n37);
   U35 : MUX2_X1 port map( A => IR_26(18), B => IR_26(13), S => n20, Z => n36);
   U36 : MUX2_X1 port map( A => IR_26(19), B => IR_26(14), S => n21, Z => n35);
   U37 : MUX2_X1 port map( A => IR_26(20), B => IR_26(15), S => n20, Z => n34);

end SYN_BEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_0;

architecture SYN_struct of MUX21_GENERIC_NBIT32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_225
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_226
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_227
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_228
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_229
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_230
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_231
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_232
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_233
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_234
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_235
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_236
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_237
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_238
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_239
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_240
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_241
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_242
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_243
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_244
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_245
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_246
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_247
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_248
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_249
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_250
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_251
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_252
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_253
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_254
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_255
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   gen1_0 : MUX21_0 port map( A => A(0), B => B(0), S => n6, Y => Y(0));
   gen1_1 : MUX21_255 port map( A => A(1), B => B(1), S => n4, Y => Y(1));
   gen1_2 : MUX21_254 port map( A => A(2), B => B(2), S => n4, Y => Y(2));
   gen1_3 : MUX21_253 port map( A => A(3), B => B(3), S => n4, Y => Y(3));
   gen1_4 : MUX21_252 port map( A => A(4), B => B(4), S => n4, Y => Y(4));
   gen1_5 : MUX21_251 port map( A => A(5), B => B(5), S => n4, Y => Y(5));
   gen1_6 : MUX21_250 port map( A => A(6), B => B(6), S => n4, Y => Y(6));
   gen1_7 : MUX21_249 port map( A => A(7), B => B(7), S => n4, Y => Y(7));
   gen1_8 : MUX21_248 port map( A => A(8), B => B(8), S => n4, Y => Y(8));
   gen1_9 : MUX21_247 port map( A => A(9), B => B(9), S => n4, Y => Y(9));
   gen1_10 : MUX21_246 port map( A => A(10), B => B(10), S => n4, Y => Y(10));
   gen1_11 : MUX21_245 port map( A => A(11), B => B(11), S => n4, Y => Y(11));
   gen1_12 : MUX21_244 port map( A => A(12), B => B(12), S => n4, Y => Y(12));
   gen1_13 : MUX21_243 port map( A => A(13), B => B(13), S => n5, Y => Y(13));
   gen1_14 : MUX21_242 port map( A => A(14), B => B(14), S => n5, Y => Y(14));
   gen1_15 : MUX21_241 port map( A => A(15), B => B(15), S => n5, Y => Y(15));
   gen1_16 : MUX21_240 port map( A => A(16), B => B(16), S => n5, Y => Y(16));
   gen1_17 : MUX21_239 port map( A => A(17), B => B(17), S => n5, Y => Y(17));
   gen1_18 : MUX21_238 port map( A => A(18), B => B(18), S => n5, Y => Y(18));
   gen1_19 : MUX21_237 port map( A => A(19), B => B(19), S => n5, Y => Y(19));
   gen1_20 : MUX21_236 port map( A => A(20), B => B(20), S => n5, Y => Y(20));
   gen1_21 : MUX21_235 port map( A => A(21), B => B(21), S => n5, Y => Y(21));
   gen1_22 : MUX21_234 port map( A => A(22), B => B(22), S => n5, Y => Y(22));
   gen1_23 : MUX21_233 port map( A => A(23), B => B(23), S => n5, Y => Y(23));
   gen1_24 : MUX21_232 port map( A => A(24), B => B(24), S => n5, Y => Y(24));
   gen1_25 : MUX21_231 port map( A => A(25), B => B(25), S => n6, Y => Y(25));
   gen1_26 : MUX21_230 port map( A => A(26), B => B(26), S => n6, Y => Y(26));
   gen1_27 : MUX21_229 port map( A => A(27), B => B(27), S => n6, Y => Y(27));
   gen1_28 : MUX21_228 port map( A => A(28), B => B(28), S => n6, Y => Y(28));
   gen1_29 : MUX21_227 port map( A => A(29), B => B(29), S => n6, Y => Y(29));
   gen1_30 : MUX21_226 port map( A => A(30), B => B(30), S => n6, Y => Y(30));
   gen1_31 : MUX21_225 port map( A => A(31), B => B(31), S => n6, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n4);
   U2 : BUF_X1 port map( A => SEL, Z => n5);
   U3 : BUF_X1 port map( A => SEL, Z => n6);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => CK, RN => n97, Q => Q(31), 
                           QN => n65);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => CK, RN => n97, Q => Q(30), 
                           QN => n66);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => CK, RN => n97, Q => Q(29), 
                           QN => n67);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => CK, RN => n97, Q => Q(28), 
                           QN => n68);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => CK, RN => n97, Q => Q(27), 
                           QN => n69);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => CK, RN => n97, Q => Q(26), 
                           QN => n70);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => CK, RN => n97, Q => Q(25), 
                           QN => n71);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => CK, RN => n97, Q => Q(24), 
                           QN => n72);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => CK, RN => n97, Q => Q(23), 
                           QN => n73);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => CK, RN => n97, Q => Q(22),
                           QN => n74);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => CK, RN => n97, Q => Q(21),
                           QN => n75);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => CK, RN => n98, Q => Q(20),
                           QN => n76);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => CK, RN => n98, Q => Q(19),
                           QN => n77);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => CK, RN => n98, Q => Q(18),
                           QN => n78);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => CK, RN => n98, Q => Q(17),
                           QN => n79);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => CK, RN => n98, Q => Q(16),
                           QN => n80);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => CK, RN => n98, Q => Q(15),
                           QN => n81);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => CK, RN => n98, Q => Q(14),
                           QN => n82);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => CK, RN => n98, Q => Q(13),
                           QN => n83);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => CK, RN => n98, Q => Q(12),
                           QN => n84);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => CK, RN => n98, Q => Q(11),
                           QN => n85);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => CK, RN => n98, Q => Q(10),
                           QN => n86);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => CK, RN => n99, Q => Q(9), 
                           QN => n87);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => CK, RN => n99, Q => Q(8), 
                           QN => n88);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => CK, RN => n99, Q => Q(7), 
                           QN => n89);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => CK, RN => n99, Q => Q(6), 
                           QN => n90);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => CK, RN => n99, Q => Q(5), 
                           QN => n91);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => CK, RN => n99, Q => Q(4), 
                           QN => n92);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => CK, RN => n99, Q => Q(3), 
                           QN => n93);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => CK, RN => n99, Q => Q(2), 
                           QN => n94);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => CK, RN => n99, Q => Q(1), 
                           QN => n95);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => CK, RN => n99, Q => Q(0), 
                           QN => n96);
   U2 : BUF_X1 port map( A => RESET, Z => n98);
   U3 : BUF_X1 port map( A => RESET, Z => n97);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n96, B2 => ENABLE, A => n39, ZN => n32);
   U6 : NAND2_X1 port map( A1 => D(0), A2 => ENABLE, ZN => n39);
   U7 : OAI21_X1 port map( B1 => n95, B2 => ENABLE, A => n40, ZN => n31);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n40);
   U9 : OAI21_X1 port map( B1 => n94, B2 => ENABLE, A => n41, ZN => n30);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n41);
   U11 : OAI21_X1 port map( B1 => n93, B2 => ENABLE, A => n43, ZN => n29);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n43);
   U13 : OAI21_X1 port map( B1 => n92, B2 => ENABLE, A => n44, ZN => n28);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n44);
   U15 : OAI21_X1 port map( B1 => n91, B2 => ENABLE, A => n45, ZN => n27);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n45);
   U17 : OAI21_X1 port map( B1 => n90, B2 => ENABLE, A => n46, ZN => n26);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n46);
   U19 : OAI21_X1 port map( B1 => n89, B2 => ENABLE, A => n47, ZN => n25);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n47);
   U21 : OAI21_X1 port map( B1 => n88, B2 => ENABLE, A => n48, ZN => n24);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n48);
   U23 : OAI21_X1 port map( B1 => n87, B2 => ENABLE, A => n49, ZN => n23);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n49);
   U25 : OAI21_X1 port map( B1 => n86, B2 => ENABLE, A => n50, ZN => n22);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n50);
   U27 : OAI21_X1 port map( B1 => n85, B2 => ENABLE, A => n51, ZN => n21);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n51);
   U29 : OAI21_X1 port map( B1 => n84, B2 => ENABLE, A => n52, ZN => n20);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n52);
   U31 : OAI21_X1 port map( B1 => n83, B2 => ENABLE, A => n54, ZN => n19);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n54);
   U33 : OAI21_X1 port map( B1 => n82, B2 => ENABLE, A => n55, ZN => n18);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n55);
   U35 : OAI21_X1 port map( B1 => n81, B2 => ENABLE, A => n56, ZN => n17);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n56);
   U37 : OAI21_X1 port map( B1 => n80, B2 => ENABLE, A => n57, ZN => n16);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n57);
   U39 : OAI21_X1 port map( B1 => n79, B2 => ENABLE, A => n58, ZN => n15);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n58);
   U41 : OAI21_X1 port map( B1 => n78, B2 => ENABLE, A => n59, ZN => n14);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n59);
   U43 : OAI21_X1 port map( B1 => n77, B2 => ENABLE, A => n60, ZN => n13);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n60);
   U45 : OAI21_X1 port map( B1 => n76, B2 => ENABLE, A => n61, ZN => n12);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n61);
   U47 : OAI21_X1 port map( B1 => n75, B2 => ENABLE, A => n62, ZN => n11);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n62);
   U49 : OAI21_X1 port map( B1 => n74, B2 => ENABLE, A => n63, ZN => n10);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n63);
   U51 : OAI21_X1 port map( B1 => n73, B2 => ENABLE, A => n33, ZN => n9);
   U52 : NAND2_X1 port map( A1 => ENABLE, A2 => D(23), ZN => n33);
   U53 : OAI21_X1 port map( B1 => n72, B2 => ENABLE, A => n34, ZN => n8);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n34);
   U55 : OAI21_X1 port map( B1 => n71, B2 => ENABLE, A => n35, ZN => n7);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n35);
   U57 : OAI21_X1 port map( B1 => n70, B2 => ENABLE, A => n36, ZN => n6);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n36);
   U59 : OAI21_X1 port map( B1 => n69, B2 => ENABLE, A => n37, ZN => n5);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n37);
   U61 : OAI21_X1 port map( B1 => n68, B2 => ENABLE, A => n38, ZN => n4);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n38);
   U63 : OAI21_X1 port map( B1 => n67, B2 => ENABLE, A => n42, ZN => n3);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n42);
   U65 : OAI21_X1 port map( B1 => n66, B2 => ENABLE, A => n53, ZN => n2);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n53);
   U67 : OAI21_X1 port map( B1 => n65, B2 => ENABLE, A => n64, ZN => n1);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n64);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DATAPTH_NBIT32_REG_BIT5 is

   port( CLK, RST : in std_logic;  PC, IR : in std_logic_vector (31 downto 0); 
         PC_OUT : out std_logic_vector (31 downto 0);  NPC_LATCH_EN, 
         ir_LATCH_EN, signed_op, trap_cs, ret_cs, RF1, RF2, WF1, 
         regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond, sb_op, RM
         , WM, EN3, S3 : in std_logic;  instruction_alu : in std_logic_vector 
         (0 to 5);  DATA_MEM_ADDR, DATA_MEM_IN : out std_logic_vector (31 
         downto 0);  DATA_MEM_OUT : in std_logic_vector (31 downto 0);  
         DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM : out std_logic);

end DATAPTH_NBIT32_REG_BIT5;

architecture SYN_STRUCTURAL of DATAPTH_NBIT32_REG_BIT5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DATAPTH_NBIT32_REG_BIT5_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_1
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FF_2
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FF_3
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_2
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_3
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component load_data
      port( data_in : in std_logic_vector (31 downto 0);  signed_val, load_op :
            in std_logic;  load_type : in std_logic_vector (1 downto 0);  
            data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT6_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 
            downto 0);  Q : out std_logic_vector (5 downto 0));
   end component;
   
   component FF_4
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_2
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_4
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_5
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT32_5
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_6
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component COND_BT_NBIT32
      port( ZERO_BIT, OPCODE_0, branch_op : in std_logic;  con_sign : out 
            std_logic);
   end component;
   
   component zero_eval_NBIT32
      port( input : in std_logic_vector (31 downto 0);  res : out std_logic);
   end component;
   
   component ALU_N32
      port( CLK : in std_logic;  FUNC : in std_logic_vector (0 to 5);  DATA1, 
            DATA2 : in std_logic_vector (31 downto 0);  OUT_ALU : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_6
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_7
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT6_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 
            downto 0);  Q : out std_logic_vector (5 downto 0));
   end component;
   
   component FF_7
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_8
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_9
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_10
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_11
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_0
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component windRF_M8_N8_F5_NBIT32
      port( CLK, RESET, ENABLE, CALL, RETRN : in std_logic;  FILL, SPILL : out 
            std_logic;  BUSin : in std_logic_vector (31 downto 0);  BUSout : 
            out std_logic_vector (31 downto 0);  RD1, RD2, WR : in std_logic;  
            ADD_WR, ADD_RD1, ADD_RD2 : in std_logic_vector (4 downto 0);  
            DATAIN : in std_logic_vector (31 downto 0);  OUT1, OUT2 : out 
            std_logic_vector (31 downto 0);  wr_signal : in std_logic);
   end component;
   
   component IR_DECODE_NBIT32_opBIT6_regBIT5
      port( CLK : in std_logic;  IR_26 : in std_logic_vector (25 downto 0);  
            OPCODE : in std_logic_vector (5 downto 0);  is_signed : in 
            std_logic;  RS1, RS2, RD : out std_logic_vector (4 downto 0);  
            IMMEDIATE : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_12
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_13
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_14
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_15
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_16
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_17
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_18
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_19
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, PC_fetch0_31_port, PC_fetch0_30_port, 
      PC_fetch0_29_port, PC_fetch0_28_port, PC_fetch0_27_port, 
      PC_fetch0_26_port, PC_fetch0_25_port, PC_fetch0_24_port, 
      PC_fetch0_23_port, PC_fetch0_22_port, PC_fetch0_21_port, 
      PC_fetch0_20_port, PC_fetch0_19_port, PC_fetch0_18_port, 
      PC_fetch0_17_port, PC_fetch0_16_port, PC_fetch0_15_port, 
      PC_fetch0_14_port, PC_fetch0_13_port, PC_fetch0_12_port, 
      PC_fetch0_11_port, PC_fetch0_10_port, PC_fetch0_9_port, PC_fetch0_8_port,
      PC_fetch0_7_port, PC_fetch0_6_port, PC_fetch0_5_port, PC_fetch0_4_port, 
      PC_fetch0_3_port, PC_fetch0_2_port, PC_fetch0_1_port, PC_fetch0_0_port, 
      NPC_31_port, NPC_30_port, NPC_29_port, NPC_28_port, NPC_27_port, 
      NPC_26_port, NPC_25_port, NPC_24_port, NPC_23_port, NPC_22_port, 
      NPC_21_port, NPC_20_port, NPC_19_port, NPC_18_port, NPC_17_port, 
      NPC_16_port, NPC_15_port, NPC_14_port, NPC_13_port, NPC_12_port, 
      NPC_11_port, NPC_10_port, NPC_9_port, NPC_8_port, NPC_7_port, NPC_6_port,
      NPC_5_port, NPC_4_port, NPC_3_port, NPC_2_port, NPC_1_port, NPC_0_port, 
      NPC_fetch1_31_port, NPC_fetch1_30_port, NPC_fetch1_29_port, 
      NPC_fetch1_28_port, NPC_fetch1_27_port, NPC_fetch1_26_port, 
      NPC_fetch1_25_port, NPC_fetch1_24_port, NPC_fetch1_23_port, 
      NPC_fetch1_22_port, NPC_fetch1_21_port, NPC_fetch1_20_port, 
      NPC_fetch1_19_port, NPC_fetch1_18_port, NPC_fetch1_17_port, 
      NPC_fetch1_16_port, NPC_fetch1_15_port, NPC_fetch1_14_port, 
      NPC_fetch1_13_port, NPC_fetch1_12_port, NPC_fetch1_11_port, 
      NPC_fetch1_10_port, NPC_fetch1_9_port, NPC_fetch1_8_port, 
      NPC_fetch1_7_port, NPC_fetch1_6_port, NPC_fetch1_5_port, 
      NPC_fetch1_4_port, NPC_fetch1_3_port, NPC_fetch1_2_port, 
      NPC_fetch1_1_port, NPC_fetch1_0_port, PC_fetch1_31_port, 
      PC_fetch1_30_port, PC_fetch1_29_port, PC_fetch1_28_port, 
      PC_fetch1_27_port, PC_fetch1_26_port, PC_fetch1_25_port, 
      PC_fetch1_24_port, PC_fetch1_23_port, PC_fetch1_22_port, 
      PC_fetch1_21_port, PC_fetch1_20_port, PC_fetch1_19_port, 
      PC_fetch1_18_port, PC_fetch1_17_port, PC_fetch1_16_port, 
      PC_fetch1_15_port, PC_fetch1_14_port, PC_fetch1_13_port, 
      PC_fetch1_12_port, PC_fetch1_11_port, PC_fetch1_10_port, PC_fetch1_9_port
      , PC_fetch1_8_port, PC_fetch1_7_port, PC_fetch1_6_port, PC_fetch1_5_port,
      PC_fetch1_4_port, PC_fetch1_3_port, PC_fetch1_2_port, PC_fetch1_1_port, 
      PC_fetch1_0_port, PC_OUT_i_31_port, PC_OUT_i_30_port, PC_OUT_i_29_port, 
      PC_OUT_i_28_port, PC_OUT_i_27_port, PC_OUT_i_26_port, PC_OUT_i_25_port, 
      PC_OUT_i_24_port, PC_OUT_i_23_port, PC_OUT_i_22_port, PC_OUT_i_21_port, 
      PC_OUT_i_20_port, PC_OUT_i_19_port, PC_OUT_i_18_port, PC_OUT_i_17_port, 
      PC_OUT_i_16_port, PC_OUT_i_15_port, PC_OUT_i_14_port, PC_OUT_i_13_port, 
      PC_OUT_i_12_port, PC_OUT_i_11_port, PC_OUT_i_10_port, PC_OUT_i_9_port, 
      PC_OUT_i_8_port, PC_OUT_i_7_port, PC_OUT_i_6_port, PC_OUT_i_5_port, 
      PC_OUT_i_4_port, PC_OUT_i_3_port, PC_OUT_i_2_port, PC_OUT_i_1_port, 
      PC_OUT_i_0_port, sel_npc, NPC_fetch_31_port, NPC_fetch_30_port, 
      NPC_fetch_29_port, NPC_fetch_28_port, NPC_fetch_27_port, 
      NPC_fetch_26_port, NPC_fetch_25_port, NPC_fetch_24_port, 
      NPC_fetch_23_port, NPC_fetch_22_port, NPC_fetch_21_port, 
      NPC_fetch_20_port, NPC_fetch_19_port, NPC_fetch_18_port, 
      NPC_fetch_17_port, NPC_fetch_16_port, NPC_fetch_15_port, 
      NPC_fetch_14_port, NPC_fetch_13_port, NPC_fetch_12_port, 
      NPC_fetch_11_port, NPC_fetch_10_port, NPC_fetch_9_port, NPC_fetch_8_port,
      NPC_fetch_7_port, NPC_fetch_6_port, NPC_fetch_5_port, NPC_fetch_4_port, 
      NPC_fetch_3_port, NPC_fetch_2_port, NPC_fetch_1_port, NPC_fetch_0_port, 
      PC_fetch_31_port, PC_fetch_30_port, PC_fetch_29_port, PC_fetch_28_port, 
      PC_fetch_27_port, PC_fetch_26_port, PC_fetch_25_port, PC_fetch_24_port, 
      PC_fetch_23_port, PC_fetch_22_port, PC_fetch_21_port, PC_fetch_20_port, 
      PC_fetch_19_port, PC_fetch_18_port, PC_fetch_17_port, PC_fetch_16_port, 
      PC_fetch_15_port, PC_fetch_14_port, PC_fetch_13_port, PC_fetch_12_port, 
      PC_fetch_11_port, PC_fetch_10_port, PC_fetch_9_port, PC_fetch_8_port, 
      PC_fetch_7_port, PC_fetch_6_port, PC_fetch_5_port, PC_fetch_4_port, 
      PC_fetch_3_port, PC_fetch_2_port, PC_fetch_1_port, PC_fetch_0_port, 
      ir_fetch_31_port, ir_fetch_30_port, ir_fetch_29_port, ir_fetch_28_port, 
      ir_fetch_27_port, ir_fetch_26_port, ir_fetch_25_port, ir_fetch_24_port, 
      ir_fetch_23_port, ir_fetch_22_port, ir_fetch_21_port, ir_fetch_20_port, 
      ir_fetch_19_port, ir_fetch_18_port, ir_fetch_17_port, ir_fetch_16_port, 
      ir_fetch_15_port, ir_fetch_14_port, ir_fetch_13_port, ir_fetch_12_port, 
      ir_fetch_11_port, ir_fetch_10_port, ir_fetch_9_port, ir_fetch_8_port, 
      ir_fetch_7_port, ir_fetch_6_port, ir_fetch_5_port, ir_fetch_4_port, 
      ir_fetch_3_port, ir_fetch_2_port, ir_fetch_1_port, ir_fetch_0_port, 
      NPC_Dec_31_port, NPC_Dec_30_port, NPC_Dec_29_port, NPC_Dec_28_port, 
      NPC_Dec_27_port, NPC_Dec_26_port, NPC_Dec_25_port, NPC_Dec_24_port, 
      NPC_Dec_23_port, NPC_Dec_22_port, NPC_Dec_21_port, NPC_Dec_20_port, 
      NPC_Dec_19_port, NPC_Dec_18_port, NPC_Dec_17_port, NPC_Dec_16_port, 
      NPC_Dec_15_port, NPC_Dec_14_port, NPC_Dec_13_port, NPC_Dec_12_port, 
      NPC_Dec_11_port, NPC_Dec_10_port, NPC_Dec_9_port, NPC_Dec_8_port, 
      NPC_Dec_7_port, NPC_Dec_6_port, NPC_Dec_5_port, NPC_Dec_4_port, 
      NPC_Dec_3_port, NPC_Dec_2_port, NPC_Dec_1_port, NPC_Dec_0_port, 
      IR_Dec_31_port, IR_Dec_30_port, IR_Dec_29_port, IR_Dec_28_port, 
      IR_Dec_27_port, IR_Dec_26_port, IR_Dec_25_port, IR_Dec_24_port, 
      IR_Dec_23_port, IR_Dec_22_port, IR_Dec_21_port, IR_Dec_20_port, 
      IR_Dec_19_port, IR_Dec_18_port, IR_Dec_17_port, IR_Dec_16_port, 
      IR_Dec_15_port, IR_Dec_14_port, IR_Dec_13_port, IR_Dec_12_port, 
      IR_Dec_11_port, IR_Dec_10_port, IR_Dec_9_port, IR_Dec_8_port, 
      IR_Dec_7_port, IR_Dec_6_port, IR_Dec_5_port, IR_Dec_4_port, IR_Dec_3_port
      , IR_Dec_2_port, IR_Dec_1_port, IR_Dec_0_port, RS1_4_port, RS1_3_port, 
      RS1_2_port, RS1_1_port, RS1_0_port, RS2_4_port, RS2_3_port, RS2_2_port, 
      RS2_1_port, RS2_0_port, RD_4_port, RD_3_port, RD_2_port, RD_1_port, 
      RD_0_port, Imm_31_port, Imm_30_port, Imm_29_port, Imm_28_port, 
      Imm_27_port, Imm_26_port, Imm_25_port, Imm_24_port, Imm_23_port, 
      Imm_22_port, Imm_21_port, Imm_20_port, Imm_19_port, Imm_18_port, 
      Imm_17_port, Imm_16_port, Imm_15_port, Imm_14_port, Imm_13_port, 
      Imm_12_port, Imm_11_port, Imm_10_port, Imm_9_port, Imm_8_port, Imm_7_port
      , Imm_6_port, Imm_5_port, Imm_4_port, Imm_3_port, Imm_2_port, Imm_1_port,
      Imm_0_port, RD_wb_4_port, RD_wb_3_port, RD_wb_2_port, RD_wb_1_port, 
      RD_wb_0_port, OUT_wb_31_port, OUT_wb_30_port, OUT_wb_29_port, 
      OUT_wb_28_port, OUT_wb_27_port, OUT_wb_26_port, OUT_wb_25_port, 
      OUT_wb_24_port, OUT_wb_23_port, OUT_wb_22_port, OUT_wb_21_port, 
      OUT_wb_20_port, OUT_wb_19_port, OUT_wb_18_port, OUT_wb_17_port, 
      OUT_wb_16_port, OUT_wb_15_port, OUT_wb_14_port, OUT_wb_13_port, 
      OUT_wb_12_port, OUT_wb_11_port, OUT_wb_10_port, OUT_wb_9_port, 
      OUT_wb_8_port, OUT_wb_7_port, OUT_wb_6_port, OUT_wb_5_port, OUT_wb_4_port
      , OUT_wb_3_port, OUT_wb_2_port, OUT_wb_1_port, OUT_wb_0_port, 
      regA_31_port, regA_30_port, regA_29_port, regA_28_port, regA_27_port, 
      regA_26_port, regA_25_port, regA_24_port, regA_23_port, regA_22_port, 
      regA_21_port, regA_20_port, regA_19_port, regA_18_port, regA_17_port, 
      regA_16_port, regA_15_port, regA_14_port, regA_13_port, regA_12_port, 
      regA_11_port, regA_10_port, regA_9_port, regA_8_port, regA_7_port, 
      regA_6_port, regA_5_port, regA_4_port, regA_3_port, regA_2_port, 
      regA_1_port, regA_0_port, regB_31_port, regB_30_port, regB_29_port, 
      regB_28_port, regB_27_port, regB_26_port, regB_25_port, regB_24_port, 
      regB_23_port, regB_22_port, regB_21_port, regB_20_port, regB_19_port, 
      regB_18_port, regB_17_port, regB_16_port, regB_15_port, regB_14_port, 
      regB_13_port, regB_12_port, regB_11_port, regB_10_port, regB_9_port, 
      regB_8_port, regB_7_port, regB_6_port, regB_5_port, regB_4_port, 
      regB_3_port, regB_2_port, regB_1_port, regB_0_port, wr_signal_wb, 
      signed_op_ex, NPC_ex_31_port, NPC_ex_30_port, NPC_ex_29_port, 
      NPC_ex_28_port, NPC_ex_27_port, NPC_ex_26_port, NPC_ex_25_port, 
      NPC_ex_24_port, NPC_ex_23_port, NPC_ex_22_port, NPC_ex_21_port, 
      NPC_ex_20_port, NPC_ex_19_port, NPC_ex_18_port, NPC_ex_17_port, 
      NPC_ex_16_port, NPC_ex_15_port, NPC_ex_14_port, NPC_ex_13_port, 
      NPC_ex_12_port, NPC_ex_11_port, NPC_ex_10_port, NPC_ex_9_port, 
      NPC_ex_8_port, NPC_ex_7_port, NPC_ex_6_port, NPC_ex_5_port, NPC_ex_4_port
      , NPC_ex_3_port, NPC_ex_2_port, NPC_ex_1_port, NPC_ex_0_port, 
      regA_ex_31_port, regA_ex_30_port, regA_ex_29_port, regA_ex_28_port, 
      regA_ex_27_port, regA_ex_26_port, regA_ex_25_port, regA_ex_24_port, 
      regA_ex_23_port, regA_ex_22_port, regA_ex_21_port, regA_ex_20_port, 
      regA_ex_19_port, regA_ex_18_port, regA_ex_17_port, regA_ex_16_port, 
      regA_ex_15_port, regA_ex_14_port, regA_ex_13_port, regA_ex_12_port, 
      regA_ex_11_port, regA_ex_10_port, regA_ex_9_port, regA_ex_8_port, 
      regA_ex_7_port, regA_ex_6_port, regA_ex_5_port, regA_ex_4_port, 
      regA_ex_3_port, regA_ex_2_port, regA_ex_1_port, regA_ex_0_port, 
      regB_ex_31_port, regB_ex_30_port, regB_ex_29_port, regB_ex_28_port, 
      regB_ex_27_port, regB_ex_26_port, regB_ex_25_port, regB_ex_24_port, 
      regB_ex_23_port, regB_ex_22_port, regB_ex_21_port, regB_ex_20_port, 
      regB_ex_19_port, regB_ex_18_port, regB_ex_17_port, regB_ex_16_port, 
      regB_ex_15_port, regB_ex_14_port, regB_ex_13_port, regB_ex_12_port, 
      regB_ex_11_port, regB_ex_10_port, regB_ex_9_port, regB_ex_8_port, 
      regB_ex_7_port, regB_ex_6_port, regB_ex_5_port, regB_ex_4_port, 
      regB_ex_3_port, regB_ex_2_port, regB_ex_1_port, regB_ex_0_port, 
      Imm_ex_31_port, Imm_ex_30_port, Imm_ex_29_port, Imm_ex_28_port, 
      Imm_ex_27_port, Imm_ex_26_port, Imm_ex_25_port, Imm_ex_24_port, 
      Imm_ex_23_port, Imm_ex_22_port, Imm_ex_21_port, Imm_ex_20_port, 
      Imm_ex_19_port, Imm_ex_18_port, Imm_ex_17_port, Imm_ex_16_port, 
      Imm_ex_15_port, Imm_ex_14_port, Imm_ex_13_port, Imm_ex_12_port, 
      Imm_ex_11_port, Imm_ex_10_port, Imm_ex_9_port, Imm_ex_8_port, 
      Imm_ex_7_port, Imm_ex_6_port, Imm_ex_5_port, Imm_ex_4_port, Imm_ex_3_port
      , Imm_ex_2_port, Imm_ex_1_port, Imm_ex_0_port, RD_ex_4_port, RD_ex_3_port
      , RD_ex_2_port, RD_ex_1_port, RD_ex_0_port, wr_signal_exe, 
      IR_26_ex_5_port, IR_26_ex_4_port, IR_26_ex_3_port, IR_26_ex_2_port, 
      IR_26_ex_1_port, IR_26_ex_0_port, LHI_ex1_31_port, LHI_ex1_30_port, 
      LHI_ex1_29_port, LHI_ex1_28_port, LHI_ex1_27_port, LHI_ex1_26_port, 
      LHI_ex1_25_port, LHI_ex1_24_port, LHI_ex1_23_port, LHI_ex1_22_port, 
      LHI_ex1_21_port, LHI_ex1_20_port, LHI_ex1_19_port, LHI_ex1_18_port, 
      LHI_ex1_17_port, LHI_ex1_16_port, LHI_ex1_15_port, LHI_ex1_14_port, 
      LHI_ex1_13_port, LHI_ex1_12_port, LHI_ex1_11_port, LHI_ex1_10_port, 
      LHI_ex1_9_port, LHI_ex1_8_port, LHI_ex1_7_port, LHI_ex1_6_port, 
      LHI_ex1_5_port, LHI_ex1_4_port, LHI_ex1_3_port, LHI_ex1_2_port, 
      LHI_ex1_1_port, LHI_ex1_0_port, LHI_ex_31_port, LHI_ex_30_port, 
      LHI_ex_29_port, LHI_ex_28_port, LHI_ex_27_port, LHI_ex_26_port, 
      LHI_ex_25_port, LHI_ex_24_port, LHI_ex_23_port, LHI_ex_22_port, 
      LHI_ex_21_port, LHI_ex_20_port, LHI_ex_19_port, LHI_ex_18_port, 
      LHI_ex_17_port, LHI_ex_16_port, LHI_ex_15_port, LHI_ex_14_port, 
      LHI_ex_13_port, LHI_ex_12_port, LHI_ex_11_port, LHI_ex_10_port, 
      LHI_ex_9_port, LHI_ex_8_port, LHI_ex_7_port, LHI_ex_6_port, LHI_ex_5_port
      , LHI_ex_4_port, LHI_ex_3_port, LHI_ex_2_port, LHI_ex_1_port, 
      LHI_ex_0_port, input1_ALU_31_port, input1_ALU_30_port, input1_ALU_29_port
      , input1_ALU_28_port, input1_ALU_27_port, input1_ALU_26_port, 
      input1_ALU_25_port, input1_ALU_24_port, input1_ALU_23_port, 
      input1_ALU_22_port, input1_ALU_21_port, input1_ALU_20_port, 
      input1_ALU_19_port, input1_ALU_18_port, input1_ALU_17_port, 
      input1_ALU_16_port, input1_ALU_15_port, input1_ALU_14_port, 
      input1_ALU_13_port, input1_ALU_12_port, input1_ALU_11_port, 
      input1_ALU_10_port, input1_ALU_9_port, input1_ALU_8_port, 
      input1_ALU_7_port, input1_ALU_6_port, input1_ALU_5_port, 
      input1_ALU_4_port, input1_ALU_3_port, input1_ALU_2_port, 
      input1_ALU_1_port, input1_ALU_0_port, input2_ALU_31_port, 
      input2_ALU_30_port, input2_ALU_29_port, input2_ALU_28_port, 
      input2_ALU_27_port, input2_ALU_26_port, input2_ALU_25_port, 
      input2_ALU_24_port, input2_ALU_23_port, input2_ALU_22_port, 
      input2_ALU_21_port, input2_ALU_20_port, input2_ALU_19_port, 
      input2_ALU_18_port, input2_ALU_17_port, input2_ALU_16_port, 
      input2_ALU_15_port, input2_ALU_14_port, input2_ALU_13_port, 
      input2_ALU_12_port, input2_ALU_11_port, input2_ALU_10_port, 
      input2_ALU_9_port, input2_ALU_8_port, input2_ALU_7_port, 
      input2_ALU_6_port, input2_ALU_5_port, input2_ALU_4_port, 
      input2_ALU_3_port, input2_ALU_2_port, input2_ALU_1_port, 
      input2_ALU_0_port, ALU_out_31_port, ALU_out_30_port, ALU_out_29_port, 
      ALU_out_28_port, ALU_out_27_port, ALU_out_26_port, ALU_out_25_port, 
      ALU_out_24_port, ALU_out_23_port, ALU_out_22_port, ALU_out_21_port, 
      ALU_out_20_port, ALU_out_19_port, ALU_out_18_port, ALU_out_17_port, 
      ALU_out_16_port, ALU_out_15_port, ALU_out_14_port, ALU_out_13_port, 
      ALU_out_12_port, ALU_out_11_port, ALU_out_10_port, ALU_out_9_port, 
      ALU_out_8_port, ALU_out_7_port, ALU_out_6_port, ALU_out_5_port, 
      ALU_out_4_port, ALU_out_3_port, ALU_out_2_port, ALU_out_1_port, 
      ALU_out_0_port, is_zero, cond, ALU_ex_31_port, ALU_ex_30_port, 
      ALU_ex_29_port, ALU_ex_28_port, ALU_ex_27_port, ALU_ex_26_port, 
      ALU_ex_25_port, ALU_ex_24_port, ALU_ex_23_port, ALU_ex_22_port, 
      ALU_ex_21_port, ALU_ex_20_port, ALU_ex_19_port, ALU_ex_18_port, 
      ALU_ex_17_port, ALU_ex_16_port, ALU_ex_15_port, ALU_ex_14_port, 
      ALU_ex_13_port, ALU_ex_12_port, ALU_ex_11_port, ALU_ex_10_port, 
      ALU_ex_9_port, ALU_ex_8_port, ALU_ex_7_port, ALU_ex_6_port, ALU_ex_5_port
      , ALU_ex_4_port, ALU_ex_3_port, ALU_ex_2_port, ALU_ex_1_port, 
      ALU_ex_0_port, signed_op_mem, NPC_mem_31_port, NPC_mem_30_port, 
      NPC_mem_29_port, NPC_mem_28_port, NPC_mem_27_port, NPC_mem_26_port, 
      NPC_mem_25_port, NPC_mem_24_port, NPC_mem_23_port, NPC_mem_22_port, 
      NPC_mem_21_port, NPC_mem_20_port, NPC_mem_19_port, NPC_mem_18_port, 
      NPC_mem_17_port, NPC_mem_16_port, NPC_mem_15_port, NPC_mem_14_port, 
      NPC_mem_13_port, NPC_mem_12_port, NPC_mem_11_port, NPC_mem_10_port, 
      NPC_mem_9_port, NPC_mem_8_port, NPC_mem_7_port, NPC_mem_6_port, 
      NPC_mem_5_port, NPC_mem_4_port, NPC_mem_3_port, NPC_mem_2_port, 
      NPC_mem_1_port, NPC_mem_0_port, cond_mem, regB_mem_31_port, 
      regB_mem_30_port, regB_mem_29_port, regB_mem_28_port, regB_mem_27_port, 
      regB_mem_26_port, regB_mem_25_port, regB_mem_24_port, regB_mem_23_port, 
      regB_mem_22_port, regB_mem_21_port, regB_mem_20_port, regB_mem_19_port, 
      regB_mem_18_port, regB_mem_17_port, regB_mem_16_port, regB_mem_15_port, 
      regB_mem_14_port, regB_mem_13_port, regB_mem_12_port, regB_mem_11_port, 
      regB_mem_10_port, regB_mem_9_port, regB_mem_8_port, RD_mem_4_port, 
      RD_mem_3_port, RD_mem_2_port, RD_mem_1_port, RD_mem_0_port, wr_signal_mem
      , IR_26_mem_5_port, IR_26_mem_4_port, IR_26_mem_3_port, IR_26_mem_2_port,
      IR_26_mem_1_port, IR_26_mem_0_port, sel_saved_reg, N13, wr_signal_mem1, 
      LMD_out_31_port, LMD_out_30_port, LMD_out_29_port, LMD_out_28_port, 
      LMD_out_27_port, LMD_out_26_port, LMD_out_25_port, LMD_out_24_port, 
      LMD_out_23_port, LMD_out_22_port, LMD_out_21_port, LMD_out_20_port, 
      LMD_out_19_port, LMD_out_18_port, LMD_out_17_port, LMD_out_16_port, 
      LMD_out_15_port, LMD_out_14_port, LMD_out_13_port, LMD_out_12_port, 
      LMD_out_11_port, LMD_out_10_port, LMD_out_9_port, LMD_out_8_port, 
      LMD_out_7_port, LMD_out_6_port, LMD_out_5_port, LMD_out_4_port, 
      LMD_out_3_port, LMD_out_2_port, LMD_out_1_port, LMD_out_0_port, 
      ALU_wb_31_port, ALU_wb_30_port, ALU_wb_29_port, ALU_wb_28_port, 
      ALU_wb_27_port, ALU_wb_26_port, ALU_wb_25_port, ALU_wb_24_port, 
      ALU_wb_23_port, ALU_wb_22_port, ALU_wb_21_port, ALU_wb_20_port, 
      ALU_wb_19_port, ALU_wb_18_port, ALU_wb_17_port, ALU_wb_16_port, 
      ALU_wb_15_port, ALU_wb_14_port, ALU_wb_13_port, ALU_wb_12_port, 
      ALU_wb_11_port, ALU_wb_10_port, ALU_wb_9_port, ALU_wb_8_port, 
      ALU_wb_7_port, ALU_wb_6_port, ALU_wb_5_port, ALU_wb_4_port, ALU_wb_3_port
      , ALU_wb_2_port, ALU_wb_1_port, ALU_wb_0_port, LMD_wb_31_port, 
      LMD_wb_30_port, LMD_wb_29_port, LMD_wb_28_port, LMD_wb_27_port, 
      LMD_wb_26_port, LMD_wb_25_port, LMD_wb_24_port, LMD_wb_23_port, 
      LMD_wb_22_port, LMD_wb_21_port, LMD_wb_20_port, LMD_wb_19_port, 
      LMD_wb_18_port, LMD_wb_17_port, LMD_wb_16_port, LMD_wb_15_port, 
      LMD_wb_14_port, LMD_wb_13_port, LMD_wb_12_port, LMD_wb_11_port, 
      LMD_wb_10_port, LMD_wb_9_port, LMD_wb_8_port, LMD_wb_7_port, 
      LMD_wb_6_port, LMD_wb_5_port, LMD_wb_4_port, LMD_wb_3_port, LMD_wb_2_port
      , LMD_wb_1_port, LMD_wb_0_port, sel_saved_reg_wb, NPC_wb_31_port, 
      NPC_wb_30_port, NPC_wb_29_port, NPC_wb_28_port, NPC_wb_27_port, 
      NPC_wb_26_port, NPC_wb_25_port, NPC_wb_24_port, NPC_wb_23_port, 
      NPC_wb_22_port, NPC_wb_21_port, NPC_wb_20_port, NPC_wb_19_port, 
      NPC_wb_18_port, NPC_wb_17_port, NPC_wb_16_port, NPC_wb_15_port, 
      NPC_wb_14_port, NPC_wb_13_port, NPC_wb_12_port, NPC_wb_11_port, 
      NPC_wb_10_port, NPC_wb_9_port, NPC_wb_8_port, NPC_wb_7_port, 
      NPC_wb_6_port, NPC_wb_5_port, NPC_wb_4_port, NPC_wb_3_port, NPC_wb_2_port
      , NPC_wb_1_port, NPC_wb_0_port, OUT_data_31_port, OUT_data_30_port, 
      OUT_data_29_port, OUT_data_28_port, OUT_data_27_port, OUT_data_26_port, 
      OUT_data_25_port, OUT_data_24_port, OUT_data_23_port, OUT_data_22_port, 
      OUT_data_21_port, OUT_data_20_port, OUT_data_19_port, OUT_data_18_port, 
      OUT_data_17_port, OUT_data_16_port, OUT_data_15_port, OUT_data_14_port, 
      OUT_data_13_port, OUT_data_12_port, OUT_data_11_port, OUT_data_10_port, 
      OUT_data_9_port, OUT_data_8_port, OUT_data_7_port, OUT_data_6_port, 
      OUT_data_5_port, OUT_data_4_port, OUT_data_3_port, OUT_data_2_port, 
      OUT_data_1_port, OUT_data_0_port, n34, n11, n12, n13_port, n14, n15, n16,
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n_3045, n_3046, n_3047, n_3048, n_3049
      , n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058,
      n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, 
      n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, 
      n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, 
      n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, 
      n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, 
      n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111 : 
      std_logic;

begin
   DATA_MEM_RM <= RM;
   DATA_MEM_WM <= WM;
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   DATA_MEM_ADDR_reg_31_inst : DLH_X1 port map( G => n43, D => ALU_ex_31_port, 
                           Q => DATA_MEM_ADDR(31));
   DATA_MEM_ADDR_reg_30_inst : DLH_X1 port map( G => n42, D => ALU_ex_30_port, 
                           Q => DATA_MEM_ADDR(30));
   DATA_MEM_ADDR_reg_29_inst : DLH_X1 port map( G => n42, D => ALU_ex_29_port, 
                           Q => DATA_MEM_ADDR(29));
   DATA_MEM_ADDR_reg_28_inst : DLH_X1 port map( G => n42, D => ALU_ex_28_port, 
                           Q => DATA_MEM_ADDR(28));
   DATA_MEM_ADDR_reg_27_inst : DLH_X1 port map( G => n42, D => ALU_ex_27_port, 
                           Q => DATA_MEM_ADDR(27));
   DATA_MEM_ADDR_reg_26_inst : DLH_X1 port map( G => n41, D => ALU_ex_26_port, 
                           Q => DATA_MEM_ADDR(26));
   DATA_MEM_ADDR_reg_25_inst : DLH_X1 port map( G => n41, D => ALU_ex_25_port, 
                           Q => DATA_MEM_ADDR(25));
   DATA_MEM_ADDR_reg_24_inst : DLH_X1 port map( G => n41, D => ALU_ex_24_port, 
                           Q => DATA_MEM_ADDR(24));
   DATA_MEM_ADDR_reg_23_inst : DLH_X1 port map( G => n42, D => ALU_ex_23_port, 
                           Q => DATA_MEM_ADDR(23));
   DATA_MEM_ADDR_reg_22_inst : DLH_X1 port map( G => n41, D => ALU_ex_22_port, 
                           Q => DATA_MEM_ADDR(22));
   DATA_MEM_ADDR_reg_21_inst : DLH_X1 port map( G => n41, D => ALU_ex_21_port, 
                           Q => DATA_MEM_ADDR(21));
   DATA_MEM_ADDR_reg_20_inst : DLH_X1 port map( G => n40, D => ALU_ex_20_port, 
                           Q => DATA_MEM_ADDR(20));
   DATA_MEM_ADDR_reg_19_inst : DLH_X1 port map( G => n42, D => ALU_ex_19_port, 
                           Q => DATA_MEM_ADDR(19));
   DATA_MEM_ADDR_reg_18_inst : DLH_X1 port map( G => n40, D => ALU_ex_18_port, 
                           Q => DATA_MEM_ADDR(18));
   DATA_MEM_ADDR_reg_17_inst : DLH_X1 port map( G => n40, D => ALU_ex_17_port, 
                           Q => DATA_MEM_ADDR(17));
   DATA_MEM_ADDR_reg_16_inst : DLH_X1 port map( G => n40, D => ALU_ex_16_port, 
                           Q => DATA_MEM_ADDR(16));
   DATA_MEM_ADDR_reg_15_inst : DLH_X1 port map( G => n42, D => ALU_ex_15_port, 
                           Q => DATA_MEM_ADDR(15));
   DATA_MEM_ADDR_reg_14_inst : DLH_X1 port map( G => n40, D => ALU_ex_14_port, 
                           Q => DATA_MEM_ADDR(14));
   DATA_MEM_ADDR_reg_13_inst : DLH_X1 port map( G => n40, D => ALU_ex_13_port, 
                           Q => DATA_MEM_ADDR(13));
   DATA_MEM_ADDR_reg_12_inst : DLH_X1 port map( G => n40, D => ALU_ex_12_port, 
                           Q => DATA_MEM_ADDR(12));
   DATA_MEM_ADDR_reg_11_inst : DLH_X1 port map( G => n41, D => ALU_ex_11_port, 
                           Q => DATA_MEM_ADDR(11));
   DATA_MEM_ADDR_reg_10_inst : DLH_X1 port map( G => n41, D => ALU_ex_10_port, 
                           Q => DATA_MEM_ADDR(10));
   DATA_MEM_ADDR_reg_9_inst : DLH_X1 port map( G => n41, D => ALU_ex_9_port, Q 
                           => DATA_MEM_ADDR(9));
   DATA_MEM_ADDR_reg_8_inst : DLH_X1 port map( G => n41, D => ALU_ex_8_port, Q 
                           => DATA_MEM_ADDR(8));
   DATA_MEM_ADDR_reg_7_inst : DLH_X1 port map( G => n42, D => ALU_ex_7_port, Q 
                           => DATA_MEM_ADDR(7));
   DATA_MEM_ADDR_reg_6_inst : DLH_X1 port map( G => n42, D => ALU_ex_6_port, Q 
                           => DATA_MEM_ADDR(6));
   DATA_MEM_ADDR_reg_5_inst : DLH_X1 port map( G => n40, D => ALU_ex_5_port, Q 
                           => DATA_MEM_ADDR(5));
   DATA_MEM_ADDR_reg_4_inst : DLH_X1 port map( G => n40, D => ALU_ex_4_port, Q 
                           => DATA_MEM_ADDR(4));
   DATA_MEM_ADDR_reg_3_inst : DLH_X1 port map( G => n42, D => ALU_ex_3_port, Q 
                           => DATA_MEM_ADDR(3));
   DATA_MEM_ADDR_reg_2_inst : DLH_X1 port map( G => n41, D => ALU_ex_2_port, Q 
                           => DATA_MEM_ADDR(2));
   DATA_MEM_ADDR_reg_1_inst : DLH_X1 port map( G => n40, D => ALU_ex_1_port, Q 
                           => DATA_MEM_ADDR(1));
   DATA_MEM_ADDR_reg_0_inst : DLH_X1 port map( G => n43, D => ALU_ex_0_port, Q 
                           => DATA_MEM_ADDR(0));
   U62 : XOR2_X1 port map( A => IR_Dec_27_port, B => IR_Dec_26_port, Z => n15);
   U63 : NAND3_X1 port map( A1 => instruction_alu(3), A2 => instruction_alu(4),
                           A3 => instruction_alu(1), ZN => n31);
   pipeline_PCING : regFFD_NBIT32_0 port map( CK => CLK, RESET => n45, ENABLE 
                           => X_Logic1_port, D(31) => PC(31), D(30) => PC(30), 
                           D(29) => PC(29), D(28) => PC(28), D(27) => PC(27), 
                           D(26) => PC(26), D(25) => PC(25), D(24) => PC(24), 
                           D(23) => PC(23), D(22) => PC(22), D(21) => PC(21), 
                           D(20) => PC(20), D(19) => PC(19), D(18) => PC(18), 
                           D(17) => PC(17), D(16) => PC(16), D(15) => PC(15), 
                           D(14) => PC(14), D(13) => PC(13), D(12) => PC(12), 
                           D(11) => PC(11), D(10) => PC(10), D(9) => PC(9), 
                           D(8) => PC(8), D(7) => PC(7), D(6) => PC(6), D(5) =>
                           PC(5), D(4) => PC(4), D(3) => PC(3), D(2) => PC(2), 
                           D(1) => PC(1), D(0) => PC(0), Q(31) => 
                           PC_fetch0_31_port, Q(30) => PC_fetch0_30_port, Q(29)
                           => PC_fetch0_29_port, Q(28) => PC_fetch0_28_port, 
                           Q(27) => PC_fetch0_27_port, Q(26) => 
                           PC_fetch0_26_port, Q(25) => PC_fetch0_25_port, Q(24)
                           => PC_fetch0_24_port, Q(23) => PC_fetch0_23_port, 
                           Q(22) => PC_fetch0_22_port, Q(21) => 
                           PC_fetch0_21_port, Q(20) => PC_fetch0_20_port, Q(19)
                           => PC_fetch0_19_port, Q(18) => PC_fetch0_18_port, 
                           Q(17) => PC_fetch0_17_port, Q(16) => 
                           PC_fetch0_16_port, Q(15) => PC_fetch0_15_port, Q(14)
                           => PC_fetch0_14_port, Q(13) => PC_fetch0_13_port, 
                           Q(12) => PC_fetch0_12_port, Q(11) => 
                           PC_fetch0_11_port, Q(10) => PC_fetch0_10_port, Q(9) 
                           => PC_fetch0_9_port, Q(8) => PC_fetch0_8_port, Q(7) 
                           => PC_fetch0_7_port, Q(6) => PC_fetch0_6_port, Q(5) 
                           => PC_fetch0_5_port, Q(4) => PC_fetch0_4_port, Q(3) 
                           => PC_fetch0_3_port, Q(2) => PC_fetch0_2_port, Q(1) 
                           => PC_fetch0_1_port, Q(0) => PC_fetch0_0_port);
   pipeline_fetch1_NPC : regFFD_NBIT32_19 port map( CK => CLK, RESET => n45, 
                           ENABLE => NPC_LATCH_EN, D(31) => NPC_31_port, D(30) 
                           => NPC_30_port, D(29) => NPC_29_port, D(28) => 
                           NPC_28_port, D(27) => NPC_27_port, D(26) => 
                           NPC_26_port, D(25) => NPC_25_port, D(24) => 
                           NPC_24_port, D(23) => NPC_23_port, D(22) => 
                           NPC_22_port, D(21) => NPC_21_port, D(20) => 
                           NPC_20_port, D(19) => NPC_19_port, D(18) => 
                           NPC_18_port, D(17) => NPC_17_port, D(16) => 
                           NPC_16_port, D(15) => NPC_15_port, D(14) => 
                           NPC_14_port, D(13) => NPC_13_port, D(12) => 
                           NPC_12_port, D(11) => NPC_11_port, D(10) => 
                           NPC_10_port, D(9) => NPC_9_port, D(8) => NPC_8_port,
                           D(7) => NPC_7_port, D(6) => NPC_6_port, D(5) => 
                           NPC_5_port, D(4) => NPC_4_port, D(3) => NPC_3_port, 
                           D(2) => NPC_2_port, D(1) => NPC_1_port, D(0) => 
                           NPC_0_port, Q(31) => NPC_fetch1_31_port, Q(30) => 
                           NPC_fetch1_30_port, Q(29) => NPC_fetch1_29_port, 
                           Q(28) => NPC_fetch1_28_port, Q(27) => 
                           NPC_fetch1_27_port, Q(26) => NPC_fetch1_26_port, 
                           Q(25) => NPC_fetch1_25_port, Q(24) => 
                           NPC_fetch1_24_port, Q(23) => NPC_fetch1_23_port, 
                           Q(22) => NPC_fetch1_22_port, Q(21) => 
                           NPC_fetch1_21_port, Q(20) => NPC_fetch1_20_port, 
                           Q(19) => NPC_fetch1_19_port, Q(18) => 
                           NPC_fetch1_18_port, Q(17) => NPC_fetch1_17_port, 
                           Q(16) => NPC_fetch1_16_port, Q(15) => 
                           NPC_fetch1_15_port, Q(14) => NPC_fetch1_14_port, 
                           Q(13) => NPC_fetch1_13_port, Q(12) => 
                           NPC_fetch1_12_port, Q(11) => NPC_fetch1_11_port, 
                           Q(10) => NPC_fetch1_10_port, Q(9) => 
                           NPC_fetch1_9_port, Q(8) => NPC_fetch1_8_port, Q(7) 
                           => NPC_fetch1_7_port, Q(6) => NPC_fetch1_6_port, 
                           Q(5) => NPC_fetch1_5_port, Q(4) => NPC_fetch1_4_port
                           , Q(3) => NPC_fetch1_3_port, Q(2) => 
                           NPC_fetch1_2_port, Q(1) => NPC_fetch1_1_port, Q(0) 
                           => NPC_fetch1_0_port);
   pipeline_fetch1_PC : regFFD_NBIT32_18 port map( CK => CLK, RESET => n45, 
                           ENABLE => ir_LATCH_EN, D(31) => PC_fetch0_31_port, 
                           D(30) => PC_fetch0_30_port, D(29) => 
                           PC_fetch0_29_port, D(28) => PC_fetch0_28_port, D(27)
                           => PC_fetch0_27_port, D(26) => PC_fetch0_26_port, 
                           D(25) => PC_fetch0_25_port, D(24) => 
                           PC_fetch0_24_port, D(23) => PC_fetch0_23_port, D(22)
                           => PC_fetch0_22_port, D(21) => PC_fetch0_21_port, 
                           D(20) => PC_fetch0_20_port, D(19) => 
                           PC_fetch0_19_port, D(18) => PC_fetch0_18_port, D(17)
                           => PC_fetch0_17_port, D(16) => PC_fetch0_16_port, 
                           D(15) => PC_fetch0_15_port, D(14) => 
                           PC_fetch0_14_port, D(13) => PC_fetch0_13_port, D(12)
                           => PC_fetch0_12_port, D(11) => PC_fetch0_11_port, 
                           D(10) => PC_fetch0_10_port, D(9) => PC_fetch0_9_port
                           , D(8) => PC_fetch0_8_port, D(7) => PC_fetch0_7_port
                           , D(6) => PC_fetch0_6_port, D(5) => PC_fetch0_5_port
                           , D(4) => PC_fetch0_4_port, D(3) => PC_fetch0_3_port
                           , D(2) => PC_fetch0_2_port, D(1) => PC_fetch0_1_port
                           , D(0) => PC_fetch0_0_port, Q(31) => 
                           PC_fetch1_31_port, Q(30) => PC_fetch1_30_port, Q(29)
                           => PC_fetch1_29_port, Q(28) => PC_fetch1_28_port, 
                           Q(27) => PC_fetch1_27_port, Q(26) => 
                           PC_fetch1_26_port, Q(25) => PC_fetch1_25_port, Q(24)
                           => PC_fetch1_24_port, Q(23) => PC_fetch1_23_port, 
                           Q(22) => PC_fetch1_22_port, Q(21) => 
                           PC_fetch1_21_port, Q(20) => PC_fetch1_20_port, Q(19)
                           => PC_fetch1_19_port, Q(18) => PC_fetch1_18_port, 
                           Q(17) => PC_fetch1_17_port, Q(16) => 
                           PC_fetch1_16_port, Q(15) => PC_fetch1_15_port, Q(14)
                           => PC_fetch1_14_port, Q(13) => PC_fetch1_13_port, 
                           Q(12) => PC_fetch1_12_port, Q(11) => 
                           PC_fetch1_11_port, Q(10) => PC_fetch1_10_port, Q(9) 
                           => PC_fetch1_9_port, Q(8) => PC_fetch1_8_port, Q(7) 
                           => PC_fetch1_7_port, Q(6) => PC_fetch1_6_port, Q(5) 
                           => PC_fetch1_5_port, Q(4) => PC_fetch1_4_port, Q(3) 
                           => PC_fetch1_3_port, Q(2) => PC_fetch1_2_port, Q(1) 
                           => PC_fetch1_1_port, Q(0) => PC_fetch1_0_port);
   MUX_PC1 : MUX21_GENERIC_NBIT32_0 port map( A(31) => PC_OUT_i_31_port, A(30) 
                           => PC_OUT_i_30_port, A(29) => PC_OUT_i_29_port, 
                           A(28) => PC_OUT_i_28_port, A(27) => PC_OUT_i_27_port
                           , A(26) => PC_OUT_i_26_port, A(25) => 
                           PC_OUT_i_25_port, A(24) => PC_OUT_i_24_port, A(23) 
                           => PC_OUT_i_23_port, A(22) => PC_OUT_i_22_port, 
                           A(21) => PC_OUT_i_21_port, A(20) => PC_OUT_i_20_port
                           , A(19) => PC_OUT_i_19_port, A(18) => 
                           PC_OUT_i_18_port, A(17) => PC_OUT_i_17_port, A(16) 
                           => PC_OUT_i_16_port, A(15) => PC_OUT_i_15_port, 
                           A(14) => PC_OUT_i_14_port, A(13) => PC_OUT_i_13_port
                           , A(12) => PC_OUT_i_12_port, A(11) => 
                           PC_OUT_i_11_port, A(10) => PC_OUT_i_10_port, A(9) =>
                           PC_OUT_i_9_port, A(8) => PC_OUT_i_8_port, A(7) => 
                           PC_OUT_i_7_port, A(6) => PC_OUT_i_6_port, A(5) => 
                           PC_OUT_i_5_port, A(4) => PC_OUT_i_4_port, A(3) => 
                           PC_OUT_i_3_port, A(2) => PC_OUT_i_2_port, A(1) => 
                           PC_OUT_i_1_port, A(0) => PC_OUT_i_0_port, B(31) => 
                           NPC_fetch1_31_port, B(30) => NPC_fetch1_30_port, 
                           B(29) => NPC_fetch1_29_port, B(28) => 
                           NPC_fetch1_28_port, B(27) => NPC_fetch1_27_port, 
                           B(26) => NPC_fetch1_26_port, B(25) => 
                           NPC_fetch1_25_port, B(24) => NPC_fetch1_24_port, 
                           B(23) => NPC_fetch1_23_port, B(22) => 
                           NPC_fetch1_22_port, B(21) => NPC_fetch1_21_port, 
                           B(20) => NPC_fetch1_20_port, B(19) => 
                           NPC_fetch1_19_port, B(18) => NPC_fetch1_18_port, 
                           B(17) => NPC_fetch1_17_port, B(16) => 
                           NPC_fetch1_16_port, B(15) => NPC_fetch1_15_port, 
                           B(14) => NPC_fetch1_14_port, B(13) => 
                           NPC_fetch1_13_port, B(12) => NPC_fetch1_12_port, 
                           B(11) => NPC_fetch1_11_port, B(10) => 
                           NPC_fetch1_10_port, B(9) => NPC_fetch1_9_port, B(8) 
                           => NPC_fetch1_8_port, B(7) => NPC_fetch1_7_port, 
                           B(6) => NPC_fetch1_6_port, B(5) => NPC_fetch1_5_port
                           , B(4) => NPC_fetch1_4_port, B(3) => 
                           NPC_fetch1_3_port, B(2) => NPC_fetch1_2_port, B(1) 
                           => NPC_fetch1_1_port, B(0) => NPC_fetch1_0_port, SEL
                           => sel_npc, Y(31) => PC_OUT(31), Y(30) => PC_OUT(30)
                           , Y(29) => PC_OUT(29), Y(28) => PC_OUT(28), Y(27) =>
                           PC_OUT(27), Y(26) => PC_OUT(26), Y(25) => PC_OUT(25)
                           , Y(24) => PC_OUT(24), Y(23) => PC_OUT(23), Y(22) =>
                           PC_OUT(22), Y(21) => PC_OUT(21), Y(20) => PC_OUT(20)
                           , Y(19) => PC_OUT(19), Y(18) => PC_OUT(18), Y(17) =>
                           PC_OUT(17), Y(16) => PC_OUT(16), Y(15) => PC_OUT(15)
                           , Y(14) => PC_OUT(14), Y(13) => PC_OUT(13), Y(12) =>
                           PC_OUT(12), Y(11) => PC_OUT(11), Y(10) => PC_OUT(10)
                           , Y(9) => PC_OUT(9), Y(8) => PC_OUT(8), Y(7) => 
                           PC_OUT(7), Y(6) => PC_OUT(6), Y(5) => PC_OUT(5), 
                           Y(4) => PC_OUT(4), Y(3) => PC_OUT(3), Y(2) => 
                           PC_OUT(2), Y(1) => PC_OUT(1), Y(0) => PC_OUT(0));
   pipeline_fetch_NPC : regFFD_NBIT32_17 port map( CK => CLK, RESET => n45, 
                           ENABLE => NPC_LATCH_EN, D(31) => NPC_fetch1_31_port,
                           D(30) => NPC_fetch1_30_port, D(29) => 
                           NPC_fetch1_29_port, D(28) => NPC_fetch1_28_port, 
                           D(27) => NPC_fetch1_27_port, D(26) => 
                           NPC_fetch1_26_port, D(25) => NPC_fetch1_25_port, 
                           D(24) => NPC_fetch1_24_port, D(23) => 
                           NPC_fetch1_23_port, D(22) => NPC_fetch1_22_port, 
                           D(21) => NPC_fetch1_21_port, D(20) => 
                           NPC_fetch1_20_port, D(19) => NPC_fetch1_19_port, 
                           D(18) => NPC_fetch1_18_port, D(17) => 
                           NPC_fetch1_17_port, D(16) => NPC_fetch1_16_port, 
                           D(15) => NPC_fetch1_15_port, D(14) => 
                           NPC_fetch1_14_port, D(13) => NPC_fetch1_13_port, 
                           D(12) => NPC_fetch1_12_port, D(11) => 
                           NPC_fetch1_11_port, D(10) => NPC_fetch1_10_port, 
                           D(9) => NPC_fetch1_9_port, D(8) => NPC_fetch1_8_port
                           , D(7) => NPC_fetch1_7_port, D(6) => 
                           NPC_fetch1_6_port, D(5) => NPC_fetch1_5_port, D(4) 
                           => NPC_fetch1_4_port, D(3) => NPC_fetch1_3_port, 
                           D(2) => NPC_fetch1_2_port, D(1) => NPC_fetch1_1_port
                           , D(0) => NPC_fetch1_0_port, Q(31) => 
                           NPC_fetch_31_port, Q(30) => NPC_fetch_30_port, Q(29)
                           => NPC_fetch_29_port, Q(28) => NPC_fetch_28_port, 
                           Q(27) => NPC_fetch_27_port, Q(26) => 
                           NPC_fetch_26_port, Q(25) => NPC_fetch_25_port, Q(24)
                           => NPC_fetch_24_port, Q(23) => NPC_fetch_23_port, 
                           Q(22) => NPC_fetch_22_port, Q(21) => 
                           NPC_fetch_21_port, Q(20) => NPC_fetch_20_port, Q(19)
                           => NPC_fetch_19_port, Q(18) => NPC_fetch_18_port, 
                           Q(17) => NPC_fetch_17_port, Q(16) => 
                           NPC_fetch_16_port, Q(15) => NPC_fetch_15_port, Q(14)
                           => NPC_fetch_14_port, Q(13) => NPC_fetch_13_port, 
                           Q(12) => NPC_fetch_12_port, Q(11) => 
                           NPC_fetch_11_port, Q(10) => NPC_fetch_10_port, Q(9) 
                           => NPC_fetch_9_port, Q(8) => NPC_fetch_8_port, Q(7) 
                           => NPC_fetch_7_port, Q(6) => NPC_fetch_6_port, Q(5) 
                           => NPC_fetch_5_port, Q(4) => NPC_fetch_4_port, Q(3) 
                           => NPC_fetch_3_port, Q(2) => NPC_fetch_2_port, Q(1) 
                           => NPC_fetch_1_port, Q(0) => NPC_fetch_0_port);
   pipeline_fetch_PC : regFFD_NBIT32_16 port map( CK => CLK, RESET => n45, 
                           ENABLE => ir_LATCH_EN, D(31) => PC_fetch1_31_port, 
                           D(30) => PC_fetch1_30_port, D(29) => 
                           PC_fetch1_29_port, D(28) => PC_fetch1_28_port, D(27)
                           => PC_fetch1_27_port, D(26) => PC_fetch1_26_port, 
                           D(25) => PC_fetch1_25_port, D(24) => 
                           PC_fetch1_24_port, D(23) => PC_fetch1_23_port, D(22)
                           => PC_fetch1_22_port, D(21) => PC_fetch1_21_port, 
                           D(20) => PC_fetch1_20_port, D(19) => 
                           PC_fetch1_19_port, D(18) => PC_fetch1_18_port, D(17)
                           => PC_fetch1_17_port, D(16) => PC_fetch1_16_port, 
                           D(15) => PC_fetch1_15_port, D(14) => 
                           PC_fetch1_14_port, D(13) => PC_fetch1_13_port, D(12)
                           => PC_fetch1_12_port, D(11) => PC_fetch1_11_port, 
                           D(10) => PC_fetch1_10_port, D(9) => PC_fetch1_9_port
                           , D(8) => PC_fetch1_8_port, D(7) => PC_fetch1_7_port
                           , D(6) => PC_fetch1_6_port, D(5) => PC_fetch1_5_port
                           , D(4) => PC_fetch1_4_port, D(3) => PC_fetch1_3_port
                           , D(2) => PC_fetch1_2_port, D(1) => PC_fetch1_1_port
                           , D(0) => PC_fetch1_0_port, Q(31) => 
                           PC_fetch_31_port, Q(30) => PC_fetch_30_port, Q(29) 
                           => PC_fetch_29_port, Q(28) => PC_fetch_28_port, 
                           Q(27) => PC_fetch_27_port, Q(26) => PC_fetch_26_port
                           , Q(25) => PC_fetch_25_port, Q(24) => 
                           PC_fetch_24_port, Q(23) => PC_fetch_23_port, Q(22) 
                           => PC_fetch_22_port, Q(21) => PC_fetch_21_port, 
                           Q(20) => PC_fetch_20_port, Q(19) => PC_fetch_19_port
                           , Q(18) => PC_fetch_18_port, Q(17) => 
                           PC_fetch_17_port, Q(16) => PC_fetch_16_port, Q(15) 
                           => PC_fetch_15_port, Q(14) => PC_fetch_14_port, 
                           Q(13) => PC_fetch_13_port, Q(12) => PC_fetch_12_port
                           , Q(11) => PC_fetch_11_port, Q(10) => 
                           PC_fetch_10_port, Q(9) => PC_fetch_9_port, Q(8) => 
                           PC_fetch_8_port, Q(7) => PC_fetch_7_port, Q(6) => 
                           PC_fetch_6_port, Q(5) => PC_fetch_5_port, Q(4) => 
                           PC_fetch_4_port, Q(3) => PC_fetch_3_port, Q(2) => 
                           PC_fetch_2_port, Q(1) => PC_fetch_1_port, Q(0) => 
                           PC_fetch_0_port);
   pipeline_fetch_ir : regFFD_NBIT32_15 port map( CK => CLK, RESET => n45, 
                           ENABLE => ir_LATCH_EN, D(31) => IR(31), D(30) => 
                           IR(30), D(29) => IR(29), D(28) => IR(28), D(27) => 
                           IR(27), D(26) => IR(26), D(25) => IR(25), D(24) => 
                           IR(24), D(23) => IR(23), D(22) => IR(22), D(21) => 
                           IR(21), D(20) => IR(20), D(19) => IR(19), D(18) => 
                           IR(18), D(17) => IR(17), D(16) => IR(16), D(15) => 
                           IR(15), D(14) => IR(14), D(13) => IR(13), D(12) => 
                           IR(12), D(11) => IR(11), D(10) => IR(10), D(9) => 
                           IR(9), D(8) => IR(8), D(7) => IR(7), D(6) => IR(6), 
                           D(5) => IR(5), D(4) => IR(4), D(3) => IR(3), D(2) =>
                           IR(2), D(1) => IR(1), D(0) => IR(0), Q(31) => 
                           ir_fetch_31_port, Q(30) => ir_fetch_30_port, Q(29) 
                           => ir_fetch_29_port, Q(28) => ir_fetch_28_port, 
                           Q(27) => ir_fetch_27_port, Q(26) => ir_fetch_26_port
                           , Q(25) => ir_fetch_25_port, Q(24) => 
                           ir_fetch_24_port, Q(23) => ir_fetch_23_port, Q(22) 
                           => ir_fetch_22_port, Q(21) => ir_fetch_21_port, 
                           Q(20) => ir_fetch_20_port, Q(19) => ir_fetch_19_port
                           , Q(18) => ir_fetch_18_port, Q(17) => 
                           ir_fetch_17_port, Q(16) => ir_fetch_16_port, Q(15) 
                           => ir_fetch_15_port, Q(14) => ir_fetch_14_port, 
                           Q(13) => ir_fetch_13_port, Q(12) => ir_fetch_12_port
                           , Q(11) => ir_fetch_11_port, Q(10) => 
                           ir_fetch_10_port, Q(9) => ir_fetch_9_port, Q(8) => 
                           ir_fetch_8_port, Q(7) => ir_fetch_7_port, Q(6) => 
                           ir_fetch_6_port, Q(5) => ir_fetch_5_port, Q(4) => 
                           ir_fetch_4_port, Q(3) => ir_fetch_3_port, Q(2) => 
                           ir_fetch_2_port, Q(1) => ir_fetch_1_port, Q(0) => 
                           ir_fetch_0_port);
   pipeline_newpc1 : regFFD_NBIT32_14 port map( CK => CLK, RESET => n45, ENABLE
                           => NPC_LATCH_EN, D(31) => NPC_fetch_31_port, D(30) 
                           => NPC_fetch_30_port, D(29) => NPC_fetch_29_port, 
                           D(28) => NPC_fetch_28_port, D(27) => 
                           NPC_fetch_27_port, D(26) => NPC_fetch_26_port, D(25)
                           => NPC_fetch_25_port, D(24) => NPC_fetch_24_port, 
                           D(23) => NPC_fetch_23_port, D(22) => 
                           NPC_fetch_22_port, D(21) => NPC_fetch_21_port, D(20)
                           => NPC_fetch_20_port, D(19) => NPC_fetch_19_port, 
                           D(18) => NPC_fetch_18_port, D(17) => 
                           NPC_fetch_17_port, D(16) => NPC_fetch_16_port, D(15)
                           => NPC_fetch_15_port, D(14) => NPC_fetch_14_port, 
                           D(13) => NPC_fetch_13_port, D(12) => 
                           NPC_fetch_12_port, D(11) => NPC_fetch_11_port, D(10)
                           => NPC_fetch_10_port, D(9) => NPC_fetch_9_port, D(8)
                           => NPC_fetch_8_port, D(7) => NPC_fetch_7_port, D(6) 
                           => NPC_fetch_6_port, D(5) => NPC_fetch_5_port, D(4) 
                           => NPC_fetch_4_port, D(3) => NPC_fetch_3_port, D(2) 
                           => NPC_fetch_2_port, D(1) => NPC_fetch_1_port, D(0) 
                           => NPC_fetch_0_port, Q(31) => NPC_Dec_31_port, Q(30)
                           => NPC_Dec_30_port, Q(29) => NPC_Dec_29_port, Q(28) 
                           => NPC_Dec_28_port, Q(27) => NPC_Dec_27_port, Q(26) 
                           => NPC_Dec_26_port, Q(25) => NPC_Dec_25_port, Q(24) 
                           => NPC_Dec_24_port, Q(23) => NPC_Dec_23_port, Q(22) 
                           => NPC_Dec_22_port, Q(21) => NPC_Dec_21_port, Q(20) 
                           => NPC_Dec_20_port, Q(19) => NPC_Dec_19_port, Q(18) 
                           => NPC_Dec_18_port, Q(17) => NPC_Dec_17_port, Q(16) 
                           => NPC_Dec_16_port, Q(15) => NPC_Dec_15_port, Q(14) 
                           => NPC_Dec_14_port, Q(13) => NPC_Dec_13_port, Q(12) 
                           => NPC_Dec_12_port, Q(11) => NPC_Dec_11_port, Q(10) 
                           => NPC_Dec_10_port, Q(9) => NPC_Dec_9_port, Q(8) => 
                           NPC_Dec_8_port, Q(7) => NPC_Dec_7_port, Q(6) => 
                           NPC_Dec_6_port, Q(5) => NPC_Dec_5_port, Q(4) => 
                           NPC_Dec_4_port, Q(3) => NPC_Dec_3_port, Q(2) => 
                           NPC_Dec_2_port, Q(1) => NPC_Dec_1_port, Q(0) => 
                           NPC_Dec_0_port);
   pipeline_pc1 : regFFD_NBIT32_13 port map( CK => CLK, RESET => n45, ENABLE =>
                           ir_LATCH_EN, D(31) => PC_fetch_31_port, D(30) => 
                           PC_fetch_30_port, D(29) => PC_fetch_29_port, D(28) 
                           => PC_fetch_28_port, D(27) => PC_fetch_27_port, 
                           D(26) => PC_fetch_26_port, D(25) => PC_fetch_25_port
                           , D(24) => PC_fetch_24_port, D(23) => 
                           PC_fetch_23_port, D(22) => PC_fetch_22_port, D(21) 
                           => PC_fetch_21_port, D(20) => PC_fetch_20_port, 
                           D(19) => PC_fetch_19_port, D(18) => PC_fetch_18_port
                           , D(17) => PC_fetch_17_port, D(16) => 
                           PC_fetch_16_port, D(15) => PC_fetch_15_port, D(14) 
                           => PC_fetch_14_port, D(13) => PC_fetch_13_port, 
                           D(12) => PC_fetch_12_port, D(11) => PC_fetch_11_port
                           , D(10) => PC_fetch_10_port, D(9) => PC_fetch_9_port
                           , D(8) => PC_fetch_8_port, D(7) => PC_fetch_7_port, 
                           D(6) => PC_fetch_6_port, D(5) => PC_fetch_5_port, 
                           D(4) => PC_fetch_4_port, D(3) => PC_fetch_3_port, 
                           D(2) => PC_fetch_2_port, D(1) => PC_fetch_1_port, 
                           D(0) => PC_fetch_0_port, Q(31) => n_3045, Q(30) => 
                           n_3046, Q(29) => n_3047, Q(28) => n_3048, Q(27) => 
                           n_3049, Q(26) => n_3050, Q(25) => n_3051, Q(24) => 
                           n_3052, Q(23) => n_3053, Q(22) => n_3054, Q(21) => 
                           n_3055, Q(20) => n_3056, Q(19) => n_3057, Q(18) => 
                           n_3058, Q(17) => n_3059, Q(16) => n_3060, Q(15) => 
                           n_3061, Q(14) => n_3062, Q(13) => n_3063, Q(12) => 
                           n_3064, Q(11) => n_3065, Q(10) => n_3066, Q(9) => 
                           n_3067, Q(8) => n_3068, Q(7) => n_3069, Q(6) => 
                           n_3070, Q(5) => n_3071, Q(4) => n_3072, Q(3) => 
                           n_3073, Q(2) => n_3074, Q(1) => n_3075, Q(0) => 
                           n_3076);
   pipeline_IR1 : regFFD_NBIT32_12 port map( CK => CLK, RESET => n45, ENABLE =>
                           ir_LATCH_EN, D(31) => ir_fetch_31_port, D(30) => 
                           ir_fetch_30_port, D(29) => ir_fetch_29_port, D(28) 
                           => ir_fetch_28_port, D(27) => ir_fetch_27_port, 
                           D(26) => ir_fetch_26_port, D(25) => ir_fetch_25_port
                           , D(24) => ir_fetch_24_port, D(23) => 
                           ir_fetch_23_port, D(22) => ir_fetch_22_port, D(21) 
                           => ir_fetch_21_port, D(20) => ir_fetch_20_port, 
                           D(19) => ir_fetch_19_port, D(18) => ir_fetch_18_port
                           , D(17) => ir_fetch_17_port, D(16) => 
                           ir_fetch_16_port, D(15) => ir_fetch_15_port, D(14) 
                           => ir_fetch_14_port, D(13) => ir_fetch_13_port, 
                           D(12) => ir_fetch_12_port, D(11) => ir_fetch_11_port
                           , D(10) => ir_fetch_10_port, D(9) => ir_fetch_9_port
                           , D(8) => ir_fetch_8_port, D(7) => ir_fetch_7_port, 
                           D(6) => ir_fetch_6_port, D(5) => ir_fetch_5_port, 
                           D(4) => ir_fetch_4_port, D(3) => ir_fetch_3_port, 
                           D(2) => ir_fetch_2_port, D(1) => ir_fetch_1_port, 
                           D(0) => ir_fetch_0_port, Q(31) => IR_Dec_31_port, 
                           Q(30) => IR_Dec_30_port, Q(29) => IR_Dec_29_port, 
                           Q(28) => IR_Dec_28_port, Q(27) => IR_Dec_27_port, 
                           Q(26) => IR_Dec_26_port, Q(25) => IR_Dec_25_port, 
                           Q(24) => IR_Dec_24_port, Q(23) => IR_Dec_23_port, 
                           Q(22) => IR_Dec_22_port, Q(21) => IR_Dec_21_port, 
                           Q(20) => IR_Dec_20_port, Q(19) => IR_Dec_19_port, 
                           Q(18) => IR_Dec_18_port, Q(17) => IR_Dec_17_port, 
                           Q(16) => IR_Dec_16_port, Q(15) => IR_Dec_15_port, 
                           Q(14) => IR_Dec_14_port, Q(13) => IR_Dec_13_port, 
                           Q(12) => IR_Dec_12_port, Q(11) => IR_Dec_11_port, 
                           Q(10) => IR_Dec_10_port, Q(9) => IR_Dec_9_port, Q(8)
                           => IR_Dec_8_port, Q(7) => IR_Dec_7_port, Q(6) => 
                           IR_Dec_6_port, Q(5) => IR_Dec_5_port, Q(4) => 
                           IR_Dec_4_port, Q(3) => IR_Dec_3_port, Q(2) => 
                           IR_Dec_2_port, Q(1) => IR_Dec_1_port, Q(0) => 
                           IR_Dec_0_port);
   IR_OP : IR_DECODE_NBIT32_opBIT6_regBIT5 port map( CLK => CLK, IR_26(25) => 
                           IR_Dec_25_port, IR_26(24) => IR_Dec_24_port, 
                           IR_26(23) => IR_Dec_23_port, IR_26(22) => 
                           IR_Dec_22_port, IR_26(21) => IR_Dec_21_port, 
                           IR_26(20) => IR_Dec_20_port, IR_26(19) => 
                           IR_Dec_19_port, IR_26(18) => IR_Dec_18_port, 
                           IR_26(17) => IR_Dec_17_port, IR_26(16) => 
                           IR_Dec_16_port, IR_26(15) => IR_Dec_15_port, 
                           IR_26(14) => IR_Dec_14_port, IR_26(13) => 
                           IR_Dec_13_port, IR_26(12) => IR_Dec_12_port, 
                           IR_26(11) => IR_Dec_11_port, IR_26(10) => 
                           IR_Dec_10_port, IR_26(9) => IR_Dec_9_port, IR_26(8) 
                           => IR_Dec_8_port, IR_26(7) => IR_Dec_7_port, 
                           IR_26(6) => IR_Dec_6_port, IR_26(5) => IR_Dec_5_port
                           , IR_26(4) => IR_Dec_4_port, IR_26(3) => 
                           IR_Dec_3_port, IR_26(2) => IR_Dec_2_port, IR_26(1) 
                           => IR_Dec_1_port, IR_26(0) => IR_Dec_0_port, 
                           OPCODE(5) => IR_Dec_31_port, OPCODE(4) => 
                           IR_Dec_30_port, OPCODE(3) => IR_Dec_29_port, 
                           OPCODE(2) => IR_Dec_28_port, OPCODE(1) => 
                           IR_Dec_27_port, OPCODE(0) => IR_Dec_26_port, 
                           is_signed => signed_op, RS1(4) => RS1_4_port, RS1(3)
                           => RS1_3_port, RS1(2) => RS1_2_port, RS1(1) => 
                           RS1_1_port, RS1(0) => RS1_0_port, RS2(4) => 
                           RS2_4_port, RS2(3) => RS2_3_port, RS2(2) => 
                           RS2_2_port, RS2(1) => RS2_1_port, RS2(0) => 
                           RS2_0_port, RD(4) => RD_4_port, RD(3) => RD_3_port, 
                           RD(2) => RD_2_port, RD(1) => RD_1_port, RD(0) => 
                           RD_0_port, IMMEDIATE(31) => Imm_31_port, 
                           IMMEDIATE(30) => Imm_30_port, IMMEDIATE(29) => 
                           Imm_29_port, IMMEDIATE(28) => Imm_28_port, 
                           IMMEDIATE(27) => Imm_27_port, IMMEDIATE(26) => 
                           Imm_26_port, IMMEDIATE(25) => Imm_25_port, 
                           IMMEDIATE(24) => Imm_24_port, IMMEDIATE(23) => 
                           Imm_23_port, IMMEDIATE(22) => Imm_22_port, 
                           IMMEDIATE(21) => Imm_21_port, IMMEDIATE(20) => 
                           Imm_20_port, IMMEDIATE(19) => Imm_19_port, 
                           IMMEDIATE(18) => Imm_18_port, IMMEDIATE(17) => 
                           Imm_17_port, IMMEDIATE(16) => Imm_16_port, 
                           IMMEDIATE(15) => Imm_15_port, IMMEDIATE(14) => 
                           Imm_14_port, IMMEDIATE(13) => Imm_13_port, 
                           IMMEDIATE(12) => Imm_12_port, IMMEDIATE(11) => 
                           Imm_11_port, IMMEDIATE(10) => Imm_10_port, 
                           IMMEDIATE(9) => Imm_9_port, IMMEDIATE(8) => 
                           Imm_8_port, IMMEDIATE(7) => Imm_7_port, IMMEDIATE(6)
                           => Imm_6_port, IMMEDIATE(5) => Imm_5_port, 
                           IMMEDIATE(4) => Imm_4_port, IMMEDIATE(3) => 
                           Imm_3_port, IMMEDIATE(2) => Imm_2_port, IMMEDIATE(1)
                           => Imm_1_port, IMMEDIATE(0) => Imm_0_port);
   RF : windRF_M8_N8_F5_NBIT32 port map( CLK => CLK, RESET => n44, ENABLE => 
                           X_Logic1_port, CALL => trap_cs, RETRN => ret_cs, 
                           FILL => n_3077, SPILL => n_3078, BUSin(31) => 
                           X_Logic0_port, BUSin(30) => X_Logic0_port, BUSin(29)
                           => X_Logic0_port, BUSin(28) => X_Logic0_port, 
                           BUSin(27) => X_Logic0_port, BUSin(26) => 
                           X_Logic0_port, BUSin(25) => X_Logic0_port, BUSin(24)
                           => X_Logic0_port, BUSin(23) => X_Logic0_port, 
                           BUSin(22) => X_Logic0_port, BUSin(21) => 
                           X_Logic0_port, BUSin(20) => X_Logic0_port, BUSin(19)
                           => X_Logic0_port, BUSin(18) => X_Logic0_port, 
                           BUSin(17) => X_Logic0_port, BUSin(16) => 
                           X_Logic0_port, BUSin(15) => X_Logic0_port, BUSin(14)
                           => X_Logic0_port, BUSin(13) => X_Logic0_port, 
                           BUSin(12) => X_Logic0_port, BUSin(11) => 
                           X_Logic0_port, BUSin(10) => X_Logic0_port, BUSin(9) 
                           => X_Logic0_port, BUSin(8) => X_Logic0_port, 
                           BUSin(7) => X_Logic0_port, BUSin(6) => X_Logic0_port
                           , BUSin(5) => X_Logic0_port, BUSin(4) => 
                           X_Logic0_port, BUSin(3) => X_Logic0_port, BUSin(2) 
                           => X_Logic0_port, BUSin(1) => X_Logic0_port, 
                           BUSin(0) => X_Logic0_port, BUSout(31) => n_3079, 
                           BUSout(30) => n_3080, BUSout(29) => n_3081, 
                           BUSout(28) => n_3082, BUSout(27) => n_3083, 
                           BUSout(26) => n_3084, BUSout(25) => n_3085, 
                           BUSout(24) => n_3086, BUSout(23) => n_3087, 
                           BUSout(22) => n_3088, BUSout(21) => n_3089, 
                           BUSout(20) => n_3090, BUSout(19) => n_3091, 
                           BUSout(18) => n_3092, BUSout(17) => n_3093, 
                           BUSout(16) => n_3094, BUSout(15) => n_3095, 
                           BUSout(14) => n_3096, BUSout(13) => n_3097, 
                           BUSout(12) => n_3098, BUSout(11) => n_3099, 
                           BUSout(10) => n_3100, BUSout(9) => n_3101, BUSout(8)
                           => n_3102, BUSout(7) => n_3103, BUSout(6) => n_3104,
                           BUSout(5) => n_3105, BUSout(4) => n_3106, BUSout(3) 
                           => n_3107, BUSout(2) => n_3108, BUSout(1) => n_3109,
                           BUSout(0) => n_3110, RD1 => RF1, RD2 => RF2, WR => 
                           WF1, ADD_WR(4) => RD_wb_4_port, ADD_WR(3) => 
                           RD_wb_3_port, ADD_WR(2) => RD_wb_2_port, ADD_WR(1) 
                           => RD_wb_1_port, ADD_WR(0) => RD_wb_0_port, 
                           ADD_RD1(4) => RS1_4_port, ADD_RD1(3) => RS1_3_port, 
                           ADD_RD1(2) => RS1_2_port, ADD_RD1(1) => RS1_1_port, 
                           ADD_RD1(0) => RS1_0_port, ADD_RD2(4) => RS2_4_port, 
                           ADD_RD2(3) => RS2_3_port, ADD_RD2(2) => RS2_2_port, 
                           ADD_RD2(1) => RS2_1_port, ADD_RD2(0) => RS2_0_port, 
                           DATAIN(31) => OUT_wb_31_port, DATAIN(30) => 
                           OUT_wb_30_port, DATAIN(29) => OUT_wb_29_port, 
                           DATAIN(28) => OUT_wb_28_port, DATAIN(27) => 
                           OUT_wb_27_port, DATAIN(26) => OUT_wb_26_port, 
                           DATAIN(25) => OUT_wb_25_port, DATAIN(24) => 
                           OUT_wb_24_port, DATAIN(23) => OUT_wb_23_port, 
                           DATAIN(22) => OUT_wb_22_port, DATAIN(21) => 
                           OUT_wb_21_port, DATAIN(20) => OUT_wb_20_port, 
                           DATAIN(19) => OUT_wb_19_port, DATAIN(18) => 
                           OUT_wb_18_port, DATAIN(17) => OUT_wb_17_port, 
                           DATAIN(16) => OUT_wb_16_port, DATAIN(15) => 
                           OUT_wb_15_port, DATAIN(14) => OUT_wb_14_port, 
                           DATAIN(13) => OUT_wb_13_port, DATAIN(12) => 
                           OUT_wb_12_port, DATAIN(11) => OUT_wb_11_port, 
                           DATAIN(10) => OUT_wb_10_port, DATAIN(9) => 
                           OUT_wb_9_port, DATAIN(8) => OUT_wb_8_port, DATAIN(7)
                           => OUT_wb_7_port, DATAIN(6) => OUT_wb_6_port, 
                           DATAIN(5) => OUT_wb_5_port, DATAIN(4) => 
                           OUT_wb_4_port, DATAIN(3) => OUT_wb_3_port, DATAIN(2)
                           => OUT_wb_2_port, DATAIN(1) => OUT_wb_1_port, 
                           DATAIN(0) => OUT_wb_0_port, OUT1(31) => regA_31_port
                           , OUT1(30) => regA_30_port, OUT1(29) => regA_29_port
                           , OUT1(28) => regA_28_port, OUT1(27) => regA_27_port
                           , OUT1(26) => regA_26_port, OUT1(25) => regA_25_port
                           , OUT1(24) => regA_24_port, OUT1(23) => regA_23_port
                           , OUT1(22) => regA_22_port, OUT1(21) => regA_21_port
                           , OUT1(20) => regA_20_port, OUT1(19) => regA_19_port
                           , OUT1(18) => regA_18_port, OUT1(17) => regA_17_port
                           , OUT1(16) => regA_16_port, OUT1(15) => regA_15_port
                           , OUT1(14) => regA_14_port, OUT1(13) => regA_13_port
                           , OUT1(12) => regA_12_port, OUT1(11) => regA_11_port
                           , OUT1(10) => regA_10_port, OUT1(9) => regA_9_port, 
                           OUT1(8) => regA_8_port, OUT1(7) => regA_7_port, 
                           OUT1(6) => regA_6_port, OUT1(5) => regA_5_port, 
                           OUT1(4) => regA_4_port, OUT1(3) => regA_3_port, 
                           OUT1(2) => regA_2_port, OUT1(1) => regA_1_port, 
                           OUT1(0) => regA_0_port, OUT2(31) => regB_31_port, 
                           OUT2(30) => regB_30_port, OUT2(29) => regB_29_port, 
                           OUT2(28) => regB_28_port, OUT2(27) => regB_27_port, 
                           OUT2(26) => regB_26_port, OUT2(25) => regB_25_port, 
                           OUT2(24) => regB_24_port, OUT2(23) => regB_23_port, 
                           OUT2(22) => regB_22_port, OUT2(21) => regB_21_port, 
                           OUT2(20) => regB_20_port, OUT2(19) => regB_19_port, 
                           OUT2(18) => regB_18_port, OUT2(17) => regB_17_port, 
                           OUT2(16) => regB_16_port, OUT2(15) => regB_15_port, 
                           OUT2(14) => regB_14_port, OUT2(13) => regB_13_port, 
                           OUT2(12) => regB_12_port, OUT2(11) => regB_11_port, 
                           OUT2(10) => regB_10_port, OUT2(9) => regB_9_port, 
                           OUT2(8) => regB_8_port, OUT2(7) => regB_7_port, 
                           OUT2(6) => regB_6_port, OUT2(5) => regB_5_port, 
                           OUT2(4) => regB_4_port, OUT2(3) => regB_3_port, 
                           OUT2(2) => regB_2_port, OUT2(1) => regB_1_port, 
                           OUT2(0) => regB_0_port, wr_signal => wr_signal_wb);
   pipeline_sign2 : FF_0 port map( CLK => CLK, RESET => n45, EN => 
                           X_Logic1_port, D => signed_op, Q => signed_op_ex);
   pipeline_newpc2 : regFFD_NBIT32_11 port map( CK => CLK, RESET => n45, ENABLE
                           => X_Logic1_port, D(31) => NPC_Dec_31_port, D(30) =>
                           NPC_Dec_30_port, D(29) => NPC_Dec_29_port, D(28) => 
                           NPC_Dec_28_port, D(27) => NPC_Dec_27_port, D(26) => 
                           NPC_Dec_26_port, D(25) => NPC_Dec_25_port, D(24) => 
                           NPC_Dec_24_port, D(23) => NPC_Dec_23_port, D(22) => 
                           NPC_Dec_22_port, D(21) => NPC_Dec_21_port, D(20) => 
                           NPC_Dec_20_port, D(19) => NPC_Dec_19_port, D(18) => 
                           NPC_Dec_18_port, D(17) => NPC_Dec_17_port, D(16) => 
                           NPC_Dec_16_port, D(15) => NPC_Dec_15_port, D(14) => 
                           NPC_Dec_14_port, D(13) => NPC_Dec_13_port, D(12) => 
                           NPC_Dec_12_port, D(11) => NPC_Dec_11_port, D(10) => 
                           NPC_Dec_10_port, D(9) => NPC_Dec_9_port, D(8) => 
                           NPC_Dec_8_port, D(7) => NPC_Dec_7_port, D(6) => 
                           NPC_Dec_6_port, D(5) => NPC_Dec_5_port, D(4) => 
                           NPC_Dec_4_port, D(3) => NPC_Dec_3_port, D(2) => 
                           NPC_Dec_2_port, D(1) => NPC_Dec_1_port, D(0) => 
                           NPC_Dec_0_port, Q(31) => NPC_ex_31_port, Q(30) => 
                           NPC_ex_30_port, Q(29) => NPC_ex_29_port, Q(28) => 
                           NPC_ex_28_port, Q(27) => NPC_ex_27_port, Q(26) => 
                           NPC_ex_26_port, Q(25) => NPC_ex_25_port, Q(24) => 
                           NPC_ex_24_port, Q(23) => NPC_ex_23_port, Q(22) => 
                           NPC_ex_22_port, Q(21) => NPC_ex_21_port, Q(20) => 
                           NPC_ex_20_port, Q(19) => NPC_ex_19_port, Q(18) => 
                           NPC_ex_18_port, Q(17) => NPC_ex_17_port, Q(16) => 
                           NPC_ex_16_port, Q(15) => NPC_ex_15_port, Q(14) => 
                           NPC_ex_14_port, Q(13) => NPC_ex_13_port, Q(12) => 
                           NPC_ex_12_port, Q(11) => NPC_ex_11_port, Q(10) => 
                           NPC_ex_10_port, Q(9) => NPC_ex_9_port, Q(8) => 
                           NPC_ex_8_port, Q(7) => NPC_ex_7_port, Q(6) => 
                           NPC_ex_6_port, Q(5) => NPC_ex_5_port, Q(4) => 
                           NPC_ex_4_port, Q(3) => NPC_ex_3_port, Q(2) => 
                           NPC_ex_2_port, Q(1) => NPC_ex_1_port, Q(0) => 
                           NPC_ex_0_port);
   pipeline_A2 : regFFD_NBIT32_10 port map( CK => CLK, RESET => n44, ENABLE => 
                           RF1, D(31) => regA_31_port, D(30) => regA_30_port, 
                           D(29) => regA_29_port, D(28) => regA_28_port, D(27) 
                           => regA_27_port, D(26) => regA_26_port, D(25) => 
                           regA_25_port, D(24) => regA_24_port, D(23) => 
                           regA_23_port, D(22) => regA_22_port, D(21) => 
                           regA_21_port, D(20) => regA_20_port, D(19) => 
                           regA_19_port, D(18) => regA_18_port, D(17) => 
                           regA_17_port, D(16) => regA_16_port, D(15) => 
                           regA_15_port, D(14) => regA_14_port, D(13) => 
                           regA_13_port, D(12) => regA_12_port, D(11) => 
                           regA_11_port, D(10) => regA_10_port, D(9) => 
                           regA_9_port, D(8) => regA_8_port, D(7) => 
                           regA_7_port, D(6) => regA_6_port, D(5) => 
                           regA_5_port, D(4) => regA_4_port, D(3) => 
                           regA_3_port, D(2) => regA_2_port, D(1) => 
                           regA_1_port, D(0) => regA_0_port, Q(31) => 
                           regA_ex_31_port, Q(30) => regA_ex_30_port, Q(29) => 
                           regA_ex_29_port, Q(28) => regA_ex_28_port, Q(27) => 
                           regA_ex_27_port, Q(26) => regA_ex_26_port, Q(25) => 
                           regA_ex_25_port, Q(24) => regA_ex_24_port, Q(23) => 
                           regA_ex_23_port, Q(22) => regA_ex_22_port, Q(21) => 
                           regA_ex_21_port, Q(20) => regA_ex_20_port, Q(19) => 
                           regA_ex_19_port, Q(18) => regA_ex_18_port, Q(17) => 
                           regA_ex_17_port, Q(16) => regA_ex_16_port, Q(15) => 
                           regA_ex_15_port, Q(14) => regA_ex_14_port, Q(13) => 
                           regA_ex_13_port, Q(12) => regA_ex_12_port, Q(11) => 
                           regA_ex_11_port, Q(10) => regA_ex_10_port, Q(9) => 
                           regA_ex_9_port, Q(8) => regA_ex_8_port, Q(7) => 
                           regA_ex_7_port, Q(6) => regA_ex_6_port, Q(5) => 
                           regA_ex_5_port, Q(4) => regA_ex_4_port, Q(3) => 
                           regA_ex_3_port, Q(2) => regA_ex_2_port, Q(1) => 
                           regA_ex_1_port, Q(0) => regA_ex_0_port);
   pipeline_B2 : regFFD_NBIT32_9 port map( CK => CLK, RESET => n44, ENABLE => 
                           RF2, D(31) => regB_31_port, D(30) => regB_30_port, 
                           D(29) => regB_29_port, D(28) => regB_28_port, D(27) 
                           => regB_27_port, D(26) => regB_26_port, D(25) => 
                           regB_25_port, D(24) => regB_24_port, D(23) => 
                           regB_23_port, D(22) => regB_22_port, D(21) => 
                           regB_21_port, D(20) => regB_20_port, D(19) => 
                           regB_19_port, D(18) => regB_18_port, D(17) => 
                           regB_17_port, D(16) => regB_16_port, D(15) => 
                           regB_15_port, D(14) => regB_14_port, D(13) => 
                           regB_13_port, D(12) => regB_12_port, D(11) => 
                           regB_11_port, D(10) => regB_10_port, D(9) => 
                           regB_9_port, D(8) => regB_8_port, D(7) => 
                           regB_7_port, D(6) => regB_6_port, D(5) => 
                           regB_5_port, D(4) => regB_4_port, D(3) => 
                           regB_3_port, D(2) => regB_2_port, D(1) => 
                           regB_1_port, D(0) => regB_0_port, Q(31) => 
                           regB_ex_31_port, Q(30) => regB_ex_30_port, Q(29) => 
                           regB_ex_29_port, Q(28) => regB_ex_28_port, Q(27) => 
                           regB_ex_27_port, Q(26) => regB_ex_26_port, Q(25) => 
                           regB_ex_25_port, Q(24) => regB_ex_24_port, Q(23) => 
                           regB_ex_23_port, Q(22) => regB_ex_22_port, Q(21) => 
                           regB_ex_21_port, Q(20) => regB_ex_20_port, Q(19) => 
                           regB_ex_19_port, Q(18) => regB_ex_18_port, Q(17) => 
                           regB_ex_17_port, Q(16) => regB_ex_16_port, Q(15) => 
                           regB_ex_15_port, Q(14) => regB_ex_14_port, Q(13) => 
                           regB_ex_13_port, Q(12) => regB_ex_12_port, Q(11) => 
                           regB_ex_11_port, Q(10) => regB_ex_10_port, Q(9) => 
                           regB_ex_9_port, Q(8) => regB_ex_8_port, Q(7) => 
                           regB_ex_7_port, Q(6) => regB_ex_6_port, Q(5) => 
                           regB_ex_5_port, Q(4) => regB_ex_4_port, Q(3) => 
                           regB_ex_3_port, Q(2) => regB_ex_2_port, Q(1) => 
                           regB_ex_1_port, Q(0) => regB_ex_0_port);
   pipeline_IMM2 : regFFD_NBIT32_8 port map( CK => CLK, RESET => n44, ENABLE =>
                           regImm_LATCH_EN, D(31) => Imm_31_port, D(30) => 
                           Imm_30_port, D(29) => Imm_29_port, D(28) => 
                           Imm_28_port, D(27) => Imm_27_port, D(26) => 
                           Imm_26_port, D(25) => Imm_25_port, D(24) => 
                           Imm_24_port, D(23) => Imm_23_port, D(22) => 
                           Imm_22_port, D(21) => Imm_21_port, D(20) => 
                           Imm_20_port, D(19) => Imm_19_port, D(18) => 
                           Imm_18_port, D(17) => Imm_17_port, D(16) => 
                           Imm_16_port, D(15) => Imm_15_port, D(14) => 
                           Imm_14_port, D(13) => Imm_13_port, D(12) => 
                           Imm_12_port, D(11) => Imm_11_port, D(10) => 
                           Imm_10_port, D(9) => Imm_9_port, D(8) => Imm_8_port,
                           D(7) => Imm_7_port, D(6) => Imm_6_port, D(5) => 
                           Imm_5_port, D(4) => Imm_4_port, D(3) => Imm_3_port, 
                           D(2) => Imm_2_port, D(1) => Imm_1_port, D(0) => 
                           Imm_0_port, Q(31) => Imm_ex_31_port, Q(30) => 
                           Imm_ex_30_port, Q(29) => Imm_ex_29_port, Q(28) => 
                           Imm_ex_28_port, Q(27) => Imm_ex_27_port, Q(26) => 
                           Imm_ex_26_port, Q(25) => Imm_ex_25_port, Q(24) => 
                           Imm_ex_24_port, Q(23) => Imm_ex_23_port, Q(22) => 
                           Imm_ex_22_port, Q(21) => Imm_ex_21_port, Q(20) => 
                           Imm_ex_20_port, Q(19) => Imm_ex_19_port, Q(18) => 
                           Imm_ex_18_port, Q(17) => Imm_ex_17_port, Q(16) => 
                           Imm_ex_16_port, Q(15) => Imm_ex_15_port, Q(14) => 
                           Imm_ex_14_port, Q(13) => Imm_ex_13_port, Q(12) => 
                           Imm_ex_12_port, Q(11) => Imm_ex_11_port, Q(10) => 
                           Imm_ex_10_port, Q(9) => Imm_ex_9_port, Q(8) => 
                           Imm_ex_8_port, Q(7) => Imm_ex_7_port, Q(6) => 
                           Imm_ex_6_port, Q(5) => Imm_ex_5_port, Q(4) => 
                           Imm_ex_4_port, Q(3) => Imm_ex_3_port, Q(2) => 
                           Imm_ex_2_port, Q(1) => Imm_ex_1_port, Q(0) => 
                           Imm_ex_0_port);
   pipeline_RD2 : regFFD_NBIT5_0 port map( CK => CLK, RESET => n44, ENABLE => 
                           X_Logic1_port, D(4) => RD_4_port, D(3) => RD_3_port,
                           D(2) => RD_2_port, D(1) => RD_1_port, D(0) => 
                           RD_0_port, Q(4) => RD_ex_4_port, Q(3) => 
                           RD_ex_3_port, Q(2) => RD_ex_2_port, Q(1) => 
                           RD_ex_1_port, Q(0) => RD_ex_0_port);
   pipeline_wr_signal : FF_7 port map( CLK => CLK, RESET => n45, EN => 
                           X_Logic1_port, D => n34, Q => wr_signal_exe);
   pipeline_IR2 : regFFD_NBIT6_0 port map( CK => CLK, RESET => n44, ENABLE => 
                           X_Logic1_port, D(5) => n36, D(4) => IR_Dec_30_port, 
                           D(3) => n35, D(2) => IR_Dec_28_port, D(1) => 
                           IR_Dec_27_port, D(0) => IR_Dec_26_port, Q(5) => 
                           IR_26_ex_5_port, Q(4) => IR_26_ex_4_port, Q(3) => 
                           IR_26_ex_3_port, Q(2) => IR_26_ex_2_port, Q(1) => 
                           IR_26_ex_1_port, Q(0) => IR_26_ex_0_port);
   pipeline_LHI2 : regFFD_NBIT32_7 port map( CK => CLK, RESET => n45, ENABLE =>
                           X_Logic1_port, D(31) => Imm_15_port, D(30) => 
                           Imm_14_port, D(29) => Imm_13_port, D(28) => 
                           Imm_12_port, D(27) => Imm_11_port, D(26) => 
                           Imm_10_port, D(25) => Imm_9_port, D(24) => 
                           Imm_8_port, D(23) => Imm_7_port, D(22) => Imm_6_port
                           , D(21) => Imm_5_port, D(20) => Imm_4_port, D(19) =>
                           Imm_3_port, D(18) => Imm_2_port, D(17) => Imm_1_port
                           , D(16) => Imm_0_port, D(15) => X_Logic0_port, D(14)
                           => X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, Q(31) => LHI_ex1_31_port, Q(30) => 
                           LHI_ex1_30_port, Q(29) => LHI_ex1_29_port, Q(28) => 
                           LHI_ex1_28_port, Q(27) => LHI_ex1_27_port, Q(26) => 
                           LHI_ex1_26_port, Q(25) => LHI_ex1_25_port, Q(24) => 
                           LHI_ex1_24_port, Q(23) => LHI_ex1_23_port, Q(22) => 
                           LHI_ex1_22_port, Q(21) => LHI_ex1_21_port, Q(20) => 
                           LHI_ex1_20_port, Q(19) => LHI_ex1_19_port, Q(18) => 
                           LHI_ex1_18_port, Q(17) => LHI_ex1_17_port, Q(16) => 
                           LHI_ex1_16_port, Q(15) => LHI_ex1_15_port, Q(14) => 
                           LHI_ex1_14_port, Q(13) => LHI_ex1_13_port, Q(12) => 
                           LHI_ex1_12_port, Q(11) => LHI_ex1_11_port, Q(10) => 
                           LHI_ex1_10_port, Q(9) => LHI_ex1_9_port, Q(8) => 
                           LHI_ex1_8_port, Q(7) => LHI_ex1_7_port, Q(6) => 
                           LHI_ex1_6_port, Q(5) => LHI_ex1_5_port, Q(4) => 
                           LHI_ex1_4_port, Q(3) => LHI_ex1_3_port, Q(2) => 
                           LHI_ex1_2_port, Q(1) => LHI_ex1_1_port, Q(0) => 
                           LHI_ex1_0_port);
   pipeline_LHI3 : regFFD_NBIT32_6 port map( CK => CLK, RESET => n45, ENABLE =>
                           X_Logic1_port, D(31) => LHI_ex1_31_port, D(30) => 
                           LHI_ex1_30_port, D(29) => LHI_ex1_29_port, D(28) => 
                           LHI_ex1_28_port, D(27) => LHI_ex1_27_port, D(26) => 
                           LHI_ex1_26_port, D(25) => LHI_ex1_25_port, D(24) => 
                           LHI_ex1_24_port, D(23) => LHI_ex1_23_port, D(22) => 
                           LHI_ex1_22_port, D(21) => LHI_ex1_21_port, D(20) => 
                           LHI_ex1_20_port, D(19) => LHI_ex1_19_port, D(18) => 
                           LHI_ex1_18_port, D(17) => LHI_ex1_17_port, D(16) => 
                           LHI_ex1_16_port, D(15) => LHI_ex1_15_port, D(14) => 
                           LHI_ex1_14_port, D(13) => LHI_ex1_13_port, D(12) => 
                           LHI_ex1_12_port, D(11) => LHI_ex1_11_port, D(10) => 
                           LHI_ex1_10_port, D(9) => LHI_ex1_9_port, D(8) => 
                           LHI_ex1_8_port, D(7) => LHI_ex1_7_port, D(6) => 
                           LHI_ex1_6_port, D(5) => LHI_ex1_5_port, D(4) => 
                           LHI_ex1_4_port, D(3) => LHI_ex1_3_port, D(2) => 
                           LHI_ex1_2_port, D(1) => LHI_ex1_1_port, D(0) => 
                           LHI_ex1_0_port, Q(31) => LHI_ex_31_port, Q(30) => 
                           LHI_ex_30_port, Q(29) => LHI_ex_29_port, Q(28) => 
                           LHI_ex_28_port, Q(27) => LHI_ex_27_port, Q(26) => 
                           LHI_ex_26_port, Q(25) => LHI_ex_25_port, Q(24) => 
                           LHI_ex_24_port, Q(23) => LHI_ex_23_port, Q(22) => 
                           LHI_ex_22_port, Q(21) => LHI_ex_21_port, Q(20) => 
                           LHI_ex_20_port, Q(19) => LHI_ex_19_port, Q(18) => 
                           LHI_ex_18_port, Q(17) => LHI_ex_17_port, Q(16) => 
                           LHI_ex_16_port, Q(15) => LHI_ex_15_port, Q(14) => 
                           LHI_ex_14_port, Q(13) => LHI_ex_13_port, Q(12) => 
                           LHI_ex_12_port, Q(11) => LHI_ex_11_port, Q(10) => 
                           LHI_ex_10_port, Q(9) => LHI_ex_9_port, Q(8) => 
                           LHI_ex_8_port, Q(7) => LHI_ex_7_port, Q(6) => 
                           LHI_ex_6_port, Q(5) => LHI_ex_5_port, Q(4) => 
                           LHI_ex_4_port, Q(3) => LHI_ex_3_port, Q(2) => 
                           LHI_ex_2_port, Q(1) => LHI_ex_1_port, Q(0) => 
                           LHI_ex_0_port);
   MUX_ALU_A : MUX21_GENERIC_NBIT32_6 port map( A(31) => NPC_ex_31_port, A(30) 
                           => NPC_ex_30_port, A(29) => NPC_ex_29_port, A(28) =>
                           NPC_ex_28_port, A(27) => NPC_ex_27_port, A(26) => 
                           NPC_ex_26_port, A(25) => NPC_ex_25_port, A(24) => 
                           NPC_ex_24_port, A(23) => NPC_ex_23_port, A(22) => 
                           NPC_ex_22_port, A(21) => NPC_ex_21_port, A(20) => 
                           NPC_ex_20_port, A(19) => NPC_ex_19_port, A(18) => 
                           NPC_ex_18_port, A(17) => NPC_ex_17_port, A(16) => 
                           NPC_ex_16_port, A(15) => NPC_ex_15_port, A(14) => 
                           NPC_ex_14_port, A(13) => NPC_ex_13_port, A(12) => 
                           NPC_ex_12_port, A(11) => NPC_ex_11_port, A(10) => 
                           NPC_ex_10_port, A(9) => NPC_ex_9_port, A(8) => 
                           NPC_ex_8_port, A(7) => NPC_ex_7_port, A(6) => 
                           NPC_ex_6_port, A(5) => NPC_ex_5_port, A(4) => 
                           NPC_ex_4_port, A(3) => NPC_ex_3_port, A(2) => 
                           NPC_ex_2_port, A(1) => NPC_ex_1_port, A(0) => 
                           NPC_ex_0_port, B(31) => regA_ex_31_port, B(30) => 
                           regA_ex_30_port, B(29) => regA_ex_29_port, B(28) => 
                           regA_ex_28_port, B(27) => regA_ex_27_port, B(26) => 
                           regA_ex_26_port, B(25) => regA_ex_25_port, B(24) => 
                           regA_ex_24_port, B(23) => regA_ex_23_port, B(22) => 
                           regA_ex_22_port, B(21) => regA_ex_21_port, B(20) => 
                           regA_ex_20_port, B(19) => regA_ex_19_port, B(18) => 
                           regA_ex_18_port, B(17) => regA_ex_17_port, B(16) => 
                           regA_ex_16_port, B(15) => regA_ex_15_port, B(14) => 
                           regA_ex_14_port, B(13) => regA_ex_13_port, B(12) => 
                           regA_ex_12_port, B(11) => regA_ex_11_port, B(10) => 
                           regA_ex_10_port, B(9) => regA_ex_9_port, B(8) => 
                           regA_ex_8_port, B(7) => regA_ex_7_port, B(6) => 
                           regA_ex_6_port, B(5) => regA_ex_5_port, B(4) => 
                           regA_ex_4_port, B(3) => regA_ex_3_port, B(2) => 
                           regA_ex_2_port, B(1) => regA_ex_1_port, B(0) => 
                           regA_ex_0_port, SEL => S1, Y(31) => 
                           input1_ALU_31_port, Y(30) => input1_ALU_30_port, 
                           Y(29) => input1_ALU_29_port, Y(28) => 
                           input1_ALU_28_port, Y(27) => input1_ALU_27_port, 
                           Y(26) => input1_ALU_26_port, Y(25) => 
                           input1_ALU_25_port, Y(24) => input1_ALU_24_port, 
                           Y(23) => input1_ALU_23_port, Y(22) => 
                           input1_ALU_22_port, Y(21) => input1_ALU_21_port, 
                           Y(20) => input1_ALU_20_port, Y(19) => 
                           input1_ALU_19_port, Y(18) => input1_ALU_18_port, 
                           Y(17) => input1_ALU_17_port, Y(16) => 
                           input1_ALU_16_port, Y(15) => input1_ALU_15_port, 
                           Y(14) => input1_ALU_14_port, Y(13) => 
                           input1_ALU_13_port, Y(12) => input1_ALU_12_port, 
                           Y(11) => input1_ALU_11_port, Y(10) => 
                           input1_ALU_10_port, Y(9) => input1_ALU_9_port, Y(8) 
                           => input1_ALU_8_port, Y(7) => input1_ALU_7_port, 
                           Y(6) => input1_ALU_6_port, Y(5) => input1_ALU_5_port
                           , Y(4) => input1_ALU_4_port, Y(3) => 
                           input1_ALU_3_port, Y(2) => input1_ALU_2_port, Y(1) 
                           => input1_ALU_1_port, Y(0) => input1_ALU_0_port);
   MUX_ALU_B : MUX21_GENERIC_NBIT32_5 port map( A(31) => Imm_ex_31_port, A(30) 
                           => Imm_ex_30_port, A(29) => Imm_ex_29_port, A(28) =>
                           Imm_ex_28_port, A(27) => Imm_ex_27_port, A(26) => 
                           Imm_ex_26_port, A(25) => Imm_ex_25_port, A(24) => 
                           Imm_ex_24_port, A(23) => Imm_ex_23_port, A(22) => 
                           Imm_ex_22_port, A(21) => Imm_ex_21_port, A(20) => 
                           Imm_ex_20_port, A(19) => Imm_ex_19_port, A(18) => 
                           Imm_ex_18_port, A(17) => Imm_ex_17_port, A(16) => 
                           Imm_ex_16_port, A(15) => Imm_ex_15_port, A(14) => 
                           Imm_ex_14_port, A(13) => Imm_ex_13_port, A(12) => 
                           Imm_ex_12_port, A(11) => Imm_ex_11_port, A(10) => 
                           Imm_ex_10_port, A(9) => Imm_ex_9_port, A(8) => 
                           Imm_ex_8_port, A(7) => Imm_ex_7_port, A(6) => 
                           Imm_ex_6_port, A(5) => Imm_ex_5_port, A(4) => 
                           Imm_ex_4_port, A(3) => Imm_ex_3_port, A(2) => 
                           Imm_ex_2_port, A(1) => Imm_ex_1_port, A(0) => 
                           Imm_ex_0_port, B(31) => regB_ex_31_port, B(30) => 
                           regB_ex_30_port, B(29) => regB_ex_29_port, B(28) => 
                           regB_ex_28_port, B(27) => regB_ex_27_port, B(26) => 
                           regB_ex_26_port, B(25) => regB_ex_25_port, B(24) => 
                           regB_ex_24_port, B(23) => regB_ex_23_port, B(22) => 
                           regB_ex_22_port, B(21) => regB_ex_21_port, B(20) => 
                           regB_ex_20_port, B(19) => regB_ex_19_port, B(18) => 
                           regB_ex_18_port, B(17) => regB_ex_17_port, B(16) => 
                           regB_ex_16_port, B(15) => regB_ex_15_port, B(14) => 
                           regB_ex_14_port, B(13) => regB_ex_13_port, B(12) => 
                           regB_ex_12_port, B(11) => regB_ex_11_port, B(10) => 
                           regB_ex_10_port, B(9) => regB_ex_9_port, B(8) => 
                           regB_ex_8_port, B(7) => regB_ex_7_port, B(6) => 
                           regB_ex_6_port, B(5) => regB_ex_5_port, B(4) => 
                           regB_ex_4_port, B(3) => regB_ex_3_port, B(2) => 
                           regB_ex_2_port, B(1) => regB_ex_1_port, B(0) => 
                           regB_ex_0_port, SEL => S2, Y(31) => 
                           input2_ALU_31_port, Y(30) => input2_ALU_30_port, 
                           Y(29) => input2_ALU_29_port, Y(28) => 
                           input2_ALU_28_port, Y(27) => input2_ALU_27_port, 
                           Y(26) => input2_ALU_26_port, Y(25) => 
                           input2_ALU_25_port, Y(24) => input2_ALU_24_port, 
                           Y(23) => input2_ALU_23_port, Y(22) => 
                           input2_ALU_22_port, Y(21) => input2_ALU_21_port, 
                           Y(20) => input2_ALU_20_port, Y(19) => 
                           input2_ALU_19_port, Y(18) => input2_ALU_18_port, 
                           Y(17) => input2_ALU_17_port, Y(16) => 
                           input2_ALU_16_port, Y(15) => input2_ALU_15_port, 
                           Y(14) => input2_ALU_14_port, Y(13) => 
                           input2_ALU_13_port, Y(12) => input2_ALU_12_port, 
                           Y(11) => input2_ALU_11_port, Y(10) => 
                           input2_ALU_10_port, Y(9) => input2_ALU_9_port, Y(8) 
                           => input2_ALU_8_port, Y(7) => input2_ALU_7_port, 
                           Y(6) => input2_ALU_6_port, Y(5) => input2_ALU_5_port
                           , Y(4) => input2_ALU_4_port, Y(3) => 
                           input2_ALU_3_port, Y(2) => input2_ALU_2_port, Y(1) 
                           => input2_ALU_1_port, Y(0) => input2_ALU_0_port);
   ALU_OP : ALU_N32 port map( CLK => CLK, FUNC(0) => instruction_alu(0), 
                           FUNC(1) => instruction_alu(1), FUNC(2) => 
                           instruction_alu(2), FUNC(3) => instruction_alu(3), 
                           FUNC(4) => instruction_alu(4), FUNC(5) => 
                           instruction_alu(5), DATA1(31) => input1_ALU_31_port,
                           DATA1(30) => input1_ALU_30_port, DATA1(29) => 
                           input1_ALU_29_port, DATA1(28) => input1_ALU_28_port,
                           DATA1(27) => input1_ALU_27_port, DATA1(26) => 
                           input1_ALU_26_port, DATA1(25) => input1_ALU_25_port,
                           DATA1(24) => input1_ALU_24_port, DATA1(23) => 
                           input1_ALU_23_port, DATA1(22) => input1_ALU_22_port,
                           DATA1(21) => input1_ALU_21_port, DATA1(20) => 
                           input1_ALU_20_port, DATA1(19) => input1_ALU_19_port,
                           DATA1(18) => input1_ALU_18_port, DATA1(17) => 
                           input1_ALU_17_port, DATA1(16) => input1_ALU_16_port,
                           DATA1(15) => input1_ALU_15_port, DATA1(14) => 
                           input1_ALU_14_port, DATA1(13) => input1_ALU_13_port,
                           DATA1(12) => input1_ALU_12_port, DATA1(11) => 
                           input1_ALU_11_port, DATA1(10) => input1_ALU_10_port,
                           DATA1(9) => input1_ALU_9_port, DATA1(8) => 
                           input1_ALU_8_port, DATA1(7) => input1_ALU_7_port, 
                           DATA1(6) => input1_ALU_6_port, DATA1(5) => 
                           input1_ALU_5_port, DATA1(4) => input1_ALU_4_port, 
                           DATA1(3) => input1_ALU_3_port, DATA1(2) => 
                           input1_ALU_2_port, DATA1(1) => input1_ALU_1_port, 
                           DATA1(0) => input1_ALU_0_port, DATA2(31) => 
                           input2_ALU_31_port, DATA2(30) => input2_ALU_30_port,
                           DATA2(29) => input2_ALU_29_port, DATA2(28) => 
                           input2_ALU_28_port, DATA2(27) => input2_ALU_27_port,
                           DATA2(26) => input2_ALU_26_port, DATA2(25) => 
                           input2_ALU_25_port, DATA2(24) => input2_ALU_24_port,
                           DATA2(23) => input2_ALU_23_port, DATA2(22) => 
                           input2_ALU_22_port, DATA2(21) => input2_ALU_21_port,
                           DATA2(20) => input2_ALU_20_port, DATA2(19) => 
                           input2_ALU_19_port, DATA2(18) => input2_ALU_18_port,
                           DATA2(17) => input2_ALU_17_port, DATA2(16) => 
                           input2_ALU_16_port, DATA2(15) => input2_ALU_15_port,
                           DATA2(14) => input2_ALU_14_port, DATA2(13) => 
                           input2_ALU_13_port, DATA2(12) => input2_ALU_12_port,
                           DATA2(11) => input2_ALU_11_port, DATA2(10) => 
                           input2_ALU_10_port, DATA2(9) => input2_ALU_9_port, 
                           DATA2(8) => input2_ALU_8_port, DATA2(7) => 
                           input2_ALU_7_port, DATA2(6) => input2_ALU_6_port, 
                           DATA2(5) => input2_ALU_5_port, DATA2(4) => 
                           input2_ALU_4_port, DATA2(3) => input2_ALU_3_port, 
                           DATA2(2) => input2_ALU_2_port, DATA2(1) => 
                           input2_ALU_1_port, DATA2(0) => input2_ALU_0_port, 
                           OUT_ALU(31) => ALU_out_31_port, OUT_ALU(30) => 
                           ALU_out_30_port, OUT_ALU(29) => ALU_out_29_port, 
                           OUT_ALU(28) => ALU_out_28_port, OUT_ALU(27) => 
                           ALU_out_27_port, OUT_ALU(26) => ALU_out_26_port, 
                           OUT_ALU(25) => ALU_out_25_port, OUT_ALU(24) => 
                           ALU_out_24_port, OUT_ALU(23) => ALU_out_23_port, 
                           OUT_ALU(22) => ALU_out_22_port, OUT_ALU(21) => 
                           ALU_out_21_port, OUT_ALU(20) => ALU_out_20_port, 
                           OUT_ALU(19) => ALU_out_19_port, OUT_ALU(18) => 
                           ALU_out_18_port, OUT_ALU(17) => ALU_out_17_port, 
                           OUT_ALU(16) => ALU_out_16_port, OUT_ALU(15) => 
                           ALU_out_15_port, OUT_ALU(14) => ALU_out_14_port, 
                           OUT_ALU(13) => ALU_out_13_port, OUT_ALU(12) => 
                           ALU_out_12_port, OUT_ALU(11) => ALU_out_11_port, 
                           OUT_ALU(10) => ALU_out_10_port, OUT_ALU(9) => 
                           ALU_out_9_port, OUT_ALU(8) => ALU_out_8_port, 
                           OUT_ALU(7) => ALU_out_7_port, OUT_ALU(6) => 
                           ALU_out_6_port, OUT_ALU(5) => ALU_out_5_port, 
                           OUT_ALU(4) => ALU_out_4_port, OUT_ALU(3) => 
                           ALU_out_3_port, OUT_ALU(2) => ALU_out_2_port, 
                           OUT_ALU(1) => ALU_out_1_port, OUT_ALU(0) => 
                           ALU_out_0_port);
   ZERO_OP : zero_eval_NBIT32 port map( input(31) => regA_ex_31_port, input(30)
                           => regA_ex_30_port, input(29) => regA_ex_29_port, 
                           input(28) => regA_ex_28_port, input(27) => 
                           regA_ex_27_port, input(26) => regA_ex_26_port, 
                           input(25) => regA_ex_25_port, input(24) => 
                           regA_ex_24_port, input(23) => regA_ex_23_port, 
                           input(22) => regA_ex_22_port, input(21) => 
                           regA_ex_21_port, input(20) => regA_ex_20_port, 
                           input(19) => regA_ex_19_port, input(18) => 
                           regA_ex_18_port, input(17) => regA_ex_17_port, 
                           input(16) => regA_ex_16_port, input(15) => 
                           regA_ex_15_port, input(14) => regA_ex_14_port, 
                           input(13) => regA_ex_13_port, input(12) => 
                           regA_ex_12_port, input(11) => regA_ex_11_port, 
                           input(10) => regA_ex_10_port, input(9) => 
                           regA_ex_9_port, input(8) => regA_ex_8_port, input(7)
                           => regA_ex_7_port, input(6) => regA_ex_6_port, 
                           input(5) => regA_ex_5_port, input(4) => 
                           regA_ex_4_port, input(3) => regA_ex_3_port, input(2)
                           => regA_ex_2_port, input(1) => regA_ex_1_port, 
                           input(0) => regA_ex_0_port, res => is_zero);
   COND_OP : COND_BT_NBIT32 port map( ZERO_BIT => is_zero, OPCODE_0 => 
                           IR_26_ex_0_port, branch_op => branch_cond, con_sign 
                           => cond);
   MUX_alu_out : MUX21_GENERIC_NBIT32_4 port map( A(31) => LHI_ex_31_port, 
                           A(30) => LHI_ex_30_port, A(29) => LHI_ex_29_port, 
                           A(28) => LHI_ex_28_port, A(27) => LHI_ex_27_port, 
                           A(26) => LHI_ex_26_port, A(25) => LHI_ex_25_port, 
                           A(24) => LHI_ex_24_port, A(23) => LHI_ex_23_port, 
                           A(22) => LHI_ex_22_port, A(21) => LHI_ex_21_port, 
                           A(20) => LHI_ex_20_port, A(19) => LHI_ex_19_port, 
                           A(18) => LHI_ex_18_port, A(17) => LHI_ex_17_port, 
                           A(16) => LHI_ex_16_port, A(15) => LHI_ex_15_port, 
                           A(14) => LHI_ex_14_port, A(13) => LHI_ex_13_port, 
                           A(12) => LHI_ex_12_port, A(11) => LHI_ex_11_port, 
                           A(10) => LHI_ex_10_port, A(9) => LHI_ex_9_port, A(8)
                           => LHI_ex_8_port, A(7) => LHI_ex_7_port, A(6) => 
                           LHI_ex_6_port, A(5) => LHI_ex_5_port, A(4) => 
                           LHI_ex_4_port, A(3) => LHI_ex_3_port, A(2) => 
                           LHI_ex_2_port, A(1) => LHI_ex_1_port, A(0) => 
                           LHI_ex_0_port, B(31) => ALU_out_31_port, B(30) => 
                           ALU_out_30_port, B(29) => ALU_out_29_port, B(28) => 
                           ALU_out_28_port, B(27) => ALU_out_27_port, B(26) => 
                           ALU_out_26_port, B(25) => ALU_out_25_port, B(24) => 
                           ALU_out_24_port, B(23) => ALU_out_23_port, B(22) => 
                           ALU_out_22_port, B(21) => ALU_out_21_port, B(20) => 
                           ALU_out_20_port, B(19) => ALU_out_19_port, B(18) => 
                           ALU_out_18_port, B(17) => ALU_out_17_port, B(16) => 
                           ALU_out_16_port, B(15) => ALU_out_15_port, B(14) => 
                           ALU_out_14_port, B(13) => ALU_out_13_port, B(12) => 
                           ALU_out_12_port, B(11) => ALU_out_11_port, B(10) => 
                           ALU_out_10_port, B(9) => ALU_out_9_port, B(8) => 
                           ALU_out_8_port, B(7) => ALU_out_7_port, B(6) => 
                           ALU_out_6_port, B(5) => ALU_out_5_port, B(4) => 
                           ALU_out_4_port, B(3) => ALU_out_3_port, B(2) => 
                           ALU_out_2_port, B(1) => ALU_out_1_port, B(0) => 
                           ALU_out_0_port, SEL => lhi_sel, Y(31) => 
                           ALU_ex_31_port, Y(30) => ALU_ex_30_port, Y(29) => 
                           ALU_ex_29_port, Y(28) => ALU_ex_28_port, Y(27) => 
                           ALU_ex_27_port, Y(26) => ALU_ex_26_port, Y(25) => 
                           ALU_ex_25_port, Y(24) => ALU_ex_24_port, Y(23) => 
                           ALU_ex_23_port, Y(22) => ALU_ex_22_port, Y(21) => 
                           ALU_ex_21_port, Y(20) => ALU_ex_20_port, Y(19) => 
                           ALU_ex_19_port, Y(18) => ALU_ex_18_port, Y(17) => 
                           ALU_ex_17_port, Y(16) => ALU_ex_16_port, Y(15) => 
                           ALU_ex_15_port, Y(14) => ALU_ex_14_port, Y(13) => 
                           ALU_ex_13_port, Y(12) => ALU_ex_12_port, Y(11) => 
                           ALU_ex_11_port, Y(10) => ALU_ex_10_port, Y(9) => 
                           ALU_ex_9_port, Y(8) => ALU_ex_8_port, Y(7) => 
                           ALU_ex_7_port, Y(6) => ALU_ex_6_port, Y(5) => 
                           ALU_ex_5_port, Y(4) => ALU_ex_4_port, Y(3) => 
                           ALU_ex_3_port, Y(2) => ALU_ex_2_port, Y(1) => 
                           ALU_ex_1_port, Y(0) => ALU_ex_0_port);
   pipeline_sign3 : FF_6 port map( CLK => CLK, RESET => n45, EN => 
                           X_Logic1_port, D => signed_op_ex, Q => signed_op_mem
                           );
   pipeline_newpc3 : regFFD_NBIT32_5 port map( CK => CLK, RESET => n45, ENABLE 
                           => X_Logic1_port, D(31) => NPC_ex_31_port, D(30) => 
                           NPC_ex_30_port, D(29) => NPC_ex_29_port, D(28) => 
                           NPC_ex_28_port, D(27) => NPC_ex_27_port, D(26) => 
                           NPC_ex_26_port, D(25) => NPC_ex_25_port, D(24) => 
                           NPC_ex_24_port, D(23) => NPC_ex_23_port, D(22) => 
                           NPC_ex_22_port, D(21) => NPC_ex_21_port, D(20) => 
                           NPC_ex_20_port, D(19) => NPC_ex_19_port, D(18) => 
                           NPC_ex_18_port, D(17) => NPC_ex_17_port, D(16) => 
                           NPC_ex_16_port, D(15) => NPC_ex_15_port, D(14) => 
                           NPC_ex_14_port, D(13) => NPC_ex_13_port, D(12) => 
                           NPC_ex_12_port, D(11) => NPC_ex_11_port, D(10) => 
                           NPC_ex_10_port, D(9) => NPC_ex_9_port, D(8) => 
                           NPC_ex_8_port, D(7) => NPC_ex_7_port, D(6) => 
                           NPC_ex_6_port, D(5) => NPC_ex_5_port, D(4) => 
                           NPC_ex_4_port, D(3) => NPC_ex_3_port, D(2) => 
                           NPC_ex_2_port, D(1) => NPC_ex_1_port, D(0) => 
                           NPC_ex_0_port, Q(31) => NPC_mem_31_port, Q(30) => 
                           NPC_mem_30_port, Q(29) => NPC_mem_29_port, Q(28) => 
                           NPC_mem_28_port, Q(27) => NPC_mem_27_port, Q(26) => 
                           NPC_mem_26_port, Q(25) => NPC_mem_25_port, Q(24) => 
                           NPC_mem_24_port, Q(23) => NPC_mem_23_port, Q(22) => 
                           NPC_mem_22_port, Q(21) => NPC_mem_21_port, Q(20) => 
                           NPC_mem_20_port, Q(19) => NPC_mem_19_port, Q(18) => 
                           NPC_mem_18_port, Q(17) => NPC_mem_17_port, Q(16) => 
                           NPC_mem_16_port, Q(15) => NPC_mem_15_port, Q(14) => 
                           NPC_mem_14_port, Q(13) => NPC_mem_13_port, Q(12) => 
                           NPC_mem_12_port, Q(11) => NPC_mem_11_port, Q(10) => 
                           NPC_mem_10_port, Q(9) => NPC_mem_9_port, Q(8) => 
                           NPC_mem_8_port, Q(7) => NPC_mem_7_port, Q(6) => 
                           NPC_mem_6_port, Q(5) => NPC_mem_5_port, Q(4) => 
                           NPC_mem_4_port, Q(3) => NPC_mem_3_port, Q(2) => 
                           NPC_mem_2_port, Q(1) => NPC_mem_1_port, Q(0) => 
                           NPC_mem_0_port);
   pipeline_cond3 : FF_5 port map( CLK => CLK, RESET => n45, EN => 
                           X_Logic1_port, D => cond, Q => cond_mem);
   pipeline_B3 : regFFD_NBIT32_4 port map( CK => CLK, RESET => n44, ENABLE => 
                           X_Logic1_port, D(31) => regB_ex_31_port, D(30) => 
                           regB_ex_30_port, D(29) => regB_ex_29_port, D(28) => 
                           regB_ex_28_port, D(27) => regB_ex_27_port, D(26) => 
                           regB_ex_26_port, D(25) => regB_ex_25_port, D(24) => 
                           regB_ex_24_port, D(23) => regB_ex_23_port, D(22) => 
                           regB_ex_22_port, D(21) => regB_ex_21_port, D(20) => 
                           regB_ex_20_port, D(19) => regB_ex_19_port, D(18) => 
                           regB_ex_18_port, D(17) => regB_ex_17_port, D(16) => 
                           regB_ex_16_port, D(15) => regB_ex_15_port, D(14) => 
                           regB_ex_14_port, D(13) => regB_ex_13_port, D(12) => 
                           regB_ex_12_port, D(11) => regB_ex_11_port, D(10) => 
                           regB_ex_10_port, D(9) => regB_ex_9_port, D(8) => 
                           regB_ex_8_port, D(7) => regB_ex_7_port, D(6) => 
                           regB_ex_6_port, D(5) => regB_ex_5_port, D(4) => 
                           regB_ex_4_port, D(3) => regB_ex_3_port, D(2) => 
                           regB_ex_2_port, D(1) => regB_ex_1_port, D(0) => 
                           regB_ex_0_port, Q(31) => regB_mem_31_port, Q(30) => 
                           regB_mem_30_port, Q(29) => regB_mem_29_port, Q(28) 
                           => regB_mem_28_port, Q(27) => regB_mem_27_port, 
                           Q(26) => regB_mem_26_port, Q(25) => regB_mem_25_port
                           , Q(24) => regB_mem_24_port, Q(23) => 
                           regB_mem_23_port, Q(22) => regB_mem_22_port, Q(21) 
                           => regB_mem_21_port, Q(20) => regB_mem_20_port, 
                           Q(19) => regB_mem_19_port, Q(18) => regB_mem_18_port
                           , Q(17) => regB_mem_17_port, Q(16) => 
                           regB_mem_16_port, Q(15) => regB_mem_15_port, Q(14) 
                           => regB_mem_14_port, Q(13) => regB_mem_13_port, 
                           Q(12) => regB_mem_12_port, Q(11) => regB_mem_11_port
                           , Q(10) => regB_mem_10_port, Q(9) => regB_mem_9_port
                           , Q(8) => regB_mem_8_port, Q(7) => DATA_MEM_IN(7), 
                           Q(6) => DATA_MEM_IN(6), Q(5) => DATA_MEM_IN(5), Q(4)
                           => DATA_MEM_IN(4), Q(3) => DATA_MEM_IN(3), Q(2) => 
                           DATA_MEM_IN(2), Q(1) => DATA_MEM_IN(1), Q(0) => 
                           DATA_MEM_IN(0));
   pipeline_RD3 : regFFD_NBIT5_2 port map( CK => CLK, RESET => n44, ENABLE => 
                           X_Logic1_port, D(4) => RD_ex_4_port, D(3) => 
                           RD_ex_3_port, D(2) => RD_ex_2_port, D(1) => 
                           RD_ex_1_port, D(0) => RD_ex_0_port, Q(4) => 
                           RD_mem_4_port, Q(3) => RD_mem_3_port, Q(2) => 
                           RD_mem_2_port, Q(1) => RD_mem_1_port, Q(0) => 
                           RD_mem_0_port);
   pipeline_wr_signal2 : FF_4 port map( CLK => CLK, RESET => n45, EN => 
                           X_Logic1_port, D => wr_signal_exe, Q => 
                           wr_signal_mem);
   pipeline_IR3 : regFFD_NBIT6_1 port map( CK => CLK, RESET => n44, ENABLE => 
                           X_Logic1_port, D(5) => IR_26_ex_5_port, D(4) => 
                           IR_26_ex_4_port, D(3) => IR_26_ex_3_port, D(2) => 
                           IR_26_ex_2_port, D(1) => IR_26_ex_1_port, D(0) => 
                           IR_26_ex_0_port, Q(5) => IR_26_mem_5_port, Q(4) => 
                           IR_26_mem_4_port, Q(3) => IR_26_mem_3_port, Q(2) => 
                           IR_26_mem_2_port, Q(1) => IR_26_mem_1_port, Q(0) => 
                           IR_26_mem_0_port);
   MUX_PC : MUX21_GENERIC_NBIT32_3 port map( A(31) => ALU_ex_31_port, A(30) => 
                           ALU_ex_30_port, A(29) => ALU_ex_29_port, A(28) => 
                           ALU_ex_28_port, A(27) => ALU_ex_27_port, A(26) => 
                           ALU_ex_26_port, A(25) => ALU_ex_25_port, A(24) => 
                           ALU_ex_24_port, A(23) => ALU_ex_23_port, A(22) => 
                           ALU_ex_22_port, A(21) => ALU_ex_21_port, A(20) => 
                           ALU_ex_20_port, A(19) => ALU_ex_19_port, A(18) => 
                           ALU_ex_18_port, A(17) => ALU_ex_17_port, A(16) => 
                           ALU_ex_16_port, A(15) => ALU_ex_15_port, A(14) => 
                           ALU_ex_14_port, A(13) => ALU_ex_13_port, A(12) => 
                           ALU_ex_12_port, A(11) => ALU_ex_11_port, A(10) => 
                           ALU_ex_10_port, A(9) => ALU_ex_9_port, A(8) => 
                           ALU_ex_8_port, A(7) => ALU_ex_7_port, A(6) => 
                           ALU_ex_6_port, A(5) => ALU_ex_5_port, A(4) => 
                           ALU_ex_4_port, A(3) => ALU_ex_3_port, A(2) => 
                           ALU_ex_2_port, A(1) => ALU_ex_1_port, A(0) => 
                           ALU_ex_0_port, B(31) => NPC_mem_31_port, B(30) => 
                           NPC_mem_30_port, B(29) => NPC_mem_29_port, B(28) => 
                           NPC_mem_28_port, B(27) => NPC_mem_27_port, B(26) => 
                           NPC_mem_26_port, B(25) => NPC_mem_25_port, B(24) => 
                           NPC_mem_24_port, B(23) => NPC_mem_23_port, B(22) => 
                           NPC_mem_22_port, B(21) => NPC_mem_21_port, B(20) => 
                           NPC_mem_20_port, B(19) => NPC_mem_19_port, B(18) => 
                           NPC_mem_18_port, B(17) => NPC_mem_17_port, B(16) => 
                           NPC_mem_16_port, B(15) => NPC_mem_15_port, B(14) => 
                           NPC_mem_14_port, B(13) => NPC_mem_13_port, B(12) => 
                           NPC_mem_12_port, B(11) => NPC_mem_11_port, B(10) => 
                           NPC_mem_10_port, B(9) => NPC_mem_9_port, B(8) => 
                           NPC_mem_8_port, B(7) => NPC_mem_7_port, B(6) => 
                           NPC_mem_6_port, B(5) => NPC_mem_5_port, B(4) => 
                           NPC_mem_4_port, B(3) => NPC_mem_3_port, B(2) => 
                           NPC_mem_2_port, B(1) => NPC_mem_1_port, B(0) => 
                           NPC_mem_0_port, SEL => sel_npc, Y(31) => 
                           PC_OUT_i_31_port, Y(30) => PC_OUT_i_30_port, Y(29) 
                           => PC_OUT_i_29_port, Y(28) => PC_OUT_i_28_port, 
                           Y(27) => PC_OUT_i_27_port, Y(26) => PC_OUT_i_26_port
                           , Y(25) => PC_OUT_i_25_port, Y(24) => 
                           PC_OUT_i_24_port, Y(23) => PC_OUT_i_23_port, Y(22) 
                           => PC_OUT_i_22_port, Y(21) => PC_OUT_i_21_port, 
                           Y(20) => PC_OUT_i_20_port, Y(19) => PC_OUT_i_19_port
                           , Y(18) => PC_OUT_i_18_port, Y(17) => 
                           PC_OUT_i_17_port, Y(16) => PC_OUT_i_16_port, Y(15) 
                           => PC_OUT_i_15_port, Y(14) => PC_OUT_i_14_port, 
                           Y(13) => PC_OUT_i_13_port, Y(12) => PC_OUT_i_12_port
                           , Y(11) => PC_OUT_i_11_port, Y(10) => 
                           PC_OUT_i_10_port, Y(9) => PC_OUT_i_9_port, Y(8) => 
                           PC_OUT_i_8_port, Y(7) => PC_OUT_i_7_port, Y(6) => 
                           PC_OUT_i_6_port, Y(5) => PC_OUT_i_5_port, Y(4) => 
                           PC_OUT_i_4_port, Y(3) => PC_OUT_i_3_port, Y(2) => 
                           PC_OUT_i_2_port, Y(1) => PC_OUT_i_1_port, Y(0) => 
                           PC_OUT_i_0_port);
   LOAD_DATA_OUT : load_data port map( data_in(31) => DATA_MEM_OUT(31), 
                           data_in(30) => DATA_MEM_OUT(30), data_in(29) => 
                           DATA_MEM_OUT(29), data_in(28) => DATA_MEM_OUT(28), 
                           data_in(27) => DATA_MEM_OUT(27), data_in(26) => 
                           DATA_MEM_OUT(26), data_in(25) => DATA_MEM_OUT(25), 
                           data_in(24) => DATA_MEM_OUT(24), data_in(23) => 
                           DATA_MEM_OUT(23), data_in(22) => DATA_MEM_OUT(22), 
                           data_in(21) => DATA_MEM_OUT(21), data_in(20) => 
                           DATA_MEM_OUT(20), data_in(19) => DATA_MEM_OUT(19), 
                           data_in(18) => DATA_MEM_OUT(18), data_in(17) => 
                           DATA_MEM_OUT(17), data_in(16) => DATA_MEM_OUT(16), 
                           data_in(15) => DATA_MEM_OUT(15), data_in(14) => 
                           DATA_MEM_OUT(14), data_in(13) => DATA_MEM_OUT(13), 
                           data_in(12) => DATA_MEM_OUT(12), data_in(11) => 
                           DATA_MEM_OUT(11), data_in(10) => DATA_MEM_OUT(10), 
                           data_in(9) => DATA_MEM_OUT(9), data_in(8) => 
                           DATA_MEM_OUT(8), data_in(7) => DATA_MEM_OUT(7), 
                           data_in(6) => DATA_MEM_OUT(6), data_in(5) => 
                           DATA_MEM_OUT(5), data_in(4) => DATA_MEM_OUT(4), 
                           data_in(3) => DATA_MEM_OUT(3), data_in(2) => 
                           DATA_MEM_OUT(2), data_in(1) => DATA_MEM_OUT(1), 
                           data_in(0) => DATA_MEM_OUT(0), signed_val => 
                           signed_op_mem, load_op => RM, load_type(1) => 
                           IR_26_mem_1_port, load_type(0) => IR_26_mem_0_port, 
                           data_out(31) => LMD_out_31_port, data_out(30) => 
                           LMD_out_30_port, data_out(29) => LMD_out_29_port, 
                           data_out(28) => LMD_out_28_port, data_out(27) => 
                           LMD_out_27_port, data_out(26) => LMD_out_26_port, 
                           data_out(25) => LMD_out_25_port, data_out(24) => 
                           LMD_out_24_port, data_out(23) => LMD_out_23_port, 
                           data_out(22) => LMD_out_22_port, data_out(21) => 
                           LMD_out_21_port, data_out(20) => LMD_out_20_port, 
                           data_out(19) => LMD_out_19_port, data_out(18) => 
                           LMD_out_18_port, data_out(17) => LMD_out_17_port, 
                           data_out(16) => LMD_out_16_port, data_out(15) => 
                           LMD_out_15_port, data_out(14) => LMD_out_14_port, 
                           data_out(13) => LMD_out_13_port, data_out(12) => 
                           LMD_out_12_port, data_out(11) => LMD_out_11_port, 
                           data_out(10) => LMD_out_10_port, data_out(9) => 
                           LMD_out_9_port, data_out(8) => LMD_out_8_port, 
                           data_out(7) => LMD_out_7_port, data_out(6) => 
                           LMD_out_6_port, data_out(5) => LMD_out_5_port, 
                           data_out(4) => LMD_out_4_port, data_out(3) => 
                           LMD_out_3_port, data_out(2) => LMD_out_2_port, 
                           data_out(1) => LMD_out_1_port, data_out(0) => 
                           LMD_out_0_port);
   pipeline_alu4 : regFFD_NBIT32_3 port map( CK => CLK, RESET => n45, ENABLE =>
                           X_Logic1_port, D(31) => ALU_ex_31_port, D(30) => 
                           ALU_ex_30_port, D(29) => ALU_ex_29_port, D(28) => 
                           ALU_ex_28_port, D(27) => ALU_ex_27_port, D(26) => 
                           ALU_ex_26_port, D(25) => ALU_ex_25_port, D(24) => 
                           ALU_ex_24_port, D(23) => ALU_ex_23_port, D(22) => 
                           ALU_ex_22_port, D(21) => ALU_ex_21_port, D(20) => 
                           ALU_ex_20_port, D(19) => ALU_ex_19_port, D(18) => 
                           ALU_ex_18_port, D(17) => ALU_ex_17_port, D(16) => 
                           ALU_ex_16_port, D(15) => ALU_ex_15_port, D(14) => 
                           ALU_ex_14_port, D(13) => ALU_ex_13_port, D(12) => 
                           ALU_ex_12_port, D(11) => ALU_ex_11_port, D(10) => 
                           ALU_ex_10_port, D(9) => ALU_ex_9_port, D(8) => 
                           ALU_ex_8_port, D(7) => ALU_ex_7_port, D(6) => 
                           ALU_ex_6_port, D(5) => ALU_ex_5_port, D(4) => 
                           ALU_ex_4_port, D(3) => ALU_ex_3_port, D(2) => 
                           ALU_ex_2_port, D(1) => ALU_ex_1_port, D(0) => 
                           ALU_ex_0_port, Q(31) => ALU_wb_31_port, Q(30) => 
                           ALU_wb_30_port, Q(29) => ALU_wb_29_port, Q(28) => 
                           ALU_wb_28_port, Q(27) => ALU_wb_27_port, Q(26) => 
                           ALU_wb_26_port, Q(25) => ALU_wb_25_port, Q(24) => 
                           ALU_wb_24_port, Q(23) => ALU_wb_23_port, Q(22) => 
                           ALU_wb_22_port, Q(21) => ALU_wb_21_port, Q(20) => 
                           ALU_wb_20_port, Q(19) => ALU_wb_19_port, Q(18) => 
                           ALU_wb_18_port, Q(17) => ALU_wb_17_port, Q(16) => 
                           ALU_wb_16_port, Q(15) => ALU_wb_15_port, Q(14) => 
                           ALU_wb_14_port, Q(13) => ALU_wb_13_port, Q(12) => 
                           ALU_wb_12_port, Q(11) => ALU_wb_11_port, Q(10) => 
                           ALU_wb_10_port, Q(9) => ALU_wb_9_port, Q(8) => 
                           ALU_wb_8_port, Q(7) => ALU_wb_7_port, Q(6) => 
                           ALU_wb_6_port, Q(5) => ALU_wb_5_port, Q(4) => 
                           ALU_wb_4_port, Q(3) => ALU_wb_3_port, Q(2) => 
                           ALU_wb_2_port, Q(1) => ALU_wb_1_port, Q(0) => 
                           ALU_wb_0_port);
   pipeline_LMD4 : regFFD_NBIT32_2 port map( CK => CLK, RESET => n45, ENABLE =>
                           RM, D(31) => LMD_out_31_port, D(30) => 
                           LMD_out_30_port, D(29) => LMD_out_29_port, D(28) => 
                           LMD_out_28_port, D(27) => LMD_out_27_port, D(26) => 
                           LMD_out_26_port, D(25) => LMD_out_25_port, D(24) => 
                           LMD_out_24_port, D(23) => LMD_out_23_port, D(22) => 
                           LMD_out_22_port, D(21) => LMD_out_21_port, D(20) => 
                           LMD_out_20_port, D(19) => LMD_out_19_port, D(18) => 
                           LMD_out_18_port, D(17) => LMD_out_17_port, D(16) => 
                           LMD_out_16_port, D(15) => LMD_out_15_port, D(14) => 
                           LMD_out_14_port, D(13) => LMD_out_13_port, D(12) => 
                           LMD_out_12_port, D(11) => LMD_out_11_port, D(10) => 
                           LMD_out_10_port, D(9) => LMD_out_9_port, D(8) => 
                           LMD_out_8_port, D(7) => LMD_out_7_port, D(6) => 
                           LMD_out_6_port, D(5) => LMD_out_5_port, D(4) => 
                           LMD_out_4_port, D(3) => LMD_out_3_port, D(2) => 
                           LMD_out_2_port, D(1) => LMD_out_1_port, D(0) => 
                           LMD_out_0_port, Q(31) => LMD_wb_31_port, Q(30) => 
                           LMD_wb_30_port, Q(29) => LMD_wb_29_port, Q(28) => 
                           LMD_wb_28_port, Q(27) => LMD_wb_27_port, Q(26) => 
                           LMD_wb_26_port, Q(25) => LMD_wb_25_port, Q(24) => 
                           LMD_wb_24_port, Q(23) => LMD_wb_23_port, Q(22) => 
                           LMD_wb_22_port, Q(21) => LMD_wb_21_port, Q(20) => 
                           LMD_wb_20_port, Q(19) => LMD_wb_19_port, Q(18) => 
                           LMD_wb_18_port, Q(17) => LMD_wb_17_port, Q(16) => 
                           LMD_wb_16_port, Q(15) => LMD_wb_15_port, Q(14) => 
                           LMD_wb_14_port, Q(13) => LMD_wb_13_port, Q(12) => 
                           LMD_wb_12_port, Q(11) => LMD_wb_11_port, Q(10) => 
                           LMD_wb_10_port, Q(9) => LMD_wb_9_port, Q(8) => 
                           LMD_wb_8_port, Q(7) => LMD_wb_7_port, Q(6) => 
                           LMD_wb_6_port, Q(5) => LMD_wb_5_port, Q(4) => 
                           LMD_wb_4_port, Q(3) => LMD_wb_3_port, Q(2) => 
                           LMD_wb_2_port, Q(1) => LMD_wb_1_port, Q(0) => 
                           LMD_wb_0_port);
   pipeline_RD4 : regFFD_NBIT5_1 port map( CK => CLK, RESET => n44, ENABLE => 
                           X_Logic1_port, D(4) => RD_mem_4_port, D(3) => 
                           RD_mem_3_port, D(2) => RD_mem_2_port, D(1) => 
                           RD_mem_1_port, D(0) => RD_mem_0_port, Q(4) => 
                           RD_wb_4_port, Q(3) => RD_wb_3_port, Q(2) => 
                           RD_wb_2_port, Q(1) => RD_wb_1_port, Q(0) => 
                           RD_wb_0_port);
   pipeline_wr_signal3 : FF_3 port map( CLK => CLK, RESET => n45, EN => 
                           X_Logic1_port, D => wr_signal_mem1, Q => 
                           wr_signal_wb);
   pipeline_WM : FF_2 port map( CLK => CLK, RESET => n45, EN => X_Logic1_port, 
                           D => WM, Q => n_3111);
   pipeline_JAL : FF_1 port map( CLK => CLK, RESET => n45, EN => X_Logic1_port,
                           D => sel_saved_reg, Q => sel_saved_reg_wb);
   pipeline_NPC_wb : regFFD_NBIT32_1 port map( CK => CLK, RESET => n45, ENABLE 
                           => X_Logic1_port, D(31) => NPC_mem_31_port, D(30) =>
                           NPC_mem_30_port, D(29) => NPC_mem_29_port, D(28) => 
                           NPC_mem_28_port, D(27) => NPC_mem_27_port, D(26) => 
                           NPC_mem_26_port, D(25) => NPC_mem_25_port, D(24) => 
                           NPC_mem_24_port, D(23) => NPC_mem_23_port, D(22) => 
                           NPC_mem_22_port, D(21) => NPC_mem_21_port, D(20) => 
                           NPC_mem_20_port, D(19) => NPC_mem_19_port, D(18) => 
                           NPC_mem_18_port, D(17) => NPC_mem_17_port, D(16) => 
                           NPC_mem_16_port, D(15) => NPC_mem_15_port, D(14) => 
                           NPC_mem_14_port, D(13) => NPC_mem_13_port, D(12) => 
                           NPC_mem_12_port, D(11) => NPC_mem_11_port, D(10) => 
                           NPC_mem_10_port, D(9) => NPC_mem_9_port, D(8) => 
                           NPC_mem_8_port, D(7) => NPC_mem_7_port, D(6) => 
                           NPC_mem_6_port, D(5) => NPC_mem_5_port, D(4) => 
                           NPC_mem_4_port, D(3) => NPC_mem_3_port, D(2) => 
                           NPC_mem_2_port, D(1) => NPC_mem_1_port, D(0) => 
                           NPC_mem_0_port, Q(31) => NPC_wb_31_port, Q(30) => 
                           NPC_wb_30_port, Q(29) => NPC_wb_29_port, Q(28) => 
                           NPC_wb_28_port, Q(27) => NPC_wb_27_port, Q(26) => 
                           NPC_wb_26_port, Q(25) => NPC_wb_25_port, Q(24) => 
                           NPC_wb_24_port, Q(23) => NPC_wb_23_port, Q(22) => 
                           NPC_wb_22_port, Q(21) => NPC_wb_21_port, Q(20) => 
                           NPC_wb_20_port, Q(19) => NPC_wb_19_port, Q(18) => 
                           NPC_wb_18_port, Q(17) => NPC_wb_17_port, Q(16) => 
                           NPC_wb_16_port, Q(15) => NPC_wb_15_port, Q(14) => 
                           NPC_wb_14_port, Q(13) => NPC_wb_13_port, Q(12) => 
                           NPC_wb_12_port, Q(11) => NPC_wb_11_port, Q(10) => 
                           NPC_wb_10_port, Q(9) => NPC_wb_9_port, Q(8) => 
                           NPC_wb_8_port, Q(7) => NPC_wb_7_port, Q(6) => 
                           NPC_wb_6_port, Q(5) => NPC_wb_5_port, Q(4) => 
                           NPC_wb_4_port, Q(3) => NPC_wb_3_port, Q(2) => 
                           NPC_wb_2_port, Q(1) => NPC_wb_1_port, Q(0) => 
                           NPC_wb_0_port);
   MUX_WB : MUX21_GENERIC_NBIT32_2 port map( A(31) => ALU_wb_31_port, A(30) => 
                           ALU_wb_30_port, A(29) => ALU_wb_29_port, A(28) => 
                           ALU_wb_28_port, A(27) => ALU_wb_27_port, A(26) => 
                           ALU_wb_26_port, A(25) => ALU_wb_25_port, A(24) => 
                           ALU_wb_24_port, A(23) => ALU_wb_23_port, A(22) => 
                           ALU_wb_22_port, A(21) => ALU_wb_21_port, A(20) => 
                           ALU_wb_20_port, A(19) => ALU_wb_19_port, A(18) => 
                           ALU_wb_18_port, A(17) => ALU_wb_17_port, A(16) => 
                           ALU_wb_16_port, A(15) => ALU_wb_15_port, A(14) => 
                           ALU_wb_14_port, A(13) => ALU_wb_13_port, A(12) => 
                           ALU_wb_12_port, A(11) => ALU_wb_11_port, A(10) => 
                           ALU_wb_10_port, A(9) => ALU_wb_9_port, A(8) => 
                           ALU_wb_8_port, A(7) => ALU_wb_7_port, A(6) => 
                           ALU_wb_6_port, A(5) => ALU_wb_5_port, A(4) => 
                           ALU_wb_4_port, A(3) => ALU_wb_3_port, A(2) => 
                           ALU_wb_2_port, A(1) => ALU_wb_1_port, A(0) => 
                           ALU_wb_0_port, B(31) => LMD_wb_31_port, B(30) => 
                           LMD_wb_30_port, B(29) => LMD_wb_29_port, B(28) => 
                           LMD_wb_28_port, B(27) => LMD_wb_27_port, B(26) => 
                           LMD_wb_26_port, B(25) => LMD_wb_25_port, B(24) => 
                           LMD_wb_24_port, B(23) => LMD_wb_23_port, B(22) => 
                           LMD_wb_22_port, B(21) => LMD_wb_21_port, B(20) => 
                           LMD_wb_20_port, B(19) => LMD_wb_19_port, B(18) => 
                           LMD_wb_18_port, B(17) => LMD_wb_17_port, B(16) => 
                           LMD_wb_16_port, B(15) => LMD_wb_15_port, B(14) => 
                           LMD_wb_14_port, B(13) => LMD_wb_13_port, B(12) => 
                           LMD_wb_12_port, B(11) => LMD_wb_11_port, B(10) => 
                           LMD_wb_10_port, B(9) => LMD_wb_9_port, B(8) => 
                           LMD_wb_8_port, B(7) => LMD_wb_7_port, B(6) => 
                           LMD_wb_6_port, B(5) => LMD_wb_5_port, B(4) => 
                           LMD_wb_4_port, B(3) => LMD_wb_3_port, B(2) => 
                           LMD_wb_2_port, B(1) => LMD_wb_1_port, B(0) => 
                           LMD_wb_0_port, SEL => S3, Y(31) => OUT_data_31_port,
                           Y(30) => OUT_data_30_port, Y(29) => OUT_data_29_port
                           , Y(28) => OUT_data_28_port, Y(27) => 
                           OUT_data_27_port, Y(26) => OUT_data_26_port, Y(25) 
                           => OUT_data_25_port, Y(24) => OUT_data_24_port, 
                           Y(23) => OUT_data_23_port, Y(22) => OUT_data_22_port
                           , Y(21) => OUT_data_21_port, Y(20) => 
                           OUT_data_20_port, Y(19) => OUT_data_19_port, Y(18) 
                           => OUT_data_18_port, Y(17) => OUT_data_17_port, 
                           Y(16) => OUT_data_16_port, Y(15) => OUT_data_15_port
                           , Y(14) => OUT_data_14_port, Y(13) => 
                           OUT_data_13_port, Y(12) => OUT_data_12_port, Y(11) 
                           => OUT_data_11_port, Y(10) => OUT_data_10_port, Y(9)
                           => OUT_data_9_port, Y(8) => OUT_data_8_port, Y(7) =>
                           OUT_data_7_port, Y(6) => OUT_data_6_port, Y(5) => 
                           OUT_data_5_port, Y(4) => OUT_data_4_port, Y(3) => 
                           OUT_data_3_port, Y(2) => OUT_data_2_port, Y(1) => 
                           OUT_data_1_port, Y(0) => OUT_data_0_port);
   MUX_jal : MUX21_GENERIC_NBIT32_1 port map( A(31) => NPC_wb_31_port, A(30) =>
                           NPC_wb_30_port, A(29) => NPC_wb_29_port, A(28) => 
                           NPC_wb_28_port, A(27) => NPC_wb_27_port, A(26) => 
                           NPC_wb_26_port, A(25) => NPC_wb_25_port, A(24) => 
                           NPC_wb_24_port, A(23) => NPC_wb_23_port, A(22) => 
                           NPC_wb_22_port, A(21) => NPC_wb_21_port, A(20) => 
                           NPC_wb_20_port, A(19) => NPC_wb_19_port, A(18) => 
                           NPC_wb_18_port, A(17) => NPC_wb_17_port, A(16) => 
                           NPC_wb_16_port, A(15) => NPC_wb_15_port, A(14) => 
                           NPC_wb_14_port, A(13) => NPC_wb_13_port, A(12) => 
                           NPC_wb_12_port, A(11) => NPC_wb_11_port, A(10) => 
                           NPC_wb_10_port, A(9) => NPC_wb_9_port, A(8) => 
                           NPC_wb_8_port, A(7) => NPC_wb_7_port, A(6) => 
                           NPC_wb_6_port, A(5) => NPC_wb_5_port, A(4) => 
                           NPC_wb_4_port, A(3) => NPC_wb_3_port, A(2) => 
                           NPC_wb_2_port, A(1) => NPC_wb_1_port, A(0) => 
                           NPC_wb_0_port, B(31) => OUT_data_31_port, B(30) => 
                           OUT_data_30_port, B(29) => OUT_data_29_port, B(28) 
                           => OUT_data_28_port, B(27) => OUT_data_27_port, 
                           B(26) => OUT_data_26_port, B(25) => OUT_data_25_port
                           , B(24) => OUT_data_24_port, B(23) => 
                           OUT_data_23_port, B(22) => OUT_data_22_port, B(21) 
                           => OUT_data_21_port, B(20) => OUT_data_20_port, 
                           B(19) => OUT_data_19_port, B(18) => OUT_data_18_port
                           , B(17) => OUT_data_17_port, B(16) => 
                           OUT_data_16_port, B(15) => OUT_data_15_port, B(14) 
                           => OUT_data_14_port, B(13) => OUT_data_13_port, 
                           B(12) => OUT_data_12_port, B(11) => OUT_data_11_port
                           , B(10) => OUT_data_10_port, B(9) => OUT_data_9_port
                           , B(8) => OUT_data_8_port, B(7) => OUT_data_7_port, 
                           B(6) => OUT_data_6_port, B(5) => OUT_data_5_port, 
                           B(4) => OUT_data_4_port, B(3) => OUT_data_3_port, 
                           B(2) => OUT_data_2_port, B(1) => OUT_data_1_port, 
                           B(0) => OUT_data_0_port, SEL => sel_saved_reg_wb, 
                           Y(31) => OUT_wb_31_port, Y(30) => OUT_wb_30_port, 
                           Y(29) => OUT_wb_29_port, Y(28) => OUT_wb_28_port, 
                           Y(27) => OUT_wb_27_port, Y(26) => OUT_wb_26_port, 
                           Y(25) => OUT_wb_25_port, Y(24) => OUT_wb_24_port, 
                           Y(23) => OUT_wb_23_port, Y(22) => OUT_wb_22_port, 
                           Y(21) => OUT_wb_21_port, Y(20) => OUT_wb_20_port, 
                           Y(19) => OUT_wb_19_port, Y(18) => OUT_wb_18_port, 
                           Y(17) => OUT_wb_17_port, Y(16) => OUT_wb_16_port, 
                           Y(15) => OUT_wb_15_port, Y(14) => OUT_wb_14_port, 
                           Y(13) => OUT_wb_13_port, Y(12) => OUT_wb_12_port, 
                           Y(11) => OUT_wb_11_port, Y(10) => OUT_wb_10_port, 
                           Y(9) => OUT_wb_9_port, Y(8) => OUT_wb_8_port, Y(7) 
                           => OUT_wb_7_port, Y(6) => OUT_wb_6_port, Y(5) => 
                           OUT_wb_5_port, Y(4) => OUT_wb_4_port, Y(3) => 
                           OUT_wb_3_port, Y(2) => OUT_wb_2_port, Y(1) => 
                           OUT_wb_1_port, Y(0) => OUT_wb_0_port);
   add_240 : DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 port map( A(31) => 
                           PC_fetch0_31_port, A(30) => PC_fetch0_30_port, A(29)
                           => PC_fetch0_29_port, A(28) => PC_fetch0_28_port, 
                           A(27) => PC_fetch0_27_port, A(26) => 
                           PC_fetch0_26_port, A(25) => PC_fetch0_25_port, A(24)
                           => PC_fetch0_24_port, A(23) => PC_fetch0_23_port, 
                           A(22) => PC_fetch0_22_port, A(21) => 
                           PC_fetch0_21_port, A(20) => PC_fetch0_20_port, A(19)
                           => PC_fetch0_19_port, A(18) => PC_fetch0_18_port, 
                           A(17) => PC_fetch0_17_port, A(16) => 
                           PC_fetch0_16_port, A(15) => PC_fetch0_15_port, A(14)
                           => PC_fetch0_14_port, A(13) => PC_fetch0_13_port, 
                           A(12) => PC_fetch0_12_port, A(11) => 
                           PC_fetch0_11_port, A(10) => PC_fetch0_10_port, A(9) 
                           => PC_fetch0_9_port, A(8) => PC_fetch0_8_port, A(7) 
                           => PC_fetch0_7_port, A(6) => PC_fetch0_6_port, A(5) 
                           => PC_fetch0_5_port, A(4) => PC_fetch0_4_port, A(3) 
                           => PC_fetch0_3_port, A(2) => PC_fetch0_2_port, A(1) 
                           => PC_fetch0_1_port, A(0) => PC_fetch0_0_port, 
                           SUM(31) => NPC_31_port, SUM(30) => NPC_30_port, 
                           SUM(29) => NPC_29_port, SUM(28) => NPC_28_port, 
                           SUM(27) => NPC_27_port, SUM(26) => NPC_26_port, 
                           SUM(25) => NPC_25_port, SUM(24) => NPC_24_port, 
                           SUM(23) => NPC_23_port, SUM(22) => NPC_22_port, 
                           SUM(21) => NPC_21_port, SUM(20) => NPC_20_port, 
                           SUM(19) => NPC_19_port, SUM(18) => NPC_18_port, 
                           SUM(17) => NPC_17_port, SUM(16) => NPC_16_port, 
                           SUM(15) => NPC_15_port, SUM(14) => NPC_14_port, 
                           SUM(13) => NPC_13_port, SUM(12) => NPC_12_port, 
                           SUM(11) => NPC_11_port, SUM(10) => NPC_10_port, 
                           SUM(9) => NPC_9_port, SUM(8) => NPC_8_port, SUM(7) 
                           => NPC_7_port, SUM(6) => NPC_6_port, SUM(5) => 
                           NPC_5_port, SUM(4) => NPC_4_port, SUM(3) => 
                           NPC_3_port, SUM(2) => NPC_2_port, SUM(1) => 
                           NPC_1_port, SUM(0) => NPC_0_port);
   U3 : INV_X1 port map( A => n49, ZN => n35);
   U4 : INV_X1 port map( A => n48, ZN => n36);
   U5 : BUF_X2 port map( A => RST, Z => n45);
   U6 : BUF_X1 port map( A => n55, Z => n38);
   U7 : BUF_X1 port map( A => n55, Z => n37);
   U8 : BUF_X1 port map( A => n55, Z => n39);
   U9 : NOR4_X1 port map( A1 => n23, A2 => IR_Dec_22_port, A3 => IR_Dec_24_port
                           , A4 => IR_Dec_23_port, ZN => n20);
   U10 : OR4_X1 port map( A1 => IR_Dec_26_port, A2 => IR_Dec_25_port, A3 => 
                           IR_Dec_2_port, A4 => IR_Dec_28_port, ZN => n23);
   U11 : OAI22_X1 port map( A1 => IR_Dec_31_port, A2 => n13_port, B1 => n14, B2
                           => n48, ZN => n34);
   U12 : INV_X1 port map( A => IR_Dec_31_port, ZN => n48);
   U13 : NOR4_X1 port map( A1 => IR_Dec_30_port, A2 => IR_Dec_28_port, A3 => 
                           n49, A4 => n15, ZN => n14);
   U14 : AOI211_X1 port map( C1 => n16, C2 => n17, A => n35, B => 
                           IR_Dec_27_port, ZN => n13_port);
   U15 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           n17);
   U16 : NOR4_X1 port map( A1 => n22, A2 => IR_Dec_3_port, A3 => IR_Dec_5_port,
                           A4 => IR_Dec_4_port, ZN => n21);
   U17 : NOR4_X1 port map( A1 => n24, A2 => IR_Dec_16_port, A3 => 
                           IR_Dec_18_port, A4 => IR_Dec_17_port, ZN => n19);
   U18 : NOR4_X1 port map( A1 => n25, A2 => IR_Dec_0_port, A3 => IR_Dec_11_port
                           , A4 => IR_Dec_10_port, ZN => n18);
   U19 : AOI21_X1 port map( B1 => jump_en, B2 => n11, A => n47, ZN => 
                           wr_signal_mem1);
   U20 : NAND4_X1 port map( A1 => IR_26_mem_1_port, A2 => IR_26_mem_0_port, A3 
                           => n12, A4 => n46, ZN => n11);
   U21 : INV_X1 port map( A => wr_signal_mem, ZN => n47);
   U22 : INV_X1 port map( A => IR_26_mem_2_port, ZN => n46);
   U23 : OR4_X1 port map( A1 => IR_Dec_13_port, A2 => IR_Dec_12_port, A3 => 
                           IR_Dec_15_port, A4 => IR_Dec_14_port, ZN => n25);
   U24 : OR4_X1 port map( A1 => IR_Dec_1_port, A2 => IR_Dec_19_port, A3 => 
                           IR_Dec_21_port, A4 => IR_Dec_20_port, ZN => n24);
   U25 : OR4_X1 port map( A1 => IR_Dec_7_port, A2 => IR_Dec_6_port, A3 => 
                           IR_Dec_9_port, A4 => IR_Dec_8_port, ZN => n22);
   U26 : OAI21_X1 port map( B1 => IR_Dec_26_port, B2 => n50, A => 
                           IR_Dec_30_port, ZN => n16);
   U27 : INV_X1 port map( A => IR_Dec_28_port, ZN => n50);
   U28 : INV_X1 port map( A => IR_Dec_29_port, ZN => n49);
   U29 : AOI22_X1 port map( A1 => n30, A2 => instruction_alu(4), B1 => 
                           instruction_alu(3), B2 => n53, ZN => n29);
   U30 : INV_X1 port map( A => instruction_alu(4), ZN => n53);
   U31 : NOR2_X1 port map( A1 => instruction_alu(3), A2 => n54, ZN => n30);
   U32 : NAND4_X1 port map( A1 => IR_26_mem_2_port, A2 => IR_26_mem_0_port, A3 
                           => IR_26_mem_4_port, A4 => n26, ZN => N13);
   U33 : NOR3_X1 port map( A1 => IR_26_mem_1_port, A2 => IR_26_mem_5_port, A3 
                           => IR_26_mem_3_port, ZN => n26);
   U34 : BUF_X2 port map( A => RST, Z => n44);
   U35 : INV_X1 port map( A => instruction_alu(2), ZN => n52);
   U36 : INV_X1 port map( A => instruction_alu(0), ZN => n51);
   U37 : OR2_X1 port map( A1 => cond_mem, A2 => jump_en, ZN => sel_npc);
   U38 : INV_X1 port map( A => instruction_alu(5), ZN => n54);
   U39 : NOR2_X1 port map( A1 => IR_26_mem_5_port, A2 => IR_26_mem_3_port, ZN 
                           => n12);
   U40 : OR4_X1 port map( A1 => n27, A2 => n28, A3 => WM, A4 => RM, ZN => 
                           DATA_MEM_ENABLE);
   U41 : NOR4_X1 port map( A1 => n31, A2 => n54, A3 => instruction_alu(0), A4 
                           => instruction_alu(2), ZN => n27);
   U42 : NOR4_X1 port map( A1 => instruction_alu(1), A2 => n29, A3 => n52, A4 
                           => n51, ZN => n28);
   U43 : AND2_X1 port map( A1 => IR_26_mem_0_port, A2 => jump_en, ZN => 
                           sel_saved_reg);
   U44 : INV_X1 port map( A => sb_op, ZN => n55);
   U45 : AND2_X1 port map( A1 => regB_mem_31_port, A2 => n37, ZN => 
                           DATA_MEM_IN(31));
   U46 : AND2_X1 port map( A1 => regB_mem_30_port, A2 => n37, ZN => 
                           DATA_MEM_IN(30));
   U47 : AND2_X1 port map( A1 => regB_mem_29_port, A2 => n37, ZN => 
                           DATA_MEM_IN(29));
   U48 : AND2_X1 port map( A1 => regB_mem_28_port, A2 => n37, ZN => 
                           DATA_MEM_IN(28));
   U49 : AND2_X1 port map( A1 => regB_mem_27_port, A2 => n37, ZN => 
                           DATA_MEM_IN(27));
   U50 : AND2_X1 port map( A1 => regB_mem_26_port, A2 => n37, ZN => 
                           DATA_MEM_IN(26));
   U51 : AND2_X1 port map( A1 => regB_mem_25_port, A2 => n37, ZN => 
                           DATA_MEM_IN(25));
   U52 : AND2_X1 port map( A1 => regB_mem_24_port, A2 => n37, ZN => 
                           DATA_MEM_IN(24));
   U53 : AND2_X1 port map( A1 => regB_mem_23_port, A2 => n37, ZN => 
                           DATA_MEM_IN(23));
   U54 : AND2_X1 port map( A1 => regB_mem_22_port, A2 => n38, ZN => 
                           DATA_MEM_IN(22));
   U55 : AND2_X1 port map( A1 => regB_mem_21_port, A2 => n38, ZN => 
                           DATA_MEM_IN(21));
   U56 : AND2_X1 port map( A1 => regB_mem_20_port, A2 => n38, ZN => 
                           DATA_MEM_IN(20));
   U57 : AND2_X1 port map( A1 => regB_mem_19_port, A2 => n38, ZN => 
                           DATA_MEM_IN(19));
   U58 : AND2_X1 port map( A1 => regB_mem_18_port, A2 => n38, ZN => 
                           DATA_MEM_IN(18));
   U59 : AND2_X1 port map( A1 => regB_mem_17_port, A2 => n38, ZN => 
                           DATA_MEM_IN(17));
   U60 : AND2_X1 port map( A1 => regB_mem_16_port, A2 => n38, ZN => 
                           DATA_MEM_IN(16));
   U61 : AND2_X1 port map( A1 => regB_mem_15_port, A2 => n38, ZN => 
                           DATA_MEM_IN(15));
   U64 : AND2_X1 port map( A1 => regB_mem_14_port, A2 => n38, ZN => 
                           DATA_MEM_IN(14));
   U65 : AND2_X1 port map( A1 => regB_mem_13_port, A2 => n38, ZN => 
                           DATA_MEM_IN(13));
   U66 : AND2_X1 port map( A1 => regB_mem_12_port, A2 => n38, ZN => 
                           DATA_MEM_IN(12));
   U67 : AND2_X1 port map( A1 => regB_mem_9_port, A2 => n37, ZN => 
                           DATA_MEM_IN(9));
   U68 : AND2_X1 port map( A1 => regB_mem_8_port, A2 => n37, ZN => 
                           DATA_MEM_IN(8));
   U69 : AND2_X1 port map( A1 => regB_mem_11_port, A2 => n39, ZN => 
                           DATA_MEM_IN(11));
   U70 : AND2_X1 port map( A1 => regB_mem_10_port, A2 => n39, ZN => 
                           DATA_MEM_IN(10));
   U71 : CLKBUF_X1 port map( A => N13, Z => n40);
   U72 : CLKBUF_X1 port map( A => N13, Z => n41);
   U73 : CLKBUF_X1 port map( A => N13, Z => n42);
   U74 : CLKBUF_X1 port map( A => N13, Z => n43);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
         std_logic;  ALU_OPCODE : out std_logic_vector (0 to 5);  
         signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
         WB_MUX_SEL, RF_WE, lhi_sel, sb_op, s_trap, s_ret : out std_logic);

end dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_7
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_6
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal aluOpcode1_5_port, aluOpcode1_4_port, aluOpcode1_3_port, 
      aluOpcode1_2_port, aluOpcode1_1_port, aluOpcode1_0_port, 
      aluOpcode2_5_port, aluOpcode2_4_port, aluOpcode2_3_port, 
      aluOpcode2_2_port, aluOpcode2_1_port, aluOpcode2_0_port, 
      iterator_trap_31_port, iterator_trap_30_port, iterator_trap_29_port, 
      iterator_trap_28_port, iterator_trap_27_port, iterator_trap_26_port, 
      iterator_trap_25_port, iterator_trap_24_port, iterator_trap_23_port, 
      iterator_trap_22_port, iterator_trap_21_port, iterator_trap_20_port, 
      iterator_trap_19_port, iterator_trap_18_port, iterator_trap_17_port, 
      iterator_trap_16_port, iterator_trap_15_port, iterator_trap_14_port, 
      iterator_trap_13_port, iterator_trap_12_port, iterator_trap_11_port, 
      iterator_trap_10_port, iterator_trap_9_port, iterator_trap_8_port, 
      iterator_trap_7_port, iterator_trap_6_port, iterator_trap_5_port, 
      iterator_trap_4_port, iterator_trap_3_port, iterator_trap_2_port, 
      iterator_trap_1_port, iterator_trap_0_port, N40, N41, N42, N43, N44, N45,
      N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60
      , N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, 
      iterator_ret_31_port, iterator_ret_30_port, iterator_ret_29_port, 
      iterator_ret_28_port, iterator_ret_27_port, iterator_ret_26_port, 
      iterator_ret_25_port, iterator_ret_24_port, iterator_ret_23_port, 
      iterator_ret_22_port, iterator_ret_21_port, iterator_ret_20_port, 
      iterator_ret_19_port, iterator_ret_18_port, iterator_ret_17_port, 
      iterator_ret_16_port, iterator_ret_15_port, iterator_ret_14_port, 
      iterator_ret_13_port, iterator_ret_12_port, iterator_ret_11_port, 
      iterator_ret_10_port, iterator_ret_9_port, iterator_ret_8_port, 
      iterator_ret_7_port, iterator_ret_6_port, iterator_ret_5_port, 
      iterator_ret_4_port, iterator_ret_3_port, iterator_ret_2_port, 
      iterator_ret_1_port, iterator_ret_0_port, N151, N152, N153, N154, N155, 
      N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, 
      N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, 
      N180, N181, N182, iterator1_31_port, iterator1_30_port, iterator1_29_port
      , iterator1_28_port, iterator1_27_port, iterator1_26_port, 
      iterator1_25_port, iterator1_24_port, iterator1_23_port, 
      iterator1_22_port, iterator1_21_port, iterator1_20_port, 
      iterator1_19_port, iterator1_18_port, iterator1_17_port, 
      iterator1_16_port, iterator1_15_port, iterator1_14_port, 
      iterator1_13_port, iterator1_12_port, iterator1_11_port, 
      iterator1_10_port, iterator1_9_port, iterator1_8_port, iterator1_7_port, 
      iterator1_6_port, iterator1_5_port, iterator1_4_port, iterator1_3_port, 
      iterator1_2_port, iterator1_1_port, iterator1_0_port, N263, N264, N265, 
      N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, 
      N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, 
      N290, N291, N292, N293, N294, iterator2_31_port, iterator2_30_port, 
      iterator2_29_port, iterator2_28_port, iterator2_27_port, 
      iterator2_26_port, iterator2_25_port, iterator2_24_port, 
      iterator2_23_port, iterator2_22_port, iterator2_21_port, 
      iterator2_20_port, iterator2_19_port, iterator2_18_port, 
      iterator2_17_port, iterator2_16_port, iterator2_15_port, 
      iterator2_14_port, iterator2_13_port, iterator2_12_port, 
      iterator2_11_port, iterator2_10_port, iterator2_9_port, iterator2_8_port,
      iterator2_7_port, iterator2_6_port, iterator2_5_port, iterator2_4_port, 
      iterator2_3_port, iterator2_2_port, iterator2_1_port, iterator2_0_port, 
      N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, 
      N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, 
      N400, N401, N402, N403, N404, N405, N406, N407, aluOpcode_i_5_port, 
      aluOpcode_i_3_port, aluOpcode_i_2_port, aluOpcode_i_1_port, 
      aluOpcode_i_0_port, signed_unsigned_i, N717, N718, n323, n324, n325, n326
      , n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
      n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
      n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
      n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, 
      n375, n376_port, n377_port, n378_port, n379_port, n380_port, n381_port, 
      n382_port, n383_port, n384_port, n385_port, n386_port, n387_port, 
      n388_port, n389_port, n390_port, n391_port, n392_port, n393_port, 
      n394_port, n395_port, n396_port, n397_port, n398_port, n399_port, 
      n400_port, n401_port, n402_port, n403_port, n404_port, n405_port, 
      n406_port, n407_port, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n424, n425, n426, n428, n429, n430, n431, n432, n433, 
      n434, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n532, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n513, n514, n515, n516, n517, n518, n519, n520, n521, 
      n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n568, n569, 
      n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, 
      n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, 
      n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, 
      n606, n607, n608, n609, n610, n611, n612, n613, n183, n184, n200, n217, 
      n218, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263_port, n264_port, n265_port, n266_port, n267_port, n268_port, 
      n269_port, n270_port, n271_port, n272_port, n273_port, n274_port, 
      n275_port, n276_port, n277_port, n278_port, n279_port, n280_port, 
      n281_port, n282_port, n283_port, n284_port, n285_port, n286_port, 
      n287_port, n288_port, n289_port, n290_port, n291_port, n292_port, 
      n293_port, n294_port, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
      n315, n316, n317, n318, n319, n320, n321, n322, n419, n420, n421, n422, 
      n423, n427, n435, n499, n500, n503, n504, n505, n506, n507, n509, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717_port, n718_port, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n773, n774, n775, n776, n777, n778, n779, n780, n781, 
      n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, 
      n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, 
      n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, 
      n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
      n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, 
      n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, 
      n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, 
      n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, 
      n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, 
      n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, 
      n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, 
      n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, 
      n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, 
      n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, 
      n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, 
      n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, 
      n974, n975, n976, n977, n978, n979, n980, n_3112, n_3113, n_3114, n_3115,
      n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, 
      n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, 
      n_3134, n_3135 : std_logic;

begin
   
   aluOpcode1_reg_5_inst : DFFR_X1 port map( D => aluOpcode_i_5_port, CK => Clk
                           , RN => n774, Q => aluOpcode1_5_port, QN => n_3112);
   aluOpcode1_reg_4_inst : DFFR_X1 port map( D => n565, CK => Clk, RN => Rst, Q
                           => aluOpcode1_4_port, QN => n_3113);
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_3_port, QN => n_3114);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_2_port, QN => n_3115);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , RN => Rst, Q => aluOpcode1_1_port, QN => n_3116);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => n774, Q => aluOpcode1_0_port, QN => n_3117);
   aluOpcode2_reg_5_inst : DFFR_X1 port map( D => aluOpcode1_5_port, CK => Clk,
                           RN => n774, Q => aluOpcode2_5_port, QN => n_3118);
   aluOpcode2_reg_4_inst : DFFR_X1 port map( D => aluOpcode1_4_port, CK => Clk,
                           RN => n774, Q => aluOpcode2_4_port, QN => n_3119);
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => aluOpcode1_3_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_3_port, QN => n_3120);
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => aluOpcode1_2_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_2_port, QN => n_3121);
   aluOpcode2_reg_1_inst : DFFR_X1 port map( D => aluOpcode1_1_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_1_port, QN => n_3122);
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => aluOpcode1_0_port, CK => Clk,
                           RN => Rst, Q => aluOpcode2_0_port, QN => n_3123);
   aluOpcode3_reg_4_inst : DFFR_X1 port map( D => aluOpcode2_4_port, CK => Clk,
                           RN => n774, Q => ALU_OPCODE(1), QN => n_3124);
   aluOpcode3_reg_3_inst : DFFR_X1 port map( D => aluOpcode2_3_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(2), QN => n_3125);
   aluOpcode3_reg_2_inst : DFFR_X1 port map( D => aluOpcode2_2_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(3), QN => n_3126);
   aluOpcode3_reg_1_inst : DFFR_X1 port map( D => aluOpcode2_1_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(4), QN => n_3127);
   aluOpcode3_reg_0_inst : DFFR_X1 port map( D => aluOpcode2_0_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(5), QN => n_3128);
   iterator_trap_reg_0_inst : DFF_X1 port map( D => n507, CK => Clk, Q => 
                           iterator_trap_0_port, QN => n323);
   s_trap_reg : DFF_X1 port map( D => n434, CK => Clk, Q => s_trap, QN => n424)
                           ;
   iterator_trap_reg_30_inst : DFF_X1 port map( D => n465, CK => Clk, Q => 
                           iterator_trap_30_port, QN => n353);
   iterator_trap_reg_29_inst : DFF_X1 port map( D => n464, CK => Clk, Q => 
                           iterator_trap_29_port, QN => n352);
   iterator_trap_reg_28_inst : DFF_X1 port map( D => n463, CK => Clk, Q => 
                           iterator_trap_28_port, QN => n351);
   iterator_trap_reg_27_inst : DFF_X1 port map( D => n462, CK => Clk, Q => 
                           iterator_trap_27_port, QN => n350);
   iterator_trap_reg_26_inst : DFF_X1 port map( D => n461, CK => Clk, Q => 
                           iterator_trap_26_port, QN => n349);
   iterator_trap_reg_25_inst : DFF_X1 port map( D => n460, CK => Clk, Q => 
                           iterator_trap_25_port, QN => n348);
   iterator_trap_reg_24_inst : DFF_X1 port map( D => n459, CK => Clk, Q => 
                           iterator_trap_24_port, QN => n347);
   iterator_trap_reg_23_inst : DFF_X1 port map( D => n458, CK => Clk, Q => 
                           iterator_trap_23_port, QN => n346);
   iterator_trap_reg_22_inst : DFF_X1 port map( D => n457, CK => Clk, Q => 
                           iterator_trap_22_port, QN => n345);
   iterator_trap_reg_21_inst : DFF_X1 port map( D => n456, CK => Clk, Q => 
                           iterator_trap_21_port, QN => n344);
   iterator_trap_reg_20_inst : DFF_X1 port map( D => n455, CK => Clk, Q => 
                           iterator_trap_20_port, QN => n343);
   iterator_trap_reg_19_inst : DFF_X1 port map( D => n454, CK => Clk, Q => 
                           iterator_trap_19_port, QN => n342);
   iterator_trap_reg_18_inst : DFF_X1 port map( D => n453, CK => Clk, Q => 
                           iterator_trap_18_port, QN => n341);
   iterator_trap_reg_17_inst : DFF_X1 port map( D => n452, CK => Clk, Q => 
                           iterator_trap_17_port, QN => n340);
   iterator_trap_reg_16_inst : DFF_X1 port map( D => n451, CK => Clk, Q => 
                           iterator_trap_16_port, QN => n339);
   iterator_trap_reg_15_inst : DFF_X1 port map( D => n450, CK => Clk, Q => 
                           iterator_trap_15_port, QN => n338);
   iterator_trap_reg_14_inst : DFF_X1 port map( D => n449, CK => Clk, Q => 
                           iterator_trap_14_port, QN => n337);
   iterator_trap_reg_13_inst : DFF_X1 port map( D => n448, CK => Clk, Q => 
                           iterator_trap_13_port, QN => n336);
   iterator_trap_reg_12_inst : DFF_X1 port map( D => n447, CK => Clk, Q => 
                           iterator_trap_12_port, QN => n335);
   iterator_trap_reg_11_inst : DFF_X1 port map( D => n446, CK => Clk, Q => 
                           iterator_trap_11_port, QN => n334);
   iterator_trap_reg_10_inst : DFF_X1 port map( D => n445, CK => Clk, Q => 
                           iterator_trap_10_port, QN => n333);
   iterator_trap_reg_9_inst : DFF_X1 port map( D => n444, CK => Clk, Q => 
                           iterator_trap_9_port, QN => n332);
   iterator_trap_reg_8_inst : DFF_X1 port map( D => n443, CK => Clk, Q => 
                           iterator_trap_8_port, QN => n331);
   iterator_trap_reg_7_inst : DFF_X1 port map( D => n442, CK => Clk, Q => 
                           iterator_trap_7_port, QN => n330);
   iterator_trap_reg_6_inst : DFF_X1 port map( D => n441, CK => Clk, Q => 
                           iterator_trap_6_port, QN => n329);
   iterator_trap_reg_5_inst : DFF_X1 port map( D => n440, CK => Clk, Q => 
                           iterator_trap_5_port, QN => n328);
   iterator_trap_reg_4_inst : DFF_X1 port map( D => n439, CK => Clk, Q => 
                           iterator_trap_4_port, QN => n327);
   iterator_trap_reg_3_inst : DFF_X1 port map( D => n438, CK => Clk, Q => 
                           iterator_trap_3_port, QN => n326);
   iterator_trap_reg_2_inst : DFF_X1 port map( D => n437, CK => Clk, Q => 
                           iterator_trap_2_port, QN => n325);
   iterator_trap_reg_1_inst : DFF_X1 port map( D => n436, CK => Clk, Q => 
                           iterator_trap_1_port, QN => n324);
   iterator_trap_reg_31_inst : DFF_X1 port map( D => n466, CK => Clk, Q => 
                           iterator_trap_31_port, QN => n354);
   iterator_ret_reg_0_inst : DFF_X1 port map( D => n467, CK => Clk, Q => 
                           iterator_ret_0_port, QN => n355);
   s_ret_reg : DFF_X1 port map( D => n433, CK => Clk, Q => s_ret, QN => n425);
   iterator_ret_reg_30_inst : DFF_X1 port map( D => n497, CK => Clk, Q => 
                           iterator_ret_30_port, QN => n385_port);
   iterator_ret_reg_29_inst : DFF_X1 port map( D => n496, CK => Clk, Q => 
                           iterator_ret_29_port, QN => n384_port);
   iterator_ret_reg_28_inst : DFF_X1 port map( D => n495, CK => Clk, Q => 
                           iterator_ret_28_port, QN => n383_port);
   iterator_ret_reg_27_inst : DFF_X1 port map( D => n494, CK => Clk, Q => 
                           iterator_ret_27_port, QN => n382_port);
   iterator_ret_reg_26_inst : DFF_X1 port map( D => n493, CK => Clk, Q => 
                           iterator_ret_26_port, QN => n381_port);
   iterator_ret_reg_25_inst : DFF_X1 port map( D => n492, CK => Clk, Q => 
                           iterator_ret_25_port, QN => n380_port);
   iterator_ret_reg_24_inst : DFF_X1 port map( D => n491, CK => Clk, Q => 
                           iterator_ret_24_port, QN => n379_port);
   iterator_ret_reg_23_inst : DFF_X1 port map( D => n490, CK => Clk, Q => 
                           iterator_ret_23_port, QN => n378_port);
   iterator_ret_reg_22_inst : DFF_X1 port map( D => n489, CK => Clk, Q => 
                           iterator_ret_22_port, QN => n377_port);
   iterator_ret_reg_21_inst : DFF_X1 port map( D => n488, CK => Clk, Q => 
                           iterator_ret_21_port, QN => n376_port);
   iterator_ret_reg_20_inst : DFF_X1 port map( D => n487, CK => Clk, Q => 
                           iterator_ret_20_port, QN => n375);
   iterator_ret_reg_19_inst : DFF_X1 port map( D => n486, CK => Clk, Q => 
                           iterator_ret_19_port, QN => n374);
   iterator_ret_reg_18_inst : DFF_X1 port map( D => n485, CK => Clk, Q => 
                           iterator_ret_18_port, QN => n373);
   iterator_ret_reg_17_inst : DFF_X1 port map( D => n484, CK => Clk, Q => 
                           iterator_ret_17_port, QN => n372);
   iterator_ret_reg_16_inst : DFF_X1 port map( D => n483, CK => Clk, Q => 
                           iterator_ret_16_port, QN => n371);
   iterator_ret_reg_15_inst : DFF_X1 port map( D => n482, CK => Clk, Q => 
                           iterator_ret_15_port, QN => n370);
   iterator_ret_reg_14_inst : DFF_X1 port map( D => n481, CK => Clk, Q => 
                           iterator_ret_14_port, QN => n369);
   iterator_ret_reg_13_inst : DFF_X1 port map( D => n480, CK => Clk, Q => 
                           iterator_ret_13_port, QN => n368);
   iterator_ret_reg_12_inst : DFF_X1 port map( D => n479, CK => Clk, Q => 
                           iterator_ret_12_port, QN => n367);
   iterator_ret_reg_11_inst : DFF_X1 port map( D => n478, CK => Clk, Q => 
                           iterator_ret_11_port, QN => n366);
   iterator_ret_reg_10_inst : DFF_X1 port map( D => n477, CK => Clk, Q => 
                           iterator_ret_10_port, QN => n365);
   iterator_ret_reg_9_inst : DFF_X1 port map( D => n476, CK => Clk, Q => 
                           iterator_ret_9_port, QN => n364);
   iterator_ret_reg_8_inst : DFF_X1 port map( D => n475, CK => Clk, Q => 
                           iterator_ret_8_port, QN => n363);
   iterator_ret_reg_7_inst : DFF_X1 port map( D => n474, CK => Clk, Q => 
                           iterator_ret_7_port, QN => n362);
   iterator_ret_reg_6_inst : DFF_X1 port map( D => n473, CK => Clk, Q => 
                           iterator_ret_6_port, QN => n361);
   iterator_ret_reg_5_inst : DFF_X1 port map( D => n472, CK => Clk, Q => 
                           iterator_ret_5_port, QN => n360);
   iterator_ret_reg_4_inst : DFF_X1 port map( D => n471, CK => Clk, Q => 
                           iterator_ret_4_port, QN => n359);
   iterator_ret_reg_3_inst : DFF_X1 port map( D => n470, CK => Clk, Q => 
                           iterator_ret_3_port, QN => n358);
   iterator_ret_reg_2_inst : DFF_X1 port map( D => n469, CK => Clk, Q => 
                           iterator_ret_2_port, QN => n357);
   iterator_ret_reg_1_inst : DFF_X1 port map( D => n468, CK => Clk, Q => 
                           iterator_ret_1_port, QN => n356);
   iterator_ret_reg_31_inst : DFF_X1 port map( D => n498, CK => Clk, Q => 
                           iterator_ret_31_port, QN => n386_port);
   iterator1_reg_0_inst : DFF_X1 port map( D => n612, CK => Clk, Q => 
                           iterator1_0_port, QN => n513);
   iterator1_reg_30_inst : DFF_X1 port map( D => n582, CK => Clk, Q => 
                           iterator1_30_port, QN => n579);
   iterator1_reg_29_inst : DFF_X1 port map( D => n583, CK => Clk, Q => 
                           iterator1_29_port, QN => n578);
   iterator1_reg_28_inst : DFF_X1 port map( D => n584, CK => Clk, Q => 
                           iterator1_28_port, QN => n577);
   iterator1_reg_27_inst : DFF_X1 port map( D => n585, CK => Clk, Q => 
                           iterator1_27_port, QN => n576);
   iterator1_reg_26_inst : DFF_X1 port map( D => n586, CK => Clk, Q => 
                           iterator1_26_port, QN => n575);
   iterator1_reg_25_inst : DFF_X1 port map( D => n587, CK => Clk, Q => 
                           iterator1_25_port, QN => n574);
   iterator1_reg_24_inst : DFF_X1 port map( D => n588, CK => Clk, Q => 
                           iterator1_24_port, QN => n573);
   iterator1_reg_23_inst : DFF_X1 port map( D => n589, CK => Clk, Q => 
                           iterator1_23_port, QN => n572);
   iterator1_reg_22_inst : DFF_X1 port map( D => n590, CK => Clk, Q => 
                           iterator1_22_port, QN => n571);
   iterator1_reg_21_inst : DFF_X1 port map( D => n591, CK => Clk, Q => 
                           iterator1_21_port, QN => n570);
   iterator1_reg_20_inst : DFF_X1 port map( D => n592, CK => Clk, Q => 
                           iterator1_20_port, QN => n569);
   iterator1_reg_19_inst : DFF_X1 port map( D => n593, CK => Clk, Q => 
                           iterator1_19_port, QN => n568);
   iterator1_reg_18_inst : DFF_X1 port map( D => n594, CK => Clk, Q => 
                           iterator1_18_port, QN => n531);
   iterator1_reg_17_inst : DFF_X1 port map( D => n595, CK => Clk, Q => 
                           iterator1_17_port, QN => n530);
   iterator1_reg_16_inst : DFF_X1 port map( D => n596, CK => Clk, Q => 
                           iterator1_16_port, QN => n529);
   iterator1_reg_15_inst : DFF_X1 port map( D => n597, CK => Clk, Q => 
                           iterator1_15_port, QN => n528);
   iterator1_reg_14_inst : DFF_X1 port map( D => n598, CK => Clk, Q => 
                           iterator1_14_port, QN => n527);
   iterator1_reg_13_inst : DFF_X1 port map( D => n599, CK => Clk, Q => 
                           iterator1_13_port, QN => n526);
   iterator1_reg_12_inst : DFF_X1 port map( D => n600, CK => Clk, Q => 
                           iterator1_12_port, QN => n525);
   iterator1_reg_11_inst : DFF_X1 port map( D => n601, CK => Clk, Q => 
                           iterator1_11_port, QN => n524);
   iterator1_reg_10_inst : DFF_X1 port map( D => n602, CK => Clk, Q => 
                           iterator1_10_port, QN => n523);
   iterator1_reg_9_inst : DFF_X1 port map( D => n603, CK => Clk, Q => 
                           iterator1_9_port, QN => n522);
   iterator1_reg_8_inst : DFF_X1 port map( D => n604, CK => Clk, Q => 
                           iterator1_8_port, QN => n521);
   iterator1_reg_7_inst : DFF_X1 port map( D => n605, CK => Clk, Q => 
                           iterator1_7_port, QN => n520);
   iterator1_reg_6_inst : DFF_X1 port map( D => n606, CK => Clk, Q => 
                           iterator1_6_port, QN => n519);
   iterator1_reg_5_inst : DFF_X1 port map( D => n607, CK => Clk, Q => 
                           iterator1_5_port, QN => n518);
   iterator1_reg_4_inst : DFF_X1 port map( D => n608, CK => Clk, Q => 
                           iterator1_4_port, QN => n517);
   iterator1_reg_3_inst : DFF_X1 port map( D => n609, CK => Clk, Q => 
                           iterator1_3_port, QN => n516);
   iterator1_reg_2_inst : DFF_X1 port map( D => n610, CK => Clk, Q => 
                           iterator1_2_port, QN => n515);
   iterator1_reg_1_inst : DFF_X1 port map( D => n611, CK => Clk, Q => 
                           iterator1_1_port, QN => n514);
   iterator1_reg_31_inst : DFF_X1 port map( D => n581, CK => Clk, Q => 
                           iterator1_31_port, QN => n580);
   iterator2_reg_0_inst : DFF_X1 port map( D => n509, CK => Clk, Q => 
                           iterator2_0_port, QN => n387_port);
   sig3_reg : DFF_X1 port map( D => n532, CK => Clk, Q => n503, QN => n_3129);
   iterator2_reg_30_inst : DFF_X1 port map( D => n563, CK => Clk, Q => 
                           iterator2_30_port, QN => n417);
   iterator2_reg_29_inst : DFF_X1 port map( D => n562, CK => Clk, Q => 
                           iterator2_29_port, QN => n416);
   iterator2_reg_28_inst : DFF_X1 port map( D => n561, CK => Clk, Q => 
                           iterator2_28_port, QN => n415);
   iterator2_reg_27_inst : DFF_X1 port map( D => n560, CK => Clk, Q => 
                           iterator2_27_port, QN => n414);
   iterator2_reg_26_inst : DFF_X1 port map( D => n559, CK => Clk, Q => 
                           iterator2_26_port, QN => n413);
   iterator2_reg_25_inst : DFF_X1 port map( D => n558, CK => Clk, Q => 
                           iterator2_25_port, QN => n412);
   iterator2_reg_24_inst : DFF_X1 port map( D => n557, CK => Clk, Q => 
                           iterator2_24_port, QN => n411);
   iterator2_reg_23_inst : DFF_X1 port map( D => n556, CK => Clk, Q => 
                           iterator2_23_port, QN => n410);
   iterator2_reg_22_inst : DFF_X1 port map( D => n555, CK => Clk, Q => 
                           iterator2_22_port, QN => n409);
   iterator2_reg_21_inst : DFF_X1 port map( D => n554, CK => Clk, Q => 
                           iterator2_21_port, QN => n408);
   iterator2_reg_20_inst : DFF_X1 port map( D => n553, CK => Clk, Q => 
                           iterator2_20_port, QN => n407_port);
   iterator2_reg_19_inst : DFF_X1 port map( D => n552, CK => Clk, Q => 
                           iterator2_19_port, QN => n406_port);
   iterator2_reg_18_inst : DFF_X1 port map( D => n551, CK => Clk, Q => 
                           iterator2_18_port, QN => n405_port);
   iterator2_reg_17_inst : DFF_X1 port map( D => n550, CK => Clk, Q => 
                           iterator2_17_port, QN => n404_port);
   iterator2_reg_16_inst : DFF_X1 port map( D => n549, CK => Clk, Q => 
                           iterator2_16_port, QN => n403_port);
   iterator2_reg_15_inst : DFF_X1 port map( D => n548, CK => Clk, Q => 
                           iterator2_15_port, QN => n402_port);
   iterator2_reg_14_inst : DFF_X1 port map( D => n547, CK => Clk, Q => 
                           iterator2_14_port, QN => n401_port);
   iterator2_reg_13_inst : DFF_X1 port map( D => n546, CK => Clk, Q => 
                           iterator2_13_port, QN => n400_port);
   iterator2_reg_12_inst : DFF_X1 port map( D => n545, CK => Clk, Q => 
                           iterator2_12_port, QN => n399_port);
   iterator2_reg_11_inst : DFF_X1 port map( D => n544, CK => Clk, Q => 
                           iterator2_11_port, QN => n398_port);
   iterator2_reg_10_inst : DFF_X1 port map( D => n543, CK => Clk, Q => 
                           iterator2_10_port, QN => n397_port);
   iterator2_reg_9_inst : DFF_X1 port map( D => n542, CK => Clk, Q => 
                           iterator2_9_port, QN => n396_port);
   iterator2_reg_8_inst : DFF_X1 port map( D => n541, CK => Clk, Q => 
                           iterator2_8_port, QN => n395_port);
   iterator2_reg_7_inst : DFF_X1 port map( D => n540, CK => Clk, Q => 
                           iterator2_7_port, QN => n394_port);
   iterator2_reg_6_inst : DFF_X1 port map( D => n539, CK => Clk, Q => 
                           iterator2_6_port, QN => n393_port);
   iterator2_reg_5_inst : DFF_X1 port map( D => n538, CK => Clk, Q => 
                           iterator2_5_port, QN => n392_port);
   iterator2_reg_4_inst : DFF_X1 port map( D => n537, CK => Clk, Q => 
                           iterator2_4_port, QN => n391_port);
   iterator2_reg_3_inst : DFF_X1 port map( D => n536, CK => Clk, Q => 
                           iterator2_3_port, QN => n390_port);
   iterator2_reg_2_inst : DFF_X1 port map( D => n535, CK => Clk, Q => 
                           iterator2_2_port, QN => n389_port);
   iterator2_reg_1_inst : DFF_X1 port map( D => n534, CK => Clk, Q => 
                           iterator2_1_port, QN => n388_port);
   sb_op_reg : DFF_X1 port map( D => n431, CK => Clk, Q => sb_op, QN => n426);
   iterator2_reg_31_inst : DFF_X1 port map( D => n564, CK => Clk, Q => 
                           iterator2_31_port, QN => n418);
   signed_unsigned_i_reg : DLH_X1 port map( G => N717, D => N718, Q => 
                           signed_unsigned_i);
   signed_unsigned_1_reg : DFF_X1 port map( D => n430, CK => Clk, Q => n_3130, 
                           QN => n504);
   signed_unsigned_2_reg : DFF_X1 port map( D => n429, CK => Clk, Q => n_3131, 
                           QN => n505);
   signed_unsigned_3_reg : DFF_X1 port map( D => n428, CK => Clk, Q => 
                           signed_unsigned, QN => n506);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   PC_LATCH_EN <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   NPC_LATCH_EN <= '0';
   IR_LATCH_EN <= '0';
   U235 : NOR4_X2 port map( A1 => n976, A2 => n980, A3 => IR_IN(29), A4 => 
                           IR_IN(31), ZN => n244);
   U277 : NOR4_X2 port map( A1 => IR_IN(6), A2 => IR_IN(10), A3 => n307, A4 => 
                           n499, ZN => n245);
   U463 : NAND3_X1 port map( A1 => n241, A2 => n242, A3 => n243, ZN => 
                           aluOpcode_i_5_port);
   U479 : NAND3_X1 port map( A1 => n263_port, A2 => n950, A3 => n264_port, ZN 
                           => aluOpcode_i_2_port);
   U480 : NAND3_X1 port map( A1 => n239, A2 => n971, A3 => n277_port, ZN => 
                           n270_port);
   U481 : NAND3_X1 port map( A1 => n291_port, A2 => n200, A3 => n217, ZN => 
                           n290_port);
   U482 : NAND3_X1 port map( A1 => n248, A2 => n954, A3 => n268_port, ZN => 
                           n299);
   U483 : NAND3_X1 port map( A1 => n217, A2 => n303, A3 => n281_port, ZN => 
                           n294_port);
   U484 : NAND3_X1 port map( A1 => n304, A2 => n963, A3 => n305, ZN => N718);
   U485 : NAND3_X1 port map( A1 => n256, A2 => n242, A3 => n314, ZN => n309);
   U486 : NAND3_X1 port map( A1 => n976, A2 => n980, A3 => n320, ZN => n255);
   U487 : NAND3_X1 port map( A1 => n955, A2 => n957, A3 => n322, ZN => 
                           n268_port);
   U488 : NAND3_X1 port map( A1 => n322, A2 => n957, A3 => IR_IN(2), ZN => n259
                           );
   U490 : NAND3_X1 port map( A1 => n976, A2 => n980, A3 => IR_IN(31), ZN => 
                           n319);
   U491 : NAND3_X1 port map( A1 => n979, A2 => n980, A3 => IR_IN(28), ZN => 
                           n292_port);
   U492 : NAND3_X1 port map( A1 => n320, A2 => n980, A3 => IR_IN(28), ZN => 
                           n217);
   U493 : NAND3_X1 port map( A1 => n322, A2 => n955, A3 => IR_IN(3), ZN => n248
                           );
   U494 : NAND3_X1 port map( A1 => n308, A2 => n980, A3 => n289_port, ZN => 
                           n307);
   U495 : NAND3_X1 port map( A1 => IR_IN(30), A2 => n976, A3 => n320, ZN => 
                           n281_port);
   add_217 : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 
                           port map( A(31) => iterator_trap_31_port, A(30) => 
                           iterator_trap_30_port, A(29) => 
                           iterator_trap_29_port, A(28) => 
                           iterator_trap_28_port, A(27) => 
                           iterator_trap_27_port, A(26) => 
                           iterator_trap_26_port, A(25) => 
                           iterator_trap_25_port, A(24) => 
                           iterator_trap_24_port, A(23) => 
                           iterator_trap_23_port, A(22) => 
                           iterator_trap_22_port, A(21) => 
                           iterator_trap_21_port, A(20) => 
                           iterator_trap_20_port, A(19) => 
                           iterator_trap_19_port, A(18) => 
                           iterator_trap_18_port, A(17) => 
                           iterator_trap_17_port, A(16) => 
                           iterator_trap_16_port, A(15) => 
                           iterator_trap_15_port, A(14) => 
                           iterator_trap_14_port, A(13) => 
                           iterator_trap_13_port, A(12) => 
                           iterator_trap_12_port, A(11) => 
                           iterator_trap_11_port, A(10) => 
                           iterator_trap_10_port, A(9) => iterator_trap_9_port,
                           A(8) => iterator_trap_8_port, A(7) => 
                           iterator_trap_7_port, A(6) => iterator_trap_6_port, 
                           A(5) => iterator_trap_5_port, A(4) => 
                           iterator_trap_4_port, A(3) => iterator_trap_3_port, 
                           A(2) => iterator_trap_2_port, A(1) => 
                           iterator_trap_1_port, A(0) => iterator_trap_0_port, 
                           SUM(31) => N71, SUM(30) => N70, SUM(29) => N69, 
                           SUM(28) => N68, SUM(27) => N67, SUM(26) => N66, 
                           SUM(25) => N65, SUM(24) => N64, SUM(23) => N63, 
                           SUM(22) => N62, SUM(21) => N61, SUM(20) => N60, 
                           SUM(19) => N59, SUM(18) => N58, SUM(17) => N57, 
                           SUM(16) => N56, SUM(15) => N55, SUM(14) => N54, 
                           SUM(13) => N53, SUM(12) => N52, SUM(11) => N51, 
                           SUM(10) => N50, SUM(9) => N49, SUM(8) => N48, SUM(7)
                           => N47, SUM(6) => N46, SUM(5) => N45, SUM(4) => N44,
                           SUM(3) => N43, SUM(2) => N42, SUM(1) => N41, SUM(0) 
                           => N40);
   add_236 : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 
                           port map( A(31) => iterator_ret_31_port, A(30) => 
                           iterator_ret_30_port, A(29) => iterator_ret_29_port,
                           A(28) => iterator_ret_28_port, A(27) => 
                           iterator_ret_27_port, A(26) => iterator_ret_26_port,
                           A(25) => iterator_ret_25_port, A(24) => 
                           iterator_ret_24_port, A(23) => iterator_ret_23_port,
                           A(22) => iterator_ret_22_port, A(21) => 
                           iterator_ret_21_port, A(20) => iterator_ret_20_port,
                           A(19) => iterator_ret_19_port, A(18) => 
                           iterator_ret_18_port, A(17) => iterator_ret_17_port,
                           A(16) => iterator_ret_16_port, A(15) => 
                           iterator_ret_15_port, A(14) => iterator_ret_14_port,
                           A(13) => iterator_ret_13_port, A(12) => 
                           iterator_ret_12_port, A(11) => iterator_ret_11_port,
                           A(10) => iterator_ret_10_port, A(9) => 
                           iterator_ret_9_port, A(8) => iterator_ret_8_port, 
                           A(7) => iterator_ret_7_port, A(6) => 
                           iterator_ret_6_port, A(5) => iterator_ret_5_port, 
                           A(4) => iterator_ret_4_port, A(3) => 
                           iterator_ret_3_port, A(2) => iterator_ret_2_port, 
                           A(1) => iterator_ret_1_port, A(0) => 
                           iterator_ret_0_port, SUM(31) => N182, SUM(30) => 
                           N181, SUM(29) => N180, SUM(28) => N179, SUM(27) => 
                           N178, SUM(26) => N177, SUM(25) => N176, SUM(24) => 
                           N175, SUM(23) => N174, SUM(22) => N173, SUM(21) => 
                           N172, SUM(20) => N171, SUM(19) => N170, SUM(18) => 
                           N169, SUM(17) => N168, SUM(16) => N167, SUM(15) => 
                           N166, SUM(14) => N165, SUM(13) => N164, SUM(12) => 
                           N163, SUM(11) => N162, SUM(10) => N161, SUM(9) => 
                           N160, SUM(8) => N159, SUM(7) => N158, SUM(6) => N157
                           , SUM(5) => N156, SUM(4) => N155, SUM(3) => N154, 
                           SUM(2) => N153, SUM(1) => N152, SUM(0) => N151);
   add_277 : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_6 
                           port map( A(31) => iterator2_31_port, A(30) => 
                           iterator2_30_port, A(29) => iterator2_29_port, A(28)
                           => iterator2_28_port, A(27) => iterator2_27_port, 
                           A(26) => iterator2_26_port, A(25) => 
                           iterator2_25_port, A(24) => iterator2_24_port, A(23)
                           => iterator2_23_port, A(22) => iterator2_22_port, 
                           A(21) => iterator2_21_port, A(20) => 
                           iterator2_20_port, A(19) => iterator2_19_port, A(18)
                           => iterator2_18_port, A(17) => iterator2_17_port, 
                           A(16) => iterator2_16_port, A(15) => 
                           iterator2_15_port, A(14) => iterator2_14_port, A(13)
                           => iterator2_13_port, A(12) => iterator2_12_port, 
                           A(11) => iterator2_11_port, A(10) => 
                           iterator2_10_port, A(9) => iterator2_9_port, A(8) =>
                           iterator2_8_port, A(7) => iterator2_7_port, A(6) => 
                           iterator2_6_port, A(5) => iterator2_5_port, A(4) => 
                           iterator2_4_port, A(3) => iterator2_3_port, A(2) => 
                           iterator2_2_port, A(1) => iterator2_1_port, A(0) => 
                           iterator2_0_port, SUM(31) => N407, SUM(30) => N406, 
                           SUM(29) => N405, SUM(28) => N404, SUM(27) => N403, 
                           SUM(26) => N402, SUM(25) => N401, SUM(24) => N400, 
                           SUM(23) => N399, SUM(22) => N398, SUM(21) => N397, 
                           SUM(20) => N396, SUM(19) => N395, SUM(18) => N394, 
                           SUM(17) => N393, SUM(16) => N392, SUM(15) => N391, 
                           SUM(14) => N390, SUM(13) => N389, SUM(12) => N388, 
                           SUM(11) => N387, SUM(10) => N386, SUM(9) => N385, 
                           SUM(8) => N384, SUM(7) => N383, SUM(6) => N382, 
                           SUM(5) => N381, SUM(4) => N380, SUM(3) => N379, 
                           SUM(2) => N378, SUM(1) => N377, SUM(0) => N376);
   add_256 : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_7 
                           port map( A(31) => iterator1_31_port, A(30) => 
                           iterator1_30_port, A(29) => iterator1_29_port, A(28)
                           => iterator1_28_port, A(27) => iterator1_27_port, 
                           A(26) => iterator1_26_port, A(25) => 
                           iterator1_25_port, A(24) => iterator1_24_port, A(23)
                           => iterator1_23_port, A(22) => iterator1_22_port, 
                           A(21) => iterator1_21_port, A(20) => 
                           iterator1_20_port, A(19) => iterator1_19_port, A(18)
                           => iterator1_18_port, A(17) => iterator1_17_port, 
                           A(16) => iterator1_16_port, A(15) => 
                           iterator1_15_port, A(14) => iterator1_14_port, A(13)
                           => iterator1_13_port, A(12) => iterator1_12_port, 
                           A(11) => iterator1_11_port, A(10) => 
                           iterator1_10_port, A(9) => iterator1_9_port, A(8) =>
                           iterator1_8_port, A(7) => iterator1_7_port, A(6) => 
                           iterator1_6_port, A(5) => iterator1_5_port, A(4) => 
                           iterator1_4_port, A(3) => iterator1_3_port, A(2) => 
                           iterator1_2_port, A(1) => iterator1_1_port, A(0) => 
                           iterator1_0_port, SUM(31) => N294, SUM(30) => N293, 
                           SUM(29) => N292, SUM(28) => N291, SUM(27) => N290, 
                           SUM(26) => N289, SUM(25) => N288, SUM(24) => N287, 
                           SUM(23) => N286, SUM(22) => N285, SUM(21) => N284, 
                           SUM(20) => N283, SUM(19) => N282, SUM(18) => N281, 
                           SUM(17) => N280, SUM(16) => N279, SUM(15) => N278, 
                           SUM(14) => N277, SUM(13) => N276, SUM(12) => N275, 
                           SUM(11) => N274, SUM(10) => N273, SUM(9) => N272, 
                           SUM(8) => N271, SUM(7) => N270, SUM(6) => N269, 
                           SUM(5) => N268, SUM(4) => N267, SUM(3) => N266, 
                           SUM(2) => N265, SUM(1) => N264, SUM(0) => N263);
   aluOpcode3_reg_5_inst : DFFR_X1 port map( D => aluOpcode2_5_port, CK => Clk,
                           RN => Rst, Q => ALU_OPCODE(0), QN => n_3132);
   sig1_reg : DFF_X1 port map( D => n567, CK => Clk, Q => n_3133, QN => n941);
   sig2_reg : DFF_X1 port map( D => n566, CK => Clk, Q => n_3134, QN => n897);
   sig4_reg : DFF_X1 port map( D => n613, CK => Clk, Q => n_3135, QN => n860);
   lhi_sel_reg : DFF_X1 port map( D => n432, CK => Clk, Q => lhi_sel, QN => 
                           n773);
   U3 : AND2_X1 port map( A1 => n826, A2 => n759, ZN => n614);
   U4 : INV_X1 port map( A => n614, ZN => n615);
   U5 : INV_X1 port map( A => n708, ZN => n616);
   U6 : INV_X1 port map( A => n705, ZN => n617);
   U7 : AND3_X1 port map( A1 => n618, A2 => n619, A3 => n620, ZN => n904);
   U8 : AND4_X1 port map( A1 => n903, A2 => n912, A3 => n911, A4 => n913, ZN =>
                           n618);
   U9 : AND4_X1 port map( A1 => n921, A2 => n920, A3 => n919, A4 => n918, ZN =>
                           n619);
   U10 : AND4_X1 port map( A1 => n925, A2 => n924, A3 => n923, A4 => n922, ZN 
                           => n620);
   U11 : AND2_X1 port map( A1 => n635, A2 => n771, ZN => n621);
   U12 : BUF_X1 port map( A => n816, Z => n755);
   U13 : INV_X1 port map( A => N389, ZN => n797);
   U14 : BUF_X1 port map( A => n816, Z => n754);
   U15 : BUF_X1 port map( A => n816, Z => n753);
   U16 : BUF_X1 port map( A => n625, Z => n758);
   U17 : BUF_X1 port map( A => n625, Z => n756);
   U18 : BUF_X2 port map( A => n899, Z => n731);
   U19 : BUF_X1 port map( A => n942, Z => n771);
   U20 : INV_X1 port map( A => N50, ZN => n918);
   U21 : BUF_X1 port map( A => n942, Z => n770);
   U22 : INV_X1 port map( A => N60, ZN => n928);
   U23 : INV_X1 port map( A => n713, ZN => n622);
   U24 : INV_X1 port map( A => n715, ZN => n623);
   U25 : INV_X1 port map( A => n747, ZN => n624);
   U26 : AND2_X1 port map( A1 => n818, A2 => n774, ZN => n625);
   U27 : AND2_X1 port map( A1 => N41, A2 => n717_port, ZN => n626);
   U28 : AND3_X1 port map( A1 => N378, A2 => N377, A3 => N376, ZN => n627);
   U29 : BUF_X1 port map( A => n942, Z => n769);
   U30 : OR2_X1 port map( A1 => N164, A2 => N167, ZN => n628);
   U31 : AND2_X1 port map( A1 => n839, A2 => n841, ZN => n629);
   U32 : MUX2_X1 port map( A => n768, B => n900, S => n639, Z => n467);
   U33 : BUF_X1 port map( A => n631, Z => n636);
   U34 : AND2_X1 port map( A1 => n908, A2 => n771, ZN => n630);
   U35 : BUF_X1 port map( A => n647, Z => n631);
   U36 : CLKBUF_X1 port map( A => N172, Z => n632);
   U37 : INV_X1 port map( A => N182, ZN => n633);
   U38 : CLKBUF_X1 port map( A => N173, Z => n634);
   U39 : NAND2_X1 port map( A1 => n744, A2 => n626, ZN => n635);
   U40 : AND4_X2 port map( A1 => n905, A2 => n904, A3 => n907, A4 => n906, ZN 
                           => n744);
   U41 : NAND3_X1 port map( A1 => n842, A2 => n840, A3 => n629, ZN => n820);
   U42 : OR2_X1 port map( A1 => N277, A2 => N279, ZN => n637);
   U43 : OR2_X1 port map( A1 => N58, A2 => N60, ZN => n638);
   U44 : INV_X1 port map( A => n355, ZN => n639);
   U45 : CLKBUF_X1 port map( A => N175, Z => n640);
   U46 : AND4_X1 port map( A1 => n641, A2 => n876, A3 => n642, A4 => n643, ZN 
                           => n864);
   U47 : INV_X1 port map( A => N160, ZN => n641);
   U48 : INV_X1 port map( A => N162, ZN => n642);
   U49 : INV_X1 port map( A => N163, ZN => n643);
   U50 : OAI22_X1 port map( A1 => n660, A2 => n797, B1 => n754, B2 => n400_port
                           , ZN => n546);
   U51 : OAI22_X1 port map( A1 => n660, A2 => n809, B1 => n753, B2 => n412, ZN 
                           => n558);
   U52 : OAI22_X1 port map( A1 => n700, A2 => n928, B1 => n769, B2 => n343, ZN 
                           => n455);
   U53 : OAI22_X1 port map( A1 => n700, A2 => n918, B1 => n770, B2 => n333, ZN 
                           => n445);
   U54 : OAI22_X1 port map( A1 => n696, A2 => n857, B1 => n756, B2 => n577, ZN 
                           => n584);
   U55 : INV_X2 port map( A => N291, ZN => n857);
   U56 : OAI22_X1 port map( A1 => n671, A2 => n837, B1 => n758, B2 => n521, ZN 
                           => n604);
   U57 : OAI22_X1 port map( A1 => n719, A2 => n786, B1 => n755, B2 => n389_port
                           , ZN => n535);
   U58 : INV_X2 port map( A => N378, ZN => n786);
   U59 : OAI22_X1 port map( A1 => n695, A2 => n909, B1 => n771, B2 => n354, ZN 
                           => n466);
   U60 : CLKBUF_X1 port map( A => N285, Z => n644);
   U61 : AND2_X1 port map( A1 => n908, A2 => n771, ZN => n645);
   U62 : BUF_X1 port map( A => n631, Z => n727);
   U63 : CLKBUF_X1 port map( A => N277, Z => n646);
   U64 : OAI21_X1 port map( B1 => n895, B2 => n639, A => n763, ZN => n647);
   U65 : CLKBUF_X1 port map( A => n883, Z => n648);
   U66 : CLKBUF_X1 port map( A => N58, Z => n649);
   U67 : OR2_X1 port map( A1 => n783, A2 => n707, ZN => n650);
   U68 : NAND4_X1 port map( A1 => n884, A2 => n648, A3 => n882, A4 => n881, ZN 
                           => n651);
   U69 : OR2_X1 port map( A1 => n783, A2 => n707, ZN => n781);
   U70 : NOR2_X1 port map( A1 => n653, A2 => n654, ZN => n652);
   U71 : NAND4_X1 port map( A1 => n673, A2 => n800, A3 => n799, A4 => n798, ZN 
                           => n653);
   U72 : OR4_X2 port map( A1 => n777, A2 => N385, A3 => N384, A4 => N383, ZN =>
                           n654);
   U73 : AND4_X1 port map( A1 => n794, A2 => n795, A3 => n796, A4 => n797, ZN 
                           => n673);
   U74 : NOR3_X1 port map( A1 => N166, A2 => N165, A3 => n628, ZN => n865);
   U75 : NOR3_X1 port map( A1 => n820, A2 => N278, A3 => n637, ZN => n824);
   U76 : INV_X1 port map( A => n658, ZN => n655);
   U77 : CLKBUF_X1 port map( A => N284, Z => n656);
   U78 : CLKBUF_X1 port map( A => N177, Z => n657);
   U79 : AND2_X1 port map( A1 => n781, A2 => n755, ZN => n658);
   U80 : AND2_X1 port map( A1 => n650, A2 => n755, ZN => n749);
   U81 : BUF_X1 port map( A => n631, Z => n728);
   U82 : CLKBUF_X1 port map( A => n744, Z => n659);
   U83 : NOR2_X1 port map( A1 => N292, A2 => N291, ZN => n720);
   U84 : INV_X1 port map( A => n704, ZN => n660);
   U85 : INV_X1 port map( A => n704, ZN => n718_port);
   U86 : CLKBUF_X1 port map( A => n690, Z => n661);
   U87 : INV_X1 port map( A => n706, ZN => n662);
   U88 : OR2_X1 port map( A1 => n763, A2 => n897, ZN => n663);
   U89 : NAND2_X1 port map( A1 => n663, A2 => n636, ZN => n566);
   U90 : INV_X1 port map( A => n768, ZN => n767);
   U91 : BUF_X1 port map( A => n899, Z => n664);
   U92 : AND3_X1 port map( A1 => n742, A2 => n859, A3 => n720, ZN => n665);
   U93 : CLKBUF_X1 port map( A => N397, Z => n666);
   U94 : OR2_X1 port map( A1 => N285, A2 => N284, ZN => n667);
   U95 : NAND2_X1 port map( A1 => n744, A2 => n626, ZN => n908);
   U96 : AND2_X1 port map( A1 => n864, A2 => n863, ZN => n668);
   U97 : AND2_X1 port map( A1 => n865, A2 => n668, ZN => n680);
   U98 : CLKBUF_X1 port map( A => n665, Z => n669);
   U99 : AND4_X1 port map( A1 => n867, A2 => N153, A3 => n894, A4 => n893, ZN 
                           => n670);
   U100 : AND4_X1 port map( A1 => n894, A2 => n633, A3 => N153, A4 => n893, ZN 
                           => n739);
   U101 : NOR3_X1 port map( A1 => n902, A2 => N59, A3 => n638, ZN => n905);
   U102 : INV_X1 port map( A => n614, ZN => n671);
   U103 : NOR2_X1 port map( A1 => N393, A2 => N396, ZN => n672);
   U104 : INV_X1 port map( A => n749, ZN => n674);
   U105 : INV_X1 port map( A => n658, ZN => n675);
   U106 : INV_X1 port map( A => n748, ZN => n676);
   U107 : CLKBUF_X1 port map( A => N398, Z => n677);
   U108 : NOR3_X1 port map( A1 => N173, A2 => N175, A3 => N172, ZN => n698);
   U109 : CLKBUF_X1 port map( A => n686, Z => n678);
   U110 : CLKBUF_X1 port map( A => N399, Z => n679);
   U111 : NAND3_X1 port map( A1 => n803, A2 => n802, A3 => n672, ZN => n778);
   U112 : NOR2_X1 port map( A1 => n661, A2 => n651, ZN => n681);
   U113 : OR2_X1 port map( A1 => n774, A2 => n773, ZN => n682);
   U114 : NAND2_X1 port map( A1 => n829, A2 => n682, ZN => n432);
   U115 : CLKBUF_X1 port map( A => n783, Z => n683);
   U116 : AND2_X1 port map( A1 => n684, A2 => n685, ZN => n779);
   U117 : AND4_X1 port map( A1 => n808, A2 => n809, A3 => n810, A4 => n811, ZN 
                           => n684);
   U118 : NOR3_X1 port map( A1 => N405, A2 => N406, A3 => N404, ZN => n685);
   U119 : AND3_X1 port map( A1 => n823, A2 => n825, A3 => n824, ZN => n686);
   U120 : INV_X1 port map( A => n748, ZN => n687);
   U121 : INV_X1 port map( A => n658, ZN => n688);
   U122 : NOR3_X1 port map( A1 => n667, A2 => N286, A3 => n821, ZN => n823);
   U123 : NOR4_X1 port map( A1 => N176, A2 => N177, A3 => N178, A4 => N179, ZN 
                           => n693);
   U124 : AND2_X1 port map( A1 => n686, A2 => n665, ZN => n689);
   U125 : NOR2_X1 port map( A1 => n690, A2 => n691, ZN => n722);
   U126 : NAND2_X1 port map( A1 => n698, A2 => n887, ZN => n690);
   U127 : NAND4_X1 port map( A1 => n884, A2 => n883, A3 => n882, A4 => n881, ZN
                           => n691);
   U128 : CLKBUF_X1 port map( A => n887, Z => n692);
   U129 : AND4_X1 port map( A1 => n891, A2 => n892, A3 => n890, A4 => n889, ZN 
                           => n738);
   U130 : INV_X1 port map( A => n747, ZN => n694);
   U131 : INV_X1 port map( A => n706, ZN => n695);
   U132 : INV_X1 port map( A => n715, ZN => n696);
   U133 : CLKBUF_X1 port map( A => N286, Z => n697);
   U134 : NAND2_X1 port map( A1 => n689, A2 => n711, ZN => n699);
   U135 : INV_X1 port map( A => n645, ZN => n700);
   U136 : NOR4_X1 port map( A1 => n778, A2 => N397, A3 => N398, A4 => N399, ZN 
                           => n780);
   U137 : AND3_X1 port map( A1 => n722, A2 => n739, A3 => n693, ZN => n701);
   U138 : INV_X1 port map( A => n714, ZN => n702);
   U139 : OR2_X1 port map( A1 => n769, A2 => n941, ZN => n703);
   U140 : NAND2_X1 port map( A1 => n734, A2 => n703, ZN => n567);
   U141 : AND2_X1 port map( A1 => n755, A2 => n650, ZN => n704);
   U142 : NAND3_X1 port map( A1 => n779, A2 => n652, A3 => n780, ZN => n783);
   U143 : AND2_X1 port map( A1 => n635, A2 => n771, ZN => n705);
   U144 : AND2_X1 port map( A1 => n908, A2 => n771, ZN => n706);
   U145 : AND2_X1 port map( A1 => n635, A2 => n771, ZN => n708);
   U146 : NAND2_X1 port map( A1 => n782, A2 => n627, ZN => n707);
   U147 : AND2_X1 port map( A1 => n862, A2 => n680, ZN => n709);
   U148 : NAND2_X1 port map( A1 => n710, A2 => n711, ZN => n826);
   U149 : AND2_X1 port map( A1 => n686, A2 => n822, ZN => n710);
   U150 : NOR2_X1 port map( A1 => n723, A2 => N294, ZN => n711);
   U151 : CLKBUF_X1 port map( A => N406, Z => n712);
   U152 : AND2_X1 port map( A1 => n699, A2 => n759, ZN => n713);
   U153 : AND2_X1 port map( A1 => n699, A2 => n759, ZN => n714);
   U154 : AND2_X1 port map( A1 => n826, A2 => n759, ZN => n715);
   U155 : INV_X1 port map( A => n713, ZN => n716);
   U156 : INV_X1 port map( A => n323, ZN => n717_port);
   U157 : INV_X1 port map( A => n704, ZN => n719);
   U158 : INV_X1 port map( A => n749, ZN => n750);
   U159 : INV_X1 port map( A => n749, ZN => n751);
   U160 : AND3_X1 port map( A1 => n742, A2 => n859, A3 => n720, ZN => n822);
   U161 : OR2_X1 port map( A1 => n756, A2 => n860, ZN => n721);
   U162 : NAND2_X1 port map( A1 => n721, A2 => n741, ZN => n613);
   U163 : AND3_X1 port map( A1 => n670, A2 => n738, A3 => n681, ZN => n862);
   U164 : NAND3_X1 port map( A1 => N265, A2 => N264, A3 => N263, ZN => n723);
   U165 : NAND2_X1 port map( A1 => n669, A2 => n678, ZN => n828);
   U166 : NAND2_X1 port map( A1 => n701, A2 => n680, ZN => n895);
   U167 : INV_X1 port map( A => n708, ZN => n724);
   U168 : INV_X1 port map( A => n630, ZN => n725);
   U169 : BUF_X1 port map( A => n898, Z => n763);
   U170 : BUF_X1 port map( A => n898, Z => n765);
   U171 : BUF_X1 port map( A => n898, Z => n764);
   U172 : OAI22_X1 port map( A1 => n962, A2 => n974, B1 => n968, B2 => n255, ZN
                           => n296);
   U173 : INV_X1 port map( A => n255, ZN => n973);
   U174 : NAND2_X1 port map( A1 => n968, A2 => n966, ZN => n184);
   U175 : INV_X1 port map( A => n303, ZN => n975);
   U176 : NAND2_X1 port map( A1 => n962, A2 => n968, ZN => n283_port);
   U177 : INV_X1 port map( A => n275_port, ZN => n962);
   U178 : NAND4_X1 port map( A1 => n963, A2 => n965, A3 => n945, A4 => n183, ZN
                           => n565);
   U179 : NAND2_X1 port map( A1 => n977, A2 => n184, ZN => n183);
   U180 : AND3_X1 port map( A1 => n965, A2 => n262, A3 => n251, ZN => n263_port
                           );
   U181 : INV_X1 port map( A => n309, ZN => n963);
   U182 : INV_X1 port map( A => n258, ZN => n948);
   U183 : INV_X1 port map( A => n271_port, ZN => n969);
   U184 : BUF_X1 port map( A => n625, Z => n757);
   U185 : AND2_X1 port map( A1 => n854, A2 => n853, ZN => n726);
   U186 : AOI211_X1 port map( C1 => n283_port, C2 => n972, A => n960, B => n423
                           , ZN => n241);
   U187 : INV_X1 port map( A => n304, ZN => n960);
   U188 : INV_X1 port map( A => n281_port, ZN => n972);
   U189 : OAI21_X1 port map( B1 => n291_port, B2 => n968, A => n239, ZN => n423
                           );
   U190 : NOR2_X1 port map( A1 => n279_port, A2 => n257, ZN => n267_port);
   U191 : INV_X1 port map( A => n775, ZN => n774);
   U192 : NOR2_X1 port map( A1 => n291_port, A2 => n218, ZN => n280_port);
   U193 : OAI21_X1 port map( B1 => n248, B2 => n302, A => n284_port, ZN => n258
                           );
   U194 : NAND2_X1 port map( A1 => n245, A2 => n435, ZN => n262);
   U195 : OAI22_X1 port map( A1 => n267_port, A2 => n248, B1 => n954, B2 => 
                           n247, ZN => n435);
   U196 : INV_X1 port map( A => n245, ZN => n959);
   U197 : AOI21_X1 port map( B1 => n289_port, B2 => n978, A => n427, ZN => n251
                           );
   U198 : INV_X1 port map( A => n280_port, ZN => n971);
   U199 : AOI22_X1 port map( A1 => n278_port, A2 => n279_port, B1 => n961, B2 
                           => n975, ZN => n277_port);
   U200 : NOR2_X1 port map( A1 => n959, A2 => n259, ZN => n278_port);
   U201 : AOI221_X1 port map( B1 => n951, B2 => n298, C1 => n257, C2 => n299, A
                           => n300, ZN => n297);
   U202 : INV_X1 port map( A => n247, ZN => n951);
   U203 : NOR4_X1 port map( A1 => n301, A2 => n958, A3 => n957, A4 => n302, ZN 
                           => n300);
   U204 : AOI211_X1 port map( C1 => n978, C2 => n266_port, A => n280_port, B =>
                           n315, ZN => n314);
   U205 : AOI21_X1 port map( B1 => n254, B2 => n968, A => n974, ZN => n315);
   U206 : NOR2_X1 port map( A1 => n292_port, A2 => n964, ZN => n427);
   U207 : INV_X1 port map( A => n184, ZN => n964);
   U208 : AOI21_X1 port map( B1 => n970, B2 => n975, A => n288_port, ZN => n242
                           );
   U209 : INV_X1 port map( A => n217, ZN => n978);
   U210 : NAND4_X1 port map( A1 => n241, A2 => n945, A3 => n251, A4 => n949, ZN
                           => aluOpcode_i_3_port);
   U211 : INV_X1 port map( A => n252, ZN => n949);
   U212 : OAI221_X1 port map( B1 => n959, B2 => n253, C1 => n254, C2 => n255, A
                           => n256, ZN => n252);
   U213 : AOI21_X1 port map( B1 => n257, B2 => n956, A => n258, ZN => n253);
   U214 : OAI21_X1 port map( B1 => n966, B2 => n292_port, A => n293_port, ZN =>
                           n287_port);
   U215 : INV_X1 port map( A => n218, ZN => n970);
   U216 : INV_X1 port map( A => n254, ZN => n961);
   U217 : AOI222_X1 port map( A1 => n244, A2 => n970, B1 => n245, B2 => n246, 
                           C1 => n977, C2 => n184, ZN => n243);
   U218 : OAI211_X1 port map( C1 => n247, C2 => n248, A => n249, B => n250, ZN 
                           => n246);
   U219 : NAND4_X1 port map( A1 => n263_port, A2 => n241, A3 => n310, A4 => 
                           n311, ZN => N717);
   U220 : AOI21_X1 port map( B1 => n245, B2 => n313, A => n309, ZN => n310);
   U221 : NOR4_X1 port map( A1 => n978, A2 => n244, A3 => n973, A4 => n312, ZN 
                           => n311);
   U222 : NAND4_X1 port map( A1 => n946, A2 => n948, A3 => n268_port, A4 => 
                           n248, ZN => n313);
   U223 : NAND2_X1 port map( A1 => n254, A2 => n966, ZN => n266_port);
   U224 : INV_X1 port map( A => n200, ZN => n977);
   U225 : NAND2_X1 port map( A1 => n944, A2 => n979, ZN => n291_port);
   U226 : NAND4_X1 port map( A1 => n271_port, A2 => n272_port, A3 => n273_port,
                           A4 => n274_port, ZN => aluOpcode_i_1_port);
   U227 : AOI22_X1 port map( A1 => n245, A2 => n282_port, B1 => n244, B2 => 
                           n283_port, ZN => n273_port);
   U228 : AOI211_X1 port map( C1 => n973, C2 => n275_port, A => n276_port, B =>
                           n270_port, ZN => n274_port);
   U229 : OAI211_X1 port map( C1 => n267_port, C2 => n248, A => n284_port, B =>
                           n947, ZN => n282_port);
   U230 : OR2_X1 port map( A1 => n259, A2 => n302, ZN => n269_port);
   U231 : INV_X1 port map( A => n259, ZN => n956);
   U232 : NAND2_X1 port map( A1 => n254, A2 => n218, ZN => n275_port);
   U233 : NAND2_X1 port map( A1 => n289_port, A2 => n290_port, ZN => n271_port)
                           ;
   U234 : INV_X1 port map( A => n298, ZN => n954);
   U236 : INV_X1 port map( A => n419, ZN => n946);
   U237 : OAI211_X1 port map( C1 => n267_port, C2 => n259, A => n250, B => n947
                           , ZN => n419);
   U238 : INV_X1 port map( A => n260, ZN => n945);
   U239 : OAI21_X1 port map( B1 => n261, B2 => n959, A => n262, ZN => n260);
   U240 : INV_X1 port map( A => n420, ZN => n947);
   U241 : OAI221_X1 port map( B1 => n268_port, B2 => n302, C1 => n267_port, C2 
                           => n954, A => n421, ZN => n420);
   U242 : AND2_X1 port map( A1 => n269_port, A2 => n249, ZN => n421);
   U243 : INV_X1 port map( A => n270_port, ZN => n950);
   U244 : AOI222_X1 port map( A1 => n244, A2 => n970, B1 => n245, B2 => 
                           n265_port, C1 => n973, C2 => n266_port, ZN => 
                           n264_port);
   U245 : OAI21_X1 port map( B1 => n267_port, B2 => n268_port, A => n269_port, 
                           ZN => n265_port);
   U246 : INV_X1 port map( A => n500, ZN => n965);
   U247 : OAI211_X1 port map( C1 => n966, C2 => n281_port, A => n293_port, B =>
                           n272_port, ZN => n500);
   U248 : AOI221_X1 port map( B1 => n978, B2 => n289_port, C1 => n961, C2 => 
                           n977, A => n306, ZN => n305);
   U249 : AOI21_X1 port map( B1 => n946, B2 => n261, A => n307, ZN => n306);
   U250 : INV_X1 port map( A => n244, ZN => n974);
   U251 : NAND2_X1 port map( A1 => n317, A2 => n976, ZN => n303);
   U252 : NAND2_X1 port map( A1 => n285_port, A2 => n286_port, ZN => 
                           aluOpcode_i_0_port);
   U253 : AOI221_X1 port map( B1 => n961, B2 => n294_port, C1 => n245, C2 => 
                           n295, A => n296, ZN => n285_port);
   U254 : NOR4_X1 port map( A1 => n287_port, A2 => n969, A3 => n288_port, A4 =>
                           n280_port, ZN => n286_port);
   U255 : NAND4_X1 port map( A1 => n261, A2 => n250, A3 => n269_port, A4 => 
                           n297, ZN => n295);
   U256 : AOI22_X1 port map( A1 => n316, A2 => n973, B1 => n318, B2 => n970, ZN
                           => n256);
   U257 : OAI21_X1 port map( B1 => n979, B2 => n319, A => n255, ZN => n318);
   U258 : OAI22_X1 port map( A1 => n218, A2 => n281_port, B1 => n966, B2 => 
                           n200, ZN => n276_port);
   U259 : OAI22_X1 port map( A1 => n505, A2 => n775, B1 => Rst, B2 => n506, ZN 
                           => n428);
   U260 : OAI22_X1 port map( A1 => n504, A2 => n775, B1 => n505, B2 => Rst, ZN 
                           => n429);
   U261 : OAI21_X1 port map( B1 => n504, B2 => Rst, A => n240, ZN => n430);
   U262 : NAND2_X1 port map( A1 => signed_unsigned_i, A2 => Rst, ZN => n240);
   U263 : OR3_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), ZN 
                           => n499);
   U264 : OAI211_X1 port map( C1 => n279_port, C2 => n321, A => n322, B => 
                           IR_IN(3), ZN => n284_port);
   U265 : NOR2_X1 port map( A1 => n955, A2 => n302, ZN => n321);
   U266 : NOR3_X1 port map( A1 => n962, A2 => IR_IN(31), A3 => IR_IN(28), ZN =>
                           n312);
   U267 : NAND4_X1 port map( A1 => n257, A2 => n301, A3 => IR_IN(3), A4 => 
                           IR_IN(5), ZN => n250);
   U268 : NAND4_X1 port map( A1 => IR_IN(28), A2 => n320, A3 => n289_port, A4 
                           => IR_IN(30), ZN => n293_port);
   U269 : NAND4_X1 port map( A1 => IR_IN(28), A2 => n320, A3 => n316, A4 => 
                           IR_IN(30), ZN => n272_port);
   U270 : NAND2_X1 port map( A1 => IR_IN(30), A2 => n308, ZN => n200);
   U271 : NAND4_X1 port map( A1 => IR_IN(4), A2 => IR_IN(3), A3 => n422, A4 => 
                           IR_IN(5), ZN => n249);
   U272 : AOI22_X1 port map( A1 => IR_IN(2), A2 => n302, B1 => n247, B2 => n955
                           , ZN => n422);
   U273 : INV_X1 port map( A => Rst, ZN => n775);
   U274 : NAND2_X1 port map( A1 => IR_IN(0), A2 => n953, ZN => n261);
   U275 : INV_X1 port map( A => n268_port, ZN => n953);
   U276 : AND3_X1 port map( A1 => IR_IN(28), A2 => n316, A3 => n317, ZN => 
                           n288_port);
   U278 : NOR2_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), ZN => n289_port);
   U279 : NAND2_X1 port map( A1 => IR_IN(0), A2 => n952, ZN => n302);
   U280 : INV_X1 port map( A => IR_IN(2), ZN => n955);
   U281 : NAND2_X1 port map( A1 => IR_IN(27), A2 => n967, ZN => n254);
   U282 : NAND2_X1 port map( A1 => IR_IN(27), A2 => IR_IN(26), ZN => n218);
   U283 : INV_X1 port map( A => IR_IN(30), ZN => n980);
   U284 : NAND2_X1 port map( A1 => IR_IN(1), A2 => IR_IN(0), ZN => n247);
   U285 : NOR2_X1 port map( A1 => n952, A2 => IR_IN(0), ZN => n257);
   U286 : INV_X1 port map( A => IR_IN(28), ZN => n976);
   U287 : NOR2_X1 port map( A1 => n979, A2 => IR_IN(31), ZN => n320);
   U288 : INV_X1 port map( A => IR_IN(29), ZN => n979);
   U289 : NOR2_X1 port map( A1 => n967, A2 => IR_IN(27), ZN => n316);
   U290 : NOR2_X1 port map( A1 => IR_IN(1), A2 => IR_IN(0), ZN => n279_port);
   U291 : NOR2_X1 port map( A1 => n958, A2 => IR_IN(4), ZN => n322);
   U292 : INV_X1 port map( A => IR_IN(3), ZN => n957);
   U293 : INV_X1 port map( A => IR_IN(26), ZN => n967);
   U294 : INV_X1 port map( A => IR_IN(1), ZN => n952);
   U295 : INV_X1 port map( A => IR_IN(5), ZN => n958);
   U296 : AND2_X1 port map( A1 => IR_IN(4), A2 => n955, ZN => n301);
   U297 : NOR4_X1 port map( A1 => n955, A2 => IR_IN(3), A3 => IR_IN(4), A4 => 
                           IR_IN(5), ZN => n298);
   U298 : NOR3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(31), A3 => IR_IN(28), 
                           ZN => n308);
   U299 : AOI22_X1 port map( A1 => n975, A2 => n961, B1 => IR_IN(31), B2 => 
                           n427, ZN => n304);
   U300 : AND3_X1 port map( A1 => IR_IN(31), A2 => IR_IN(30), A3 => IR_IN(29), 
                           ZN => n317);
   U301 : BUF_X1 port map( A => n899, Z => n729);
   U302 : BUF_X1 port map( A => n899, Z => n730);
   U303 : INV_X1 port map( A => n630, ZN => n732);
   U304 : INV_X1 port map( A => n708, ZN => n733);
   U305 : INV_X1 port map( A => n645, ZN => n734);
   U306 : INV_X1 port map( A => n705, ZN => n735);
   U307 : INV_X1 port map( A => n705, ZN => n736);
   U308 : INV_X1 port map( A => n621, ZN => n737);
   U309 : AND4_X1 port map( A1 => n937, A2 => n938, A3 => n909, A4 => N42, ZN 
                           => n907);
   U310 : INV_X1 port map( A => n714, ZN => n740);
   U311 : INV_X1 port map( A => n715, ZN => n741);
   U312 : INV_X1 port map( A => n614, ZN => n743);
   U313 : INV_X1 port map( A => n745, ZN => n760);
   U314 : INV_X1 port map( A => n713, ZN => n761);
   U315 : INV_X1 port map( A => n745, ZN => n762);
   U316 : AND2_X1 port map( A1 => n826, A2 => n759, ZN => n747);
   U317 : AND4_X1 port map( A1 => n933, A2 => n934, A3 => n935, A4 => n936, ZN 
                           => n906);
   U318 : AND3_X1 port map( A1 => n856, A2 => n855, A3 => n726, ZN => n742);
   U319 : AND2_X1 port map( A1 => n826, A2 => n759, ZN => n745);
   U320 : INV_X1 port map( A => n513, ZN => n746);
   U321 : INV_X1 port map( A => n658, ZN => n752);
   U322 : AND2_X1 port map( A1 => n781, A2 => n755, ZN => n748);
   U323 : INV_X1 port map( A => n647, ZN => n768);
   U324 : CLKBUF_X1 port map( A => n625, Z => n759);
   U325 : CLKBUF_X1 port map( A => n898, Z => n766);
   U326 : INV_X1 port map( A => n319, ZN => n944);
   U327 : NAND3_X1 port map( A1 => IR_IN(29), A2 => n289_port, A3 => n944, ZN 
                           => n239);
   U328 : INV_X1 port map( A => n316, ZN => n966);
   U329 : INV_X1 port map( A => n289_port, ZN => n968);
   U330 : INV_X1 port map( A => n239, ZN => n776);
   U331 : OAI21_X1 port map( B1 => n503, B2 => n776, A => n774, ZN => n817);
   U332 : INV_X1 port map( A => n817, ZN => n816);
   U333 : INV_X1 port map( A => N379, ZN => n787);
   U334 : INV_X1 port map( A => N380, ZN => n788);
   U335 : INV_X1 port map( A => N381, ZN => n789);
   U336 : INV_X1 port map( A => N382, ZN => n790);
   U337 : NAND4_X1 port map( A1 => n787, A2 => n788, A3 => n789, A4 => n790, ZN
                           => n777);
   U338 : INV_X1 port map( A => N386, ZN => n794);
   U339 : INV_X1 port map( A => N387, ZN => n795);
   U340 : INV_X1 port map( A => N388, ZN => n796);
   U341 : INV_X1 port map( A => N393, ZN => n801);
   U342 : INV_X1 port map( A => N394, ZN => n802);
   U343 : INV_X1 port map( A => N395, ZN => n803);
   U344 : INV_X1 port map( A => N396, ZN => n804);
   U345 : INV_X1 port map( A => N400, ZN => n808);
   U346 : INV_X1 port map( A => N401, ZN => n809);
   U347 : INV_X1 port map( A => N402, ZN => n810);
   U348 : INV_X1 port map( A => N403, ZN => n811);
   U349 : INV_X1 port map( A => N407, ZN => n782);
   U350 : OAI22_X1 port map( A1 => n676, A2 => n782, B1 => n418, B2 => n755, ZN
                           => n564);
   U351 : OAI211_X1 port map( C1 => N378, C2 => n683, A => n748, B => n782, ZN 
                           => n784);
   U352 : OAI21_X1 port map( B1 => n426, B2 => n774, A => n784, ZN => n431);
   U353 : INV_X1 port map( A => N377, ZN => n785);
   U354 : OAI22_X1 port map( A1 => n785, A2 => n750, B1 => n388_port, B2 => 
                           n755, ZN => n534);
   U355 : OAI22_X1 port map( A1 => n750, A2 => n787, B1 => n390_port, B2 => 
                           n755, ZN => n536);
   U356 : OAI22_X1 port map( A1 => n660, A2 => n788, B1 => n391_port, B2 => 
                           n755, ZN => n537);
   U357 : OAI22_X1 port map( A1 => n687, A2 => n789, B1 => n392_port, B2 => 
                           n755, ZN => n538);
   U358 : OAI22_X1 port map( A1 => n687, A2 => n790, B1 => n393_port, B2 => 
                           n755, ZN => n539);
   U359 : INV_X1 port map( A => N383, ZN => n791);
   U360 : OAI22_X1 port map( A1 => n718_port, A2 => n791, B1 => n394_port, B2 
                           => n755, ZN => n540);
   U361 : INV_X1 port map( A => N384, ZN => n792);
   U362 : OAI22_X1 port map( A1 => n688, A2 => n792, B1 => n395_port, B2 => 
                           n755, ZN => n541);
   U363 : INV_X1 port map( A => N385, ZN => n793);
   U364 : OAI22_X1 port map( A1 => n751, A2 => n793, B1 => n396_port, B2 => 
                           n755, ZN => n542);
   U365 : OAI22_X1 port map( A1 => n687, A2 => n794, B1 => n397_port, B2 => 
                           n754, ZN => n543);
   U366 : OAI22_X1 port map( A1 => n676, A2 => n795, B1 => n398_port, B2 => 
                           n754, ZN => n544);
   U367 : OAI22_X1 port map( A1 => n688, A2 => n796, B1 => n399_port, B2 => 
                           n754, ZN => n545);
   U368 : INV_X1 port map( A => N390, ZN => n798);
   U369 : OAI22_X1 port map( A1 => n655, A2 => n798, B1 => n401_port, B2 => 
                           n754, ZN => n547);
   U370 : INV_X1 port map( A => N391, ZN => n799);
   U371 : OAI22_X1 port map( A1 => n751, A2 => n799, B1 => n402_port, B2 => 
                           n754, ZN => n548);
   U372 : INV_X1 port map( A => N392, ZN => n800);
   U373 : OAI22_X1 port map( A1 => n719, A2 => n800, B1 => n403_port, B2 => 
                           n754, ZN => n549);
   U374 : OAI22_X1 port map( A1 => n752, A2 => n801, B1 => n404_port, B2 => 
                           n754, ZN => n550);
   U375 : OAI22_X1 port map( A1 => n718_port, A2 => n802, B1 => n405_port, B2 
                           => n754, ZN => n551);
   U376 : OAI22_X1 port map( A1 => n750, A2 => n803, B1 => n406_port, B2 => 
                           n754, ZN => n552);
   U377 : OAI22_X1 port map( A1 => n655, A2 => n804, B1 => n407_port, B2 => 
                           n754, ZN => n553);
   U378 : INV_X1 port map( A => n666, ZN => n805);
   U379 : OAI22_X1 port map( A1 => n675, A2 => n805, B1 => n408, B2 => n753, ZN
                           => n554);
   U380 : INV_X1 port map( A => n677, ZN => n806);
   U381 : OAI22_X1 port map( A1 => n806, A2 => n674, B1 => n409, B2 => n753, ZN
                           => n555);
   U382 : INV_X1 port map( A => n679, ZN => n807);
   U383 : OAI22_X1 port map( A1 => n752, A2 => n807, B1 => n410, B2 => n753, ZN
                           => n556);
   U384 : OAI22_X1 port map( A1 => n751, A2 => n808, B1 => n411, B2 => n753, ZN
                           => n557);
   U385 : OAI22_X1 port map( A1 => n675, A2 => n810, B1 => n413, B2 => n753, ZN
                           => n559);
   U386 : OAI22_X1 port map( A1 => n718_port, A2 => n811, B1 => n414, B2 => 
                           n753, ZN => n560);
   U387 : INV_X1 port map( A => N404, ZN => n812);
   U388 : OAI22_X1 port map( A1 => n812, A2 => n674, B1 => n415, B2 => n753, ZN
                           => n561);
   U389 : INV_X1 port map( A => N405, ZN => n813);
   U390 : OAI22_X1 port map( A1 => n676, A2 => n813, B1 => n416, B2 => n753, ZN
                           => n562);
   U391 : INV_X1 port map( A => n712, ZN => n814);
   U392 : OAI22_X1 port map( A1 => n719, A2 => n814, B1 => n417, B2 => n753, ZN
                           => n563);
   U393 : INV_X1 port map( A => n503, ZN => n815);
   U394 : OAI21_X1 port map( B1 => n753, B2 => n815, A => n674, ZN => n532);
   U395 : MUX2_X1 port map( A => n817, B => n658, S => n387_port, Z => n509);
   U396 : OAI21_X1 port map( B1 => n218, B2 => n217, A => n860, ZN => n818);
   U397 : INV_X1 port map( A => N266, ZN => n832);
   U398 : INV_X1 port map( A => N267, ZN => n833);
   U399 : INV_X1 port map( A => N268, ZN => n834);
   U400 : INV_X1 port map( A => N269, ZN => n835);
   U401 : NAND4_X1 port map( A1 => n832, A2 => n833, A3 => n834, A4 => n835, ZN
                           => n819);
   U402 : NOR4_X1 port map( A1 => n819, A2 => N272, A3 => N271, A4 => N270, ZN 
                           => n825);
   U403 : INV_X1 port map( A => N273, ZN => n839);
   U404 : INV_X1 port map( A => N274, ZN => n840);
   U405 : INV_X1 port map( A => N275, ZN => n841);
   U406 : INV_X1 port map( A => N276, ZN => n842);
   U407 : INV_X1 port map( A => N280, ZN => n846);
   U408 : INV_X1 port map( A => N281, ZN => n847);
   U409 : INV_X1 port map( A => N282, ZN => n848);
   U410 : INV_X1 port map( A => N283, ZN => n849);
   U411 : NAND4_X1 port map( A1 => n849, A2 => n847, A3 => n848, A4 => n846, ZN
                           => n821);
   U412 : INV_X1 port map( A => N287, ZN => n853);
   U413 : INV_X1 port map( A => N288, ZN => n854);
   U414 : INV_X1 port map( A => N289, ZN => n855);
   U415 : INV_X1 port map( A => N290, ZN => n856);
   U416 : INV_X1 port map( A => N294, ZN => n827);
   U417 : OAI22_X1 port map( A1 => n622, A2 => n827, B1 => n580, B2 => n758, ZN
                           => n581);
   U418 : OAI211_X1 port map( C1 => N265, C2 => n828, A => n747, B => n827, ZN 
                           => n829);
   U419 : INV_X1 port map( A => N264, ZN => n830);
   U420 : OAI22_X1 port map( A1 => n830, A2 => n760, B1 => n514, B2 => n758, ZN
                           => n611);
   U421 : INV_X1 port map( A => N265, ZN => n831);
   U422 : OAI22_X1 port map( A1 => n831, A2 => n761, B1 => n515, B2 => n758, ZN
                           => n610);
   U423 : OAI22_X1 port map( A1 => n623, A2 => n832, B1 => n516, B2 => n758, ZN
                           => n609);
   U424 : OAI22_X1 port map( A1 => n694, A2 => n833, B1 => n517, B2 => n758, ZN
                           => n608);
   U425 : OAI22_X1 port map( A1 => n743, A2 => n834, B1 => n518, B2 => n758, ZN
                           => n607);
   U426 : OAI22_X1 port map( A1 => n716, A2 => n835, B1 => n519, B2 => n758, ZN
                           => n606);
   U427 : INV_X1 port map( A => N270, ZN => n836);
   U428 : OAI22_X1 port map( A1 => n624, A2 => n836, B1 => n520, B2 => n758, ZN
                           => n605);
   U429 : INV_X1 port map( A => N271, ZN => n837);
   U430 : INV_X1 port map( A => N272, ZN => n838);
   U431 : OAI22_X1 port map( A1 => n762, A2 => n838, B1 => n522, B2 => n758, ZN
                           => n603);
   U432 : OAI22_X1 port map( A1 => n694, A2 => n839, B1 => n523, B2 => n758, ZN
                           => n602);
   U433 : OAI22_X1 port map( A1 => n702, A2 => n840, B1 => n524, B2 => n757, ZN
                           => n601);
   U434 : OAI22_X1 port map( A1 => n702, A2 => n841, B1 => n525, B2 => n757, ZN
                           => n600);
   U435 : OAI22_X1 port map( A1 => n696, A2 => n842, B1 => n526, B2 => n757, ZN
                           => n599);
   U436 : INV_X1 port map( A => n646, ZN => n843);
   U437 : OAI22_X1 port map( A1 => n716, A2 => n843, B1 => n527, B2 => n757, ZN
                           => n598);
   U438 : INV_X1 port map( A => N278, ZN => n844);
   U439 : OAI22_X1 port map( A1 => n761, A2 => n844, B1 => n528, B2 => n757, ZN
                           => n597);
   U440 : INV_X1 port map( A => N279, ZN => n845);
   U441 : OAI22_X1 port map( A1 => n740, A2 => n845, B1 => n529, B2 => n757, ZN
                           => n596);
   U442 : OAI22_X1 port map( A1 => n741, A2 => n846, B1 => n530, B2 => n757, ZN
                           => n595);
   U443 : OAI22_X1 port map( A1 => n716, A2 => n847, B1 => n531, B2 => n757, ZN
                           => n594);
   U444 : OAI22_X1 port map( A1 => n671, A2 => n848, B1 => n568, B2 => n757, ZN
                           => n593);
   U445 : OAI22_X1 port map( A1 => n740, A2 => n849, B1 => n569, B2 => n757, ZN
                           => n592);
   U446 : INV_X1 port map( A => n656, ZN => n850);
   U447 : OAI22_X1 port map( A1 => n762, A2 => n850, B1 => n570, B2 => n756, ZN
                           => n591);
   U448 : INV_X1 port map( A => n644, ZN => n851);
   U449 : OAI22_X1 port map( A1 => n624, A2 => n851, B1 => n571, B2 => n756, ZN
                           => n590);
   U450 : INV_X1 port map( A => n697, ZN => n852);
   U451 : OAI22_X1 port map( A1 => n760, A2 => n852, B1 => n572, B2 => n756, ZN
                           => n589);
   U452 : OAI22_X1 port map( A1 => n702, A2 => n853, B1 => n573, B2 => n756, ZN
                           => n588);
   U453 : OAI22_X1 port map( A1 => n622, A2 => n854, B1 => n574, B2 => n756, ZN
                           => n587);
   U454 : OAI22_X1 port map( A1 => n743, A2 => n855, B1 => n575, B2 => n756, ZN
                           => n586);
   U455 : OAI22_X1 port map( A1 => n702, A2 => n856, B1 => n576, B2 => n756, ZN
                           => n585);
   U456 : INV_X1 port map( A => N292, ZN => n858);
   U457 : OAI22_X1 port map( A1 => n615, A2 => n858, B1 => n578, B2 => n756, ZN
                           => n583);
   U458 : INV_X1 port map( A => N293, ZN => n859);
   U459 : OAI22_X1 port map( A1 => n615, A2 => n859, B1 => n579, B2 => n756, ZN
                           => n582);
   U460 : OAI22_X1 port map( A1 => n746, A2 => n740, B1 => n513, B2 => n757, ZN
                           => n612);
   U461 : INV_X1 port map( A => N159, ZN => n875);
   U462 : INV_X1 port map( A => N158, ZN => n874);
   U489 : INV_X1 port map( A => N157, ZN => n873);
   U496 : INV_X1 port map( A => N156, ZN => n872);
   U497 : NAND4_X1 port map( A1 => n875, A2 => n874, A3 => n873, A4 => n872, ZN
                           => n861);
   U498 : NOR4_X1 port map( A1 => n861, A2 => N152, A3 => N154, A4 => N155, ZN 
                           => n863);
   U499 : INV_X1 port map( A => N171, ZN => n884);
   U500 : INV_X1 port map( A => N170, ZN => n883);
   U501 : INV_X1 port map( A => N169, ZN => n882);
   U502 : INV_X1 port map( A => N168, ZN => n881);
   U503 : INV_X1 port map( A => n640, ZN => n888);
   U504 : INV_X1 port map( A => N174, ZN => n887);
   U505 : INV_X1 port map( A => n634, ZN => n886);
   U506 : INV_X1 port map( A => n632, ZN => n885);
   U507 : INV_X1 port map( A => N179, ZN => n892);
   U508 : INV_X1 port map( A => N178, ZN => n891);
   U509 : INV_X1 port map( A => n657, ZN => n890);
   U510 : INV_X1 port map( A => N176, ZN => n889);
   U511 : INV_X1 port map( A => N182, ZN => n867);
   U512 : INV_X1 port map( A => N181, ZN => n894);
   U513 : INV_X1 port map( A => N180, ZN => n893);
   U514 : OAI21_X1 port map( B1 => n200, B2 => n968, A => n897, ZN => n866);
   U515 : NAND2_X1 port map( A1 => n866, A2 => n774, ZN => n900);
   U516 : INV_X1 port map( A => n900, ZN => n898);
   U517 : OAI21_X1 port map( B1 => n639, B2 => n895, A => n763, ZN => n899);
   U518 : OAI22_X1 port map( A1 => n730, A2 => n867, B1 => n386_port, B2 => 
                           n763, ZN => n498);
   U519 : INV_X1 port map( A => N152, ZN => n868);
   U520 : OAI22_X1 port map( A1 => n636, A2 => n868, B1 => n356, B2 => n766, ZN
                           => n468);
   U521 : INV_X1 port map( A => N153, ZN => n869);
   U522 : OAI22_X1 port map( A1 => n869, A2 => n728, B1 => n357, B2 => n765, ZN
                           => n469);
   U523 : INV_X1 port map( A => N154, ZN => n870);
   U524 : OAI22_X1 port map( A1 => n767, A2 => n870, B1 => n358, B2 => n765, ZN
                           => n470);
   U525 : INV_X1 port map( A => N155, ZN => n871);
   U526 : OAI22_X1 port map( A1 => n728, A2 => n871, B1 => n359, B2 => n765, ZN
                           => n471);
   U527 : OAI22_X1 port map( A1 => n731, A2 => n872, B1 => n360, B2 => n765, ZN
                           => n472);
   U528 : OAI22_X1 port map( A1 => n731, A2 => n873, B1 => n361, B2 => n765, ZN
                           => n473);
   U529 : OAI22_X1 port map( A1 => n767, A2 => n874, B1 => n362, B2 => n765, ZN
                           => n474);
   U530 : OAI22_X1 port map( A1 => n767, A2 => n875, B1 => n363, B2 => n765, ZN
                           => n475);
   U531 : OAI22_X1 port map( A1 => n767, A2 => n641, B1 => n364, B2 => n765, ZN
                           => n476);
   U532 : INV_X1 port map( A => N161, ZN => n876);
   U533 : OAI22_X1 port map( A1 => n727, A2 => n876, B1 => n365, B2 => n765, ZN
                           => n477);
   U534 : OAI22_X1 port map( A1 => n767, A2 => n642, B1 => n366, B2 => n765, ZN
                           => n478);
   U535 : OAI22_X1 port map( A1 => n727, A2 => n643, B1 => n367, B2 => n765, ZN
                           => n479);
   U536 : INV_X1 port map( A => N164, ZN => n877);
   U537 : OAI22_X1 port map( A1 => n731, A2 => n877, B1 => n368, B2 => n764, ZN
                           => n480);
   U538 : INV_X1 port map( A => N165, ZN => n878);
   U539 : OAI22_X1 port map( A1 => n729, A2 => n878, B1 => n369, B2 => n764, ZN
                           => n481);
   U540 : INV_X1 port map( A => N166, ZN => n879);
   U541 : OAI22_X1 port map( A1 => n731, A2 => n879, B1 => n370, B2 => n764, ZN
                           => n482);
   U542 : INV_X1 port map( A => N167, ZN => n880);
   U543 : OAI22_X1 port map( A1 => n730, A2 => n880, B1 => n371, B2 => n764, ZN
                           => n483);
   U544 : OAI22_X1 port map( A1 => n728, A2 => n881, B1 => n372, B2 => n764, ZN
                           => n484);
   U545 : OAI22_X1 port map( A1 => n664, A2 => n882, B1 => n373, B2 => n764, ZN
                           => n485);
   U546 : OAI22_X1 port map( A1 => n636, A2 => n648, B1 => n374, B2 => n764, ZN
                           => n486);
   U547 : OAI22_X1 port map( A1 => n664, A2 => n884, B1 => n375, B2 => n764, ZN
                           => n487);
   U548 : OAI22_X1 port map( A1 => n731, A2 => n885, B1 => n376_port, B2 => 
                           n764, ZN => n488);
   U549 : OAI22_X1 port map( A1 => n730, A2 => n886, B1 => n377_port, B2 => 
                           n764, ZN => n489);
   U550 : OAI22_X1 port map( A1 => n727, A2 => n692, B1 => n378_port, B2 => 
                           n763, ZN => n490);
   U551 : OAI22_X1 port map( A1 => n729, A2 => n888, B1 => n379_port, B2 => 
                           n764, ZN => n491);
   U552 : OAI22_X1 port map( A1 => n729, A2 => n889, B1 => n380_port, B2 => 
                           n763, ZN => n492);
   U553 : OAI22_X1 port map( A1 => n730, A2 => n890, B1 => n381_port, B2 => 
                           n763, ZN => n493);
   U554 : OAI22_X1 port map( A1 => n729, A2 => n891, B1 => n382_port, B2 => 
                           n763, ZN => n494);
   U555 : OAI22_X1 port map( A1 => n731, A2 => n892, B1 => n383_port, B2 => 
                           n763, ZN => n495);
   U556 : OAI22_X1 port map( A1 => n664, A2 => n893, B1 => n384_port, B2 => 
                           n763, ZN => n496);
   U557 : OAI22_X1 port map( A1 => n664, A2 => n894, B1 => n385_port, B2 => 
                           n763, ZN => n497);
   U558 : NAND2_X1 port map( A1 => n709, A2 => n763, ZN => n896);
   U559 : OAI22_X1 port map( A1 => N151, A2 => n896, B1 => n425, B2 => n774, ZN
                           => n433);
   U560 : OAI21_X1 port map( B1 => n200, B2 => n966, A => n941, ZN => n901);
   U561 : NAND2_X1 port map( A1 => n901, A2 => n774, ZN => n943);
   U562 : INV_X1 port map( A => n943, ZN => n942);
   U563 : INV_X1 port map( A => N42, ZN => n910);
   U564 : INV_X1 port map( A => N64, ZN => n932);
   U565 : INV_X1 port map( A => N63, ZN => n931);
   U566 : INV_X1 port map( A => N62, ZN => n930);
   U567 : INV_X1 port map( A => N61, ZN => n929);
   U568 : NAND4_X1 port map( A1 => n932, A2 => n931, A3 => n930, A4 => n929, ZN
                           => n902);
   U569 : INV_X1 port map( A => N45, ZN => n913);
   U570 : INV_X1 port map( A => N44, ZN => n912);
   U571 : INV_X1 port map( A => N43, ZN => n911);
   U572 : NOR4_X1 port map( A1 => N46, A2 => N47, A3 => N48, A4 => N49, ZN => 
                           n903);
   U573 : INV_X1 port map( A => N53, ZN => n921);
   U574 : INV_X1 port map( A => N52, ZN => n920);
   U575 : INV_X1 port map( A => N51, ZN => n919);
   U576 : INV_X1 port map( A => N57, ZN => n925);
   U577 : INV_X1 port map( A => N56, ZN => n924);
   U578 : INV_X1 port map( A => N55, ZN => n923);
   U579 : INV_X1 port map( A => N54, ZN => n922);
   U580 : INV_X1 port map( A => N71, ZN => n909);
   U581 : INV_X1 port map( A => N41, ZN => n939);
   U582 : OAI22_X1 port map( A1 => n939, A2 => n725, B1 => n324, B2 => n771, ZN
                           => n436);
   U583 : OAI22_X1 port map( A1 => n910, A2 => n725, B1 => n325, B2 => n771, ZN
                           => n437);
   U584 : OAI22_X1 port map( A1 => n735, A2 => n911, B1 => n326, B2 => n771, ZN
                           => n438);
   U585 : OAI22_X1 port map( A1 => n736, A2 => n912, B1 => n327, B2 => n771, ZN
                           => n439);
   U586 : OAI22_X1 port map( A1 => n734, A2 => n913, B1 => n328, B2 => n771, ZN
                           => n440);
   U587 : INV_X1 port map( A => N46, ZN => n914);
   U588 : OAI22_X1 port map( A1 => n733, A2 => n914, B1 => n329, B2 => n771, ZN
                           => n441);
   U589 : INV_X1 port map( A => N47, ZN => n915);
   U590 : OAI22_X1 port map( A1 => n732, A2 => n915, B1 => n330, B2 => n771, ZN
                           => n442);
   U591 : INV_X1 port map( A => N48, ZN => n916);
   U592 : OAI22_X1 port map( A1 => n662, A2 => n916, B1 => n331, B2 => n771, ZN
                           => n443);
   U593 : INV_X1 port map( A => N49, ZN => n917);
   U594 : OAI22_X1 port map( A1 => n724, A2 => n917, B1 => n332, B2 => n771, ZN
                           => n444);
   U595 : OAI22_X1 port map( A1 => n735, A2 => n919, B1 => n334, B2 => n770, ZN
                           => n446);
   U596 : OAI22_X1 port map( A1 => n662, A2 => n920, B1 => n335, B2 => n770, ZN
                           => n447);
   U597 : OAI22_X1 port map( A1 => n736, A2 => n921, B1 => n336, B2 => n770, ZN
                           => n448);
   U598 : OAI22_X1 port map( A1 => n737, A2 => n922, B1 => n337, B2 => n770, ZN
                           => n449);
   U599 : OAI22_X1 port map( A1 => n734, A2 => n923, B1 => n338, B2 => n770, ZN
                           => n450);
   U600 : OAI22_X1 port map( A1 => n617, A2 => n924, B1 => n339, B2 => n770, ZN
                           => n451);
   U601 : OAI22_X1 port map( A1 => n700, A2 => n925, B1 => n340, B2 => n770, ZN
                           => n452);
   U602 : INV_X1 port map( A => n649, ZN => n926);
   U603 : OAI22_X1 port map( A1 => n737, A2 => n926, B1 => n341, B2 => n770, ZN
                           => n453);
   U604 : INV_X1 port map( A => N59, ZN => n927);
   U605 : OAI22_X1 port map( A1 => n733, A2 => n927, B1 => n342, B2 => n770, ZN
                           => n454);
   U606 : OAI22_X1 port map( A1 => n662, A2 => n929, B1 => n344, B2 => n769, ZN
                           => n456);
   U607 : OAI22_X1 port map( A1 => n616, A2 => n930, B1 => n345, B2 => n769, ZN
                           => n457);
   U608 : OAI22_X1 port map( A1 => n695, A2 => n931, B1 => n346, B2 => n769, ZN
                           => n458);
   U609 : OAI22_X1 port map( A1 => n616, A2 => n932, B1 => n347, B2 => n770, ZN
                           => n459);
   U610 : INV_X1 port map( A => N65, ZN => n933);
   U611 : OAI22_X1 port map( A1 => n732, A2 => n933, B1 => n348, B2 => n769, ZN
                           => n460);
   U612 : INV_X1 port map( A => N66, ZN => n934);
   U613 : OAI22_X1 port map( A1 => n695, A2 => n934, B1 => n349, B2 => n769, ZN
                           => n461);
   U614 : INV_X1 port map( A => N67, ZN => n935);
   U615 : OAI22_X1 port map( A1 => n737, A2 => n935, B1 => n350, B2 => n769, ZN
                           => n462);
   U616 : INV_X1 port map( A => N68, ZN => n936);
   U617 : OAI22_X1 port map( A1 => n732, A2 => n936, B1 => n351, B2 => n769, ZN
                           => n463);
   U618 : INV_X1 port map( A => N69, ZN => n937);
   U619 : OAI22_X1 port map( A1 => n724, A2 => n937, B1 => n352, B2 => n769, ZN
                           => n464);
   U620 : INV_X1 port map( A => N70, ZN => n938);
   U621 : OAI22_X1 port map( A1 => n617, A2 => n938, B1 => n353, B2 => n769, ZN
                           => n465);
   U622 : NAND4_X1 port map( A1 => N40, A2 => n769, A3 => n659, A4 => n939, ZN 
                           => n940);
   U623 : OAI21_X1 port map( B1 => n424, B2 => n774, A => n940, ZN => n434);
   U624 : MUX2_X1 port map( A => n943, B => n621, S => n323, Z => n507);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ISSUE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (63 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ISSUE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (63 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DATAPTH_NBIT32_REG_BIT5
      port( CLK, RST : in std_logic;  PC, IR : in std_logic_vector (31 downto 
            0);  PC_OUT : out std_logic_vector (31 downto 0);  NPC_LATCH_EN, 
            ir_LATCH_EN, signed_op, trap_cs, ret_cs, RF1, RF2, WF1, 
            regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond, sb_op,
            RM, WM, EN3, S3 : in std_logic;  instruction_alu : in 
            std_logic_vector (0 to 5);  DATA_MEM_ADDR, DATA_MEM_IN : out 
            std_logic_vector (31 downto 0);  DATA_MEM_OUT : in std_logic_vector
            (31 downto 0);  DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM : out 
            std_logic);
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
            std_logic;  ALU_OPCODE : out std_logic_vector (0 to 5);  
            signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
            WB_MUX_SEL, RF_WE, lhi_sel, sb_op, s_trap, s_ret : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_25_port, IR_24_port, IR_23_port, IR_22_port, IR_21_port, 
      IR_20_port, IR_19_port, IR_18_port, IR_17_port, IR_16_port, IR_15_port, 
      IR_14_port, IR_13_port, IR_12_port, IR_11_port, IR_10_port, IR_9_port, 
      IR_8_port, IR_7_port, IR_6_port, IR_5_port, IR_4_port, IR_3_port, 
      IR_2_port, IR_1_port, IR_0_port, IR_LATCH_EN_i, PC_31_port, PC_30_port, 
      PC_29_port, PC_28_port, PC_27_port, PC_26_port, PC_25_port, PC_24_port, 
      PC_23_port, PC_22_port, PC_21_port, PC_20_port, PC_19_port, PC_18_port, 
      PC_17_port, PC_16_port, PC_15_port, PC_14_port, PC_13_port, PC_12_port, 
      PC_11_port, PC_10_port, PC_9_port, PC_8_port, PC_7_port, PC_6_port, 
      PC_5_port, PC_4_port, PC_3_port, PC_2_port, PC_1_port, PC_0_port, 
      PC_LATCH_EN_i, NPC_LATCH_EN_i, RegA_LATCH_EN_i, RegB_LATCH_EN_i, 
      RegIMM_LATCH_EN_i, MUXA_SEL_i, MUXB_SEL_i, ALU_OUTREG_EN_i, EQ_COND_i, 
      ALU_OPCODE_i_5_port, ALU_OPCODE_i_4_port, ALU_OPCODE_i_3_port, 
      ALU_OPCODE_i_2_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_0_port, 
      signed_unsigned_i, DRAM_WE_i, LMD_LATCH_EN_i, JUMP_EN_i, WB_MUX_SEL_i, 
      RF_WE_i, lhi_sel_i, sb_op_i, trap_cs_i, ret_cs_i, DATA_MEM_IN_i_31_port, 
      DATA_MEM_IN_i_30_port, DATA_MEM_IN_i_29_port, DATA_MEM_IN_i_28_port, 
      DATA_MEM_IN_i_27_port, DATA_MEM_IN_i_26_port, DATA_MEM_IN_i_25_port, 
      DATA_MEM_IN_i_24_port, DATA_MEM_IN_i_23_port, DATA_MEM_IN_i_22_port, 
      DATA_MEM_IN_i_21_port, DATA_MEM_IN_i_20_port, DATA_MEM_IN_i_19_port, 
      DATA_MEM_IN_i_18_port, DATA_MEM_IN_i_17_port, DATA_MEM_IN_i_16_port, 
      DATA_MEM_IN_i_15_port, DATA_MEM_IN_i_14_port, DATA_MEM_IN_i_13_port, 
      DATA_MEM_IN_i_12_port, DATA_MEM_IN_i_11_port, DATA_MEM_IN_i_10_port, 
      DATA_MEM_IN_i_9_port, DATA_MEM_IN_i_8_port, DATA_MEM_IN_i_7_port, 
      DATA_MEM_IN_i_6_port, DATA_MEM_IN_i_5_port, DATA_MEM_IN_i_4_port, 
      DATA_MEM_IN_i_3_port, DATA_MEM_IN_i_2_port, DATA_MEM_IN_i_1_port, 
      DATA_MEM_IN_i_0_port, dram_data_i_31_port, dram_data_i_30_port, 
      dram_data_i_29_port, dram_data_i_28_port, dram_data_i_27_port, 
      dram_data_i_26_port, dram_data_i_25_port, dram_data_i_24_port, 
      dram_data_i_23_port, dram_data_i_22_port, dram_data_i_21_port, 
      dram_data_i_20_port, dram_data_i_19_port, dram_data_i_18_port, 
      dram_data_i_17_port, dram_data_i_16_port, dram_data_i_15_port, 
      dram_data_i_14_port, dram_data_i_13_port, dram_data_i_12_port, 
      dram_data_i_11_port, dram_data_i_10_port, dram_data_i_9_port, 
      dram_data_i_8_port, dram_data_i_7_port, dram_data_i_6_port, 
      dram_data_i_5_port, dram_data_i_4_port, dram_data_i_3_port, 
      dram_data_i_2_port, dram_data_i_1_port, dram_data_i_0_port, DATA_MEM_WM_i
      , n1, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, 
      n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, 
      n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, 
      n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, 
      n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, 
      n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, 
      n_3214, n_3215, n_3216, n_3217 : std_logic;

begin
   
   DRAM_READNOTWRITE_reg : DFF_X1 port map( D => n271, CK => CLK, Q => 
                           DRAM_READNOTWRITE, QN => n_3169);
   n1 <= '0';
   IR_0_port <= '0';
   IR_1_port <= '0';
   IR_2_port <= '0';
   IR_3_port <= '0';
   IR_4_port <= '0';
   IR_5_port <= '0';
   IR_6_port <= '0';
   IR_7_port <= '0';
   IR_8_port <= '0';
   IR_9_port <= '0';
   IR_10_port <= '0';
   IR_11_port <= '0';
   IR_12_port <= '0';
   IR_13_port <= '0';
   IR_14_port <= '0';
   IR_15_port <= '0';
   IR_16_port <= '0';
   IR_17_port <= '0';
   IR_18_port <= '0';
   IR_19_port <= '0';
   IR_20_port <= '0';
   IR_21_port <= '0';
   IR_22_port <= '0';
   IR_23_port <= '0';
   IR_24_port <= '0';
   IR_25_port <= '0';
   IR_26_port <= '0';
   IR_27_port <= '0';
   IR_28_port <= '0';
   IR_29_port <= '0';
   IR_30_port <= '0';
   IR_31_port <= '0';
   PC_0_port <= '0';
   IRAM_ADDRESS(0) <= '0';
   PC_1_port <= '0';
   IRAM_ADDRESS(1) <= '0';
   PC_2_port <= '0';
   IRAM_ADDRESS(2) <= '0';
   PC_3_port <= '0';
   IRAM_ADDRESS(3) <= '0';
   PC_4_port <= '0';
   IRAM_ADDRESS(4) <= '0';
   PC_5_port <= '0';
   IRAM_ADDRESS(5) <= '0';
   PC_6_port <= '0';
   IRAM_ADDRESS(6) <= '0';
   PC_7_port <= '0';
   IRAM_ADDRESS(7) <= '0';
   PC_8_port <= '0';
   IRAM_ADDRESS(8) <= '0';
   PC_9_port <= '0';
   IRAM_ADDRESS(9) <= '0';
   PC_10_port <= '0';
   IRAM_ADDRESS(10) <= '0';
   PC_11_port <= '0';
   IRAM_ADDRESS(11) <= '0';
   PC_12_port <= '0';
   IRAM_ADDRESS(12) <= '0';
   PC_13_port <= '0';
   IRAM_ADDRESS(13) <= '0';
   PC_14_port <= '0';
   IRAM_ADDRESS(14) <= '0';
   PC_15_port <= '0';
   IRAM_ADDRESS(15) <= '0';
   PC_16_port <= '0';
   IRAM_ADDRESS(16) <= '0';
   PC_17_port <= '0';
   IRAM_ADDRESS(17) <= '0';
   PC_18_port <= '0';
   IRAM_ADDRESS(18) <= '0';
   PC_19_port <= '0';
   IRAM_ADDRESS(19) <= '0';
   PC_20_port <= '0';
   IRAM_ADDRESS(20) <= '0';
   PC_21_port <= '0';
   IRAM_ADDRESS(21) <= '0';
   PC_22_port <= '0';
   IRAM_ADDRESS(22) <= '0';
   PC_23_port <= '0';
   IRAM_ADDRESS(23) <= '0';
   PC_24_port <= '0';
   IRAM_ADDRESS(24) <= '0';
   PC_25_port <= '0';
   IRAM_ADDRESS(25) <= '0';
   PC_26_port <= '0';
   IRAM_ADDRESS(26) <= '0';
   PC_27_port <= '0';
   IRAM_ADDRESS(27) <= '0';
   PC_28_port <= '0';
   IRAM_ADDRESS(28) <= '0';
   PC_29_port <= '0';
   IRAM_ADDRESS(29) <= '0';
   PC_30_port <= '0';
   IRAM_ADDRESS(30) <= '0';
   PC_31_port <= '0';
   IRAM_ADDRESS(31) <= '0';
   RF_WE_i <= '0';
   WB_MUX_SEL_i <= '0';
   PC_LATCH_EN_i <= '0';
   JUMP_EN_i <= '0';
   LMD_LATCH_EN_i <= '0';
   DRAM_WE_i <= '0';
   EQ_COND_i <= '0';
   ALU_OUTREG_EN_i <= '0';
   MUXB_SEL_i <= '0';
   MUXA_SEL_i <= '0';
   RegIMM_LATCH_EN_i <= '0';
   RegB_LATCH_EN_i <= '0';
   RegA_LATCH_EN_i <= '0';
   NPC_LATCH_EN_i <= '0';
   IR_LATCH_EN_i <= '0';
   CU_I : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 
                           port map( Clk => CLK, Rst => RST, IR_IN(31) => 
                           IR_31_port, IR_IN(30) => IR_30_port, IR_IN(29) => 
                           IR_29_port, IR_IN(28) => IR_28_port, IR_IN(27) => 
                           IR_27_port, IR_IN(26) => IR_26_port, IR_IN(25) => 
                           IR_25_port, IR_IN(24) => IR_24_port, IR_IN(23) => 
                           IR_23_port, IR_IN(22) => IR_22_port, IR_IN(21) => 
                           IR_21_port, IR_IN(20) => IR_20_port, IR_IN(19) => 
                           IR_19_port, IR_IN(18) => IR_18_port, IR_IN(17) => 
                           IR_17_port, IR_IN(16) => IR_16_port, IR_IN(15) => 
                           IR_15_port, IR_IN(14) => IR_14_port, IR_IN(13) => 
                           IR_13_port, IR_IN(12) => IR_12_port, IR_IN(11) => 
                           IR_11_port, IR_IN(10) => IR_10_port, IR_IN(9) => 
                           IR_9_port, IR_IN(8) => IR_8_port, IR_IN(7) => 
                           IR_7_port, IR_IN(6) => IR_6_port, IR_IN(5) => 
                           IR_5_port, IR_IN(4) => IR_4_port, IR_IN(3) => 
                           IR_3_port, IR_IN(2) => IR_2_port, IR_IN(1) => 
                           IR_1_port, IR_IN(0) => IR_0_port, IR_LATCH_EN => 
                           n_3170, NPC_LATCH_EN => n_3171, RegA_LATCH_EN => 
                           n_3172, RegB_LATCH_EN => n_3173, RegIMM_LATCH_EN => 
                           n_3174, MUXA_SEL => n_3175, MUXB_SEL => n_3176, 
                           ALU_OUTREG_EN => n_3177, EQ_COND => n_3178, 
                           ALU_OPCODE(0) => ALU_OPCODE_i_5_port, ALU_OPCODE(1) 
                           => ALU_OPCODE_i_4_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_i_0_port, signed_unsigned => 
                           signed_unsigned_i, DRAM_WE => n_3179, LMD_LATCH_EN 
                           => n_3180, JUMP_EN => n_3181, PC_LATCH_EN => n_3182,
                           WB_MUX_SEL => n_3183, RF_WE => n_3184, lhi_sel => 
                           lhi_sel_i, sb_op => sb_op_i, s_trap => trap_cs_i, 
                           s_ret => ret_cs_i);
   DTPTH_I : DATAPTH_NBIT32_REG_BIT5 port map( CLK => CLK, RST => RST, PC(31) 
                           => PC_31_port, PC(30) => PC_30_port, PC(29) => 
                           PC_29_port, PC(28) => PC_28_port, PC(27) => 
                           PC_27_port, PC(26) => PC_26_port, PC(25) => 
                           PC_25_port, PC(24) => PC_24_port, PC(23) => 
                           PC_23_port, PC(22) => PC_22_port, PC(21) => 
                           PC_21_port, PC(20) => PC_20_port, PC(19) => 
                           PC_19_port, PC(18) => PC_18_port, PC(17) => 
                           PC_17_port, PC(16) => PC_16_port, PC(15) => 
                           PC_15_port, PC(14) => PC_14_port, PC(13) => 
                           PC_13_port, PC(12) => PC_12_port, PC(11) => 
                           PC_11_port, PC(10) => PC_10_port, PC(9) => PC_9_port
                           , PC(8) => PC_8_port, PC(7) => PC_7_port, PC(6) => 
                           PC_6_port, PC(5) => PC_5_port, PC(4) => PC_4_port, 
                           PC(3) => PC_3_port, PC(2) => PC_2_port, PC(1) => 
                           PC_1_port, PC(0) => PC_0_port, IR(31) => IR_31_port,
                           IR(30) => IR_30_port, IR(29) => IR_29_port, IR(28) 
                           => IR_28_port, IR(27) => IR_27_port, IR(26) => 
                           IR_26_port, IR(25) => IR_25_port, IR(24) => 
                           IR_24_port, IR(23) => IR_23_port, IR(22) => 
                           IR_22_port, IR(21) => IR_21_port, IR(20) => 
                           IR_20_port, IR(19) => IR_19_port, IR(18) => 
                           IR_18_port, IR(17) => IR_17_port, IR(16) => 
                           IR_16_port, IR(15) => IR_15_port, IR(14) => 
                           IR_14_port, IR(13) => IR_13_port, IR(12) => 
                           IR_12_port, IR(11) => IR_11_port, IR(10) => 
                           IR_10_port, IR(9) => IR_9_port, IR(8) => IR_8_port, 
                           IR(7) => IR_7_port, IR(6) => IR_6_port, IR(5) => 
                           IR_5_port, IR(4) => IR_4_port, IR(3) => IR_3_port, 
                           IR(2) => IR_2_port, IR(1) => IR_1_port, IR(0) => 
                           IR_0_port, PC_OUT(31) => n_3185, PC_OUT(30) => 
                           n_3186, PC_OUT(29) => n_3187, PC_OUT(28) => n_3188, 
                           PC_OUT(27) => n_3189, PC_OUT(26) => n_3190, 
                           PC_OUT(25) => n_3191, PC_OUT(24) => n_3192, 
                           PC_OUT(23) => n_3193, PC_OUT(22) => n_3194, 
                           PC_OUT(21) => n_3195, PC_OUT(20) => n_3196, 
                           PC_OUT(19) => n_3197, PC_OUT(18) => n_3198, 
                           PC_OUT(17) => n_3199, PC_OUT(16) => n_3200, 
                           PC_OUT(15) => n_3201, PC_OUT(14) => n_3202, 
                           PC_OUT(13) => n_3203, PC_OUT(12) => n_3204, 
                           PC_OUT(11) => n_3205, PC_OUT(10) => n_3206, 
                           PC_OUT(9) => n_3207, PC_OUT(8) => n_3208, PC_OUT(7) 
                           => n_3209, PC_OUT(6) => n_3210, PC_OUT(5) => n_3211,
                           PC_OUT(4) => n_3212, PC_OUT(3) => n_3213, PC_OUT(2) 
                           => n_3214, PC_OUT(1) => n_3215, PC_OUT(0) => n_3216,
                           NPC_LATCH_EN => NPC_LATCH_EN_i, ir_LATCH_EN => 
                           IR_LATCH_EN_i, signed_op => signed_unsigned_i, 
                           trap_cs => trap_cs_i, ret_cs => ret_cs_i, RF1 => 
                           RegA_LATCH_EN_i, RF2 => RegB_LATCH_EN_i, WF1 => 
                           RF_WE_i, regImm_LATCH_EN => RegIMM_LATCH_EN_i, S1 =>
                           MUXA_SEL_i, S2 => MUXB_SEL_i, EN2 => ALU_OUTREG_EN_i
                           , lhi_sel => lhi_sel_i, jump_en => JUMP_EN_i, 
                           branch_cond => EQ_COND_i, sb_op => sb_op_i, RM => 
                           LMD_LATCH_EN_i, WM => DRAM_WE_i, EN3 => 
                           PC_LATCH_EN_i, S3 => WB_MUX_SEL_i, 
                           instruction_alu(0) => ALU_OPCODE_i_5_port, 
                           instruction_alu(1) => ALU_OPCODE_i_4_port, 
                           instruction_alu(2) => ALU_OPCODE_i_3_port, 
                           instruction_alu(3) => ALU_OPCODE_i_2_port, 
                           instruction_alu(4) => ALU_OPCODE_i_1_port, 
                           instruction_alu(5) => ALU_OPCODE_i_0_port, 
                           DATA_MEM_ADDR(31) => DRAM_ADDRESS(31), 
                           DATA_MEM_ADDR(30) => DRAM_ADDRESS(30), 
                           DATA_MEM_ADDR(29) => DRAM_ADDRESS(29), 
                           DATA_MEM_ADDR(28) => DRAM_ADDRESS(28), 
                           DATA_MEM_ADDR(27) => DRAM_ADDRESS(27), 
                           DATA_MEM_ADDR(26) => DRAM_ADDRESS(26), 
                           DATA_MEM_ADDR(25) => DRAM_ADDRESS(25), 
                           DATA_MEM_ADDR(24) => DRAM_ADDRESS(24), 
                           DATA_MEM_ADDR(23) => DRAM_ADDRESS(23), 
                           DATA_MEM_ADDR(22) => DRAM_ADDRESS(22), 
                           DATA_MEM_ADDR(21) => DRAM_ADDRESS(21), 
                           DATA_MEM_ADDR(20) => DRAM_ADDRESS(20), 
                           DATA_MEM_ADDR(19) => DRAM_ADDRESS(19), 
                           DATA_MEM_ADDR(18) => DRAM_ADDRESS(18), 
                           DATA_MEM_ADDR(17) => DRAM_ADDRESS(17), 
                           DATA_MEM_ADDR(16) => DRAM_ADDRESS(16), 
                           DATA_MEM_ADDR(15) => DRAM_ADDRESS(15), 
                           DATA_MEM_ADDR(14) => DRAM_ADDRESS(14), 
                           DATA_MEM_ADDR(13) => DRAM_ADDRESS(13), 
                           DATA_MEM_ADDR(12) => DRAM_ADDRESS(12), 
                           DATA_MEM_ADDR(11) => DRAM_ADDRESS(11), 
                           DATA_MEM_ADDR(10) => DRAM_ADDRESS(10), 
                           DATA_MEM_ADDR(9) => DRAM_ADDRESS(9), 
                           DATA_MEM_ADDR(8) => DRAM_ADDRESS(8), 
                           DATA_MEM_ADDR(7) => DRAM_ADDRESS(7), 
                           DATA_MEM_ADDR(6) => DRAM_ADDRESS(6), 
                           DATA_MEM_ADDR(5) => DRAM_ADDRESS(5), 
                           DATA_MEM_ADDR(4) => DRAM_ADDRESS(4), 
                           DATA_MEM_ADDR(3) => DRAM_ADDRESS(3), 
                           DATA_MEM_ADDR(2) => DRAM_ADDRESS(2), 
                           DATA_MEM_ADDR(1) => DRAM_ADDRESS(1), 
                           DATA_MEM_ADDR(0) => DRAM_ADDRESS(0), DATA_MEM_IN(31)
                           => DATA_MEM_IN_i_31_port, DATA_MEM_IN(30) => 
                           DATA_MEM_IN_i_30_port, DATA_MEM_IN(29) => 
                           DATA_MEM_IN_i_29_port, DATA_MEM_IN(28) => 
                           DATA_MEM_IN_i_28_port, DATA_MEM_IN(27) => 
                           DATA_MEM_IN_i_27_port, DATA_MEM_IN(26) => 
                           DATA_MEM_IN_i_26_port, DATA_MEM_IN(25) => 
                           DATA_MEM_IN_i_25_port, DATA_MEM_IN(24) => 
                           DATA_MEM_IN_i_24_port, DATA_MEM_IN(23) => 
                           DATA_MEM_IN_i_23_port, DATA_MEM_IN(22) => 
                           DATA_MEM_IN_i_22_port, DATA_MEM_IN(21) => 
                           DATA_MEM_IN_i_21_port, DATA_MEM_IN(20) => 
                           DATA_MEM_IN_i_20_port, DATA_MEM_IN(19) => 
                           DATA_MEM_IN_i_19_port, DATA_MEM_IN(18) => 
                           DATA_MEM_IN_i_18_port, DATA_MEM_IN(17) => 
                           DATA_MEM_IN_i_17_port, DATA_MEM_IN(16) => 
                           DATA_MEM_IN_i_16_port, DATA_MEM_IN(15) => 
                           DATA_MEM_IN_i_15_port, DATA_MEM_IN(14) => 
                           DATA_MEM_IN_i_14_port, DATA_MEM_IN(13) => 
                           DATA_MEM_IN_i_13_port, DATA_MEM_IN(12) => 
                           DATA_MEM_IN_i_12_port, DATA_MEM_IN(11) => 
                           DATA_MEM_IN_i_11_port, DATA_MEM_IN(10) => 
                           DATA_MEM_IN_i_10_port, DATA_MEM_IN(9) => 
                           DATA_MEM_IN_i_9_port, DATA_MEM_IN(8) => 
                           DATA_MEM_IN_i_8_port, DATA_MEM_IN(7) => 
                           DATA_MEM_IN_i_7_port, DATA_MEM_IN(6) => 
                           DATA_MEM_IN_i_6_port, DATA_MEM_IN(5) => 
                           DATA_MEM_IN_i_5_port, DATA_MEM_IN(4) => 
                           DATA_MEM_IN_i_4_port, DATA_MEM_IN(3) => 
                           DATA_MEM_IN_i_3_port, DATA_MEM_IN(2) => 
                           DATA_MEM_IN_i_2_port, DATA_MEM_IN(1) => 
                           DATA_MEM_IN_i_1_port, DATA_MEM_IN(0) => 
                           DATA_MEM_IN_i_0_port, DATA_MEM_OUT(31) => 
                           dram_data_i_31_port, DATA_MEM_OUT(30) => 
                           dram_data_i_30_port, DATA_MEM_OUT(29) => 
                           dram_data_i_29_port, DATA_MEM_OUT(28) => 
                           dram_data_i_28_port, DATA_MEM_OUT(27) => 
                           dram_data_i_27_port, DATA_MEM_OUT(26) => 
                           dram_data_i_26_port, DATA_MEM_OUT(25) => 
                           dram_data_i_25_port, DATA_MEM_OUT(24) => 
                           dram_data_i_24_port, DATA_MEM_OUT(23) => 
                           dram_data_i_23_port, DATA_MEM_OUT(22) => 
                           dram_data_i_22_port, DATA_MEM_OUT(21) => 
                           dram_data_i_21_port, DATA_MEM_OUT(20) => 
                           dram_data_i_20_port, DATA_MEM_OUT(19) => 
                           dram_data_i_19_port, DATA_MEM_OUT(18) => 
                           dram_data_i_18_port, DATA_MEM_OUT(17) => 
                           dram_data_i_17_port, DATA_MEM_OUT(16) => 
                           dram_data_i_16_port, DATA_MEM_OUT(15) => 
                           dram_data_i_15_port, DATA_MEM_OUT(14) => 
                           dram_data_i_14_port, DATA_MEM_OUT(13) => 
                           dram_data_i_13_port, DATA_MEM_OUT(12) => 
                           dram_data_i_12_port, DATA_MEM_OUT(11) => 
                           dram_data_i_11_port, DATA_MEM_OUT(10) => 
                           dram_data_i_10_port, DATA_MEM_OUT(9) => 
                           dram_data_i_9_port, DATA_MEM_OUT(8) => 
                           dram_data_i_8_port, DATA_MEM_OUT(7) => 
                           dram_data_i_7_port, DATA_MEM_OUT(6) => 
                           dram_data_i_6_port, DATA_MEM_OUT(5) => 
                           dram_data_i_5_port, DATA_MEM_OUT(4) => 
                           dram_data_i_4_port, DATA_MEM_OUT(3) => 
                           dram_data_i_3_port, DATA_MEM_OUT(2) => 
                           dram_data_i_2_port, DATA_MEM_OUT(1) => 
                           dram_data_i_1_port, DATA_MEM_OUT(0) => 
                           dram_data_i_0_port, DATA_MEM_ENABLE => DRAM_ISSUE, 
                           DATA_MEM_RM => n_3217, DATA_MEM_WM => DATA_MEM_WM_i)
                           ;
   DRAM_DATA_tri_32_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(32));
   DRAM_DATA_tri_33_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(33));
   DRAM_DATA_tri_34_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(34));
   DRAM_DATA_tri_35_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(35));
   DRAM_DATA_tri_36_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(36));
   DRAM_DATA_tri_37_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(37));
   DRAM_DATA_tri_38_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(38));
   DRAM_DATA_tri_39_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(39));
   DRAM_DATA_tri_40_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(40));
   DRAM_DATA_tri_41_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(41));
   DRAM_DATA_tri_42_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(42));
   DRAM_DATA_tri_43_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(43));
   DRAM_DATA_tri_44_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(44));
   DRAM_DATA_tri_45_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(45));
   DRAM_DATA_tri_46_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(46));
   DRAM_DATA_tri_47_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(47));
   DRAM_DATA_tri_48_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(48));
   DRAM_DATA_tri_49_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(49));
   DRAM_DATA_tri_50_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(50));
   DRAM_DATA_tri_51_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(51));
   DRAM_DATA_tri_52_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(52));
   DRAM_DATA_tri_53_inst : TBUF_X1 port map( A => n1, EN => n265, Z => 
                           DRAM_DATA(53));
   DRAM_DATA_tri_54_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(54));
   DRAM_DATA_tri_55_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(55));
   DRAM_DATA_tri_56_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(56));
   DRAM_DATA_tri_57_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(57));
   DRAM_DATA_tri_58_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(58));
   DRAM_DATA_tri_59_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(59));
   DRAM_DATA_tri_60_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(60));
   DRAM_DATA_tri_61_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(61));
   DRAM_DATA_tri_62_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(62));
   DRAM_DATA_tri_63_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(63));
   DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_8_port, EN => 
                           n267, Z => DRAM_DATA(8));
   DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_9_port, EN => 
                           n267, Z => DRAM_DATA(9));
   DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_10_port, EN => 
                           n267, Z => DRAM_DATA(10));
   DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_11_port, EN => 
                           n267, Z => DRAM_DATA(11));
   DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_12_port, EN => 
                           n268, Z => DRAM_DATA(12));
   DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_13_port, EN => 
                           n268, Z => DRAM_DATA(13));
   DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_14_port, EN => 
                           n268, Z => DRAM_DATA(14));
   DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_15_port, EN => 
                           n268, Z => DRAM_DATA(15));
   DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_16_port, EN => 
                           n268, Z => DRAM_DATA(16));
   DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_17_port, EN => 
                           n268, Z => DRAM_DATA(17));
   DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_18_port, EN => 
                           n268, Z => DRAM_DATA(18));
   DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_19_port, EN => 
                           n268, Z => DRAM_DATA(19));
   DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_20_port, EN => 
                           n268, Z => DRAM_DATA(20));
   DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_21_port, EN => 
                           n268, Z => DRAM_DATA(21));
   DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_22_port, EN => 
                           n268, Z => DRAM_DATA(22));
   DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_23_port, EN => 
                           n269, Z => DRAM_DATA(23));
   DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_24_port, EN => 
                           n269, Z => DRAM_DATA(24));
   DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_25_port, EN => 
                           n269, Z => DRAM_DATA(25));
   DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_26_port, EN => 
                           n269, Z => DRAM_DATA(26));
   DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_27_port, EN => 
                           n269, Z => DRAM_DATA(27));
   DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_28_port, EN => 
                           n269, Z => DRAM_DATA(28));
   DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_29_port, EN => 
                           n269, Z => DRAM_DATA(29));
   DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_30_port, EN => 
                           n269, Z => DRAM_DATA(30));
   DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_31_port, EN => 
                           n269, Z => DRAM_DATA(31));
   DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_0_port, EN => 
                           n266, Z => DRAM_DATA(0));
   DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_1_port, EN => 
                           n267, Z => DRAM_DATA(1));
   DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_2_port, EN => 
                           n267, Z => DRAM_DATA(2));
   DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_3_port, EN => 
                           n267, Z => DRAM_DATA(3));
   DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_4_port, EN => 
                           n267, Z => DRAM_DATA(4));
   DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_5_port, EN => 
                           n267, Z => DRAM_DATA(5));
   DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_6_port, EN => 
                           n267, Z => DRAM_DATA(6));
   DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_7_port, EN => 
                           n267, Z => DRAM_DATA(7));
   U342 : BUF_X1 port map( A => n263, Z => n270);
   U343 : BUF_X1 port map( A => n263, Z => n269);
   U344 : BUF_X1 port map( A => n263, Z => n268);
   U345 : BUF_X1 port map( A => n262, Z => n267);
   U346 : BUF_X1 port map( A => n262, Z => n266);
   U347 : BUF_X1 port map( A => n262, Z => n265);
   U348 : BUF_X1 port map( A => n262, Z => n264);
   U349 : BUF_X1 port map( A => n263, Z => n271);
   U350 : BUF_X1 port map( A => n272, Z => n262);
   U351 : BUF_X1 port map( A => n272, Z => n263);
   U352 : AND2_X1 port map( A1 => DRAM_DATA(63), A2 => n271, ZN => 
                           dram_data_i_31_port);
   U353 : AND2_X1 port map( A1 => DRAM_DATA(40), A2 => n271, ZN => 
                           dram_data_i_8_port);
   U354 : AND2_X1 port map( A1 => DRAM_DATA(41), A2 => n271, ZN => 
                           dram_data_i_9_port);
   U355 : AND2_X1 port map( A1 => DRAM_DATA(42), A2 => n269, ZN => 
                           dram_data_i_10_port);
   U356 : AND2_X1 port map( A1 => DRAM_DATA(43), A2 => n269, ZN => 
                           dram_data_i_11_port);
   U357 : AND2_X1 port map( A1 => DRAM_DATA(44), A2 => n270, ZN => 
                           dram_data_i_12_port);
   U358 : AND2_X1 port map( A1 => DRAM_DATA(45), A2 => n270, ZN => 
                           dram_data_i_13_port);
   U359 : AND2_X1 port map( A1 => DRAM_DATA(46), A2 => n270, ZN => 
                           dram_data_i_14_port);
   U360 : AND2_X1 port map( A1 => DRAM_DATA(47), A2 => n270, ZN => 
                           dram_data_i_15_port);
   U361 : AND2_X1 port map( A1 => DRAM_DATA(52), A2 => n270, ZN => 
                           dram_data_i_20_port);
   U362 : AND2_X1 port map( A1 => DRAM_DATA(53), A2 => n270, ZN => 
                           dram_data_i_21_port);
   U363 : AND2_X1 port map( A1 => DRAM_DATA(54), A2 => n270, ZN => 
                           dram_data_i_22_port);
   U364 : AND2_X1 port map( A1 => DRAM_DATA(55), A2 => n270, ZN => 
                           dram_data_i_23_port);
   U365 : AND2_X1 port map( A1 => DRAM_DATA(56), A2 => n270, ZN => 
                           dram_data_i_24_port);
   U366 : AND2_X1 port map( A1 => DRAM_DATA(57), A2 => n270, ZN => 
                           dram_data_i_25_port);
   U367 : AND2_X1 port map( A1 => DRAM_DATA(58), A2 => n270, ZN => 
                           dram_data_i_26_port);
   U368 : AND2_X1 port map( A1 => DRAM_DATA(59), A2 => n271, ZN => 
                           dram_data_i_27_port);
   U369 : AND2_X1 port map( A1 => DRAM_DATA(60), A2 => n271, ZN => 
                           dram_data_i_28_port);
   U370 : AND2_X1 port map( A1 => DRAM_DATA(61), A2 => n271, ZN => 
                           dram_data_i_29_port);
   U371 : AND2_X1 port map( A1 => DRAM_DATA(62), A2 => n271, ZN => 
                           dram_data_i_30_port);
   U372 : AND2_X1 port map( A1 => DRAM_DATA(48), A2 => n270, ZN => 
                           dram_data_i_16_port);
   U373 : AND2_X1 port map( A1 => DRAM_DATA(49), A2 => n270, ZN => 
                           dram_data_i_17_port);
   U374 : AND2_X1 port map( A1 => DRAM_DATA(50), A2 => n270, ZN => 
                           dram_data_i_18_port);
   U375 : AND2_X1 port map( A1 => DRAM_DATA(51), A2 => n270, ZN => 
                           dram_data_i_19_port);
   U376 : AND2_X1 port map( A1 => DRAM_DATA(32), A2 => n269, ZN => 
                           dram_data_i_0_port);
   U377 : AND2_X1 port map( A1 => DRAM_DATA(33), A2 => n270, ZN => 
                           dram_data_i_1_port);
   U378 : AND2_X1 port map( A1 => DRAM_DATA(34), A2 => n271, ZN => 
                           dram_data_i_2_port);
   U379 : AND2_X1 port map( A1 => DRAM_DATA(35), A2 => n271, ZN => 
                           dram_data_i_3_port);
   U380 : AND2_X1 port map( A1 => DRAM_DATA(36), A2 => n271, ZN => 
                           dram_data_i_4_port);
   U381 : AND2_X1 port map( A1 => DRAM_DATA(37), A2 => n271, ZN => 
                           dram_data_i_5_port);
   U382 : AND2_X1 port map( A1 => DRAM_DATA(38), A2 => n271, ZN => 
                           dram_data_i_6_port);
   U383 : AND2_X1 port map( A1 => DRAM_DATA(39), A2 => n271, ZN => 
                           dram_data_i_7_port);
   U384 : INV_X1 port map( A => DATA_MEM_WM_i, ZN => n272);

end SYN_dlx_rtl;



    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 ( 
        Clk, Rst, IR_IN, IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, 
        RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
        EQ_COND, .ALU_OPCODE({\ALU_OPCODE[5] , \ALU_OPCODE[4] , 
        \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), 
        signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
        WB_MUX_SEL, RF_WE, lhi_sel, sb_op );
  input [31:0] IR_IN;
  input Clk, Rst;
  output IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN,
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND,
         \ALU_OPCODE[5] , \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] ,
         \ALU_OPCODE[1] , \ALU_OPCODE[0] , signed_unsigned, DRAM_WE,
         LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE, lhi_sel, sb_op;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26, n3,
         signed_unsigned_i, N393, N394, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n146, n147, n148, n149, n150, n1;
  wire   [5:0] ALU_OPCODE;
  wire   [5:0] aluOpcode1;
  wire   [5:0] aluOpcode2;
  wire   [5:0] aluOpcode_i;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];
  assign IR_LATCH_EN = 1'b0;
  assign NPC_LATCH_EN = 1'b0;
  assign RegA_LATCH_EN = 1'b0;
  assign RegB_LATCH_EN = 1'b0;
  assign RegIMM_LATCH_EN = 1'b0;
  assign MUXA_SEL = 1'b0;
  assign MUXB_SEL = 1'b0;
  assign ALU_OUTREG_EN = 1'b0;
  assign EQ_COND = 1'b0;
  assign DRAM_WE = 1'b0;
  assign LMD_LATCH_EN = 1'b0;
  assign JUMP_EN = 1'b0;
  assign PC_LATCH_EN = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign RF_WE = 1'b0;

  DFFR_X1 \aluOpcode1_reg[5]  ( .D(aluOpcode_i[5]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[5]) );
  DFFR_X1 \aluOpcode1_reg[4]  ( .D(aluOpcode_i[4]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[4]) );
  DFFR_X1 \aluOpcode1_reg[3]  ( .D(aluOpcode_i[3]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[3]) );
  DFFR_X1 \aluOpcode1_reg[2]  ( .D(aluOpcode_i[2]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[2]) );
  DFFR_X1 \aluOpcode1_reg[1]  ( .D(aluOpcode_i[1]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[1]) );
  DFFR_X1 \aluOpcode1_reg[0]  ( .D(aluOpcode_i[0]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[0]) );
  DFFR_X1 \aluOpcode2_reg[5]  ( .D(aluOpcode1[5]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[5]) );
  DFFR_X1 \aluOpcode2_reg[4]  ( .D(aluOpcode1[4]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[4]) );
  DFFR_X1 \aluOpcode2_reg[3]  ( .D(aluOpcode1[3]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[3]) );
  DFFR_X1 \aluOpcode2_reg[2]  ( .D(aluOpcode1[2]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[2]) );
  DFFR_X1 \aluOpcode2_reg[1]  ( .D(aluOpcode1[1]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[1]) );
  DFFR_X1 \aluOpcode2_reg[0]  ( .D(aluOpcode1[0]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[0]) );
  DFFR_X1 \aluOpcode3_reg[5]  ( .D(aluOpcode2[5]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[5]) );
  DFFR_X1 \aluOpcode3_reg[4]  ( .D(aluOpcode2[4]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[4]) );
  DFFR_X1 \aluOpcode3_reg[3]  ( .D(aluOpcode2[3]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[3]) );
  DFFR_X1 \aluOpcode3_reg[2]  ( .D(aluOpcode2[2]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[2]) );
  DFFR_X1 \aluOpcode3_reg[1]  ( .D(aluOpcode2[1]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[1]) );
  DFFR_X1 \aluOpcode3_reg[0]  ( .D(aluOpcode2[0]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[0]) );
  DLH_X1 signed_unsigned_i_reg ( .G(N393), .D(N394), .Q(signed_unsigned_i) );
  DFF_X1 signed_unsigned_2_reg ( .D(n149), .CK(Clk), .Q(signed_unsigned), .QN(
        n145) );
  DFF_X1 lhi_sel_reg ( .D(n148), .CK(Clk), .Q(n3), .QN(n143) );
  DFF_X1 sb_op_reg ( .D(n147), .CK(Clk), .Q(sb_op), .QN(n146) );
  NOR2_X1 U3 ( .A1(Rst), .A2(n146), .ZN(n147) );
  NOR2_X1 U4 ( .A1(n143), .A2(Rst), .ZN(n148) );
  OAI22_X1 U5 ( .A1(n9), .A2(n10), .B1(Rst), .B2(n145), .ZN(n149) );
  INV_X1 U6 ( .A(Rst), .ZN(n9) );
  OAI21_X1 U7 ( .B1(Rst), .B2(n10), .A(n11), .ZN(n150) );
  NAND2_X1 U8 ( .A1(signed_unsigned_i), .A2(Rst), .ZN(n11) );
  OAI211_X1 U10 ( .C1(n12), .C2(n13), .A(n14), .B(n15), .ZN(aluOpcode_i[5]) );
  INV_X1 U11 ( .A(n16), .ZN(n15) );
  OAI211_X1 U12 ( .C1(n17), .C2(n18), .A(n19), .B(n20), .ZN(n16) );
  AND3_X1 U13 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n18) );
  NAND3_X1 U14 ( .A1(IR_IN[0]), .A2(n24), .A3(IR_IN[1]), .ZN(n22) );
  OAI211_X1 U15 ( .C1(n25), .C2(n17), .A(n26), .B(n27), .ZN(aluOpcode_i[4]) );
  OAI211_X1 U16 ( .C1(n28), .C2(n17), .A(n14), .B(n29), .ZN(aluOpcode_i[3]) );
  NOR2_X1 U17 ( .A1(n30), .A2(n31), .ZN(n29) );
  NOR3_X1 U18 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n28) );
  INV_X1 U19 ( .A(n25), .ZN(n33) );
  NOR2_X1 U20 ( .A1(n35), .A2(n36), .ZN(n25) );
  INV_X1 U21 ( .A(n37), .ZN(n36) );
  OAI21_X1 U22 ( .B1(n38), .B2(n39), .A(n40), .ZN(n32) );
  NAND3_X1 U23 ( .A1(n41), .A2(n42), .A3(n43), .ZN(aluOpcode_i[2]) );
  AOI221_X1 U24 ( .B1(n44), .B2(n45), .C1(n46), .C2(n47), .A(n48), .ZN(n43) );
  NAND2_X1 U25 ( .A1(n49), .A2(n50), .ZN(n47) );
  AOI21_X1 U26 ( .B1(n51), .B2(n52), .A(n53), .ZN(n41) );
  OAI211_X1 U27 ( .C1(n54), .C2(n17), .A(n55), .B(n56), .ZN(aluOpcode_i[1]) );
  AOI221_X1 U28 ( .B1(n51), .B2(n57), .C1(n58), .C2(n59), .A(n60), .ZN(n56) );
  NOR2_X1 U29 ( .A1(n61), .A2(n62), .ZN(n55) );
  AOI21_X1 U30 ( .B1(n13), .B2(n63), .A(n64), .ZN(n62) );
  AND3_X1 U31 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n54) );
  NAND3_X1 U32 ( .A1(n68), .A2(n69), .A3(n70), .ZN(aluOpcode_i[0]) );
  AOI211_X1 U33 ( .C1(n51), .C2(n45), .A(n60), .B(n71), .ZN(n70) );
  OAI211_X1 U34 ( .C1(n72), .C2(n13), .A(n73), .B(n74), .ZN(n60) );
  NOR2_X1 U35 ( .A1(n48), .A2(n75), .ZN(n74) );
  NOR3_X1 U36 ( .A1(n76), .A2(IR_IN_29), .A3(n64), .ZN(n75) );
  INV_X1 U37 ( .A(n57), .ZN(n72) );
  INV_X1 U38 ( .A(n77), .ZN(n51) );
  AOI21_X1 U39 ( .B1(n46), .B2(n78), .A(n79), .ZN(n69) );
  NAND4_X1 U40 ( .A1(n80), .A2(n81), .A3(n82), .A4(n83), .ZN(n78) );
  AND4_X1 U41 ( .A1(n21), .A2(n84), .A3(n37), .A4(n85), .ZN(n83) );
  OAI21_X1 U42 ( .B1(n86), .B2(n87), .A(n88), .ZN(n82) );
  OAI21_X1 U43 ( .B1(n89), .B2(n87), .A(n90), .ZN(n80) );
  INV_X1 U44 ( .A(n38), .ZN(n87) );
  NOR2_X1 U45 ( .A1(n91), .A2(n24), .ZN(n38) );
  AOI22_X1 U46 ( .A1(n92), .A2(n52), .B1(n58), .B2(n93), .ZN(n68) );
  INV_X1 U47 ( .A(n94), .ZN(n92) );
  OAI211_X1 U48 ( .C1(n95), .C2(n96), .A(n27), .B(n73), .ZN(N394) );
  INV_X1 U49 ( .A(n97), .ZN(n73) );
  OAI21_X1 U50 ( .B1(n64), .B2(n98), .A(n99), .ZN(n97) );
  AOI22_X1 U51 ( .A1(n100), .A2(n45), .B1(n93), .B2(IR_IN_30), .ZN(n95) );
  NOR2_X1 U52 ( .A1(IR_IN_30), .A2(n101), .ZN(n100) );
  NAND4_X1 U53 ( .A1(n42), .A2(n27), .A3(n102), .A4(n103), .ZN(N393) );
  AOI211_X1 U54 ( .C1(n104), .C2(n57), .A(n105), .B(n106), .ZN(n103) );
  NAND2_X1 U55 ( .A1(n77), .A2(n13), .ZN(n105) );
  AOI21_X1 U56 ( .B1(n46), .B2(n107), .A(n108), .ZN(n102) );
  INV_X1 U57 ( .A(n14), .ZN(n108) );
  AOI211_X1 U58 ( .C1(n57), .C2(n58), .A(n109), .B(n53), .ZN(n14) );
  NAND2_X1 U59 ( .A1(n99), .A2(n110), .ZN(n53) );
  OR3_X1 U60 ( .A1(n111), .A2(n112), .A3(n94), .ZN(n110) );
  NAND3_X1 U61 ( .A1(n113), .A2(n114), .A3(n93), .ZN(n99) );
  AOI21_X1 U62 ( .B1(n76), .B2(n115), .A(n64), .ZN(n109) );
  NAND2_X1 U63 ( .A1(n12), .A2(n116), .ZN(n57) );
  NAND4_X1 U64 ( .A1(n101), .A2(n49), .A3(n67), .A4(n117), .ZN(n107) );
  INV_X1 U65 ( .A(n24), .ZN(n117) );
  INV_X1 U66 ( .A(n34), .ZN(n67) );
  NAND2_X1 U67 ( .A1(n81), .A2(n118), .ZN(n34) );
  NAND3_X1 U68 ( .A1(n119), .A2(IR_IN[3]), .A3(n120), .ZN(n118) );
  NAND3_X1 U69 ( .A1(n90), .A2(IR_IN[3]), .A3(n119), .ZN(n81) );
  AOI21_X1 U70 ( .B1(n121), .B2(n91), .A(n35), .ZN(n49) );
  NAND2_X1 U71 ( .A1(n85), .A2(n66), .ZN(n35) );
  OAI21_X1 U72 ( .B1(n120), .B2(n88), .A(n24), .ZN(n66) );
  NOR4_X1 U73 ( .A1(n122), .A2(n123), .A3(IR_IN[2]), .A4(IR_IN[4]), .ZN(n24)
         );
  NAND3_X1 U74 ( .A1(IR_IN[1]), .A2(IR_IN[0]), .A3(n86), .ZN(n85) );
  AND4_X1 U75 ( .A1(n65), .A2(n40), .A3(n37), .A4(n21), .ZN(n101) );
  NAND3_X1 U76 ( .A1(n124), .A2(n125), .A3(n88), .ZN(n21) );
  NAND2_X1 U77 ( .A1(n91), .A2(IR_IN[0]), .ZN(n37) );
  NAND2_X1 U78 ( .A1(n89), .A2(n88), .ZN(n40) );
  AOI211_X1 U79 ( .C1(n121), .C2(n86), .A(n126), .B(n127), .ZN(n65) );
  OAI21_X1 U80 ( .B1(n128), .B2(n39), .A(n23), .ZN(n127) );
  AND2_X1 U81 ( .A1(n84), .A2(n129), .ZN(n23) );
  NAND4_X1 U82 ( .A1(n124), .A2(IR_IN[1]), .A3(IR_IN[0]), .A4(n125), .ZN(n129)
         );
  NAND3_X1 U83 ( .A1(n90), .A2(n124), .A3(IR_IN[2]), .ZN(n84) );
  AND3_X1 U84 ( .A1(IR_IN[5]), .A2(IR_IN[3]), .A3(IR_IN[4]), .ZN(n124) );
  INV_X1 U85 ( .A(n91), .ZN(n128) );
  NOR4_X1 U86 ( .A1(n122), .A2(IR_IN[2]), .A3(IR_IN[3]), .A4(IR_IN[4]), .ZN(
        n91) );
  INV_X1 U87 ( .A(n50), .ZN(n126) );
  OAI21_X1 U88 ( .B1(n120), .B2(n90), .A(n89), .ZN(n50) );
  AND2_X1 U89 ( .A1(n119), .A2(n123), .ZN(n89) );
  INV_X1 U90 ( .A(IR_IN[3]), .ZN(n123) );
  NOR3_X1 U91 ( .A1(n122), .A2(IR_IN[4]), .A3(n125), .ZN(n119) );
  INV_X1 U92 ( .A(IR_IN[5]), .ZN(n122) );
  INV_X1 U93 ( .A(n39), .ZN(n90) );
  NAND2_X1 U94 ( .A1(IR_IN[0]), .A2(n130), .ZN(n39) );
  NOR4_X1 U95 ( .A1(n125), .A2(IR_IN[3]), .A3(IR_IN[4]), .A4(IR_IN[5]), .ZN(
        n86) );
  INV_X1 U96 ( .A(IR_IN[2]), .ZN(n125) );
  OR2_X1 U97 ( .A1(n88), .A2(n120), .ZN(n121) );
  NOR2_X1 U98 ( .A1(IR_IN[0]), .A2(IR_IN[1]), .ZN(n120) );
  NOR2_X1 U99 ( .A1(n130), .A2(IR_IN[0]), .ZN(n88) );
  INV_X1 U100 ( .A(IR_IN[1]), .ZN(n130) );
  INV_X1 U101 ( .A(n17), .ZN(n46) );
  NAND4_X1 U102 ( .A1(n104), .A2(n45), .A3(n131), .A4(n132), .ZN(n17) );
  NOR4_X1 U103 ( .A1(IR_IN_30), .A2(IR_IN[9]), .A3(IR_IN[8]), .A4(IR_IN[7]), 
        .ZN(n132) );
  NOR2_X1 U104 ( .A1(IR_IN[6]), .A2(IR_IN[10]), .ZN(n131) );
  INV_X1 U105 ( .A(n96), .ZN(n104) );
  NAND3_X1 U106 ( .A1(n133), .A2(n111), .A3(n114), .ZN(n96) );
  AND4_X1 U107 ( .A1(n134), .A2(n19), .A3(n135), .A4(n136), .ZN(n27) );
  AOI211_X1 U108 ( .C1(n106), .C2(n52), .A(n71), .B(n30), .ZN(n136) );
  OAI22_X1 U109 ( .A1(n12), .A2(n63), .B1(n137), .B2(n77), .ZN(n30) );
  NOR2_X1 U110 ( .A1(n52), .A2(n59), .ZN(n137) );
  INV_X1 U111 ( .A(n44), .ZN(n63) );
  NOR2_X1 U112 ( .A1(n76), .A2(n133), .ZN(n44) );
  OAI21_X1 U113 ( .B1(n116), .B2(n98), .A(n20), .ZN(n71) );
  NAND3_X1 U114 ( .A1(n52), .A2(n113), .A3(IR_IN_28), .ZN(n20) );
  INV_X1 U115 ( .A(n98), .ZN(n106) );
  OAI21_X1 U116 ( .B1(n93), .B2(n45), .A(n138), .ZN(n135) );
  INV_X1 U117 ( .A(n116), .ZN(n93) );
  NAND3_X1 U118 ( .A1(n59), .A2(n114), .A3(n113), .ZN(n19) );
  NOR3_X1 U119 ( .A1(n139), .A2(n133), .A3(n111), .ZN(n113) );
  INV_X1 U120 ( .A(n48), .ZN(n134) );
  NOR3_X1 U121 ( .A1(n12), .A2(IR_IN_29), .A3(n76), .ZN(n48) );
  NAND3_X1 U122 ( .A1(n114), .A2(n139), .A3(IR_IN_31), .ZN(n76) );
  AOI211_X1 U123 ( .C1(n59), .C2(n138), .A(n140), .B(n31), .ZN(n42) );
  OAI222_X1 U124 ( .A1(n116), .A2(n77), .B1(n112), .B2(n94), .C1(n64), .C2(n98), .ZN(n31) );
  NAND3_X1 U125 ( .A1(IR_IN_28), .A2(n139), .A3(n141), .ZN(n98) );
  INV_X1 U126 ( .A(n45), .ZN(n64) );
  NAND3_X1 U127 ( .A1(n133), .A2(n139), .A3(IR_IN_28), .ZN(n94) );
  NOR2_X1 U128 ( .A1(n45), .A2(n52), .ZN(n112) );
  NAND3_X1 U129 ( .A1(n114), .A2(n139), .A3(n141), .ZN(n77) );
  INV_X1 U130 ( .A(IR_IN_30), .ZN(n139) );
  NAND2_X1 U131 ( .A1(IR_IN_27), .A2(n142), .ZN(n116) );
  INV_X1 U132 ( .A(n26), .ZN(n140) );
  AOI211_X1 U133 ( .C1(n52), .C2(n58), .A(n79), .B(n61), .ZN(n26) );
  AND4_X1 U134 ( .A1(n141), .A2(IR_IN_28), .A3(n52), .A4(IR_IN_30), .ZN(n61)
         );
  AND4_X1 U135 ( .A1(n45), .A2(n141), .A3(IR_IN_28), .A4(IR_IN_30), .ZN(n79)
         );
  NOR2_X1 U136 ( .A1(IR_IN_26), .A2(IR_IN_27), .ZN(n45) );
  INV_X1 U137 ( .A(n115), .ZN(n58) );
  NAND3_X1 U138 ( .A1(IR_IN_30), .A2(n114), .A3(n141), .ZN(n115) );
  NOR2_X1 U139 ( .A1(n133), .A2(IR_IN_31), .ZN(n141) );
  INV_X1 U140 ( .A(IR_IN_28), .ZN(n114) );
  NOR2_X1 U141 ( .A1(n142), .A2(IR_IN_27), .ZN(n52) );
  INV_X1 U142 ( .A(IR_IN_26), .ZN(n142) );
  INV_X1 U143 ( .A(n13), .ZN(n138) );
  NAND4_X1 U144 ( .A1(IR_IN_28), .A2(IR_IN_30), .A3(n133), .A4(n111), .ZN(n13)
         );
  INV_X1 U145 ( .A(IR_IN_31), .ZN(n111) );
  INV_X1 U146 ( .A(IR_IN_29), .ZN(n133) );
  INV_X1 U147 ( .A(n12), .ZN(n59) );
  NAND2_X1 U148 ( .A1(IR_IN_27), .A2(IR_IN_26), .ZN(n12) );
  DFF_X1 signed_unsigned_1_reg ( .D(n150), .CK(Clk), .QN(n10) );
  INV_X1 U9 ( .A(n3), .ZN(n1) );
  INV_X4 U164 ( .A(n1), .ZN(lhi_sel) );
endmodule


module regFFD_NBIT32_0 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96;

  DFFR_X1 \Q_reg[31]  ( .D(n96), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n64) );
  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n63) );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n62) );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n61) );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n60) );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n59) );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n58) );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n57) );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n56) );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n55) );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n54) );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n53) );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n52) );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n51) );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n50) );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n49) );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n48) );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n47) );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n46) );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n45) );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n44) );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n43) );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n42) );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n41) );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n40) );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n39) );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n38) );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n37) );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n36) );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n35) );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n34) );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n33) );
  OAI21_X1 U2 ( .B1(n33), .B2(ENABLE), .A(n1), .ZN(n65) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n34), .B2(ENABLE), .A(n2), .ZN(n66) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n2) );
  OAI21_X1 U6 ( .B1(n35), .B2(ENABLE), .A(n3), .ZN(n67) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n3) );
  OAI21_X1 U8 ( .B1(n36), .B2(ENABLE), .A(n4), .ZN(n68) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n4) );
  OAI21_X1 U10 ( .B1(n37), .B2(ENABLE), .A(n5), .ZN(n69) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n5) );
  OAI21_X1 U12 ( .B1(n38), .B2(ENABLE), .A(n6), .ZN(n70) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n6) );
  OAI21_X1 U14 ( .B1(n39), .B2(ENABLE), .A(n7), .ZN(n71) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n7) );
  OAI21_X1 U16 ( .B1(n40), .B2(ENABLE), .A(n8), .ZN(n72) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n8) );
  OAI21_X1 U18 ( .B1(n41), .B2(ENABLE), .A(n9), .ZN(n73) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n9) );
  OAI21_X1 U20 ( .B1(n42), .B2(ENABLE), .A(n10), .ZN(n74) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n10) );
  OAI21_X1 U22 ( .B1(n43), .B2(ENABLE), .A(n11), .ZN(n75) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n11) );
  OAI21_X1 U24 ( .B1(n44), .B2(ENABLE), .A(n12), .ZN(n76) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n12) );
  OAI21_X1 U26 ( .B1(n45), .B2(ENABLE), .A(n13), .ZN(n77) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n13) );
  OAI21_X1 U28 ( .B1(n46), .B2(ENABLE), .A(n14), .ZN(n78) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n14) );
  OAI21_X1 U30 ( .B1(n47), .B2(ENABLE), .A(n15), .ZN(n79) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n15) );
  OAI21_X1 U32 ( .B1(n48), .B2(ENABLE), .A(n16), .ZN(n80) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n16) );
  OAI21_X1 U34 ( .B1(n49), .B2(ENABLE), .A(n17), .ZN(n81) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n17) );
  OAI21_X1 U36 ( .B1(n50), .B2(ENABLE), .A(n18), .ZN(n82) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n18) );
  OAI21_X1 U38 ( .B1(n51), .B2(ENABLE), .A(n19), .ZN(n83) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n19) );
  OAI21_X1 U40 ( .B1(n52), .B2(ENABLE), .A(n20), .ZN(n84) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n20) );
  OAI21_X1 U42 ( .B1(n53), .B2(ENABLE), .A(n21), .ZN(n85) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n21) );
  OAI21_X1 U44 ( .B1(n54), .B2(ENABLE), .A(n22), .ZN(n86) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n22) );
  OAI21_X1 U46 ( .B1(n55), .B2(ENABLE), .A(n23), .ZN(n87) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n23) );
  OAI21_X1 U48 ( .B1(n56), .B2(ENABLE), .A(n24), .ZN(n88) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n24) );
  OAI21_X1 U50 ( .B1(n57), .B2(ENABLE), .A(n25), .ZN(n89) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n25) );
  OAI21_X1 U52 ( .B1(n58), .B2(ENABLE), .A(n26), .ZN(n90) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n26) );
  OAI21_X1 U54 ( .B1(n59), .B2(ENABLE), .A(n27), .ZN(n91) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n27) );
  OAI21_X1 U56 ( .B1(n60), .B2(ENABLE), .A(n28), .ZN(n92) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n28) );
  OAI21_X1 U58 ( .B1(n61), .B2(ENABLE), .A(n29), .ZN(n93) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n29) );
  OAI21_X1 U60 ( .B1(n62), .B2(ENABLE), .A(n30), .ZN(n94) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n30) );
  OAI21_X1 U62 ( .B1(n63), .B2(ENABLE), .A(n31), .ZN(n95) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n31) );
  OAI21_X1 U64 ( .B1(n64), .B2(ENABLE), .A(n32), .ZN(n96) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n32) );
endmodule


module regFFD_NBIT32_18 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_17 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_767 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_766 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0 UIV ( .A(S), .Y(SB) );
  ND2_0 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_767 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_766 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_255 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_765 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_764 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_763 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_255 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_255 UIV ( .A(S), .Y(SB) );
  ND2_765 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_764 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_763 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_254 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_762 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_761 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_760 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_254 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_254 UIV ( .A(S), .Y(SB) );
  ND2_762 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_761 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_760 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_253 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_759 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_758 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_757 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_253 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_253 UIV ( .A(S), .Y(SB) );
  ND2_759 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_758 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_757 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_252 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_756 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_755 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_754 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_252 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_252 UIV ( .A(S), .Y(SB) );
  ND2_756 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_755 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_754 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_251 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_753 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_752 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_751 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_251 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_251 UIV ( .A(S), .Y(SB) );
  ND2_753 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_752 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_751 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_250 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_750 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_749 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_748 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_250 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_250 UIV ( .A(S), .Y(SB) );
  ND2_750 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_749 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_748 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_249 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_747 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_746 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_745 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_249 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_249 UIV ( .A(S), .Y(SB) );
  ND2_747 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_746 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_745 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_248 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_744 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_743 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_742 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_248 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_248 UIV ( .A(S), .Y(SB) );
  ND2_744 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_743 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_742 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_247 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_741 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_740 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_739 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_247 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_247 UIV ( .A(S), .Y(SB) );
  ND2_741 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_740 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_739 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_246 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_738 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_737 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_736 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_246 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_246 UIV ( .A(S), .Y(SB) );
  ND2_738 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_737 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_736 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_245 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_735 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_734 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_733 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_245 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_245 UIV ( .A(S), .Y(SB) );
  ND2_735 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_734 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_733 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_244 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_732 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_731 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_730 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_244 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_244 UIV ( .A(S), .Y(SB) );
  ND2_732 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_731 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_730 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_243 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_729 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_728 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_727 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_243 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_243 UIV ( .A(S), .Y(SB) );
  ND2_729 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_728 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_727 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_242 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_726 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_725 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_724 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_242 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_242 UIV ( .A(S), .Y(SB) );
  ND2_726 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_725 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_724 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_241 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_723 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_722 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_721 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_241 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_241 UIV ( .A(S), .Y(SB) );
  ND2_723 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_722 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_721 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_240 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_720 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_719 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_718 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_240 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_240 UIV ( .A(S), .Y(SB) );
  ND2_720 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_719 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_718 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_239 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_717 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_716 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_715 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_239 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_239 UIV ( .A(S), .Y(SB) );
  ND2_717 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_716 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_715 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_238 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_714 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_713 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_712 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_238 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_238 UIV ( .A(S), .Y(SB) );
  ND2_714 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_713 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_712 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_237 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_711 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_710 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_709 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_237 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_237 UIV ( .A(S), .Y(SB) );
  ND2_711 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_710 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_709 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_236 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_708 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_707 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_706 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_236 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_236 UIV ( .A(S), .Y(SB) );
  ND2_708 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_707 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_706 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_235 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_705 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_704 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_703 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_235 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_235 UIV ( .A(S), .Y(SB) );
  ND2_705 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_704 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_703 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_234 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_702 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_701 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_700 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_234 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_234 UIV ( .A(S), .Y(SB) );
  ND2_702 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_701 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_700 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_233 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_699 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_698 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_697 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_233 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_233 UIV ( .A(S), .Y(SB) );
  ND2_699 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_698 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_697 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_232 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_696 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_695 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_694 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_232 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_232 UIV ( .A(S), .Y(SB) );
  ND2_696 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_695 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_694 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_231 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_693 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_692 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_691 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_231 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_231 UIV ( .A(S), .Y(SB) );
  ND2_693 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_692 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_691 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_230 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_690 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_689 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_688 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_230 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_230 UIV ( .A(S), .Y(SB) );
  ND2_690 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_689 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_688 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_229 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_687 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_686 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_685 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_229 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_229 UIV ( .A(S), .Y(SB) );
  ND2_687 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_686 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_685 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_228 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_684 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_683 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_682 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_228 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_228 UIV ( .A(S), .Y(SB) );
  ND2_684 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_683 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_682 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_227 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_681 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_680 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_679 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_227 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_227 UIV ( .A(S), .Y(SB) );
  ND2_681 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_680 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_679 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_226 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_678 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_677 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_676 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_226 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_226 UIV ( .A(S), .Y(SB) );
  ND2_678 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_677 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_676 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_225 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_675 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_674 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_673 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_225 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_225 UIV ( .A(S), .Y(SB) );
  ND2_675 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_674 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_673 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_0 gen1_0 ( .A(A[0]), .B(B[0]), .S(n3), .Y(Y[0]) );
  MUX21_255 gen1_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_254 gen1_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_253 gen1_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_252 gen1_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_251 gen1_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_250 gen1_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_249 gen1_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_248 gen1_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_247 gen1_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_246 gen1_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_245 gen1_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_244 gen1_12 ( .A(A[12]), .B(B[12]), .S(n1), .Y(Y[12]) );
  MUX21_243 gen1_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_242 gen1_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_241 gen1_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_240 gen1_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_239 gen1_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_238 gen1_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_237 gen1_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_236 gen1_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_235 gen1_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_234 gen1_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_233 gen1_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_232 gen1_24 ( .A(A[24]), .B(B[24]), .S(n2), .Y(Y[24]) );
  MUX21_231 gen1_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_230 gen1_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_229 gen1_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_228 gen1_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_227 gen1_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_226 gen1_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_225 gen1_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  CLKBUF_X3 U1 ( .A(SEL), .Z(n1) );
  CLKBUF_X3 U2 ( .A(SEL), .Z(n2) );
  CLKBUF_X3 U3 ( .A(SEL), .Z(n3) );
endmodule


module regFFD_NBIT32_16 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_15 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_14 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_13 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_12 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_11 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n163) );
  OAI21_X1 U2 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U4 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U6 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U8 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U10 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U12 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U14 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U16 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U18 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U20 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U22 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U24 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U26 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U28 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U30 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U32 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U34 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U36 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U38 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U40 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U42 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U44 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U46 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U48 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U50 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U52 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U54 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U56 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U58 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U60 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U62 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U64 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
  SDFFR_X1 \Q_reg[31]  ( .D(1'b1), .SI(1'b0), .SE(n97), .CK(CK), .RN(RESET), 
        .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n135) );
  INV_X1 U66 ( .A(n100), .ZN(n97) );
endmodule


module sign_eval_N_in5_N_out32 ( IR_out, signed_val, Immediate );
  input [4:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   Immediate_31, n1;
  assign Immediate[5] = Immediate_31;
  assign Immediate[6] = Immediate_31;
  assign Immediate[7] = Immediate_31;
  assign Immediate[8] = Immediate_31;
  assign Immediate[9] = Immediate_31;
  assign Immediate[10] = Immediate_31;
  assign Immediate[11] = Immediate_31;
  assign Immediate[12] = Immediate_31;
  assign Immediate[13] = Immediate_31;
  assign Immediate[14] = Immediate_31;
  assign Immediate[15] = Immediate_31;
  assign Immediate[16] = Immediate_31;
  assign Immediate[17] = Immediate_31;
  assign Immediate[18] = Immediate_31;
  assign Immediate[19] = Immediate_31;
  assign Immediate[20] = Immediate_31;
  assign Immediate[21] = Immediate_31;
  assign Immediate[22] = Immediate_31;
  assign Immediate[23] = Immediate_31;
  assign Immediate[24] = Immediate_31;
  assign Immediate[25] = Immediate_31;
  assign Immediate[26] = Immediate_31;
  assign Immediate[27] = Immediate_31;
  assign Immediate[28] = Immediate_31;
  assign Immediate[29] = Immediate_31;
  assign Immediate[30] = Immediate_31;
  assign Immediate[31] = Immediate_31;
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];

  NOR2_X1 U1 ( .A1(signed_val), .A2(n1), .ZN(Immediate_31) );
  INV_X1 U2 ( .A(IR_out[4]), .ZN(n1) );
endmodule


module sign_eval_N_in16_N_out32 ( IR_out, signed_val, Immediate );
  input [15:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   Immediate_31, n1;
  assign Immediate[16] = Immediate_31;
  assign Immediate[17] = Immediate_31;
  assign Immediate[18] = Immediate_31;
  assign Immediate[19] = Immediate_31;
  assign Immediate[20] = Immediate_31;
  assign Immediate[21] = Immediate_31;
  assign Immediate[22] = Immediate_31;
  assign Immediate[23] = Immediate_31;
  assign Immediate[24] = Immediate_31;
  assign Immediate[25] = Immediate_31;
  assign Immediate[26] = Immediate_31;
  assign Immediate[27] = Immediate_31;
  assign Immediate[28] = Immediate_31;
  assign Immediate[29] = Immediate_31;
  assign Immediate[30] = Immediate_31;
  assign Immediate[31] = Immediate_31;
  assign Immediate[15] = IR_out[15];
  assign Immediate[14] = IR_out[14];
  assign Immediate[13] = IR_out[13];
  assign Immediate[12] = IR_out[12];
  assign Immediate[11] = IR_out[11];
  assign Immediate[10] = IR_out[10];
  assign Immediate[9] = IR_out[9];
  assign Immediate[8] = IR_out[8];
  assign Immediate[7] = IR_out[7];
  assign Immediate[6] = IR_out[6];
  assign Immediate[5] = IR_out[5];
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];

  NOR2_X1 U1 ( .A1(signed_val), .A2(n1), .ZN(Immediate_31) );
  INV_X1 U2 ( .A(IR_out[15]), .ZN(n1) );
endmodule


module sign_eval_N_in26_N_out32 ( IR_out, signed_val, Immediate );
  input [25:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   Immediate_31, n1;
  assign Immediate[26] = Immediate_31;
  assign Immediate[27] = Immediate_31;
  assign Immediate[28] = Immediate_31;
  assign Immediate[29] = Immediate_31;
  assign Immediate[30] = Immediate_31;
  assign Immediate[31] = Immediate_31;
  assign Immediate[25] = IR_out[25];
  assign Immediate[24] = IR_out[24];
  assign Immediate[23] = IR_out[23];
  assign Immediate[22] = IR_out[22];
  assign Immediate[21] = IR_out[21];
  assign Immediate[20] = IR_out[20];
  assign Immediate[19] = IR_out[19];
  assign Immediate[18] = IR_out[18];
  assign Immediate[17] = IR_out[17];
  assign Immediate[16] = IR_out[16];
  assign Immediate[15] = IR_out[15];
  assign Immediate[14] = IR_out[14];
  assign Immediate[13] = IR_out[13];
  assign Immediate[12] = IR_out[12];
  assign Immediate[11] = IR_out[11];
  assign Immediate[10] = IR_out[10];
  assign Immediate[9] = IR_out[9];
  assign Immediate[8] = IR_out[8];
  assign Immediate[7] = IR_out[7];
  assign Immediate[6] = IR_out[6];
  assign Immediate[5] = IR_out[5];
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];

  NOR2_X1 U1 ( .A1(signed_val), .A2(n1), .ZN(Immediate_31) );
  INV_X1 U2 ( .A(IR_out[25]), .ZN(n1) );
endmodule


module IR_DECODE_NBIT32_opBIT6_regBIT5 ( CLK, IR_26, OPCODE, is_signed, RS1, 
        RS2, RD, IMMEDIATE );
  input [25:0] IR_26;
  input [5:0] OPCODE;
  output [4:0] RS1;
  output [4:0] RS2;
  output [4:0] RD;
  output [31:0] IMMEDIATE;
  input CLK, is_signed;
  wire   N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38;
  wire   [31:0] IMMEDIATE_16;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;
  assign N133 = IR_26[21];
  assign N134 = IR_26[22];
  assign N135 = IR_26[23];
  assign N136 = IR_26[24];
  assign N137 = IR_26[25];
  assign N138 = IR_26[16];
  assign N139 = IR_26[17];
  assign N140 = IR_26[18];
  assign N141 = IR_26[19];
  assign N142 = IR_26[20];

  DLH_X1 \RD_reg[4]  ( .G(CLK), .D(N147), .Q(RD[4]) );
  DLH_X1 \RD_reg[3]  ( .G(CLK), .D(N146), .Q(RD[3]) );
  DLH_X1 \RD_reg[2]  ( .G(CLK), .D(N145), .Q(RD[2]) );
  DLH_X1 \RD_reg[1]  ( .G(CLK), .D(N144), .Q(RD[1]) );
  DLH_X1 \RD_reg[0]  ( .G(CLK), .D(N143), .Q(RD[0]) );
  DLH_X1 \IMMEDIATE_reg[31]  ( .G(CLK), .D(n36), .Q(IMMEDIATE[31]) );
  DLH_X1 \IMMEDIATE_reg[30]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[30]) );
  DLH_X1 \IMMEDIATE_reg[29]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[29]) );
  DLH_X1 \IMMEDIATE_reg[28]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[28]) );
  DLH_X1 \IMMEDIATE_reg[27]  ( .G(CLK), .D(n36), .Q(IMMEDIATE[27]) );
  DLH_X1 \IMMEDIATE_reg[26]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[26]) );
  DLH_X1 \IMMEDIATE_reg[25]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[25]) );
  DLH_X1 \IMMEDIATE_reg[24]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[24]) );
  DLH_X1 \IMMEDIATE_reg[23]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[23]) );
  DLH_X1 \IMMEDIATE_reg[22]  ( .G(CLK), .D(n36), .Q(IMMEDIATE[22]) );
  DLH_X1 \IMMEDIATE_reg[21]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[21]) );
  DLH_X1 \IMMEDIATE_reg[20]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[20]) );
  DLH_X1 \IMMEDIATE_reg[19]  ( .G(CLK), .D(n36), .Q(IMMEDIATE[19]) );
  DLH_X1 \IMMEDIATE_reg[18]  ( .G(CLK), .D(n36), .Q(IMMEDIATE[18]) );
  DLH_X1 \IMMEDIATE_reg[17]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[17]) );
  DLH_X1 \IMMEDIATE_reg[16]  ( .G(CLK), .D(n32), .Q(IMMEDIATE[16]) );
  DLH_X1 \IMMEDIATE_reg[15]  ( .G(CLK), .D(N163), .Q(IMMEDIATE[15]) );
  DLH_X1 \IMMEDIATE_reg[14]  ( .G(CLK), .D(N162), .Q(IMMEDIATE[14]) );
  DLH_X1 \IMMEDIATE_reg[13]  ( .G(CLK), .D(N161), .Q(IMMEDIATE[13]) );
  DLH_X1 \IMMEDIATE_reg[12]  ( .G(CLK), .D(N160), .Q(IMMEDIATE[12]) );
  DLH_X1 \IMMEDIATE_reg[11]  ( .G(CLK), .D(N159), .Q(IMMEDIATE[11]) );
  DLH_X1 \IMMEDIATE_reg[10]  ( .G(CLK), .D(N158), .Q(IMMEDIATE[10]) );
  DLH_X1 \IMMEDIATE_reg[9]  ( .G(CLK), .D(N157), .Q(IMMEDIATE[9]) );
  DLH_X1 \IMMEDIATE_reg[8]  ( .G(CLK), .D(N156), .Q(IMMEDIATE[8]) );
  DLH_X1 \IMMEDIATE_reg[7]  ( .G(CLK), .D(N155), .Q(IMMEDIATE[7]) );
  DLH_X1 \IMMEDIATE_reg[6]  ( .G(CLK), .D(N154), .Q(IMMEDIATE[6]) );
  DLH_X1 \IMMEDIATE_reg[5]  ( .G(CLK), .D(N153), .Q(IMMEDIATE[5]) );
  DLH_X1 \IMMEDIATE_reg[4]  ( .G(CLK), .D(N152), .Q(IMMEDIATE[4]) );
  DLH_X1 \IMMEDIATE_reg[3]  ( .G(CLK), .D(N151), .Q(IMMEDIATE[3]) );
  DLH_X1 \IMMEDIATE_reg[2]  ( .G(CLK), .D(N150), .Q(IMMEDIATE[2]) );
  DLH_X1 \IMMEDIATE_reg[1]  ( .G(CLK), .D(N149), .Q(IMMEDIATE[1]) );
  DLH_X1 \IMMEDIATE_reg[0]  ( .G(CLK), .D(N148), .Q(IMMEDIATE[0]) );
  DLH_X1 \RS1_reg[4]  ( .G(CLK), .D(N137), .Q(RS1[4]) );
  DLH_X1 \RS1_reg[3]  ( .G(CLK), .D(N136), .Q(RS1[3]) );
  DLH_X1 \RS1_reg[2]  ( .G(CLK), .D(N135), .Q(RS1[2]) );
  DLH_X1 \RS1_reg[1]  ( .G(CLK), .D(N134), .Q(RS1[1]) );
  DLH_X1 \RS1_reg[0]  ( .G(CLK), .D(N133), .Q(RS1[0]) );
  DLH_X1 \RS2_reg[4]  ( .G(CLK), .D(N142), .Q(RS2[4]) );
  DLH_X1 \RS2_reg[3]  ( .G(CLK), .D(N141), .Q(RS2[3]) );
  DLH_X1 \RS2_reg[2]  ( .G(CLK), .D(N140), .Q(RS2[2]) );
  DLH_X1 \RS2_reg[1]  ( .G(CLK), .D(N139), .Q(RS2[1]) );
  DLH_X1 \RS2_reg[0]  ( .G(CLK), .D(N138), .Q(RS2[0]) );
  sign_eval_N_in5_N_out32 SIGN_EXTENSION_imm5 ( .IR_out(IR_26[15:11]), 
        .signed_val(is_signed) );
  sign_eval_N_in16_N_out32 SIGN_EXTENSION_imm16 ( .IR_out(IR_26[15:0]), 
        .signed_val(is_signed), .Immediate({IMMEDIATE_16[31], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, IMMEDIATE_16[15:0]}) );
  sign_eval_N_in26_N_out32 SIGN_EXTENSION_imm26 ( .IR_out({N137, N136, N135, 
        N134, N133, N142, N141, N140, N139, N138, IR_26[15:0]}), .signed_val(
        1'b0) );
  NAND4_X1 U3 ( .A1(n8), .A2(n21), .A3(n22), .A4(n23), .ZN(n1) );
  NAND4_X1 U4 ( .A1(n8), .A2(n21), .A3(n22), .A4(n23), .ZN(n38) );
  NAND4_X1 U5 ( .A1(n7), .A2(n24), .A3(n25), .A4(n26), .ZN(n2) );
  INV_X1 U6 ( .A(OPCODE[3]), .ZN(n3) );
  AND3_X2 U7 ( .A1(n3), .A2(n28), .A3(n27), .ZN(n8) );
  MUX2_X1 U8 ( .A(IR_26[15]), .B(N142), .S(n4), .Z(N147) );
  NAND4_X1 U9 ( .A1(n8), .A2(n19), .A3(n20), .A4(n23), .ZN(n4) );
  AND3_X1 U10 ( .A1(n11), .A2(n12), .A3(n29), .ZN(n5) );
  AND3_X1 U11 ( .A1(n11), .A2(n12), .A3(n3), .ZN(n7) );
  MUX2_X1 U12 ( .A(IR_26[14]), .B(N141), .S(n35), .Z(N146) );
  AND3_X2 U13 ( .A1(n11), .A2(n29), .A3(n12), .ZN(n6) );
  AND2_X2 U14 ( .A1(n34), .A2(IMMEDIATE_16[31]), .ZN(n32) );
  NAND3_X1 U15 ( .A1(n28), .A2(n13), .A3(n27), .ZN(n9) );
  NAND4_X1 U16 ( .A1(n6), .A2(n24), .A3(n25), .A4(n15), .ZN(n33) );
  NAND4_X1 U17 ( .A1(n6), .A2(n16), .A3(n14), .A4(n15), .ZN(n10) );
  INV_X1 U18 ( .A(OPCODE[5]), .ZN(n11) );
  INV_X1 U19 ( .A(OPCODE[4]), .ZN(n12) );
  INV_X1 U20 ( .A(OPCODE[3]), .ZN(n13) );
  NAND4_X1 U21 ( .A1(n6), .A2(n21), .A3(n14), .A4(n15), .ZN(n34) );
  INV_X1 U22 ( .A(OPCODE[0]), .ZN(n14) );
  INV_X1 U23 ( .A(OPCODE[2]), .ZN(n15) );
  NAND4_X1 U24 ( .A1(n5), .A2(n16), .A3(n17), .A4(n18), .ZN(n35) );
  INV_X1 U25 ( .A(OPCODE[1]), .ZN(n16) );
  INV_X1 U26 ( .A(OPCODE[2]), .ZN(n17) );
  INV_X1 U27 ( .A(OPCODE[0]), .ZN(n18) );
  NAND4_X1 U28 ( .A1(n17), .A2(n19), .A3(n20), .A4(n6), .ZN(n30) );
  INV_X1 U29 ( .A(OPCODE[1]), .ZN(n19) );
  INV_X1 U30 ( .A(OPCODE[0]), .ZN(n20) );
  INV_X1 U31 ( .A(OPCODE[1]), .ZN(n21) );
  INV_X1 U32 ( .A(OPCODE[0]), .ZN(n22) );
  INV_X1 U33 ( .A(OPCODE[2]), .ZN(n23) );
  NAND4_X1 U34 ( .A1(n7), .A2(n24), .A3(n25), .A4(n26), .ZN(n37) );
  INV_X1 U35 ( .A(OPCODE[1]), .ZN(n24) );
  INV_X1 U36 ( .A(OPCODE[0]), .ZN(n25) );
  INV_X1 U37 ( .A(OPCODE[2]), .ZN(n26) );
  INV_X1 U38 ( .A(OPCODE[5]), .ZN(n27) );
  INV_X1 U39 ( .A(OPCODE[4]), .ZN(n28) );
  INV_X1 U40 ( .A(OPCODE[3]), .ZN(n29) );
  MUX2_X1 U41 ( .A(N140), .B(IR_26[13]), .S(n31), .Z(N145) );
  NOR4_X1 U42 ( .A1(n9), .A2(OPCODE[1]), .A3(OPCODE[0]), .A4(OPCODE[2]), .ZN(
        n31) );
  AND2_X1 U43 ( .A1(n33), .A2(IMMEDIATE_16[31]), .ZN(n36) );
  AND2_X1 U44 ( .A1(n1), .A2(IMMEDIATE_16[15]), .ZN(N163) );
  AND2_X1 U45 ( .A1(n10), .A2(IMMEDIATE_16[14]), .ZN(N162) );
  AND2_X1 U46 ( .A1(n33), .A2(IMMEDIATE_16[13]), .ZN(N161) );
  AND2_X1 U47 ( .A1(n1), .A2(IMMEDIATE_16[12]), .ZN(N160) );
  AND2_X1 U48 ( .A1(n38), .A2(IMMEDIATE_16[11]), .ZN(N159) );
  AND2_X1 U49 ( .A1(n1), .A2(IMMEDIATE_16[10]), .ZN(N158) );
  AND2_X1 U50 ( .A1(n10), .A2(IMMEDIATE_16[9]), .ZN(N157) );
  AND2_X1 U51 ( .A1(n1), .A2(IMMEDIATE_16[8]), .ZN(N156) );
  AND2_X1 U52 ( .A1(n38), .A2(IMMEDIATE_16[7]), .ZN(N155) );
  AND2_X1 U53 ( .A1(n30), .A2(IMMEDIATE_16[6]), .ZN(N154) );
  AND2_X1 U54 ( .A1(n30), .A2(IMMEDIATE_16[5]), .ZN(N153) );
  AND2_X1 U55 ( .A1(n38), .A2(IMMEDIATE_16[4]), .ZN(N152) );
  AND2_X1 U56 ( .A1(n38), .A2(IMMEDIATE_16[3]), .ZN(N151) );
  AND2_X1 U57 ( .A1(n10), .A2(IMMEDIATE_16[2]), .ZN(N150) );
  AND2_X1 U58 ( .A1(n10), .A2(IMMEDIATE_16[1]), .ZN(N149) );
  AND2_X1 U59 ( .A1(n30), .A2(IMMEDIATE_16[0]), .ZN(N148) );
  MUX2_X1 U60 ( .A(IR_26[12]), .B(N139), .S(n2), .Z(N144) );
  MUX2_X1 U61 ( .A(IR_26[11]), .B(N138), .S(n37), .Z(N143) );
endmodule


module register_file ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, 
        ADD_RD2, DATAIN, OUT1, OUT2, wr_signal );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR, wr_signal;
  wire   \REGISTERS[2][31] , \REGISTERS[2][30] , \REGISTERS[2][29] ,
         \REGISTERS[2][28] , \REGISTERS[2][27] , \REGISTERS[2][26] ,
         \REGISTERS[2][25] , \REGISTERS[2][24] , \REGISTERS[2][23] ,
         \REGISTERS[2][22] , \REGISTERS[2][21] , \REGISTERS[2][20] ,
         \REGISTERS[2][19] , \REGISTERS[2][18] , \REGISTERS[2][17] ,
         \REGISTERS[2][16] , \REGISTERS[2][15] , \REGISTERS[2][14] ,
         \REGISTERS[2][13] , \REGISTERS[2][12] , \REGISTERS[2][11] ,
         \REGISTERS[2][10] , \REGISTERS[2][9] , \REGISTERS[2][8] ,
         \REGISTERS[2][7] , \REGISTERS[2][6] , \REGISTERS[2][5] ,
         \REGISTERS[2][4] , \REGISTERS[2][3] , \REGISTERS[2][2] ,
         \REGISTERS[2][1] , \REGISTERS[2][0] , \REGISTERS[3][31] ,
         \REGISTERS[3][30] , \REGISTERS[3][29] , \REGISTERS[3][28] ,
         \REGISTERS[3][27] , \REGISTERS[3][26] , \REGISTERS[3][25] ,
         \REGISTERS[3][24] , \REGISTERS[3][23] , \REGISTERS[3][22] ,
         \REGISTERS[3][21] , \REGISTERS[3][20] , \REGISTERS[3][19] ,
         \REGISTERS[3][18] , \REGISTERS[3][17] , \REGISTERS[3][16] ,
         \REGISTERS[3][15] , \REGISTERS[3][14] , \REGISTERS[3][13] ,
         \REGISTERS[3][12] , \REGISTERS[3][11] , \REGISTERS[3][10] ,
         \REGISTERS[3][9] , \REGISTERS[3][8] , \REGISTERS[3][7] ,
         \REGISTERS[3][6] , \REGISTERS[3][5] , \REGISTERS[3][4] ,
         \REGISTERS[3][3] , \REGISTERS[3][2] , \REGISTERS[3][1] ,
         \REGISTERS[3][0] , \REGISTERS[6][31] , \REGISTERS[6][30] ,
         \REGISTERS[6][29] , \REGISTERS[6][28] , \REGISTERS[6][27] ,
         \REGISTERS[6][26] , \REGISTERS[6][25] , \REGISTERS[6][24] ,
         \REGISTERS[6][23] , \REGISTERS[6][22] , \REGISTERS[6][21] ,
         \REGISTERS[6][20] , \REGISTERS[6][19] , \REGISTERS[6][18] ,
         \REGISTERS[6][17] , \REGISTERS[6][16] , \REGISTERS[6][15] ,
         \REGISTERS[6][14] , \REGISTERS[6][13] , \REGISTERS[6][12] ,
         \REGISTERS[6][11] , \REGISTERS[6][10] , \REGISTERS[6][9] ,
         \REGISTERS[6][8] , \REGISTERS[6][7] , \REGISTERS[6][6] ,
         \REGISTERS[6][5] , \REGISTERS[6][4] , \REGISTERS[6][3] ,
         \REGISTERS[6][2] , \REGISTERS[6][1] , \REGISTERS[6][0] ,
         \REGISTERS[7][31] , \REGISTERS[7][30] , \REGISTERS[7][29] ,
         \REGISTERS[7][28] , \REGISTERS[7][27] , \REGISTERS[7][26] ,
         \REGISTERS[7][25] , \REGISTERS[7][24] , \REGISTERS[7][23] ,
         \REGISTERS[7][22] , \REGISTERS[7][21] , \REGISTERS[7][20] ,
         \REGISTERS[7][19] , \REGISTERS[7][18] , \REGISTERS[7][17] ,
         \REGISTERS[7][16] , \REGISTERS[7][15] , \REGISTERS[7][14] ,
         \REGISTERS[7][13] , \REGISTERS[7][12] , \REGISTERS[7][11] ,
         \REGISTERS[7][10] , \REGISTERS[7][9] , \REGISTERS[7][8] ,
         \REGISTERS[7][7] , \REGISTERS[7][6] , \REGISTERS[7][5] ,
         \REGISTERS[7][4] , \REGISTERS[7][3] , \REGISTERS[7][2] ,
         \REGISTERS[7][1] , \REGISTERS[7][0] , \REGISTERS[10][31] ,
         \REGISTERS[10][30] , \REGISTERS[10][29] , \REGISTERS[10][28] ,
         \REGISTERS[10][27] , \REGISTERS[10][26] , \REGISTERS[10][25] ,
         \REGISTERS[10][24] , \REGISTERS[10][23] , \REGISTERS[10][22] ,
         \REGISTERS[10][21] , \REGISTERS[10][20] , \REGISTERS[10][19] ,
         \REGISTERS[10][18] , \REGISTERS[10][17] , \REGISTERS[10][16] ,
         \REGISTERS[10][15] , \REGISTERS[10][14] , \REGISTERS[10][13] ,
         \REGISTERS[10][12] , \REGISTERS[10][11] , \REGISTERS[10][10] ,
         \REGISTERS[10][9] , \REGISTERS[10][8] , \REGISTERS[10][7] ,
         \REGISTERS[10][6] , \REGISTERS[10][5] , \REGISTERS[10][4] ,
         \REGISTERS[10][3] , \REGISTERS[10][2] , \REGISTERS[10][1] ,
         \REGISTERS[10][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[14][31] , \REGISTERS[14][30] , \REGISTERS[14][29] ,
         \REGISTERS[14][28] , \REGISTERS[14][27] , \REGISTERS[14][26] ,
         \REGISTERS[14][25] , \REGISTERS[14][24] , \REGISTERS[14][23] ,
         \REGISTERS[14][22] , \REGISTERS[14][21] , \REGISTERS[14][20] ,
         \REGISTERS[14][19] , \REGISTERS[14][18] , \REGISTERS[14][17] ,
         \REGISTERS[14][16] , \REGISTERS[14][15] , \REGISTERS[14][14] ,
         \REGISTERS[14][13] , \REGISTERS[14][12] , \REGISTERS[14][11] ,
         \REGISTERS[14][10] , \REGISTERS[14][9] , \REGISTERS[14][8] ,
         \REGISTERS[14][7] , \REGISTERS[14][6] , \REGISTERS[14][5] ,
         \REGISTERS[14][4] , \REGISTERS[14][3] , \REGISTERS[14][2] ,
         \REGISTERS[14][1] , \REGISTERS[14][0] , \REGISTERS[15][31] ,
         \REGISTERS[15][30] , \REGISTERS[15][29] , \REGISTERS[15][28] ,
         \REGISTERS[15][27] , \REGISTERS[15][26] , \REGISTERS[15][25] ,
         \REGISTERS[15][24] , \REGISTERS[15][23] , \REGISTERS[15][22] ,
         \REGISTERS[15][21] , \REGISTERS[15][20] , \REGISTERS[15][19] ,
         \REGISTERS[15][18] , \REGISTERS[15][17] , \REGISTERS[15][16] ,
         \REGISTERS[15][15] , \REGISTERS[15][14] , \REGISTERS[15][13] ,
         \REGISTERS[15][12] , \REGISTERS[15][11] , \REGISTERS[15][10] ,
         \REGISTERS[15][9] , \REGISTERS[15][8] , \REGISTERS[15][7] ,
         \REGISTERS[15][6] , \REGISTERS[15][5] , \REGISTERS[15][4] ,
         \REGISTERS[15][3] , \REGISTERS[15][2] , \REGISTERS[15][1] ,
         \REGISTERS[15][0] , \REGISTERS[18][31] , \REGISTERS[18][30] ,
         \REGISTERS[18][29] , \REGISTERS[18][28] , \REGISTERS[18][27] ,
         \REGISTERS[18][26] , \REGISTERS[18][25] , \REGISTERS[18][24] ,
         \REGISTERS[18][23] , \REGISTERS[18][22] , \REGISTERS[18][21] ,
         \REGISTERS[18][20] , \REGISTERS[18][19] , \REGISTERS[18][18] ,
         \REGISTERS[18][17] , \REGISTERS[18][16] , \REGISTERS[18][15] ,
         \REGISTERS[18][14] , \REGISTERS[18][13] , \REGISTERS[18][12] ,
         \REGISTERS[18][11] , \REGISTERS[18][10] , \REGISTERS[18][9] ,
         \REGISTERS[18][8] , \REGISTERS[18][7] , \REGISTERS[18][6] ,
         \REGISTERS[18][5] , \REGISTERS[18][4] , \REGISTERS[18][3] ,
         \REGISTERS[18][2] , \REGISTERS[18][1] , \REGISTERS[18][0] ,
         \REGISTERS[19][31] , \REGISTERS[19][30] , \REGISTERS[19][29] ,
         \REGISTERS[19][28] , \REGISTERS[19][27] , \REGISTERS[19][26] ,
         \REGISTERS[19][25] , \REGISTERS[19][24] , \REGISTERS[19][23] ,
         \REGISTERS[19][22] , \REGISTERS[19][21] , \REGISTERS[19][20] ,
         \REGISTERS[19][19] , \REGISTERS[19][18] , \REGISTERS[19][17] ,
         \REGISTERS[19][16] , \REGISTERS[19][15] , \REGISTERS[19][14] ,
         \REGISTERS[19][13] , \REGISTERS[19][12] , \REGISTERS[19][11] ,
         \REGISTERS[19][10] , \REGISTERS[19][9] , \REGISTERS[19][8] ,
         \REGISTERS[19][7] , \REGISTERS[19][6] , \REGISTERS[19][5] ,
         \REGISTERS[19][4] , \REGISTERS[19][3] , \REGISTERS[19][2] ,
         \REGISTERS[19][1] , \REGISTERS[19][0] , \REGISTERS[22][31] ,
         \REGISTERS[22][30] , \REGISTERS[22][29] , \REGISTERS[22][28] ,
         \REGISTERS[22][27] , \REGISTERS[22][26] , \REGISTERS[22][25] ,
         \REGISTERS[22][24] , \REGISTERS[22][23] , \REGISTERS[22][22] ,
         \REGISTERS[22][21] , \REGISTERS[22][20] , \REGISTERS[22][19] ,
         \REGISTERS[22][18] , \REGISTERS[22][17] , \REGISTERS[22][16] ,
         \REGISTERS[22][15] , \REGISTERS[22][14] , \REGISTERS[22][13] ,
         \REGISTERS[22][12] , \REGISTERS[22][11] , \REGISTERS[22][10] ,
         \REGISTERS[22][9] , \REGISTERS[22][8] , \REGISTERS[22][7] ,
         \REGISTERS[22][6] , \REGISTERS[22][5] , \REGISTERS[22][4] ,
         \REGISTERS[22][3] , \REGISTERS[22][2] , \REGISTERS[22][1] ,
         \REGISTERS[22][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[26][31] , \REGISTERS[26][30] , \REGISTERS[26][29] ,
         \REGISTERS[26][28] , \REGISTERS[26][27] , \REGISTERS[26][26] ,
         \REGISTERS[26][25] , \REGISTERS[26][24] , \REGISTERS[26][23] ,
         \REGISTERS[26][22] , \REGISTERS[26][21] , \REGISTERS[26][20] ,
         \REGISTERS[26][19] , \REGISTERS[26][18] , \REGISTERS[26][17] ,
         \REGISTERS[26][16] , \REGISTERS[26][15] , \REGISTERS[26][14] ,
         \REGISTERS[26][13] , \REGISTERS[26][12] , \REGISTERS[26][11] ,
         \REGISTERS[26][10] , \REGISTERS[26][9] , \REGISTERS[26][8] ,
         \REGISTERS[26][7] , \REGISTERS[26][6] , \REGISTERS[26][5] ,
         \REGISTERS[26][4] , \REGISTERS[26][3] , \REGISTERS[26][2] ,
         \REGISTERS[26][1] , \REGISTERS[26][0] , \REGISTERS[27][31] ,
         \REGISTERS[27][30] , \REGISTERS[27][29] , \REGISTERS[27][28] ,
         \REGISTERS[27][27] , \REGISTERS[27][26] , \REGISTERS[27][25] ,
         \REGISTERS[27][24] , \REGISTERS[27][23] , \REGISTERS[27][22] ,
         \REGISTERS[27][21] , \REGISTERS[27][20] , \REGISTERS[27][19] ,
         \REGISTERS[27][18] , \REGISTERS[27][17] , \REGISTERS[27][16] ,
         \REGISTERS[27][15] , \REGISTERS[27][14] , \REGISTERS[27][13] ,
         \REGISTERS[27][12] , \REGISTERS[27][11] , \REGISTERS[27][10] ,
         \REGISTERS[27][9] , \REGISTERS[27][8] , \REGISTERS[27][7] ,
         \REGISTERS[27][6] , \REGISTERS[27][5] , \REGISTERS[27][4] ,
         \REGISTERS[27][3] , \REGISTERS[27][2] , \REGISTERS[27][1] ,
         \REGISTERS[27][0] , \REGISTERS[28][31] , \REGISTERS[28][30] ,
         \REGISTERS[28][29] , \REGISTERS[28][28] , \REGISTERS[28][27] ,
         \REGISTERS[28][26] , \REGISTERS[28][25] , \REGISTERS[28][24] ,
         \REGISTERS[28][23] , \REGISTERS[28][22] , \REGISTERS[28][21] ,
         \REGISTERS[28][20] , \REGISTERS[28][19] , \REGISTERS[28][18] ,
         \REGISTERS[28][17] , \REGISTERS[28][16] , \REGISTERS[28][15] ,
         \REGISTERS[28][14] , \REGISTERS[28][13] , \REGISTERS[28][12] ,
         \REGISTERS[28][11] , \REGISTERS[28][10] , \REGISTERS[28][9] ,
         \REGISTERS[28][8] , \REGISTERS[28][7] , \REGISTERS[28][6] ,
         \REGISTERS[28][5] , \REGISTERS[28][4] , \REGISTERS[28][3] ,
         \REGISTERS[28][2] , \REGISTERS[28][1] , \REGISTERS[28][0] ,
         \REGISTERS[29][31] , \REGISTERS[29][30] , \REGISTERS[29][29] ,
         \REGISTERS[29][28] , \REGISTERS[29][27] , \REGISTERS[29][26] ,
         \REGISTERS[29][25] , \REGISTERS[29][24] , \REGISTERS[29][23] ,
         \REGISTERS[29][22] , \REGISTERS[29][21] , \REGISTERS[29][20] ,
         \REGISTERS[29][19] , \REGISTERS[29][18] , \REGISTERS[29][17] ,
         \REGISTERS[29][16] , \REGISTERS[29][15] , \REGISTERS[29][14] ,
         \REGISTERS[29][13] , \REGISTERS[29][12] , \REGISTERS[29][11] ,
         \REGISTERS[29][10] , \REGISTERS[29][9] , \REGISTERS[29][8] ,
         \REGISTERS[29][7] , \REGISTERS[29][6] , \REGISTERS[29][5] ,
         \REGISTERS[29][4] , \REGISTERS[29][3] , \REGISTERS[29][2] ,
         \REGISTERS[29][1] , \REGISTERS[29][0] , N286, N287, N288, N289, N290,
         N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301,
         N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312,
         N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323,
         N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334,
         N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345,
         N346, N347, N348, N349, N350, N351, N352, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420;

  DFFR_X1 \REGISTERS_reg[0][31]  ( .D(n3420), .CK(CLK), .RN(RESET), .QN(n1138)
         );
  DFFR_X1 \REGISTERS_reg[0][30]  ( .D(n3419), .CK(CLK), .RN(RESET), .QN(n1137)
         );
  DFFR_X1 \REGISTERS_reg[0][29]  ( .D(n3418), .CK(CLK), .RN(RESET), .QN(n1136)
         );
  DFFR_X1 \REGISTERS_reg[0][28]  ( .D(n3417), .CK(CLK), .RN(RESET), .QN(n1135)
         );
  DFFR_X1 \REGISTERS_reg[0][27]  ( .D(n3416), .CK(CLK), .RN(RESET), .QN(n1134)
         );
  DFFR_X1 \REGISTERS_reg[0][26]  ( .D(n3415), .CK(CLK), .RN(RESET), .QN(n1133)
         );
  DFFR_X1 \REGISTERS_reg[0][25]  ( .D(n3414), .CK(CLK), .RN(RESET), .QN(n1132)
         );
  DFFR_X1 \REGISTERS_reg[0][24]  ( .D(n3413), .CK(CLK), .RN(RESET), .QN(n1131)
         );
  DFFR_X1 \REGISTERS_reg[0][23]  ( .D(n3412), .CK(CLK), .RN(RESET), .QN(n1130)
         );
  DFFR_X1 \REGISTERS_reg[0][22]  ( .D(n3411), .CK(CLK), .RN(RESET), .QN(n1129)
         );
  DFFR_X1 \REGISTERS_reg[0][21]  ( .D(n3410), .CK(CLK), .RN(RESET), .QN(n1128)
         );
  DFFR_X1 \REGISTERS_reg[0][20]  ( .D(n3409), .CK(CLK), .RN(RESET), .QN(n1127)
         );
  DFFR_X1 \REGISTERS_reg[0][19]  ( .D(n3408), .CK(CLK), .RN(RESET), .QN(n1126)
         );
  DFFR_X1 \REGISTERS_reg[0][18]  ( .D(n3407), .CK(CLK), .RN(RESET), .QN(n1125)
         );
  DFFR_X1 \REGISTERS_reg[0][17]  ( .D(n3406), .CK(CLK), .RN(RESET), .QN(n1124)
         );
  DFFR_X1 \REGISTERS_reg[0][16]  ( .D(n3405), .CK(CLK), .RN(RESET), .QN(n1123)
         );
  DFFR_X1 \REGISTERS_reg[0][15]  ( .D(n3404), .CK(CLK), .RN(RESET), .QN(n1122)
         );
  DFFR_X1 \REGISTERS_reg[0][14]  ( .D(n3403), .CK(CLK), .RN(RESET), .QN(n1121)
         );
  DFFR_X1 \REGISTERS_reg[0][13]  ( .D(n3402), .CK(CLK), .RN(RESET), .QN(n1120)
         );
  DFFR_X1 \REGISTERS_reg[0][12]  ( .D(n3401), .CK(CLK), .RN(RESET), .QN(n1119)
         );
  DFFR_X1 \REGISTERS_reg[0][11]  ( .D(n3400), .CK(CLK), .RN(RESET), .QN(n1118)
         );
  DFFR_X1 \REGISTERS_reg[0][10]  ( .D(n3399), .CK(CLK), .RN(RESET), .QN(n1117)
         );
  DFFR_X1 \REGISTERS_reg[0][9]  ( .D(n3398), .CK(CLK), .RN(RESET), .QN(n1116)
         );
  DFFR_X1 \REGISTERS_reg[0][8]  ( .D(n3397), .CK(CLK), .RN(RESET), .QN(n1115)
         );
  DFFR_X1 \REGISTERS_reg[0][7]  ( .D(n3396), .CK(CLK), .RN(RESET), .QN(n1114)
         );
  DFFR_X1 \REGISTERS_reg[0][6]  ( .D(n3395), .CK(CLK), .RN(RESET), .QN(n1113)
         );
  DFFR_X1 \REGISTERS_reg[0][5]  ( .D(n3394), .CK(CLK), .RN(RESET), .QN(n1112)
         );
  DFFR_X1 \REGISTERS_reg[0][4]  ( .D(n3393), .CK(CLK), .RN(RESET), .QN(n1111)
         );
  DFFR_X1 \REGISTERS_reg[0][3]  ( .D(n3392), .CK(CLK), .RN(RESET), .QN(n1110)
         );
  DFFR_X1 \REGISTERS_reg[0][2]  ( .D(n3391), .CK(CLK), .RN(RESET), .QN(n1109)
         );
  DFFR_X1 \REGISTERS_reg[0][1]  ( .D(n3390), .CK(CLK), .RN(RESET), .QN(n1108)
         );
  DFFR_X1 \REGISTERS_reg[0][0]  ( .D(n3389), .CK(CLK), .RN(RESET), .QN(n1107)
         );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n3388), .CK(CLK), .RN(RESET), .QN(n1104)
         );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n3387), .CK(CLK), .RN(RESET), .QN(n1103)
         );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n3386), .CK(CLK), .RN(RESET), .QN(n1102)
         );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n3385), .CK(CLK), .RN(RESET), .QN(n1101)
         );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n3384), .CK(CLK), .RN(RESET), .QN(n1100)
         );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n3383), .CK(CLK), .RN(RESET), .QN(n1099)
         );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n3382), .CK(CLK), .RN(RESET), .QN(n1098)
         );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n3381), .CK(CLK), .RN(RESET), .QN(n1097)
         );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n3380), .CK(CLK), .RN(RESET), .QN(n1096)
         );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n3379), .CK(CLK), .RN(RESET), .QN(n1095)
         );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n3378), .CK(CLK), .RN(RESET), .QN(n1094)
         );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n3377), .CK(CLK), .RN(RESET), .QN(n1093)
         );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n3376), .CK(CLK), .RN(RESET), .QN(n1092)
         );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n3375), .CK(CLK), .RN(RESET), .QN(n1091)
         );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n3374), .CK(CLK), .RN(RESET), .QN(n1090)
         );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n3373), .CK(CLK), .RN(RESET), .QN(n1089)
         );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n3372), .CK(CLK), .RN(RESET), .QN(n1088)
         );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n3371), .CK(CLK), .RN(RESET), .QN(n1087)
         );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n3370), .CK(CLK), .RN(RESET), .QN(n1086)
         );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n3369), .CK(CLK), .RN(RESET), .QN(n1085)
         );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n3368), .CK(CLK), .RN(RESET), .QN(n1084)
         );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n3367), .CK(CLK), .RN(RESET), .QN(n1083)
         );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n3366), .CK(CLK), .RN(RESET), .QN(n1082)
         );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n3365), .CK(CLK), .RN(RESET), .QN(n1081)
         );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n3364), .CK(CLK), .RN(RESET), .QN(n1080)
         );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n3363), .CK(CLK), .RN(RESET), .QN(n1079)
         );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n3362), .CK(CLK), .RN(RESET), .QN(n1078)
         );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n3361), .CK(CLK), .RN(RESET), .QN(n1077)
         );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n3360), .CK(CLK), .RN(RESET), .QN(n1076)
         );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n3359), .CK(CLK), .RN(RESET), .QN(n1075)
         );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n3358), .CK(CLK), .RN(RESET), .QN(n1074)
         );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n3357), .CK(CLK), .RN(RESET), .QN(n1073)
         );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n3356), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][31] ) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n3355), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][30] ) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n3354), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][29] ) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n3353), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][28] ) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n3352), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][27] ) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n3351), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][26] ) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n3350), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][25] ) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n3349), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][24] ) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n3348), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][23] ) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n3347), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][22] ) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n3346), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][21] ) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n3345), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][20] ) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n3344), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][19] ) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n3343), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][18] ) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n3342), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][17] ) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n3341), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][16] ) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n3340), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][15] ) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n3339), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][14] ) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n3338), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][13] ) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n3337), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][12] ) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n3336), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][11] ) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n3335), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][10] ) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n3334), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][9] ) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n3333), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][8] ) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n3332), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][7] ) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n3331), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][6] ) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n3330), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][5] ) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n3329), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][4] ) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n3328), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][3] ) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n3327), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][2] ) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n3326), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][1] ) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n3325), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[2][0] ) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n3324), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][31] ) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n3323), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][30] ) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n3322), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][29] ) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n3321), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][28] ) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n3320), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][27] ) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n3319), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][26] ) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n3318), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][25] ) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n3317), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][24] ) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n3316), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][23] ) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n3315), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][22] ) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n3314), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][21] ) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n3313), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][20] ) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n3312), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][19] ) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n3311), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][18] ) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n3310), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][17] ) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n3309), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][16] ) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n3308), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][15] ) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n3307), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][14] ) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n3306), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][13] ) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n3305), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][12] ) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n3304), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][11] ) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n3303), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][10] ) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n3302), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][9] ) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n3301), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][8] ) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n3300), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][7] ) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n3299), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][6] ) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n3298), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][5] ) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n3297), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][4] ) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n3296), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][3] ) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n3295), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][2] ) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n3294), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][1] ) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n3293), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[3][0] ) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n3292), .CK(CLK), .RN(RESET), .QN(n1002)
         );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n3291), .CK(CLK), .RN(RESET), .QN(n1001)
         );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n3290), .CK(CLK), .RN(RESET), .QN(n1000)
         );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n3289), .CK(CLK), .RN(RESET), .QN(n999)
         );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n3288), .CK(CLK), .RN(RESET), .QN(n998)
         );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n3287), .CK(CLK), .RN(RESET), .QN(n997)
         );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n3286), .CK(CLK), .RN(RESET), .QN(n996)
         );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n3285), .CK(CLK), .RN(RESET), .QN(n995)
         );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n3284), .CK(CLK), .RN(RESET), .QN(n994)
         );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n3283), .CK(CLK), .RN(RESET), .QN(n993)
         );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n3282), .CK(CLK), .RN(RESET), .QN(n992)
         );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n3281), .CK(CLK), .RN(RESET), .QN(n991)
         );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n3280), .CK(CLK), .RN(RESET), .QN(n990)
         );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n3279), .CK(CLK), .RN(RESET), .QN(n989)
         );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n3278), .CK(CLK), .RN(RESET), .QN(n988)
         );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n3277), .CK(CLK), .RN(RESET), .QN(n987)
         );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n3276), .CK(CLK), .RN(RESET), .QN(n986)
         );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n3275), .CK(CLK), .RN(RESET), .QN(n985)
         );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n3274), .CK(CLK), .RN(RESET), .QN(n984)
         );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n3273), .CK(CLK), .RN(RESET), .QN(n983)
         );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n3272), .CK(CLK), .RN(RESET), .QN(n982)
         );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n3271), .CK(CLK), .RN(RESET), .QN(n981)
         );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n3270), .CK(CLK), .RN(RESET), .QN(n980)
         );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n3269), .CK(CLK), .RN(RESET), .QN(n979)
         );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n3268), .CK(CLK), .RN(RESET), .QN(n978)
         );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n3267), .CK(CLK), .RN(RESET), .QN(n977)
         );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n3266), .CK(CLK), .RN(RESET), .QN(n976)
         );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n3265), .CK(CLK), .RN(RESET), .QN(n975)
         );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n3264), .CK(CLK), .RN(RESET), .QN(n974)
         );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n3263), .CK(CLK), .RN(RESET), .QN(n973)
         );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n3262), .CK(CLK), .RN(RESET), .QN(n972)
         );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n3261), .CK(CLK), .RN(RESET), .QN(n971)
         );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n3260), .CK(CLK), .RN(RESET), .QN(n968)
         );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n3259), .CK(CLK), .RN(RESET), .QN(n967)
         );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n3258), .CK(CLK), .RN(RESET), .QN(n966)
         );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n3257), .CK(CLK), .RN(RESET), .QN(n965)
         );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n3256), .CK(CLK), .RN(RESET), .QN(n964)
         );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n3255), .CK(CLK), .RN(RESET), .QN(n963)
         );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n3254), .CK(CLK), .RN(RESET), .QN(n962)
         );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n3253), .CK(CLK), .RN(RESET), .QN(n961)
         );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n3252), .CK(CLK), .RN(RESET), .QN(n960)
         );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n3251), .CK(CLK), .RN(RESET), .QN(n959)
         );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n3250), .CK(CLK), .RN(RESET), .QN(n958)
         );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n3249), .CK(CLK), .RN(RESET), .QN(n957)
         );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n3248), .CK(CLK), .RN(RESET), .QN(n956)
         );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n3247), .CK(CLK), .RN(RESET), .QN(n955)
         );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n3246), .CK(CLK), .RN(RESET), .QN(n954)
         );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n3245), .CK(CLK), .RN(RESET), .QN(n953)
         );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n3244), .CK(CLK), .RN(RESET), .QN(n952)
         );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n3243), .CK(CLK), .RN(RESET), .QN(n951)
         );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n3242), .CK(CLK), .RN(RESET), .QN(n950)
         );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n3241), .CK(CLK), .RN(RESET), .QN(n949)
         );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n3240), .CK(CLK), .RN(RESET), .QN(n948)
         );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n3239), .CK(CLK), .RN(RESET), .QN(n947)
         );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n3238), .CK(CLK), .RN(RESET), .QN(n946)
         );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n3237), .CK(CLK), .RN(RESET), .QN(n945)
         );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n3236), .CK(CLK), .RN(RESET), .QN(n944)
         );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n3235), .CK(CLK), .RN(RESET), .QN(n943)
         );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n3234), .CK(CLK), .RN(RESET), .QN(n942)
         );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n3233), .CK(CLK), .RN(RESET), .QN(n941)
         );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n3232), .CK(CLK), .RN(RESET), .QN(n940)
         );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n3231), .CK(CLK), .RN(RESET), .QN(n939)
         );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n3230), .CK(CLK), .RN(RESET), .QN(n938)
         );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n3229), .CK(CLK), .RN(RESET), .QN(n937)
         );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n3228), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][31] ) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n3227), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][30] ) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n3226), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][29] ) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n3225), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][28] ) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n3224), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][27] ) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n3223), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][26] ) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n3222), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][25] ) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n3221), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][24] ) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n3220), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][23] ) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n3219), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][22] ) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n3218), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][21] ) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n3217), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][20] ) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n3216), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][19] ) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n3215), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][18] ) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n3214), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][17] ) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n3213), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][16] ) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n3212), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][15] ) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n3211), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][14] ) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n3210), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][13] ) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n3209), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][12] ) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n3208), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][11] ) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n3207), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][10] ) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n3206), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][9] ) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n3205), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][8] ) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n3204), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][7] ) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n3203), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][6] ) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n3202), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][5] ) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n3201), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][4] ) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n3200), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][3] ) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n3199), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][2] ) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n3198), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][1] ) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n3197), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[6][0] ) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n3196), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][31] ) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n3195), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][30] ) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n3194), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][29] ) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n3193), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][28] ) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n3192), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][27] ) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n3191), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][26] ) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n3190), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][25] ) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n3189), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][24] ) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n3188), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][23] ) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n3187), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][22] ) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n3186), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][21] ) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n3185), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][20] ) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n3184), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][19] ) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n3183), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][18] ) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n3182), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][17] ) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n3181), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][16] ) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n3180), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][15] ) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n3179), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][14] ) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n3178), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][13] ) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n3177), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][12] ) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n3176), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][11] ) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n3175), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][10] ) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n3174), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][9] ) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n3173), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][8] ) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n3172), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][7] ) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n3171), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][6] ) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n3170), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][5] ) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n3169), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][4] ) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n3168), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][3] ) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n3167), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][2] ) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n3166), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][1] ) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n3165), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[7][0] ) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n3164), .CK(CLK), .RN(RESET), .QN(n861)
         );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n3163), .CK(CLK), .RN(RESET), .QN(n860)
         );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n3162), .CK(CLK), .RN(RESET), .QN(n859)
         );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n3161), .CK(CLK), .RN(RESET), .QN(n858)
         );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n3160), .CK(CLK), .RN(RESET), .QN(n857)
         );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n3159), .CK(CLK), .RN(RESET), .QN(n856)
         );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n3158), .CK(CLK), .RN(RESET), .QN(n855)
         );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n3157), .CK(CLK), .RN(RESET), .QN(n854)
         );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n3156), .CK(CLK), .RN(RESET), .QN(n853)
         );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n3155), .CK(CLK), .RN(RESET), .QN(n852)
         );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n3154), .CK(CLK), .RN(RESET), .QN(n851)
         );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n3153), .CK(CLK), .RN(RESET), .QN(n850)
         );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n3152), .CK(CLK), .RN(RESET), .QN(n849)
         );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n3151), .CK(CLK), .RN(RESET), .QN(n848)
         );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n3150), .CK(CLK), .RN(RESET), .QN(n847)
         );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n3149), .CK(CLK), .RN(RESET), .QN(n846)
         );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n3148), .CK(CLK), .RN(RESET), .QN(n845)
         );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n3147), .CK(CLK), .RN(RESET), .QN(n844)
         );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n3146), .CK(CLK), .RN(RESET), .QN(n843)
         );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n3145), .CK(CLK), .RN(RESET), .QN(n842)
         );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n3144), .CK(CLK), .RN(RESET), .QN(n841)
         );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n3143), .CK(CLK), .RN(RESET), .QN(n840)
         );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n3142), .CK(CLK), .RN(RESET), .QN(n839)
         );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n3141), .CK(CLK), .RN(RESET), .QN(n838)
         );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n3140), .CK(CLK), .RN(RESET), .QN(n837)
         );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n3139), .CK(CLK), .RN(RESET), .QN(n836)
         );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n3138), .CK(CLK), .RN(RESET), .QN(n835)
         );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n3137), .CK(CLK), .RN(RESET), .QN(n834)
         );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n3136), .CK(CLK), .RN(RESET), .QN(n833)
         );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n3135), .CK(CLK), .RN(RESET), .QN(n832)
         );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n3134), .CK(CLK), .RN(RESET), .QN(n831)
         );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n3133), .CK(CLK), .RN(RESET), .QN(n830)
         );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n3132), .CK(CLK), .RN(RESET), .QN(n827)
         );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n3131), .CK(CLK), .RN(RESET), .QN(n826)
         );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n3130), .CK(CLK), .RN(RESET), .QN(n825)
         );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n3129), .CK(CLK), .RN(RESET), .QN(n824)
         );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n3128), .CK(CLK), .RN(RESET), .QN(n823)
         );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n3127), .CK(CLK), .RN(RESET), .QN(n822)
         );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n3126), .CK(CLK), .RN(RESET), .QN(n821)
         );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n3125), .CK(CLK), .RN(RESET), .QN(n820)
         );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n3124), .CK(CLK), .RN(RESET), .QN(n819)
         );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n3123), .CK(CLK), .RN(RESET), .QN(n818)
         );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n3122), .CK(CLK), .RN(RESET), .QN(n817)
         );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n3121), .CK(CLK), .RN(RESET), .QN(n816)
         );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n3120), .CK(CLK), .RN(RESET), .QN(n815)
         );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n3119), .CK(CLK), .RN(RESET), .QN(n814)
         );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n3118), .CK(CLK), .RN(RESET), .QN(n813)
         );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n3117), .CK(CLK), .RN(RESET), .QN(n812)
         );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n3116), .CK(CLK), .RN(RESET), .QN(n811)
         );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n3115), .CK(CLK), .RN(RESET), .QN(n810)
         );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n3114), .CK(CLK), .RN(RESET), .QN(n809)
         );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n3113), .CK(CLK), .RN(RESET), .QN(n808)
         );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n3112), .CK(CLK), .RN(RESET), .QN(n807)
         );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n3111), .CK(CLK), .RN(RESET), .QN(n806)
         );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n3110), .CK(CLK), .RN(RESET), .QN(n805)
         );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n3109), .CK(CLK), .RN(RESET), .QN(n804)
         );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n3108), .CK(CLK), .RN(RESET), .QN(n803)
         );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n3107), .CK(CLK), .RN(RESET), .QN(n802)
         );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n3106), .CK(CLK), .RN(RESET), .QN(n801)
         );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n3105), .CK(CLK), .RN(RESET), .QN(n800)
         );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n3104), .CK(CLK), .RN(RESET), .QN(n799)
         );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n3103), .CK(CLK), .RN(RESET), .QN(n798)
         );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n3102), .CK(CLK), .RN(RESET), .QN(n797)
         );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n3101), .CK(CLK), .RN(RESET), .QN(n796)
         );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n3100), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][31] ) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n3099), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][30] ) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n3098), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][29] ) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n3097), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][28] ) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n3096), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][27] ) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n3095), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][26] ) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n3094), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][25] ) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n3093), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][24] ) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n3092), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][23] ) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n3091), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][22] ) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n3090), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][21] ) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n3089), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][20] ) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n3088), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][19] ) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n3087), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][18] ) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n3086), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][17] ) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n3085), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][16] ) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n3084), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][15] ) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n3083), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][14] ) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n3082), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][13] ) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n3081), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][12] ) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n3080), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][11] ) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n3079), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][10] ) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n3078), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][9] ) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n3077), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][8] ) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n3076), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][7] ) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n3075), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][6] ) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n3074), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][5] ) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n3073), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][4] ) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n3072), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][3] ) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n3071), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][2] ) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n3070), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][1] ) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n3069), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[10][0] ) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n3068), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][31] ) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n3067), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][30] ) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n3066), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][29] ) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n3065), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][28] ) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n3064), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][27] ) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n3063), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][26] ) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n3062), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][25] ) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n3061), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][24] ) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n3060), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][23] ) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n3059), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][22] ) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n3058), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][21] ) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n3057), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][20] ) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n3056), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][19] ) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n3055), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][18] ) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n3054), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][17] ) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n3053), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][16] ) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n3052), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][15] ) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n3051), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][14] ) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n3050), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][13] ) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n3049), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][12] ) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n3048), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][11] ) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n3047), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][10] ) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n3046), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][9] ) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n3045), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][8] ) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n3044), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][7] ) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n3043), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][6] ) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n3042), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][5] ) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n3041), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][4] ) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n3040), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][3] ) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n3039), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][2] ) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n3038), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][1] ) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n3037), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[11][0] ) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n3036), .CK(CLK), .RN(RESET), .QN(n725)
         );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n3035), .CK(CLK), .RN(RESET), .QN(n724)
         );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n3034), .CK(CLK), .RN(RESET), .QN(n723)
         );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n3033), .CK(CLK), .RN(RESET), .QN(n722)
         );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n3032), .CK(CLK), .RN(RESET), .QN(n721)
         );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n3031), .CK(CLK), .RN(RESET), .QN(n720)
         );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n3030), .CK(CLK), .RN(RESET), .QN(n719)
         );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n3029), .CK(CLK), .RN(RESET), .QN(n718)
         );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n3028), .CK(CLK), .RN(RESET), .QN(n717)
         );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n3027), .CK(CLK), .RN(RESET), .QN(n716)
         );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n3026), .CK(CLK), .RN(RESET), .QN(n715)
         );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n3025), .CK(CLK), .RN(RESET), .QN(n714)
         );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n3024), .CK(CLK), .RN(RESET), .QN(n713)
         );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n3023), .CK(CLK), .RN(RESET), .QN(n712)
         );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n3022), .CK(CLK), .RN(RESET), .QN(n711)
         );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n3021), .CK(CLK), .RN(RESET), .QN(n710)
         );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n3020), .CK(CLK), .RN(RESET), .QN(n709)
         );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n3019), .CK(CLK), .RN(RESET), .QN(n708)
         );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n3018), .CK(CLK), .RN(RESET), .QN(n707)
         );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n3017), .CK(CLK), .RN(RESET), .QN(n706)
         );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n3016), .CK(CLK), .RN(RESET), .QN(n705)
         );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n3015), .CK(CLK), .RN(RESET), .QN(n704)
         );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n3014), .CK(CLK), .RN(RESET), .QN(n703)
         );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n3013), .CK(CLK), .RN(RESET), .QN(n702)
         );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n3012), .CK(CLK), .RN(RESET), .QN(n701)
         );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n3011), .CK(CLK), .RN(RESET), .QN(n700)
         );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n3010), .CK(CLK), .RN(RESET), .QN(n699)
         );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n3009), .CK(CLK), .RN(RESET), .QN(n698)
         );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n3008), .CK(CLK), .RN(RESET), .QN(n697)
         );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n3007), .CK(CLK), .RN(RESET), .QN(n696)
         );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n3006), .CK(CLK), .RN(RESET), .QN(n695)
         );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n3005), .CK(CLK), .RN(RESET), .QN(n694)
         );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n3004), .CK(CLK), .RN(RESET), .QN(n691)
         );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n3003), .CK(CLK), .RN(RESET), .QN(n690)
         );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n3002), .CK(CLK), .RN(RESET), .QN(n689)
         );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n3001), .CK(CLK), .RN(RESET), .QN(n688)
         );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n3000), .CK(CLK), .RN(RESET), .QN(n687)
         );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n2999), .CK(CLK), .RN(RESET), .QN(n686)
         );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n2998), .CK(CLK), .RN(RESET), .QN(n685)
         );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n2997), .CK(CLK), .RN(RESET), .QN(n684)
         );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n2996), .CK(CLK), .RN(RESET), .QN(n683)
         );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n2995), .CK(CLK), .RN(RESET), .QN(n682)
         );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n2994), .CK(CLK), .RN(RESET), .QN(n681)
         );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n2993), .CK(CLK), .RN(RESET), .QN(n680)
         );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n2992), .CK(CLK), .RN(RESET), .QN(n679)
         );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n2991), .CK(CLK), .RN(RESET), .QN(n678)
         );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n2990), .CK(CLK), .RN(RESET), .QN(n677)
         );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n2989), .CK(CLK), .RN(RESET), .QN(n676)
         );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n2988), .CK(CLK), .RN(RESET), .QN(n675)
         );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n2987), .CK(CLK), .RN(RESET), .QN(n674)
         );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n2986), .CK(CLK), .RN(RESET), .QN(n673)
         );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n2985), .CK(CLK), .RN(RESET), .QN(n672)
         );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n2984), .CK(CLK), .RN(RESET), .QN(n671)
         );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n2983), .CK(CLK), .RN(RESET), .QN(n670)
         );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n2982), .CK(CLK), .RN(RESET), .QN(n669)
         );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n2981), .CK(CLK), .RN(RESET), .QN(n668)
         );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n2980), .CK(CLK), .RN(RESET), .QN(n667)
         );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n2979), .CK(CLK), .RN(RESET), .QN(n666)
         );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n2978), .CK(CLK), .RN(RESET), .QN(n665)
         );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n2977), .CK(CLK), .RN(RESET), .QN(n664)
         );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n2976), .CK(CLK), .RN(RESET), .QN(n663)
         );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n2975), .CK(CLK), .RN(RESET), .QN(n662)
         );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n2974), .CK(CLK), .RN(RESET), .QN(n661)
         );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n2973), .CK(CLK), .RN(RESET), .QN(n660)
         );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n2972), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][31] ) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n2971), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][30] ) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n2970), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][29] ) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n2969), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][28] ) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n2968), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][27] ) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n2967), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][26] ) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n2966), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][25] ) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n2965), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][24] ) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n2964), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][23] ) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n2963), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][22] ) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n2962), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][21] ) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n2961), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][20] ) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n2960), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][19] ) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n2959), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][18] ) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n2958), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][17] ) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n2957), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][16] ) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n2956), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][15] ) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n2955), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][14] ) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n2954), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][13] ) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n2953), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][12] ) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n2952), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][11] ) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n2951), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][10] ) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n2950), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][9] ) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n2949), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][8] ) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n2948), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][7] ) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n2947), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][6] ) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n2946), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][5] ) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n2945), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][4] ) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n2944), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][3] ) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n2943), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][2] ) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n2942), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][1] ) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n2941), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[14][0] ) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n2940), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][31] ) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n2939), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][30] ) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n2938), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][29] ) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n2937), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][28] ) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n2936), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][27] ) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n2935), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][26] ) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n2934), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][25] ) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n2933), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][24] ) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n2932), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][23] ) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n2931), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][22] ) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n2930), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][21] ) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n2929), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][20] ) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n2928), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][19] ) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n2927), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][18] ) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n2926), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][17] ) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n2925), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][16] ) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n2924), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][15] ) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n2923), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][14] ) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n2922), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][13] ) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n2921), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][12] ) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n2920), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][11] ) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n2919), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][10] ) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n2918), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][9] ) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n2917), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][8] ) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n2916), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][7] ) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n2915), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][6] ) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n2914), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][5] ) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n2913), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][4] ) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n2912), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][3] ) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n2911), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][2] ) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n2910), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][1] ) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n2909), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[15][0] ) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n2908), .CK(CLK), .RN(RESET), .QN(n587)
         );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n2907), .CK(CLK), .RN(RESET), .QN(n586)
         );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n2906), .CK(CLK), .RN(RESET), .QN(n585)
         );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n2905), .CK(CLK), .RN(RESET), .QN(n584)
         );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n2904), .CK(CLK), .RN(RESET), .QN(n583)
         );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n2903), .CK(CLK), .RN(RESET), .QN(n582)
         );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n2902), .CK(CLK), .RN(RESET), .QN(n581)
         );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n2901), .CK(CLK), .RN(RESET), .QN(n580)
         );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n2900), .CK(CLK), .RN(RESET), .QN(n579)
         );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n2899), .CK(CLK), .RN(RESET), .QN(n578)
         );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n2898), .CK(CLK), .RN(RESET), .QN(n577)
         );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n2897), .CK(CLK), .RN(RESET), .QN(n576)
         );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n2896), .CK(CLK), .RN(RESET), .QN(n575)
         );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n2895), .CK(CLK), .RN(RESET), .QN(n574)
         );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n2894), .CK(CLK), .RN(RESET), .QN(n573)
         );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n2893), .CK(CLK), .RN(RESET), .QN(n572)
         );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n2892), .CK(CLK), .RN(RESET), .QN(n571)
         );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n2891), .CK(CLK), .RN(RESET), .QN(n570)
         );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n2890), .CK(CLK), .RN(RESET), .QN(n569)
         );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n2889), .CK(CLK), .RN(RESET), .QN(n568)
         );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n2888), .CK(CLK), .RN(RESET), .QN(n567)
         );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n2887), .CK(CLK), .RN(RESET), .QN(n566)
         );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n2886), .CK(CLK), .RN(RESET), .QN(n565)
         );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n2885), .CK(CLK), .RN(RESET), .QN(n564)
         );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n2884), .CK(CLK), .RN(RESET), .QN(n563)
         );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n2883), .CK(CLK), .RN(RESET), .QN(n562)
         );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n2882), .CK(CLK), .RN(RESET), .QN(n561)
         );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n2881), .CK(CLK), .RN(RESET), .QN(n560)
         );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n2880), .CK(CLK), .RN(RESET), .QN(n559)
         );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n2879), .CK(CLK), .RN(RESET), .QN(n558)
         );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n2878), .CK(CLK), .RN(RESET), .QN(n557)
         );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n2877), .CK(CLK), .RN(RESET), .QN(n556)
         );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n2876), .CK(CLK), .RN(RESET), .QN(n553)
         );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n2875), .CK(CLK), .RN(RESET), .QN(n552)
         );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n2874), .CK(CLK), .RN(RESET), .QN(n551)
         );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n2873), .CK(CLK), .RN(RESET), .QN(n550)
         );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n2872), .CK(CLK), .RN(RESET), .QN(n549)
         );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n2871), .CK(CLK), .RN(RESET), .QN(n548)
         );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n2870), .CK(CLK), .RN(RESET), .QN(n547)
         );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n2869), .CK(CLK), .RN(RESET), .QN(n546)
         );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n2868), .CK(CLK), .RN(RESET), .QN(n545)
         );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n2867), .CK(CLK), .RN(RESET), .QN(n544)
         );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n2866), .CK(CLK), .RN(RESET), .QN(n543)
         );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n2865), .CK(CLK), .RN(RESET), .QN(n542)
         );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n2864), .CK(CLK), .RN(RESET), .QN(n541)
         );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n2863), .CK(CLK), .RN(RESET), .QN(n540)
         );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n2862), .CK(CLK), .RN(RESET), .QN(n539)
         );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n2861), .CK(CLK), .RN(RESET), .QN(n538)
         );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n2860), .CK(CLK), .RN(RESET), .QN(n537)
         );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n2859), .CK(CLK), .RN(RESET), .QN(n536)
         );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n2858), .CK(CLK), .RN(RESET), .QN(n535)
         );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n2857), .CK(CLK), .RN(RESET), .QN(n534)
         );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n2856), .CK(CLK), .RN(RESET), .QN(n533)
         );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n2855), .CK(CLK), .RN(RESET), .QN(n532)
         );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n2854), .CK(CLK), .RN(RESET), .QN(n531)
         );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n2853), .CK(CLK), .RN(RESET), .QN(n530)
         );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n2852), .CK(CLK), .RN(RESET), .QN(n529)
         );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n2851), .CK(CLK), .RN(RESET), .QN(n528)
         );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n2850), .CK(CLK), .RN(RESET), .QN(n527)
         );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n2849), .CK(CLK), .RN(RESET), .QN(n526)
         );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n2848), .CK(CLK), .RN(RESET), .QN(n525)
         );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n2847), .CK(CLK), .RN(RESET), .QN(n524)
         );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n2846), .CK(CLK), .RN(RESET), .QN(n523)
         );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n2845), .CK(CLK), .RN(RESET), .QN(n522)
         );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n2844), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][31] ) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n2843), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][30] ) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n2842), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][29] ) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n2841), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][28] ) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n2840), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][27] ) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n2839), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][26] ) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n2838), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][25] ) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n2837), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][24] ) );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n2836), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][23] ) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n2835), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][22] ) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n2834), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][21] ) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n2833), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][20] ) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n2832), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][19] ) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n2831), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][18] ) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n2830), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][17] ) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n2829), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][16] ) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n2828), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][15] ) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n2827), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][14] ) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n2826), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][13] ) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n2825), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][12] ) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n2824), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][11] ) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n2823), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][10] ) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n2822), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][9] ) );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n2821), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][8] ) );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n2820), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][7] ) );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n2819), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][6] ) );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n2818), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][5] ) );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n2817), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][4] ) );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n2816), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][3] ) );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n2815), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][2] ) );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n2814), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][1] ) );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n2813), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[18][0] ) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n2812), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][31] ) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n2811), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][30] ) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n2810), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][29] ) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n2809), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][28] ) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n2808), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][27] ) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n2807), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][26] ) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n2806), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][25] ) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n2805), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][24] ) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n2804), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][23] ) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n2803), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][22] ) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n2802), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][21] ) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n2801), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][20] ) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n2800), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][19] ) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n2799), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][18] ) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n2798), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][17] ) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n2797), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][16] ) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n2796), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][15] ) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n2795), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][14] ) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n2794), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][13] ) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n2793), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][12] ) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n2792), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][11] ) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n2791), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][10] ) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n2790), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][9] ) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n2789), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][8] ) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n2788), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][7] ) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n2787), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][6] ) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n2786), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][5] ) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n2785), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][4] ) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n2784), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][3] ) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n2783), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][2] ) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n2782), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][1] ) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n2781), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[19][0] ) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n2780), .CK(CLK), .RN(RESET), .QN(n451)
         );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n2779), .CK(CLK), .RN(RESET), .QN(n450)
         );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n2778), .CK(CLK), .RN(RESET), .QN(n449)
         );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n2777), .CK(CLK), .RN(RESET), .QN(n448)
         );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n2776), .CK(CLK), .RN(RESET), .QN(n447)
         );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n2775), .CK(CLK), .RN(RESET), .QN(n446)
         );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n2774), .CK(CLK), .RN(RESET), .QN(n445)
         );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n2773), .CK(CLK), .RN(RESET), .QN(n444)
         );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n2772), .CK(CLK), .RN(RESET), .QN(n443)
         );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n2771), .CK(CLK), .RN(RESET), .QN(n442)
         );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n2770), .CK(CLK), .RN(RESET), .QN(n441)
         );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n2769), .CK(CLK), .RN(RESET), .QN(n440)
         );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n2768), .CK(CLK), .RN(RESET), .QN(n439)
         );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n2767), .CK(CLK), .RN(RESET), .QN(n438)
         );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n2766), .CK(CLK), .RN(RESET), .QN(n437)
         );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n2765), .CK(CLK), .RN(RESET), .QN(n436)
         );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n2764), .CK(CLK), .RN(RESET), .QN(n435)
         );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n2763), .CK(CLK), .RN(RESET), .QN(n434)
         );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n2762), .CK(CLK), .RN(RESET), .QN(n433)
         );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n2761), .CK(CLK), .RN(RESET), .QN(n432)
         );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n2760), .CK(CLK), .RN(RESET), .QN(n431)
         );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n2759), .CK(CLK), .RN(RESET), .QN(n430)
         );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n2758), .CK(CLK), .RN(RESET), .QN(n429)
         );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n2757), .CK(CLK), .RN(RESET), .QN(n428)
         );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n2756), .CK(CLK), .RN(RESET), .QN(n427)
         );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n2755), .CK(CLK), .RN(RESET), .QN(n426)
         );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n2754), .CK(CLK), .RN(RESET), .QN(n425)
         );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n2753), .CK(CLK), .RN(RESET), .QN(n424)
         );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n2752), .CK(CLK), .RN(RESET), .QN(n423)
         );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n2751), .CK(CLK), .RN(RESET), .QN(n422)
         );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n2750), .CK(CLK), .RN(RESET), .QN(n421)
         );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n2749), .CK(CLK), .RN(RESET), .QN(n420)
         );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n2748), .CK(CLK), .RN(RESET), .QN(n417)
         );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n2747), .CK(CLK), .RN(RESET), .QN(n416)
         );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n2746), .CK(CLK), .RN(RESET), .QN(n415)
         );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n2745), .CK(CLK), .RN(RESET), .QN(n414)
         );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n2744), .CK(CLK), .RN(RESET), .QN(n413)
         );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n2743), .CK(CLK), .RN(RESET), .QN(n412)
         );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n2742), .CK(CLK), .RN(RESET), .QN(n411)
         );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n2741), .CK(CLK), .RN(RESET), .QN(n410)
         );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n2740), .CK(CLK), .RN(RESET), .QN(n409)
         );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n2739), .CK(CLK), .RN(RESET), .QN(n408)
         );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n2738), .CK(CLK), .RN(RESET), .QN(n407)
         );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n2737), .CK(CLK), .RN(RESET), .QN(n406)
         );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n2736), .CK(CLK), .RN(RESET), .QN(n405)
         );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n2735), .CK(CLK), .RN(RESET), .QN(n404)
         );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n2734), .CK(CLK), .RN(RESET), .QN(n403)
         );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n2733), .CK(CLK), .RN(RESET), .QN(n402)
         );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n2732), .CK(CLK), .RN(RESET), .QN(n401)
         );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n2731), .CK(CLK), .RN(RESET), .QN(n400)
         );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n2730), .CK(CLK), .RN(RESET), .QN(n399)
         );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n2729), .CK(CLK), .RN(RESET), .QN(n398)
         );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n2728), .CK(CLK), .RN(RESET), .QN(n397)
         );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n2727), .CK(CLK), .RN(RESET), .QN(n396)
         );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n2726), .CK(CLK), .RN(RESET), .QN(n395)
         );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n2725), .CK(CLK), .RN(RESET), .QN(n394)
         );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n2724), .CK(CLK), .RN(RESET), .QN(n393)
         );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n2723), .CK(CLK), .RN(RESET), .QN(n392)
         );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n2722), .CK(CLK), .RN(RESET), .QN(n391)
         );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n2721), .CK(CLK), .RN(RESET), .QN(n390)
         );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n2720), .CK(CLK), .RN(RESET), .QN(n389)
         );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n2719), .CK(CLK), .RN(RESET), .QN(n388)
         );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n2718), .CK(CLK), .RN(RESET), .QN(n387)
         );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n2717), .CK(CLK), .RN(RESET), .QN(n386)
         );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n2716), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][31] ) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n2715), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][30] ) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n2714), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][29] ) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n2713), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][28] ) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n2712), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][27] ) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n2711), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][26] ) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n2710), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][25] ) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n2709), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][24] ) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n2708), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][23] ) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n2707), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][22] ) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n2706), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][21] ) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n2705), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][20] ) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n2704), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][19] ) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n2703), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][18] ) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n2702), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][17] ) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n2701), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][16] ) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n2700), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][15] ) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n2699), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][14] ) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n2698), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][13] ) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n2697), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][12] ) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n2696), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][11] ) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n2695), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][10] ) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n2694), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][9] ) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n2693), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][8] ) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n2692), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][7] ) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n2691), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][6] ) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n2690), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][5] ) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n2689), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][4] ) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n2688), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][3] ) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n2687), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][2] ) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n2686), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][1] ) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n2685), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[22][0] ) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n2684), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][31] ) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n2683), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][30] ) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n2682), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][29] ) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n2681), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][28] ) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n2680), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][27] ) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n2679), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][26] ) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n2678), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][25] ) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n2677), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][24] ) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n2676), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][23] ) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n2675), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][22] ) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n2674), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][21] ) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n2673), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][20] ) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n2672), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][19] ) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n2671), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][18] ) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n2670), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][17] ) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n2669), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][16] ) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n2668), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][15] ) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n2667), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][14] ) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n2666), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][13] ) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n2665), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][12] ) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n2664), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][11] ) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n2663), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][10] ) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n2662), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][9] ) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n2661), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][8] ) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n2660), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][7] ) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n2659), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][6] ) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n2658), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][5] ) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n2657), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][4] ) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n2656), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][3] ) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n2655), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][2] ) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n2654), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][1] ) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n2653), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[23][0] ) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n2652), .CK(CLK), .RN(RESET), .QN(n312)
         );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n2651), .CK(CLK), .RN(RESET), .QN(n311)
         );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n2650), .CK(CLK), .RN(RESET), .QN(n310)
         );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n2649), .CK(CLK), .RN(RESET), .QN(n309)
         );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n2648), .CK(CLK), .RN(RESET), .QN(n308)
         );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n2647), .CK(CLK), .RN(RESET), .QN(n307)
         );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n2646), .CK(CLK), .RN(RESET), .QN(n306)
         );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n2645), .CK(CLK), .RN(RESET), .QN(n305)
         );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n2644), .CK(CLK), .RN(RESET), .QN(n304)
         );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n2643), .CK(CLK), .RN(RESET), .QN(n303)
         );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n2642), .CK(CLK), .RN(RESET), .QN(n302)
         );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n2641), .CK(CLK), .RN(RESET), .QN(n301)
         );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n2640), .CK(CLK), .RN(RESET), .QN(n300)
         );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n2639), .CK(CLK), .RN(RESET), .QN(n299)
         );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n2638), .CK(CLK), .RN(RESET), .QN(n298)
         );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n2637), .CK(CLK), .RN(RESET), .QN(n297)
         );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n2636), .CK(CLK), .RN(RESET), .QN(n296)
         );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n2635), .CK(CLK), .RN(RESET), .QN(n295)
         );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n2634), .CK(CLK), .RN(RESET), .QN(n294)
         );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n2633), .CK(CLK), .RN(RESET), .QN(n293)
         );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n2632), .CK(CLK), .RN(RESET), .QN(n292)
         );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n2631), .CK(CLK), .RN(RESET), .QN(n291)
         );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n2630), .CK(CLK), .RN(RESET), .QN(n290)
         );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n2629), .CK(CLK), .RN(RESET), .QN(n289)
         );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n2628), .CK(CLK), .RN(RESET), .QN(n288)
         );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n2627), .CK(CLK), .RN(RESET), .QN(n287)
         );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n2626), .CK(CLK), .RN(RESET), .QN(n286)
         );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n2625), .CK(CLK), .RN(RESET), .QN(n285)
         );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n2624), .CK(CLK), .RN(RESET), .QN(n284)
         );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n2623), .CK(CLK), .RN(RESET), .QN(n283)
         );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n2622), .CK(CLK), .RN(RESET), .QN(n282)
         );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n2621), .CK(CLK), .RN(RESET), .QN(n281)
         );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n2620), .CK(CLK), .RN(RESET), .QN(n277)
         );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n2619), .CK(CLK), .RN(RESET), .QN(n276)
         );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n2618), .CK(CLK), .RN(RESET), .QN(n275)
         );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n2617), .CK(CLK), .RN(RESET), .QN(n274)
         );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n2616), .CK(CLK), .RN(RESET), .QN(n273)
         );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n2615), .CK(CLK), .RN(RESET), .QN(n272)
         );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n2614), .CK(CLK), .RN(RESET), .QN(n271)
         );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n2613), .CK(CLK), .RN(RESET), .QN(n270)
         );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n2612), .CK(CLK), .RN(RESET), .QN(n269)
         );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n2611), .CK(CLK), .RN(RESET), .QN(n268)
         );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n2610), .CK(CLK), .RN(RESET), .QN(n267)
         );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n2609), .CK(CLK), .RN(RESET), .QN(n266)
         );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n2608), .CK(CLK), .RN(RESET), .QN(n265)
         );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n2607), .CK(CLK), .RN(RESET), .QN(n264)
         );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n2606), .CK(CLK), .RN(RESET), .QN(n263)
         );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n2605), .CK(CLK), .RN(RESET), .QN(n262)
         );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n2604), .CK(CLK), .RN(RESET), .QN(n261)
         );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n2603), .CK(CLK), .RN(RESET), .QN(n260)
         );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n2602), .CK(CLK), .RN(RESET), .QN(n259)
         );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n2601), .CK(CLK), .RN(RESET), .QN(n258)
         );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n2600), .CK(CLK), .RN(RESET), .QN(n257)
         );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n2599), .CK(CLK), .RN(RESET), .QN(n256)
         );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n2598), .CK(CLK), .RN(RESET), .QN(n255)
         );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n2597), .CK(CLK), .RN(RESET), .QN(n254)
         );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n2596), .CK(CLK), .RN(RESET), .QN(n253)
         );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n2595), .CK(CLK), .RN(RESET), .QN(n252)
         );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n2594), .CK(CLK), .RN(RESET), .QN(n251)
         );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n2593), .CK(CLK), .RN(RESET), .QN(n250)
         );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n2592), .CK(CLK), .RN(RESET), .QN(n249)
         );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n2591), .CK(CLK), .RN(RESET), .QN(n248)
         );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n2590), .CK(CLK), .RN(RESET), .QN(n247)
         );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n2589), .CK(CLK), .RN(RESET), .QN(n246)
         );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n2588), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][31] ) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n2587), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][30] ) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n2586), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][29] ) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n2585), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][28] ) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n2584), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][27] ) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n2583), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][26] ) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n2582), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][25] ) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n2581), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][24] ) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n2580), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][23] ) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n2579), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][22] ) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n2578), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][21] ) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n2577), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][20] ) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n2576), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][19] ) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n2575), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][18] ) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n2574), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][17] ) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n2573), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][16] ) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n2572), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][15] ) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n2571), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][14] ) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n2570), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][13] ) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n2569), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][12] ) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n2568), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][11] ) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n2567), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][10] ) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n2566), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][9] ) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n2565), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][8] ) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n2564), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][7] ) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n2563), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][6] ) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n2562), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][5] ) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n2561), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][4] ) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n2560), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][3] ) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n2559), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][2] ) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n2558), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][1] ) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n2557), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[26][0] ) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n2556), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][31] ) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n2555), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][30] ) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n2554), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][29] ) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n2553), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][28] ) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n2552), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][27] ) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n2551), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][26] ) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n2550), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][25] ) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n2549), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][24] ) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n2548), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][23] ) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n2547), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][22] ) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n2546), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][21] ) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n2545), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][20] ) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n2544), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][19] ) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n2543), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][18] ) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n2542), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][17] ) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n2541), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][16] ) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n2540), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][15] ) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n2539), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][14] ) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n2538), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][13] ) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n2537), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][12] ) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n2536), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][11] ) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n2535), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][10] ) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n2534), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][9] ) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n2533), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][8] ) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n2532), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][7] ) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n2531), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][6] ) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n2530), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][5] ) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n2529), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][4] ) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n2528), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][3] ) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n2527), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][2] ) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n2526), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][1] ) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n2525), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[27][0] ) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n2524), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][31] ) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n2523), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][30] ) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n2522), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][29] ) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n2521), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][28] ) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n2520), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][27] ) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n2519), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][26] ) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n2518), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][25] ) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n2517), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][24] ) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n2516), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][23] ) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n2515), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][22] ) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n2514), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][21] ) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n2513), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][20] ) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n2512), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][19] ) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n2511), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][18] ) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n2510), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][17] ) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n2509), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][16] ) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n2508), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][15] ) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n2507), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][14] ) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n2506), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][13] ) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n2505), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][12] ) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n2504), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][11] ) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n2503), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][10] ) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n2502), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][9] ) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n2501), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][8] ) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n2500), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][7] ) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n2499), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][6] ) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n2498), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][5] ) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n2497), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][4] ) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n2496), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][3] ) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n2495), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][2] ) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n2494), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][1] ) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n2493), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[28][0] ) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n2492), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][31] ) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n2491), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][30] ) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n2490), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][29] ) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n2489), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][28] ) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n2488), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][27] ) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n2487), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][26] ) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n2486), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][25] ) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n2485), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][24] ) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n2484), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][23] ) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n2483), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][22] ) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n2482), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][21] ) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n2481), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][20] ) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n2480), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][19] ) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n2479), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][18] ) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n2478), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][17] ) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n2477), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][16] ) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n2476), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][15] ) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n2475), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][14] ) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n2474), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][13] ) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n2473), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][12] ) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n2472), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][11] ) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n2471), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][10] ) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n2470), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][9] ) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n2469), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][8] ) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n2468), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][7] ) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n2467), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][6] ) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n2466), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][5] ) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n2465), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][4] ) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n2464), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][3] ) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n2463), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][2] ) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n2462), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][1] ) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n2461), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[29][0] ) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n2460), .CK(CLK), .RN(RESET), .QN(n102)
         );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n2459), .CK(CLK), .RN(RESET), .QN(n101)
         );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n2458), .CK(CLK), .RN(RESET), .QN(n100)
         );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n2457), .CK(CLK), .RN(RESET), .QN(n99)
         );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n2456), .CK(CLK), .RN(RESET), .QN(n98)
         );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n2455), .CK(CLK), .RN(RESET), .QN(n97)
         );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n2454), .CK(CLK), .RN(RESET), .QN(n96)
         );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n2453), .CK(CLK), .RN(RESET), .QN(n95)
         );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n2452), .CK(CLK), .RN(RESET), .QN(n94)
         );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n2451), .CK(CLK), .RN(RESET), .QN(n93)
         );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n2450), .CK(CLK), .RN(RESET), .QN(n92)
         );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n2449), .CK(CLK), .RN(RESET), .QN(n91)
         );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n2448), .CK(CLK), .RN(RESET), .QN(n90)
         );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n2447), .CK(CLK), .RN(RESET), .QN(n89)
         );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n2446), .CK(CLK), .RN(RESET), .QN(n88)
         );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n2445), .CK(CLK), .RN(RESET), .QN(n87)
         );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n2444), .CK(CLK), .RN(RESET), .QN(n86)
         );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n2443), .CK(CLK), .RN(RESET), .QN(n85)
         );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n2442), .CK(CLK), .RN(RESET), .QN(n84)
         );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n2441), .CK(CLK), .RN(RESET), .QN(n83)
         );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n2440), .CK(CLK), .RN(RESET), .QN(n82)
         );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n2439), .CK(CLK), .RN(RESET), .QN(n81)
         );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n2438), .CK(CLK), .RN(RESET), .QN(n80)
         );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n2437), .CK(CLK), .RN(RESET), .QN(n79)
         );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n2436), .CK(CLK), .RN(RESET), .QN(n78)
         );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n2435), .CK(CLK), .RN(RESET), .QN(n77)
         );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n2434), .CK(CLK), .RN(RESET), .QN(n76)
         );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n2433), .CK(CLK), .RN(RESET), .QN(n75)
         );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n2432), .CK(CLK), .RN(RESET), .QN(n74)
         );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n2431), .CK(CLK), .RN(RESET), .QN(n73)
         );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n2430), .CK(CLK), .RN(RESET), .QN(n72)
         );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n2429), .CK(CLK), .RN(RESET), .QN(n71)
         );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n2428), .CK(CLK), .RN(RESET), .QN(n66)
         );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n2427), .CK(CLK), .RN(RESET), .QN(n64)
         );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n2426), .CK(CLK), .RN(RESET), .QN(n62)
         );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n2425), .CK(CLK), .RN(RESET), .QN(n60)
         );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n2424), .CK(CLK), .RN(RESET), .QN(n58)
         );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n2423), .CK(CLK), .RN(RESET), .QN(n56)
         );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n2422), .CK(CLK), .RN(RESET), .QN(n54)
         );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n2421), .CK(CLK), .RN(RESET), .QN(n52)
         );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n2420), .CK(CLK), .RN(RESET), .QN(n50)
         );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n2419), .CK(CLK), .RN(RESET), .QN(n48)
         );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n2418), .CK(CLK), .RN(RESET), .QN(n46)
         );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n2417), .CK(CLK), .RN(RESET), .QN(n44)
         );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n2416), .CK(CLK), .RN(RESET), .QN(n42)
         );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n2415), .CK(CLK), .RN(RESET), .QN(n40)
         );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n2414), .CK(CLK), .RN(RESET), .QN(n38)
         );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n2413), .CK(CLK), .RN(RESET), .QN(n36)
         );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n2412), .CK(CLK), .RN(RESET), .QN(n34)
         );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n2411), .CK(CLK), .RN(RESET), .QN(n32)
         );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n2410), .CK(CLK), .RN(RESET), .QN(n30)
         );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n2409), .CK(CLK), .RN(RESET), .QN(n28)
         );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n2408), .CK(CLK), .RN(RESET), .QN(n26)
         );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n2407), .CK(CLK), .RN(RESET), .QN(n24)
         );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n2406), .CK(CLK), .RN(RESET), .QN(n22)
         );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n2405), .CK(CLK), .RN(RESET), .QN(n20)
         );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n2404), .CK(CLK), .RN(RESET), .QN(n18)
         );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n2403), .CK(CLK), .RN(RESET), .QN(n16)
         );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n2402), .CK(CLK), .RN(RESET), .QN(n14)
         );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n2401), .CK(CLK), .RN(RESET), .QN(n12)
         );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n2400), .CK(CLK), .RN(RESET), .QN(n10)
         );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n2399), .CK(CLK), .RN(RESET), .QN(n8) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n2398), .CK(CLK), .RN(RESET), .QN(n6) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n2397), .CK(CLK), .RN(RESET), .QN(n4) );
  DLH_X1 \OUT1_reg[31]  ( .G(N286), .D(N318), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(N286), .D(N317), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(N286), .D(N316), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(N286), .D(N315), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(N286), .D(N314), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(N286), .D(N313), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(N286), .D(N312), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(N286), .D(N311), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(N286), .D(N310), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(N286), .D(N309), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(N286), .D(N308), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(N286), .D(N307), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(N286), .D(N306), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(N286), .D(N305), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(N286), .D(N304), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(N286), .D(N303), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(N286), .D(N302), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(N286), .D(N301), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(N286), .D(N300), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(N286), .D(N299), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(N286), .D(N298), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(N286), .D(N297), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(N286), .D(N296), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(N286), .D(N295), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(N286), .D(N294), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(N286), .D(N293), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(N286), .D(N292), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(N286), .D(N291), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(N286), .D(N290), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(N286), .D(N289), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(N286), .D(N288), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(N286), .D(N287), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(N319), .D(N351), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(N319), .D(N350), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(N319), .D(N349), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(N319), .D(N348), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(N319), .D(N347), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(N319), .D(N346), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(N319), .D(N345), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(N319), .D(N344), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(N319), .D(N343), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(N319), .D(N342), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(N319), .D(N341), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(N319), .D(N340), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(N319), .D(N339), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(N319), .D(N338), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(N319), .D(N337), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(N319), .D(N336), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(N319), .D(N335), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(N319), .D(N334), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(N319), .D(N333), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(N319), .D(N332), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(N319), .D(N331), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(N319), .D(N330), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(N319), .D(N329), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(N319), .D(N328), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(N319), .D(N327), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(N319), .D(N326), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(N319), .D(N325), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(N319), .D(N324), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(N319), .D(N323), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(N319), .D(N322), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(N319), .D(N321), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(N319), .D(N320), .Q(OUT2[0]) );
  OAI22_X1 U3 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(n2397) );
  OAI22_X1 U4 ( .A1(n1), .A2(n5), .B1(n3), .B2(n6), .ZN(n2398) );
  OAI22_X1 U5 ( .A1(n1), .A2(n7), .B1(n3), .B2(n8), .ZN(n2399) );
  OAI22_X1 U6 ( .A1(n1), .A2(n9), .B1(n3), .B2(n10), .ZN(n2400) );
  OAI22_X1 U7 ( .A1(n1), .A2(n11), .B1(n3), .B2(n12), .ZN(n2401) );
  OAI22_X1 U8 ( .A1(n1), .A2(n13), .B1(n3), .B2(n14), .ZN(n2402) );
  OAI22_X1 U9 ( .A1(n1), .A2(n15), .B1(n3), .B2(n16), .ZN(n2403) );
  OAI22_X1 U10 ( .A1(n1), .A2(n17), .B1(n3), .B2(n18), .ZN(n2404) );
  OAI22_X1 U11 ( .A1(n1), .A2(n19), .B1(n3), .B2(n20), .ZN(n2405) );
  OAI22_X1 U12 ( .A1(n1), .A2(n21), .B1(n3), .B2(n22), .ZN(n2406) );
  OAI22_X1 U13 ( .A1(n1), .A2(n23), .B1(n3), .B2(n24), .ZN(n2407) );
  OAI22_X1 U14 ( .A1(n1), .A2(n25), .B1(n3), .B2(n26), .ZN(n2408) );
  OAI22_X1 U15 ( .A1(n1), .A2(n27), .B1(n3), .B2(n28), .ZN(n2409) );
  OAI22_X1 U16 ( .A1(n1), .A2(n29), .B1(n3), .B2(n30), .ZN(n2410) );
  OAI22_X1 U17 ( .A1(n1), .A2(n31), .B1(n3), .B2(n32), .ZN(n2411) );
  OAI22_X1 U18 ( .A1(n1), .A2(n33), .B1(n3), .B2(n34), .ZN(n2412) );
  OAI22_X1 U19 ( .A1(n1), .A2(n35), .B1(n3), .B2(n36), .ZN(n2413) );
  OAI22_X1 U20 ( .A1(n1), .A2(n37), .B1(n3), .B2(n38), .ZN(n2414) );
  OAI22_X1 U21 ( .A1(n1), .A2(n39), .B1(n3), .B2(n40), .ZN(n2415) );
  OAI22_X1 U22 ( .A1(n1), .A2(n41), .B1(n3), .B2(n42), .ZN(n2416) );
  OAI22_X1 U23 ( .A1(n1), .A2(n43), .B1(n3), .B2(n44), .ZN(n2417) );
  OAI22_X1 U24 ( .A1(n1), .A2(n45), .B1(n3), .B2(n46), .ZN(n2418) );
  OAI22_X1 U25 ( .A1(n1), .A2(n47), .B1(n3), .B2(n48), .ZN(n2419) );
  OAI22_X1 U26 ( .A1(n1), .A2(n49), .B1(n3), .B2(n50), .ZN(n2420) );
  OAI22_X1 U27 ( .A1(n1), .A2(n51), .B1(n3), .B2(n52), .ZN(n2421) );
  OAI22_X1 U28 ( .A1(n1), .A2(n53), .B1(n3), .B2(n54), .ZN(n2422) );
  OAI22_X1 U29 ( .A1(n1), .A2(n55), .B1(n3), .B2(n56), .ZN(n2423) );
  OAI22_X1 U30 ( .A1(n1), .A2(n57), .B1(n3), .B2(n58), .ZN(n2424) );
  OAI22_X1 U31 ( .A1(n1), .A2(n59), .B1(n3), .B2(n60), .ZN(n2425) );
  OAI22_X1 U32 ( .A1(n1), .A2(n61), .B1(n3), .B2(n62), .ZN(n2426) );
  OAI22_X1 U33 ( .A1(n1), .A2(n63), .B1(n3), .B2(n64), .ZN(n2427) );
  OAI22_X1 U34 ( .A1(n1), .A2(n65), .B1(n3), .B2(n66), .ZN(n2428) );
  OAI22_X1 U37 ( .A1(n2), .A2(n69), .B1(n70), .B2(n71), .ZN(n2429) );
  OAI22_X1 U38 ( .A1(n5), .A2(n69), .B1(n70), .B2(n72), .ZN(n2430) );
  OAI22_X1 U39 ( .A1(n7), .A2(n69), .B1(n70), .B2(n73), .ZN(n2431) );
  OAI22_X1 U40 ( .A1(n9), .A2(n69), .B1(n70), .B2(n74), .ZN(n2432) );
  OAI22_X1 U41 ( .A1(n11), .A2(n69), .B1(n70), .B2(n75), .ZN(n2433) );
  OAI22_X1 U42 ( .A1(n13), .A2(n69), .B1(n70), .B2(n76), .ZN(n2434) );
  OAI22_X1 U43 ( .A1(n15), .A2(n69), .B1(n70), .B2(n77), .ZN(n2435) );
  OAI22_X1 U44 ( .A1(n17), .A2(n69), .B1(n70), .B2(n78), .ZN(n2436) );
  OAI22_X1 U45 ( .A1(n19), .A2(n69), .B1(n70), .B2(n79), .ZN(n2437) );
  OAI22_X1 U46 ( .A1(n21), .A2(n69), .B1(n70), .B2(n80), .ZN(n2438) );
  OAI22_X1 U47 ( .A1(n23), .A2(n69), .B1(n70), .B2(n81), .ZN(n2439) );
  OAI22_X1 U48 ( .A1(n25), .A2(n69), .B1(n70), .B2(n82), .ZN(n2440) );
  OAI22_X1 U49 ( .A1(n27), .A2(n69), .B1(n70), .B2(n83), .ZN(n2441) );
  OAI22_X1 U50 ( .A1(n29), .A2(n69), .B1(n70), .B2(n84), .ZN(n2442) );
  OAI22_X1 U51 ( .A1(n31), .A2(n69), .B1(n70), .B2(n85), .ZN(n2443) );
  OAI22_X1 U52 ( .A1(n33), .A2(n69), .B1(n70), .B2(n86), .ZN(n2444) );
  OAI22_X1 U53 ( .A1(n35), .A2(n69), .B1(n70), .B2(n87), .ZN(n2445) );
  OAI22_X1 U54 ( .A1(n37), .A2(n69), .B1(n70), .B2(n88), .ZN(n2446) );
  OAI22_X1 U55 ( .A1(n39), .A2(n69), .B1(n70), .B2(n89), .ZN(n2447) );
  OAI22_X1 U56 ( .A1(n41), .A2(n69), .B1(n70), .B2(n90), .ZN(n2448) );
  OAI22_X1 U57 ( .A1(n43), .A2(n69), .B1(n70), .B2(n91), .ZN(n2449) );
  OAI22_X1 U58 ( .A1(n45), .A2(n69), .B1(n70), .B2(n92), .ZN(n2450) );
  OAI22_X1 U59 ( .A1(n47), .A2(n69), .B1(n70), .B2(n93), .ZN(n2451) );
  OAI22_X1 U60 ( .A1(n49), .A2(n69), .B1(n70), .B2(n94), .ZN(n2452) );
  OAI22_X1 U61 ( .A1(n51), .A2(n69), .B1(n70), .B2(n95), .ZN(n2453) );
  OAI22_X1 U62 ( .A1(n53), .A2(n69), .B1(n70), .B2(n96), .ZN(n2454) );
  OAI22_X1 U63 ( .A1(n55), .A2(n69), .B1(n70), .B2(n97), .ZN(n2455) );
  OAI22_X1 U64 ( .A1(n57), .A2(n69), .B1(n70), .B2(n98), .ZN(n2456) );
  OAI22_X1 U65 ( .A1(n59), .A2(n69), .B1(n70), .B2(n99), .ZN(n2457) );
  OAI22_X1 U66 ( .A1(n61), .A2(n69), .B1(n70), .B2(n100), .ZN(n2458) );
  OAI22_X1 U67 ( .A1(n63), .A2(n69), .B1(n70), .B2(n101), .ZN(n2459) );
  OAI22_X1 U68 ( .A1(n65), .A2(n69), .B1(n70), .B2(n102), .ZN(n2460) );
  INV_X1 U71 ( .A(n104), .ZN(n2461) );
  AOI22_X1 U72 ( .A1(DATAIN[0]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][0] ), 
        .ZN(n104) );
  INV_X1 U73 ( .A(n107), .ZN(n2462) );
  AOI22_X1 U74 ( .A1(DATAIN[1]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][1] ), 
        .ZN(n107) );
  INV_X1 U75 ( .A(n108), .ZN(n2463) );
  AOI22_X1 U76 ( .A1(DATAIN[2]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][2] ), 
        .ZN(n108) );
  INV_X1 U77 ( .A(n109), .ZN(n2464) );
  AOI22_X1 U78 ( .A1(DATAIN[3]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][3] ), 
        .ZN(n109) );
  INV_X1 U79 ( .A(n110), .ZN(n2465) );
  AOI22_X1 U80 ( .A1(DATAIN[4]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][4] ), 
        .ZN(n110) );
  INV_X1 U81 ( .A(n111), .ZN(n2466) );
  AOI22_X1 U82 ( .A1(DATAIN[5]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][5] ), 
        .ZN(n111) );
  INV_X1 U83 ( .A(n112), .ZN(n2467) );
  AOI22_X1 U84 ( .A1(DATAIN[6]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][6] ), 
        .ZN(n112) );
  INV_X1 U85 ( .A(n113), .ZN(n2468) );
  AOI22_X1 U86 ( .A1(DATAIN[7]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][7] ), 
        .ZN(n113) );
  INV_X1 U87 ( .A(n114), .ZN(n2469) );
  AOI22_X1 U88 ( .A1(DATAIN[8]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][8] ), 
        .ZN(n114) );
  INV_X1 U89 ( .A(n115), .ZN(n2470) );
  AOI22_X1 U90 ( .A1(DATAIN[9]), .A2(n105), .B1(n106), .B2(\REGISTERS[29][9] ), 
        .ZN(n115) );
  INV_X1 U91 ( .A(n116), .ZN(n2471) );
  AOI22_X1 U92 ( .A1(DATAIN[10]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][10] ), .ZN(n116) );
  INV_X1 U93 ( .A(n117), .ZN(n2472) );
  AOI22_X1 U94 ( .A1(DATAIN[11]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][11] ), .ZN(n117) );
  INV_X1 U95 ( .A(n118), .ZN(n2473) );
  AOI22_X1 U96 ( .A1(DATAIN[12]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][12] ), .ZN(n118) );
  INV_X1 U97 ( .A(n119), .ZN(n2474) );
  AOI22_X1 U98 ( .A1(DATAIN[13]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][13] ), .ZN(n119) );
  INV_X1 U99 ( .A(n120), .ZN(n2475) );
  AOI22_X1 U100 ( .A1(DATAIN[14]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][14] ), .ZN(n120) );
  INV_X1 U101 ( .A(n121), .ZN(n2476) );
  AOI22_X1 U102 ( .A1(DATAIN[15]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][15] ), .ZN(n121) );
  INV_X1 U103 ( .A(n122), .ZN(n2477) );
  AOI22_X1 U104 ( .A1(DATAIN[16]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][16] ), .ZN(n122) );
  INV_X1 U105 ( .A(n123), .ZN(n2478) );
  AOI22_X1 U106 ( .A1(DATAIN[17]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][17] ), .ZN(n123) );
  INV_X1 U107 ( .A(n124), .ZN(n2479) );
  AOI22_X1 U108 ( .A1(DATAIN[18]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][18] ), .ZN(n124) );
  INV_X1 U109 ( .A(n125), .ZN(n2480) );
  AOI22_X1 U110 ( .A1(DATAIN[19]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][19] ), .ZN(n125) );
  INV_X1 U111 ( .A(n126), .ZN(n2481) );
  AOI22_X1 U112 ( .A1(DATAIN[20]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][20] ), .ZN(n126) );
  INV_X1 U113 ( .A(n127), .ZN(n2482) );
  AOI22_X1 U114 ( .A1(DATAIN[21]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][21] ), .ZN(n127) );
  INV_X1 U115 ( .A(n128), .ZN(n2483) );
  AOI22_X1 U116 ( .A1(DATAIN[22]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][22] ), .ZN(n128) );
  INV_X1 U117 ( .A(n129), .ZN(n2484) );
  AOI22_X1 U118 ( .A1(DATAIN[23]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][23] ), .ZN(n129) );
  INV_X1 U119 ( .A(n130), .ZN(n2485) );
  AOI22_X1 U120 ( .A1(DATAIN[24]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][24] ), .ZN(n130) );
  INV_X1 U121 ( .A(n131), .ZN(n2486) );
  AOI22_X1 U122 ( .A1(DATAIN[25]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][25] ), .ZN(n131) );
  INV_X1 U123 ( .A(n132), .ZN(n2487) );
  AOI22_X1 U124 ( .A1(DATAIN[26]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][26] ), .ZN(n132) );
  INV_X1 U125 ( .A(n133), .ZN(n2488) );
  AOI22_X1 U126 ( .A1(DATAIN[27]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][27] ), .ZN(n133) );
  INV_X1 U127 ( .A(n134), .ZN(n2489) );
  AOI22_X1 U128 ( .A1(DATAIN[28]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][28] ), .ZN(n134) );
  INV_X1 U129 ( .A(n135), .ZN(n2490) );
  AOI22_X1 U130 ( .A1(DATAIN[29]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][29] ), .ZN(n135) );
  INV_X1 U131 ( .A(n136), .ZN(n2491) );
  AOI22_X1 U132 ( .A1(DATAIN[30]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][30] ), .ZN(n136) );
  INV_X1 U133 ( .A(n137), .ZN(n2492) );
  AOI22_X1 U134 ( .A1(DATAIN[31]), .A2(n105), .B1(n106), .B2(
        \REGISTERS[29][31] ), .ZN(n137) );
  INV_X1 U137 ( .A(n139), .ZN(n2493) );
  AOI22_X1 U138 ( .A1(DATAIN[0]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][0] ), .ZN(n139) );
  INV_X1 U139 ( .A(n142), .ZN(n2494) );
  AOI22_X1 U140 ( .A1(DATAIN[1]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][1] ), .ZN(n142) );
  INV_X1 U141 ( .A(n143), .ZN(n2495) );
  AOI22_X1 U142 ( .A1(DATAIN[2]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][2] ), .ZN(n143) );
  INV_X1 U143 ( .A(n144), .ZN(n2496) );
  AOI22_X1 U144 ( .A1(DATAIN[3]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][3] ), .ZN(n144) );
  INV_X1 U145 ( .A(n145), .ZN(n2497) );
  AOI22_X1 U146 ( .A1(DATAIN[4]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][4] ), .ZN(n145) );
  INV_X1 U147 ( .A(n146), .ZN(n2498) );
  AOI22_X1 U148 ( .A1(DATAIN[5]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][5] ), .ZN(n146) );
  INV_X1 U149 ( .A(n147), .ZN(n2499) );
  AOI22_X1 U150 ( .A1(DATAIN[6]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][6] ), .ZN(n147) );
  INV_X1 U151 ( .A(n148), .ZN(n2500) );
  AOI22_X1 U152 ( .A1(DATAIN[7]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][7] ), .ZN(n148) );
  INV_X1 U153 ( .A(n149), .ZN(n2501) );
  AOI22_X1 U154 ( .A1(DATAIN[8]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][8] ), .ZN(n149) );
  INV_X1 U155 ( .A(n150), .ZN(n2502) );
  AOI22_X1 U156 ( .A1(DATAIN[9]), .A2(n140), .B1(n141), .B2(\REGISTERS[28][9] ), .ZN(n150) );
  INV_X1 U157 ( .A(n151), .ZN(n2503) );
  AOI22_X1 U158 ( .A1(DATAIN[10]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][10] ), .ZN(n151) );
  INV_X1 U159 ( .A(n152), .ZN(n2504) );
  AOI22_X1 U160 ( .A1(DATAIN[11]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][11] ), .ZN(n152) );
  INV_X1 U161 ( .A(n153), .ZN(n2505) );
  AOI22_X1 U162 ( .A1(DATAIN[12]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][12] ), .ZN(n153) );
  INV_X1 U163 ( .A(n154), .ZN(n2506) );
  AOI22_X1 U164 ( .A1(DATAIN[13]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][13] ), .ZN(n154) );
  INV_X1 U165 ( .A(n155), .ZN(n2507) );
  AOI22_X1 U166 ( .A1(DATAIN[14]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][14] ), .ZN(n155) );
  INV_X1 U167 ( .A(n156), .ZN(n2508) );
  AOI22_X1 U168 ( .A1(DATAIN[15]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][15] ), .ZN(n156) );
  INV_X1 U169 ( .A(n157), .ZN(n2509) );
  AOI22_X1 U170 ( .A1(DATAIN[16]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][16] ), .ZN(n157) );
  INV_X1 U171 ( .A(n158), .ZN(n2510) );
  AOI22_X1 U172 ( .A1(DATAIN[17]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][17] ), .ZN(n158) );
  INV_X1 U173 ( .A(n159), .ZN(n2511) );
  AOI22_X1 U174 ( .A1(DATAIN[18]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][18] ), .ZN(n159) );
  INV_X1 U175 ( .A(n160), .ZN(n2512) );
  AOI22_X1 U176 ( .A1(DATAIN[19]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][19] ), .ZN(n160) );
  INV_X1 U177 ( .A(n161), .ZN(n2513) );
  AOI22_X1 U178 ( .A1(DATAIN[20]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][20] ), .ZN(n161) );
  INV_X1 U179 ( .A(n162), .ZN(n2514) );
  AOI22_X1 U180 ( .A1(DATAIN[21]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][21] ), .ZN(n162) );
  INV_X1 U181 ( .A(n163), .ZN(n2515) );
  AOI22_X1 U182 ( .A1(DATAIN[22]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][22] ), .ZN(n163) );
  INV_X1 U183 ( .A(n164), .ZN(n2516) );
  AOI22_X1 U184 ( .A1(DATAIN[23]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][23] ), .ZN(n164) );
  INV_X1 U185 ( .A(n165), .ZN(n2517) );
  AOI22_X1 U186 ( .A1(DATAIN[24]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][24] ), .ZN(n165) );
  INV_X1 U187 ( .A(n166), .ZN(n2518) );
  AOI22_X1 U188 ( .A1(DATAIN[25]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][25] ), .ZN(n166) );
  INV_X1 U189 ( .A(n167), .ZN(n2519) );
  AOI22_X1 U190 ( .A1(DATAIN[26]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][26] ), .ZN(n167) );
  INV_X1 U191 ( .A(n168), .ZN(n2520) );
  AOI22_X1 U192 ( .A1(DATAIN[27]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][27] ), .ZN(n168) );
  INV_X1 U193 ( .A(n169), .ZN(n2521) );
  AOI22_X1 U194 ( .A1(DATAIN[28]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][28] ), .ZN(n169) );
  INV_X1 U195 ( .A(n170), .ZN(n2522) );
  AOI22_X1 U196 ( .A1(DATAIN[29]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][29] ), .ZN(n170) );
  INV_X1 U197 ( .A(n171), .ZN(n2523) );
  AOI22_X1 U198 ( .A1(DATAIN[30]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][30] ), .ZN(n171) );
  INV_X1 U199 ( .A(n172), .ZN(n2524) );
  AOI22_X1 U200 ( .A1(DATAIN[31]), .A2(n140), .B1(n141), .B2(
        \REGISTERS[28][31] ), .ZN(n172) );
  INV_X1 U203 ( .A(n174), .ZN(n2525) );
  AOI22_X1 U204 ( .A1(DATAIN[0]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][0] ), .ZN(n174) );
  INV_X1 U205 ( .A(n177), .ZN(n2526) );
  AOI22_X1 U206 ( .A1(DATAIN[1]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][1] ), .ZN(n177) );
  INV_X1 U207 ( .A(n178), .ZN(n2527) );
  AOI22_X1 U208 ( .A1(DATAIN[2]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][2] ), .ZN(n178) );
  INV_X1 U209 ( .A(n179), .ZN(n2528) );
  AOI22_X1 U210 ( .A1(DATAIN[3]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][3] ), .ZN(n179) );
  INV_X1 U211 ( .A(n180), .ZN(n2529) );
  AOI22_X1 U212 ( .A1(DATAIN[4]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][4] ), .ZN(n180) );
  INV_X1 U213 ( .A(n181), .ZN(n2530) );
  AOI22_X1 U214 ( .A1(DATAIN[5]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][5] ), .ZN(n181) );
  INV_X1 U215 ( .A(n182), .ZN(n2531) );
  AOI22_X1 U216 ( .A1(DATAIN[6]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][6] ), .ZN(n182) );
  INV_X1 U217 ( .A(n183), .ZN(n2532) );
  AOI22_X1 U218 ( .A1(DATAIN[7]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][7] ), .ZN(n183) );
  INV_X1 U219 ( .A(n184), .ZN(n2533) );
  AOI22_X1 U220 ( .A1(DATAIN[8]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][8] ), .ZN(n184) );
  INV_X1 U221 ( .A(n185), .ZN(n2534) );
  AOI22_X1 U222 ( .A1(DATAIN[9]), .A2(n175), .B1(n176), .B2(\REGISTERS[27][9] ), .ZN(n185) );
  INV_X1 U223 ( .A(n186), .ZN(n2535) );
  AOI22_X1 U224 ( .A1(DATAIN[10]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][10] ), .ZN(n186) );
  INV_X1 U225 ( .A(n187), .ZN(n2536) );
  AOI22_X1 U226 ( .A1(DATAIN[11]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][11] ), .ZN(n187) );
  INV_X1 U227 ( .A(n188), .ZN(n2537) );
  AOI22_X1 U228 ( .A1(DATAIN[12]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][12] ), .ZN(n188) );
  INV_X1 U229 ( .A(n189), .ZN(n2538) );
  AOI22_X1 U230 ( .A1(DATAIN[13]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][13] ), .ZN(n189) );
  INV_X1 U231 ( .A(n190), .ZN(n2539) );
  AOI22_X1 U232 ( .A1(DATAIN[14]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][14] ), .ZN(n190) );
  INV_X1 U233 ( .A(n191), .ZN(n2540) );
  AOI22_X1 U234 ( .A1(DATAIN[15]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][15] ), .ZN(n191) );
  INV_X1 U235 ( .A(n192), .ZN(n2541) );
  AOI22_X1 U236 ( .A1(DATAIN[16]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][16] ), .ZN(n192) );
  INV_X1 U237 ( .A(n193), .ZN(n2542) );
  AOI22_X1 U238 ( .A1(DATAIN[17]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][17] ), .ZN(n193) );
  INV_X1 U239 ( .A(n194), .ZN(n2543) );
  AOI22_X1 U240 ( .A1(DATAIN[18]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][18] ), .ZN(n194) );
  INV_X1 U241 ( .A(n195), .ZN(n2544) );
  AOI22_X1 U242 ( .A1(DATAIN[19]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][19] ), .ZN(n195) );
  INV_X1 U243 ( .A(n196), .ZN(n2545) );
  AOI22_X1 U244 ( .A1(DATAIN[20]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][20] ), .ZN(n196) );
  INV_X1 U245 ( .A(n197), .ZN(n2546) );
  AOI22_X1 U246 ( .A1(DATAIN[21]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][21] ), .ZN(n197) );
  INV_X1 U247 ( .A(n198), .ZN(n2547) );
  AOI22_X1 U248 ( .A1(DATAIN[22]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][22] ), .ZN(n198) );
  INV_X1 U249 ( .A(n199), .ZN(n2548) );
  AOI22_X1 U250 ( .A1(DATAIN[23]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][23] ), .ZN(n199) );
  INV_X1 U251 ( .A(n200), .ZN(n2549) );
  AOI22_X1 U252 ( .A1(DATAIN[24]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][24] ), .ZN(n200) );
  INV_X1 U253 ( .A(n201), .ZN(n2550) );
  AOI22_X1 U254 ( .A1(DATAIN[25]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][25] ), .ZN(n201) );
  INV_X1 U255 ( .A(n202), .ZN(n2551) );
  AOI22_X1 U256 ( .A1(DATAIN[26]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][26] ), .ZN(n202) );
  INV_X1 U257 ( .A(n203), .ZN(n2552) );
  AOI22_X1 U258 ( .A1(DATAIN[27]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][27] ), .ZN(n203) );
  INV_X1 U259 ( .A(n204), .ZN(n2553) );
  AOI22_X1 U260 ( .A1(DATAIN[28]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][28] ), .ZN(n204) );
  INV_X1 U261 ( .A(n205), .ZN(n2554) );
  AOI22_X1 U262 ( .A1(DATAIN[29]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][29] ), .ZN(n205) );
  INV_X1 U263 ( .A(n206), .ZN(n2555) );
  AOI22_X1 U264 ( .A1(DATAIN[30]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][30] ), .ZN(n206) );
  INV_X1 U265 ( .A(n207), .ZN(n2556) );
  AOI22_X1 U266 ( .A1(DATAIN[31]), .A2(n175), .B1(n176), .B2(
        \REGISTERS[27][31] ), .ZN(n207) );
  INV_X1 U269 ( .A(n209), .ZN(n2557) );
  AOI22_X1 U270 ( .A1(DATAIN[0]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][0] ), .ZN(n209) );
  INV_X1 U271 ( .A(n212), .ZN(n2558) );
  AOI22_X1 U272 ( .A1(DATAIN[1]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][1] ), .ZN(n212) );
  INV_X1 U273 ( .A(n213), .ZN(n2559) );
  AOI22_X1 U274 ( .A1(DATAIN[2]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][2] ), .ZN(n213) );
  INV_X1 U275 ( .A(n214), .ZN(n2560) );
  AOI22_X1 U276 ( .A1(DATAIN[3]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][3] ), .ZN(n214) );
  INV_X1 U277 ( .A(n215), .ZN(n2561) );
  AOI22_X1 U278 ( .A1(DATAIN[4]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][4] ), .ZN(n215) );
  INV_X1 U279 ( .A(n216), .ZN(n2562) );
  AOI22_X1 U280 ( .A1(DATAIN[5]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][5] ), .ZN(n216) );
  INV_X1 U281 ( .A(n217), .ZN(n2563) );
  AOI22_X1 U282 ( .A1(DATAIN[6]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][6] ), .ZN(n217) );
  INV_X1 U283 ( .A(n218), .ZN(n2564) );
  AOI22_X1 U284 ( .A1(DATAIN[7]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][7] ), .ZN(n218) );
  INV_X1 U285 ( .A(n219), .ZN(n2565) );
  AOI22_X1 U286 ( .A1(DATAIN[8]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][8] ), .ZN(n219) );
  INV_X1 U287 ( .A(n220), .ZN(n2566) );
  AOI22_X1 U288 ( .A1(DATAIN[9]), .A2(n210), .B1(n211), .B2(\REGISTERS[26][9] ), .ZN(n220) );
  INV_X1 U289 ( .A(n221), .ZN(n2567) );
  AOI22_X1 U290 ( .A1(DATAIN[10]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][10] ), .ZN(n221) );
  INV_X1 U291 ( .A(n222), .ZN(n2568) );
  AOI22_X1 U292 ( .A1(DATAIN[11]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][11] ), .ZN(n222) );
  INV_X1 U293 ( .A(n223), .ZN(n2569) );
  AOI22_X1 U294 ( .A1(DATAIN[12]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][12] ), .ZN(n223) );
  INV_X1 U295 ( .A(n224), .ZN(n2570) );
  AOI22_X1 U296 ( .A1(DATAIN[13]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][13] ), .ZN(n224) );
  INV_X1 U297 ( .A(n225), .ZN(n2571) );
  AOI22_X1 U298 ( .A1(DATAIN[14]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][14] ), .ZN(n225) );
  INV_X1 U299 ( .A(n226), .ZN(n2572) );
  AOI22_X1 U300 ( .A1(DATAIN[15]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][15] ), .ZN(n226) );
  INV_X1 U301 ( .A(n227), .ZN(n2573) );
  AOI22_X1 U302 ( .A1(DATAIN[16]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][16] ), .ZN(n227) );
  INV_X1 U303 ( .A(n228), .ZN(n2574) );
  AOI22_X1 U304 ( .A1(DATAIN[17]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][17] ), .ZN(n228) );
  INV_X1 U305 ( .A(n229), .ZN(n2575) );
  AOI22_X1 U306 ( .A1(DATAIN[18]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][18] ), .ZN(n229) );
  INV_X1 U307 ( .A(n230), .ZN(n2576) );
  AOI22_X1 U308 ( .A1(DATAIN[19]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][19] ), .ZN(n230) );
  INV_X1 U309 ( .A(n231), .ZN(n2577) );
  AOI22_X1 U310 ( .A1(DATAIN[20]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][20] ), .ZN(n231) );
  INV_X1 U311 ( .A(n232), .ZN(n2578) );
  AOI22_X1 U312 ( .A1(DATAIN[21]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][21] ), .ZN(n232) );
  INV_X1 U313 ( .A(n233), .ZN(n2579) );
  AOI22_X1 U314 ( .A1(DATAIN[22]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][22] ), .ZN(n233) );
  INV_X1 U315 ( .A(n234), .ZN(n2580) );
  AOI22_X1 U316 ( .A1(DATAIN[23]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][23] ), .ZN(n234) );
  INV_X1 U317 ( .A(n235), .ZN(n2581) );
  AOI22_X1 U318 ( .A1(DATAIN[24]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][24] ), .ZN(n235) );
  INV_X1 U319 ( .A(n236), .ZN(n2582) );
  AOI22_X1 U320 ( .A1(DATAIN[25]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][25] ), .ZN(n236) );
  INV_X1 U321 ( .A(n237), .ZN(n2583) );
  AOI22_X1 U322 ( .A1(DATAIN[26]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][26] ), .ZN(n237) );
  INV_X1 U323 ( .A(n238), .ZN(n2584) );
  AOI22_X1 U324 ( .A1(DATAIN[27]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][27] ), .ZN(n238) );
  INV_X1 U325 ( .A(n239), .ZN(n2585) );
  AOI22_X1 U326 ( .A1(DATAIN[28]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][28] ), .ZN(n239) );
  INV_X1 U327 ( .A(n240), .ZN(n2586) );
  AOI22_X1 U328 ( .A1(DATAIN[29]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][29] ), .ZN(n240) );
  INV_X1 U329 ( .A(n241), .ZN(n2587) );
  AOI22_X1 U330 ( .A1(DATAIN[30]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][30] ), .ZN(n241) );
  INV_X1 U331 ( .A(n242), .ZN(n2588) );
  AOI22_X1 U332 ( .A1(DATAIN[31]), .A2(n210), .B1(n211), .B2(
        \REGISTERS[26][31] ), .ZN(n242) );
  OAI22_X1 U335 ( .A1(n2), .A2(n244), .B1(n245), .B2(n246), .ZN(n2589) );
  OAI22_X1 U336 ( .A1(n5), .A2(n244), .B1(n245), .B2(n247), .ZN(n2590) );
  OAI22_X1 U337 ( .A1(n7), .A2(n244), .B1(n245), .B2(n248), .ZN(n2591) );
  OAI22_X1 U338 ( .A1(n9), .A2(n244), .B1(n245), .B2(n249), .ZN(n2592) );
  OAI22_X1 U339 ( .A1(n11), .A2(n244), .B1(n245), .B2(n250), .ZN(n2593) );
  OAI22_X1 U340 ( .A1(n13), .A2(n244), .B1(n245), .B2(n251), .ZN(n2594) );
  OAI22_X1 U341 ( .A1(n15), .A2(n244), .B1(n245), .B2(n252), .ZN(n2595) );
  OAI22_X1 U342 ( .A1(n17), .A2(n244), .B1(n245), .B2(n253), .ZN(n2596) );
  OAI22_X1 U343 ( .A1(n19), .A2(n244), .B1(n245), .B2(n254), .ZN(n2597) );
  OAI22_X1 U344 ( .A1(n21), .A2(n244), .B1(n245), .B2(n255), .ZN(n2598) );
  OAI22_X1 U345 ( .A1(n23), .A2(n244), .B1(n245), .B2(n256), .ZN(n2599) );
  OAI22_X1 U346 ( .A1(n25), .A2(n244), .B1(n245), .B2(n257), .ZN(n2600) );
  OAI22_X1 U347 ( .A1(n27), .A2(n244), .B1(n245), .B2(n258), .ZN(n2601) );
  OAI22_X1 U348 ( .A1(n29), .A2(n244), .B1(n245), .B2(n259), .ZN(n2602) );
  OAI22_X1 U349 ( .A1(n31), .A2(n244), .B1(n245), .B2(n260), .ZN(n2603) );
  OAI22_X1 U350 ( .A1(n33), .A2(n244), .B1(n245), .B2(n261), .ZN(n2604) );
  OAI22_X1 U351 ( .A1(n35), .A2(n244), .B1(n245), .B2(n262), .ZN(n2605) );
  OAI22_X1 U352 ( .A1(n37), .A2(n244), .B1(n245), .B2(n263), .ZN(n2606) );
  OAI22_X1 U353 ( .A1(n39), .A2(n244), .B1(n245), .B2(n264), .ZN(n2607) );
  OAI22_X1 U354 ( .A1(n41), .A2(n244), .B1(n245), .B2(n265), .ZN(n2608) );
  OAI22_X1 U355 ( .A1(n43), .A2(n244), .B1(n245), .B2(n266), .ZN(n2609) );
  OAI22_X1 U356 ( .A1(n45), .A2(n244), .B1(n245), .B2(n267), .ZN(n2610) );
  OAI22_X1 U357 ( .A1(n47), .A2(n244), .B1(n245), .B2(n268), .ZN(n2611) );
  OAI22_X1 U358 ( .A1(n49), .A2(n244), .B1(n245), .B2(n269), .ZN(n2612) );
  OAI22_X1 U359 ( .A1(n51), .A2(n244), .B1(n245), .B2(n270), .ZN(n2613) );
  OAI22_X1 U360 ( .A1(n53), .A2(n244), .B1(n245), .B2(n271), .ZN(n2614) );
  OAI22_X1 U361 ( .A1(n55), .A2(n244), .B1(n245), .B2(n272), .ZN(n2615) );
  OAI22_X1 U362 ( .A1(n57), .A2(n244), .B1(n245), .B2(n273), .ZN(n2616) );
  OAI22_X1 U363 ( .A1(n59), .A2(n244), .B1(n245), .B2(n274), .ZN(n2617) );
  OAI22_X1 U364 ( .A1(n61), .A2(n244), .B1(n245), .B2(n275), .ZN(n2618) );
  OAI22_X1 U365 ( .A1(n63), .A2(n244), .B1(n245), .B2(n276), .ZN(n2619) );
  OAI22_X1 U366 ( .A1(n65), .A2(n244), .B1(n245), .B2(n277), .ZN(n2620) );
  OAI22_X1 U369 ( .A1(n2), .A2(n279), .B1(n280), .B2(n281), .ZN(n2621) );
  OAI22_X1 U370 ( .A1(n5), .A2(n279), .B1(n280), .B2(n282), .ZN(n2622) );
  OAI22_X1 U371 ( .A1(n7), .A2(n279), .B1(n280), .B2(n283), .ZN(n2623) );
  OAI22_X1 U372 ( .A1(n9), .A2(n279), .B1(n280), .B2(n284), .ZN(n2624) );
  OAI22_X1 U373 ( .A1(n11), .A2(n279), .B1(n280), .B2(n285), .ZN(n2625) );
  OAI22_X1 U374 ( .A1(n13), .A2(n279), .B1(n280), .B2(n286), .ZN(n2626) );
  OAI22_X1 U375 ( .A1(n15), .A2(n279), .B1(n280), .B2(n287), .ZN(n2627) );
  OAI22_X1 U376 ( .A1(n17), .A2(n279), .B1(n280), .B2(n288), .ZN(n2628) );
  OAI22_X1 U377 ( .A1(n19), .A2(n279), .B1(n280), .B2(n289), .ZN(n2629) );
  OAI22_X1 U378 ( .A1(n21), .A2(n279), .B1(n280), .B2(n290), .ZN(n2630) );
  OAI22_X1 U379 ( .A1(n23), .A2(n279), .B1(n280), .B2(n291), .ZN(n2631) );
  OAI22_X1 U380 ( .A1(n25), .A2(n279), .B1(n280), .B2(n292), .ZN(n2632) );
  OAI22_X1 U381 ( .A1(n27), .A2(n279), .B1(n280), .B2(n293), .ZN(n2633) );
  OAI22_X1 U382 ( .A1(n29), .A2(n279), .B1(n280), .B2(n294), .ZN(n2634) );
  OAI22_X1 U383 ( .A1(n31), .A2(n279), .B1(n280), .B2(n295), .ZN(n2635) );
  OAI22_X1 U384 ( .A1(n33), .A2(n279), .B1(n280), .B2(n296), .ZN(n2636) );
  OAI22_X1 U385 ( .A1(n35), .A2(n279), .B1(n280), .B2(n297), .ZN(n2637) );
  OAI22_X1 U386 ( .A1(n37), .A2(n279), .B1(n280), .B2(n298), .ZN(n2638) );
  OAI22_X1 U387 ( .A1(n39), .A2(n279), .B1(n280), .B2(n299), .ZN(n2639) );
  OAI22_X1 U388 ( .A1(n41), .A2(n279), .B1(n280), .B2(n300), .ZN(n2640) );
  OAI22_X1 U389 ( .A1(n43), .A2(n279), .B1(n280), .B2(n301), .ZN(n2641) );
  OAI22_X1 U390 ( .A1(n45), .A2(n279), .B1(n280), .B2(n302), .ZN(n2642) );
  OAI22_X1 U391 ( .A1(n47), .A2(n279), .B1(n280), .B2(n303), .ZN(n2643) );
  OAI22_X1 U392 ( .A1(n49), .A2(n279), .B1(n280), .B2(n304), .ZN(n2644) );
  OAI22_X1 U393 ( .A1(n51), .A2(n279), .B1(n280), .B2(n305), .ZN(n2645) );
  OAI22_X1 U394 ( .A1(n53), .A2(n279), .B1(n280), .B2(n306), .ZN(n2646) );
  OAI22_X1 U395 ( .A1(n55), .A2(n279), .B1(n280), .B2(n307), .ZN(n2647) );
  OAI22_X1 U396 ( .A1(n57), .A2(n279), .B1(n280), .B2(n308), .ZN(n2648) );
  OAI22_X1 U397 ( .A1(n59), .A2(n279), .B1(n280), .B2(n309), .ZN(n2649) );
  OAI22_X1 U398 ( .A1(n61), .A2(n279), .B1(n280), .B2(n310), .ZN(n2650) );
  OAI22_X1 U399 ( .A1(n63), .A2(n279), .B1(n280), .B2(n311), .ZN(n2651) );
  OAI22_X1 U400 ( .A1(n65), .A2(n279), .B1(n280), .B2(n312), .ZN(n2652) );
  AND3_X1 U403 ( .A1(ADD_WR[3]), .A2(n314), .A3(ADD_WR[4]), .ZN(n68) );
  INV_X1 U404 ( .A(n315), .ZN(n2653) );
  AOI22_X1 U405 ( .A1(DATAIN[0]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][0] ), .ZN(n315) );
  INV_X1 U406 ( .A(n318), .ZN(n2654) );
  AOI22_X1 U407 ( .A1(DATAIN[1]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][1] ), .ZN(n318) );
  INV_X1 U408 ( .A(n319), .ZN(n2655) );
  AOI22_X1 U409 ( .A1(DATAIN[2]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][2] ), .ZN(n319) );
  INV_X1 U410 ( .A(n320), .ZN(n2656) );
  AOI22_X1 U411 ( .A1(DATAIN[3]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][3] ), .ZN(n320) );
  INV_X1 U412 ( .A(n321), .ZN(n2657) );
  AOI22_X1 U413 ( .A1(DATAIN[4]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][4] ), .ZN(n321) );
  INV_X1 U414 ( .A(n322), .ZN(n2658) );
  AOI22_X1 U415 ( .A1(DATAIN[5]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][5] ), .ZN(n322) );
  INV_X1 U416 ( .A(n323), .ZN(n2659) );
  AOI22_X1 U417 ( .A1(DATAIN[6]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][6] ), .ZN(n323) );
  INV_X1 U418 ( .A(n324), .ZN(n2660) );
  AOI22_X1 U419 ( .A1(DATAIN[7]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][7] ), .ZN(n324) );
  INV_X1 U420 ( .A(n325), .ZN(n2661) );
  AOI22_X1 U421 ( .A1(DATAIN[8]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][8] ), .ZN(n325) );
  INV_X1 U422 ( .A(n326), .ZN(n2662) );
  AOI22_X1 U423 ( .A1(DATAIN[9]), .A2(n316), .B1(n317), .B2(\REGISTERS[23][9] ), .ZN(n326) );
  INV_X1 U424 ( .A(n327), .ZN(n2663) );
  AOI22_X1 U425 ( .A1(DATAIN[10]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][10] ), .ZN(n327) );
  INV_X1 U426 ( .A(n328), .ZN(n2664) );
  AOI22_X1 U427 ( .A1(DATAIN[11]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][11] ), .ZN(n328) );
  INV_X1 U428 ( .A(n329), .ZN(n2665) );
  AOI22_X1 U429 ( .A1(DATAIN[12]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][12] ), .ZN(n329) );
  INV_X1 U430 ( .A(n330), .ZN(n2666) );
  AOI22_X1 U431 ( .A1(DATAIN[13]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][13] ), .ZN(n330) );
  INV_X1 U432 ( .A(n331), .ZN(n2667) );
  AOI22_X1 U433 ( .A1(DATAIN[14]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][14] ), .ZN(n331) );
  INV_X1 U434 ( .A(n332), .ZN(n2668) );
  AOI22_X1 U435 ( .A1(DATAIN[15]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][15] ), .ZN(n332) );
  INV_X1 U436 ( .A(n333), .ZN(n2669) );
  AOI22_X1 U437 ( .A1(DATAIN[16]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][16] ), .ZN(n333) );
  INV_X1 U438 ( .A(n334), .ZN(n2670) );
  AOI22_X1 U439 ( .A1(DATAIN[17]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][17] ), .ZN(n334) );
  INV_X1 U440 ( .A(n335), .ZN(n2671) );
  AOI22_X1 U441 ( .A1(DATAIN[18]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][18] ), .ZN(n335) );
  INV_X1 U442 ( .A(n336), .ZN(n2672) );
  AOI22_X1 U443 ( .A1(DATAIN[19]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][19] ), .ZN(n336) );
  INV_X1 U444 ( .A(n337), .ZN(n2673) );
  AOI22_X1 U445 ( .A1(DATAIN[20]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][20] ), .ZN(n337) );
  INV_X1 U446 ( .A(n338), .ZN(n2674) );
  AOI22_X1 U447 ( .A1(DATAIN[21]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][21] ), .ZN(n338) );
  INV_X1 U448 ( .A(n339), .ZN(n2675) );
  AOI22_X1 U449 ( .A1(DATAIN[22]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][22] ), .ZN(n339) );
  INV_X1 U450 ( .A(n340), .ZN(n2676) );
  AOI22_X1 U451 ( .A1(DATAIN[23]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][23] ), .ZN(n340) );
  INV_X1 U452 ( .A(n341), .ZN(n2677) );
  AOI22_X1 U453 ( .A1(DATAIN[24]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][24] ), .ZN(n341) );
  INV_X1 U454 ( .A(n342), .ZN(n2678) );
  AOI22_X1 U455 ( .A1(DATAIN[25]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][25] ), .ZN(n342) );
  INV_X1 U456 ( .A(n343), .ZN(n2679) );
  AOI22_X1 U457 ( .A1(DATAIN[26]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][26] ), .ZN(n343) );
  INV_X1 U458 ( .A(n344), .ZN(n2680) );
  AOI22_X1 U459 ( .A1(DATAIN[27]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][27] ), .ZN(n344) );
  INV_X1 U460 ( .A(n345), .ZN(n2681) );
  AOI22_X1 U461 ( .A1(DATAIN[28]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][28] ), .ZN(n345) );
  INV_X1 U462 ( .A(n346), .ZN(n2682) );
  AOI22_X1 U463 ( .A1(DATAIN[29]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][29] ), .ZN(n346) );
  INV_X1 U464 ( .A(n347), .ZN(n2683) );
  AOI22_X1 U465 ( .A1(DATAIN[30]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][30] ), .ZN(n347) );
  INV_X1 U466 ( .A(n348), .ZN(n2684) );
  AOI22_X1 U467 ( .A1(DATAIN[31]), .A2(n316), .B1(n317), .B2(
        \REGISTERS[23][31] ), .ZN(n348) );
  INV_X1 U470 ( .A(n350), .ZN(n2685) );
  AOI22_X1 U471 ( .A1(DATAIN[0]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][0] ), .ZN(n350) );
  INV_X1 U472 ( .A(n353), .ZN(n2686) );
  AOI22_X1 U473 ( .A1(DATAIN[1]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][1] ), .ZN(n353) );
  INV_X1 U474 ( .A(n354), .ZN(n2687) );
  AOI22_X1 U475 ( .A1(DATAIN[2]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][2] ), .ZN(n354) );
  INV_X1 U476 ( .A(n355), .ZN(n2688) );
  AOI22_X1 U477 ( .A1(DATAIN[3]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][3] ), .ZN(n355) );
  INV_X1 U478 ( .A(n356), .ZN(n2689) );
  AOI22_X1 U479 ( .A1(DATAIN[4]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][4] ), .ZN(n356) );
  INV_X1 U480 ( .A(n357), .ZN(n2690) );
  AOI22_X1 U481 ( .A1(DATAIN[5]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][5] ), .ZN(n357) );
  INV_X1 U482 ( .A(n358), .ZN(n2691) );
  AOI22_X1 U483 ( .A1(DATAIN[6]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][6] ), .ZN(n358) );
  INV_X1 U484 ( .A(n359), .ZN(n2692) );
  AOI22_X1 U485 ( .A1(DATAIN[7]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][7] ), .ZN(n359) );
  INV_X1 U486 ( .A(n360), .ZN(n2693) );
  AOI22_X1 U487 ( .A1(DATAIN[8]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][8] ), .ZN(n360) );
  INV_X1 U488 ( .A(n361), .ZN(n2694) );
  AOI22_X1 U489 ( .A1(DATAIN[9]), .A2(n351), .B1(n352), .B2(\REGISTERS[22][9] ), .ZN(n361) );
  INV_X1 U490 ( .A(n362), .ZN(n2695) );
  AOI22_X1 U491 ( .A1(DATAIN[10]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][10] ), .ZN(n362) );
  INV_X1 U492 ( .A(n363), .ZN(n2696) );
  AOI22_X1 U493 ( .A1(DATAIN[11]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][11] ), .ZN(n363) );
  INV_X1 U494 ( .A(n364), .ZN(n2697) );
  AOI22_X1 U495 ( .A1(DATAIN[12]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][12] ), .ZN(n364) );
  INV_X1 U496 ( .A(n365), .ZN(n2698) );
  AOI22_X1 U497 ( .A1(DATAIN[13]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][13] ), .ZN(n365) );
  INV_X1 U498 ( .A(n366), .ZN(n2699) );
  AOI22_X1 U499 ( .A1(DATAIN[14]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][14] ), .ZN(n366) );
  INV_X1 U500 ( .A(n367), .ZN(n2700) );
  AOI22_X1 U501 ( .A1(DATAIN[15]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][15] ), .ZN(n367) );
  INV_X1 U502 ( .A(n368), .ZN(n2701) );
  AOI22_X1 U503 ( .A1(DATAIN[16]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][16] ), .ZN(n368) );
  INV_X1 U504 ( .A(n369), .ZN(n2702) );
  AOI22_X1 U505 ( .A1(DATAIN[17]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][17] ), .ZN(n369) );
  INV_X1 U506 ( .A(n370), .ZN(n2703) );
  AOI22_X1 U507 ( .A1(DATAIN[18]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][18] ), .ZN(n370) );
  INV_X1 U508 ( .A(n371), .ZN(n2704) );
  AOI22_X1 U509 ( .A1(DATAIN[19]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][19] ), .ZN(n371) );
  INV_X1 U510 ( .A(n372), .ZN(n2705) );
  AOI22_X1 U511 ( .A1(DATAIN[20]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][20] ), .ZN(n372) );
  INV_X1 U512 ( .A(n373), .ZN(n2706) );
  AOI22_X1 U513 ( .A1(DATAIN[21]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][21] ), .ZN(n373) );
  INV_X1 U514 ( .A(n374), .ZN(n2707) );
  AOI22_X1 U515 ( .A1(DATAIN[22]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][22] ), .ZN(n374) );
  INV_X1 U516 ( .A(n375), .ZN(n2708) );
  AOI22_X1 U517 ( .A1(DATAIN[23]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][23] ), .ZN(n375) );
  INV_X1 U518 ( .A(n376), .ZN(n2709) );
  AOI22_X1 U519 ( .A1(DATAIN[24]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][24] ), .ZN(n376) );
  INV_X1 U520 ( .A(n377), .ZN(n2710) );
  AOI22_X1 U521 ( .A1(DATAIN[25]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][25] ), .ZN(n377) );
  INV_X1 U522 ( .A(n378), .ZN(n2711) );
  AOI22_X1 U523 ( .A1(DATAIN[26]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][26] ), .ZN(n378) );
  INV_X1 U524 ( .A(n379), .ZN(n2712) );
  AOI22_X1 U525 ( .A1(DATAIN[27]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][27] ), .ZN(n379) );
  INV_X1 U526 ( .A(n380), .ZN(n2713) );
  AOI22_X1 U527 ( .A1(DATAIN[28]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][28] ), .ZN(n380) );
  INV_X1 U528 ( .A(n381), .ZN(n2714) );
  AOI22_X1 U529 ( .A1(DATAIN[29]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][29] ), .ZN(n381) );
  INV_X1 U530 ( .A(n382), .ZN(n2715) );
  AOI22_X1 U531 ( .A1(DATAIN[30]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][30] ), .ZN(n382) );
  INV_X1 U532 ( .A(n383), .ZN(n2716) );
  AOI22_X1 U533 ( .A1(DATAIN[31]), .A2(n351), .B1(n352), .B2(
        \REGISTERS[22][31] ), .ZN(n383) );
  OAI22_X1 U536 ( .A1(n2), .A2(n384), .B1(n385), .B2(n386), .ZN(n2717) );
  OAI22_X1 U537 ( .A1(n5), .A2(n384), .B1(n385), .B2(n387), .ZN(n2718) );
  OAI22_X1 U538 ( .A1(n7), .A2(n384), .B1(n385), .B2(n388), .ZN(n2719) );
  OAI22_X1 U539 ( .A1(n9), .A2(n384), .B1(n385), .B2(n389), .ZN(n2720) );
  OAI22_X1 U540 ( .A1(n11), .A2(n384), .B1(n385), .B2(n390), .ZN(n2721) );
  OAI22_X1 U541 ( .A1(n13), .A2(n384), .B1(n385), .B2(n391), .ZN(n2722) );
  OAI22_X1 U542 ( .A1(n15), .A2(n384), .B1(n385), .B2(n392), .ZN(n2723) );
  OAI22_X1 U543 ( .A1(n17), .A2(n384), .B1(n385), .B2(n393), .ZN(n2724) );
  OAI22_X1 U544 ( .A1(n19), .A2(n384), .B1(n385), .B2(n394), .ZN(n2725) );
  OAI22_X1 U545 ( .A1(n21), .A2(n384), .B1(n385), .B2(n395), .ZN(n2726) );
  OAI22_X1 U546 ( .A1(n23), .A2(n384), .B1(n385), .B2(n396), .ZN(n2727) );
  OAI22_X1 U547 ( .A1(n25), .A2(n384), .B1(n385), .B2(n397), .ZN(n2728) );
  OAI22_X1 U548 ( .A1(n27), .A2(n384), .B1(n385), .B2(n398), .ZN(n2729) );
  OAI22_X1 U549 ( .A1(n29), .A2(n384), .B1(n385), .B2(n399), .ZN(n2730) );
  OAI22_X1 U550 ( .A1(n31), .A2(n384), .B1(n385), .B2(n400), .ZN(n2731) );
  OAI22_X1 U551 ( .A1(n33), .A2(n384), .B1(n385), .B2(n401), .ZN(n2732) );
  OAI22_X1 U552 ( .A1(n35), .A2(n384), .B1(n385), .B2(n402), .ZN(n2733) );
  OAI22_X1 U553 ( .A1(n37), .A2(n384), .B1(n385), .B2(n403), .ZN(n2734) );
  OAI22_X1 U554 ( .A1(n39), .A2(n384), .B1(n385), .B2(n404), .ZN(n2735) );
  OAI22_X1 U555 ( .A1(n41), .A2(n384), .B1(n385), .B2(n405), .ZN(n2736) );
  OAI22_X1 U556 ( .A1(n43), .A2(n384), .B1(n385), .B2(n406), .ZN(n2737) );
  OAI22_X1 U557 ( .A1(n45), .A2(n384), .B1(n385), .B2(n407), .ZN(n2738) );
  OAI22_X1 U558 ( .A1(n47), .A2(n384), .B1(n385), .B2(n408), .ZN(n2739) );
  OAI22_X1 U559 ( .A1(n49), .A2(n384), .B1(n385), .B2(n409), .ZN(n2740) );
  OAI22_X1 U560 ( .A1(n51), .A2(n384), .B1(n385), .B2(n410), .ZN(n2741) );
  OAI22_X1 U561 ( .A1(n53), .A2(n384), .B1(n385), .B2(n411), .ZN(n2742) );
  OAI22_X1 U562 ( .A1(n55), .A2(n384), .B1(n385), .B2(n412), .ZN(n2743) );
  OAI22_X1 U563 ( .A1(n57), .A2(n384), .B1(n385), .B2(n413), .ZN(n2744) );
  OAI22_X1 U564 ( .A1(n59), .A2(n384), .B1(n385), .B2(n414), .ZN(n2745) );
  OAI22_X1 U565 ( .A1(n61), .A2(n384), .B1(n385), .B2(n415), .ZN(n2746) );
  OAI22_X1 U566 ( .A1(n63), .A2(n384), .B1(n385), .B2(n416), .ZN(n2747) );
  OAI22_X1 U567 ( .A1(n65), .A2(n384), .B1(n385), .B2(n417), .ZN(n2748) );
  OAI22_X1 U570 ( .A1(n2), .A2(n418), .B1(n419), .B2(n420), .ZN(n2749) );
  OAI22_X1 U571 ( .A1(n5), .A2(n418), .B1(n419), .B2(n421), .ZN(n2750) );
  OAI22_X1 U572 ( .A1(n7), .A2(n418), .B1(n419), .B2(n422), .ZN(n2751) );
  OAI22_X1 U573 ( .A1(n9), .A2(n418), .B1(n419), .B2(n423), .ZN(n2752) );
  OAI22_X1 U574 ( .A1(n11), .A2(n418), .B1(n419), .B2(n424), .ZN(n2753) );
  OAI22_X1 U575 ( .A1(n13), .A2(n418), .B1(n419), .B2(n425), .ZN(n2754) );
  OAI22_X1 U576 ( .A1(n15), .A2(n418), .B1(n419), .B2(n426), .ZN(n2755) );
  OAI22_X1 U577 ( .A1(n17), .A2(n418), .B1(n419), .B2(n427), .ZN(n2756) );
  OAI22_X1 U578 ( .A1(n19), .A2(n418), .B1(n419), .B2(n428), .ZN(n2757) );
  OAI22_X1 U579 ( .A1(n21), .A2(n418), .B1(n419), .B2(n429), .ZN(n2758) );
  OAI22_X1 U580 ( .A1(n23), .A2(n418), .B1(n419), .B2(n430), .ZN(n2759) );
  OAI22_X1 U581 ( .A1(n25), .A2(n418), .B1(n419), .B2(n431), .ZN(n2760) );
  OAI22_X1 U582 ( .A1(n27), .A2(n418), .B1(n419), .B2(n432), .ZN(n2761) );
  OAI22_X1 U583 ( .A1(n29), .A2(n418), .B1(n419), .B2(n433), .ZN(n2762) );
  OAI22_X1 U584 ( .A1(n31), .A2(n418), .B1(n419), .B2(n434), .ZN(n2763) );
  OAI22_X1 U585 ( .A1(n33), .A2(n418), .B1(n419), .B2(n435), .ZN(n2764) );
  OAI22_X1 U586 ( .A1(n35), .A2(n418), .B1(n419), .B2(n436), .ZN(n2765) );
  OAI22_X1 U587 ( .A1(n37), .A2(n418), .B1(n419), .B2(n437), .ZN(n2766) );
  OAI22_X1 U588 ( .A1(n39), .A2(n418), .B1(n419), .B2(n438), .ZN(n2767) );
  OAI22_X1 U589 ( .A1(n41), .A2(n418), .B1(n419), .B2(n439), .ZN(n2768) );
  OAI22_X1 U590 ( .A1(n43), .A2(n418), .B1(n419), .B2(n440), .ZN(n2769) );
  OAI22_X1 U591 ( .A1(n45), .A2(n418), .B1(n419), .B2(n441), .ZN(n2770) );
  OAI22_X1 U592 ( .A1(n47), .A2(n418), .B1(n419), .B2(n442), .ZN(n2771) );
  OAI22_X1 U593 ( .A1(n49), .A2(n418), .B1(n419), .B2(n443), .ZN(n2772) );
  OAI22_X1 U594 ( .A1(n51), .A2(n418), .B1(n419), .B2(n444), .ZN(n2773) );
  OAI22_X1 U595 ( .A1(n53), .A2(n418), .B1(n419), .B2(n445), .ZN(n2774) );
  OAI22_X1 U596 ( .A1(n55), .A2(n418), .B1(n419), .B2(n446), .ZN(n2775) );
  OAI22_X1 U597 ( .A1(n57), .A2(n418), .B1(n419), .B2(n447), .ZN(n2776) );
  OAI22_X1 U598 ( .A1(n59), .A2(n418), .B1(n419), .B2(n448), .ZN(n2777) );
  OAI22_X1 U599 ( .A1(n61), .A2(n418), .B1(n419), .B2(n449), .ZN(n2778) );
  OAI22_X1 U600 ( .A1(n63), .A2(n418), .B1(n419), .B2(n450), .ZN(n2779) );
  OAI22_X1 U601 ( .A1(n65), .A2(n418), .B1(n419), .B2(n451), .ZN(n2780) );
  INV_X1 U604 ( .A(n452), .ZN(n2781) );
  AOI22_X1 U605 ( .A1(DATAIN[0]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][0] ), .ZN(n452) );
  INV_X1 U606 ( .A(n455), .ZN(n2782) );
  AOI22_X1 U607 ( .A1(DATAIN[1]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][1] ), .ZN(n455) );
  INV_X1 U608 ( .A(n456), .ZN(n2783) );
  AOI22_X1 U609 ( .A1(DATAIN[2]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][2] ), .ZN(n456) );
  INV_X1 U610 ( .A(n457), .ZN(n2784) );
  AOI22_X1 U611 ( .A1(DATAIN[3]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][3] ), .ZN(n457) );
  INV_X1 U612 ( .A(n458), .ZN(n2785) );
  AOI22_X1 U613 ( .A1(DATAIN[4]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][4] ), .ZN(n458) );
  INV_X1 U614 ( .A(n459), .ZN(n2786) );
  AOI22_X1 U615 ( .A1(DATAIN[5]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][5] ), .ZN(n459) );
  INV_X1 U616 ( .A(n460), .ZN(n2787) );
  AOI22_X1 U617 ( .A1(DATAIN[6]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][6] ), .ZN(n460) );
  INV_X1 U618 ( .A(n461), .ZN(n2788) );
  AOI22_X1 U619 ( .A1(DATAIN[7]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][7] ), .ZN(n461) );
  INV_X1 U620 ( .A(n462), .ZN(n2789) );
  AOI22_X1 U621 ( .A1(DATAIN[8]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][8] ), .ZN(n462) );
  INV_X1 U622 ( .A(n463), .ZN(n2790) );
  AOI22_X1 U623 ( .A1(DATAIN[9]), .A2(n453), .B1(n454), .B2(\REGISTERS[19][9] ), .ZN(n463) );
  INV_X1 U624 ( .A(n464), .ZN(n2791) );
  AOI22_X1 U625 ( .A1(DATAIN[10]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][10] ), .ZN(n464) );
  INV_X1 U626 ( .A(n465), .ZN(n2792) );
  AOI22_X1 U627 ( .A1(DATAIN[11]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][11] ), .ZN(n465) );
  INV_X1 U628 ( .A(n466), .ZN(n2793) );
  AOI22_X1 U629 ( .A1(DATAIN[12]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][12] ), .ZN(n466) );
  INV_X1 U630 ( .A(n467), .ZN(n2794) );
  AOI22_X1 U631 ( .A1(DATAIN[13]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][13] ), .ZN(n467) );
  INV_X1 U632 ( .A(n468), .ZN(n2795) );
  AOI22_X1 U633 ( .A1(DATAIN[14]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][14] ), .ZN(n468) );
  INV_X1 U634 ( .A(n469), .ZN(n2796) );
  AOI22_X1 U635 ( .A1(DATAIN[15]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][15] ), .ZN(n469) );
  INV_X1 U636 ( .A(n470), .ZN(n2797) );
  AOI22_X1 U637 ( .A1(DATAIN[16]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][16] ), .ZN(n470) );
  INV_X1 U638 ( .A(n471), .ZN(n2798) );
  AOI22_X1 U639 ( .A1(DATAIN[17]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][17] ), .ZN(n471) );
  INV_X1 U640 ( .A(n472), .ZN(n2799) );
  AOI22_X1 U641 ( .A1(DATAIN[18]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][18] ), .ZN(n472) );
  INV_X1 U642 ( .A(n473), .ZN(n2800) );
  AOI22_X1 U643 ( .A1(DATAIN[19]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][19] ), .ZN(n473) );
  INV_X1 U644 ( .A(n474), .ZN(n2801) );
  AOI22_X1 U645 ( .A1(DATAIN[20]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][20] ), .ZN(n474) );
  INV_X1 U646 ( .A(n475), .ZN(n2802) );
  AOI22_X1 U647 ( .A1(DATAIN[21]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][21] ), .ZN(n475) );
  INV_X1 U648 ( .A(n476), .ZN(n2803) );
  AOI22_X1 U649 ( .A1(DATAIN[22]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][22] ), .ZN(n476) );
  INV_X1 U650 ( .A(n477), .ZN(n2804) );
  AOI22_X1 U651 ( .A1(DATAIN[23]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][23] ), .ZN(n477) );
  INV_X1 U652 ( .A(n478), .ZN(n2805) );
  AOI22_X1 U653 ( .A1(DATAIN[24]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][24] ), .ZN(n478) );
  INV_X1 U654 ( .A(n479), .ZN(n2806) );
  AOI22_X1 U655 ( .A1(DATAIN[25]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][25] ), .ZN(n479) );
  INV_X1 U656 ( .A(n480), .ZN(n2807) );
  AOI22_X1 U657 ( .A1(DATAIN[26]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][26] ), .ZN(n480) );
  INV_X1 U658 ( .A(n481), .ZN(n2808) );
  AOI22_X1 U659 ( .A1(DATAIN[27]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][27] ), .ZN(n481) );
  INV_X1 U660 ( .A(n482), .ZN(n2809) );
  AOI22_X1 U661 ( .A1(DATAIN[28]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][28] ), .ZN(n482) );
  INV_X1 U662 ( .A(n483), .ZN(n2810) );
  AOI22_X1 U663 ( .A1(DATAIN[29]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][29] ), .ZN(n483) );
  INV_X1 U664 ( .A(n484), .ZN(n2811) );
  AOI22_X1 U665 ( .A1(DATAIN[30]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][30] ), .ZN(n484) );
  INV_X1 U666 ( .A(n485), .ZN(n2812) );
  AOI22_X1 U667 ( .A1(DATAIN[31]), .A2(n453), .B1(n454), .B2(
        \REGISTERS[19][31] ), .ZN(n485) );
  INV_X1 U670 ( .A(n486), .ZN(n2813) );
  AOI22_X1 U671 ( .A1(DATAIN[0]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][0] ), .ZN(n486) );
  INV_X1 U672 ( .A(n489), .ZN(n2814) );
  AOI22_X1 U673 ( .A1(DATAIN[1]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][1] ), .ZN(n489) );
  INV_X1 U674 ( .A(n490), .ZN(n2815) );
  AOI22_X1 U675 ( .A1(DATAIN[2]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][2] ), .ZN(n490) );
  INV_X1 U676 ( .A(n491), .ZN(n2816) );
  AOI22_X1 U677 ( .A1(DATAIN[3]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][3] ), .ZN(n491) );
  INV_X1 U678 ( .A(n492), .ZN(n2817) );
  AOI22_X1 U679 ( .A1(DATAIN[4]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][4] ), .ZN(n492) );
  INV_X1 U680 ( .A(n493), .ZN(n2818) );
  AOI22_X1 U681 ( .A1(DATAIN[5]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][5] ), .ZN(n493) );
  INV_X1 U682 ( .A(n494), .ZN(n2819) );
  AOI22_X1 U683 ( .A1(DATAIN[6]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][6] ), .ZN(n494) );
  INV_X1 U684 ( .A(n495), .ZN(n2820) );
  AOI22_X1 U685 ( .A1(DATAIN[7]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][7] ), .ZN(n495) );
  INV_X1 U686 ( .A(n496), .ZN(n2821) );
  AOI22_X1 U687 ( .A1(DATAIN[8]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][8] ), .ZN(n496) );
  INV_X1 U688 ( .A(n497), .ZN(n2822) );
  AOI22_X1 U689 ( .A1(DATAIN[9]), .A2(n487), .B1(n488), .B2(\REGISTERS[18][9] ), .ZN(n497) );
  INV_X1 U690 ( .A(n498), .ZN(n2823) );
  AOI22_X1 U691 ( .A1(DATAIN[10]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][10] ), .ZN(n498) );
  INV_X1 U692 ( .A(n499), .ZN(n2824) );
  AOI22_X1 U693 ( .A1(DATAIN[11]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][11] ), .ZN(n499) );
  INV_X1 U694 ( .A(n500), .ZN(n2825) );
  AOI22_X1 U695 ( .A1(DATAIN[12]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][12] ), .ZN(n500) );
  INV_X1 U696 ( .A(n501), .ZN(n2826) );
  AOI22_X1 U697 ( .A1(DATAIN[13]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][13] ), .ZN(n501) );
  INV_X1 U698 ( .A(n502), .ZN(n2827) );
  AOI22_X1 U699 ( .A1(DATAIN[14]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][14] ), .ZN(n502) );
  INV_X1 U700 ( .A(n503), .ZN(n2828) );
  AOI22_X1 U701 ( .A1(DATAIN[15]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][15] ), .ZN(n503) );
  INV_X1 U702 ( .A(n504), .ZN(n2829) );
  AOI22_X1 U703 ( .A1(DATAIN[16]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][16] ), .ZN(n504) );
  INV_X1 U704 ( .A(n505), .ZN(n2830) );
  AOI22_X1 U705 ( .A1(DATAIN[17]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][17] ), .ZN(n505) );
  INV_X1 U706 ( .A(n506), .ZN(n2831) );
  AOI22_X1 U707 ( .A1(DATAIN[18]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][18] ), .ZN(n506) );
  INV_X1 U708 ( .A(n507), .ZN(n2832) );
  AOI22_X1 U709 ( .A1(DATAIN[19]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][19] ), .ZN(n507) );
  INV_X1 U710 ( .A(n508), .ZN(n2833) );
  AOI22_X1 U711 ( .A1(DATAIN[20]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][20] ), .ZN(n508) );
  INV_X1 U712 ( .A(n509), .ZN(n2834) );
  AOI22_X1 U713 ( .A1(DATAIN[21]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][21] ), .ZN(n509) );
  INV_X1 U714 ( .A(n510), .ZN(n2835) );
  AOI22_X1 U715 ( .A1(DATAIN[22]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][22] ), .ZN(n510) );
  INV_X1 U716 ( .A(n511), .ZN(n2836) );
  AOI22_X1 U717 ( .A1(DATAIN[23]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][23] ), .ZN(n511) );
  INV_X1 U718 ( .A(n512), .ZN(n2837) );
  AOI22_X1 U719 ( .A1(DATAIN[24]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][24] ), .ZN(n512) );
  INV_X1 U720 ( .A(n513), .ZN(n2838) );
  AOI22_X1 U721 ( .A1(DATAIN[25]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][25] ), .ZN(n513) );
  INV_X1 U722 ( .A(n514), .ZN(n2839) );
  AOI22_X1 U723 ( .A1(DATAIN[26]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][26] ), .ZN(n514) );
  INV_X1 U724 ( .A(n515), .ZN(n2840) );
  AOI22_X1 U725 ( .A1(DATAIN[27]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][27] ), .ZN(n515) );
  INV_X1 U726 ( .A(n516), .ZN(n2841) );
  AOI22_X1 U727 ( .A1(DATAIN[28]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][28] ), .ZN(n516) );
  INV_X1 U728 ( .A(n517), .ZN(n2842) );
  AOI22_X1 U729 ( .A1(DATAIN[29]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][29] ), .ZN(n517) );
  INV_X1 U730 ( .A(n518), .ZN(n2843) );
  AOI22_X1 U731 ( .A1(DATAIN[30]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][30] ), .ZN(n518) );
  INV_X1 U732 ( .A(n519), .ZN(n2844) );
  AOI22_X1 U733 ( .A1(DATAIN[31]), .A2(n487), .B1(n488), .B2(
        \REGISTERS[18][31] ), .ZN(n519) );
  OAI22_X1 U736 ( .A1(n2), .A2(n520), .B1(n521), .B2(n522), .ZN(n2845) );
  OAI22_X1 U737 ( .A1(n5), .A2(n520), .B1(n521), .B2(n523), .ZN(n2846) );
  OAI22_X1 U738 ( .A1(n7), .A2(n520), .B1(n521), .B2(n524), .ZN(n2847) );
  OAI22_X1 U739 ( .A1(n9), .A2(n520), .B1(n521), .B2(n525), .ZN(n2848) );
  OAI22_X1 U740 ( .A1(n11), .A2(n520), .B1(n521), .B2(n526), .ZN(n2849) );
  OAI22_X1 U741 ( .A1(n13), .A2(n520), .B1(n521), .B2(n527), .ZN(n2850) );
  OAI22_X1 U742 ( .A1(n15), .A2(n520), .B1(n521), .B2(n528), .ZN(n2851) );
  OAI22_X1 U743 ( .A1(n17), .A2(n520), .B1(n521), .B2(n529), .ZN(n2852) );
  OAI22_X1 U744 ( .A1(n19), .A2(n520), .B1(n521), .B2(n530), .ZN(n2853) );
  OAI22_X1 U745 ( .A1(n21), .A2(n520), .B1(n521), .B2(n531), .ZN(n2854) );
  OAI22_X1 U746 ( .A1(n23), .A2(n520), .B1(n521), .B2(n532), .ZN(n2855) );
  OAI22_X1 U747 ( .A1(n25), .A2(n520), .B1(n521), .B2(n533), .ZN(n2856) );
  OAI22_X1 U748 ( .A1(n27), .A2(n520), .B1(n521), .B2(n534), .ZN(n2857) );
  OAI22_X1 U749 ( .A1(n29), .A2(n520), .B1(n521), .B2(n535), .ZN(n2858) );
  OAI22_X1 U750 ( .A1(n31), .A2(n520), .B1(n521), .B2(n536), .ZN(n2859) );
  OAI22_X1 U751 ( .A1(n33), .A2(n520), .B1(n521), .B2(n537), .ZN(n2860) );
  OAI22_X1 U752 ( .A1(n35), .A2(n520), .B1(n521), .B2(n538), .ZN(n2861) );
  OAI22_X1 U753 ( .A1(n37), .A2(n520), .B1(n521), .B2(n539), .ZN(n2862) );
  OAI22_X1 U754 ( .A1(n39), .A2(n520), .B1(n521), .B2(n540), .ZN(n2863) );
  OAI22_X1 U755 ( .A1(n41), .A2(n520), .B1(n521), .B2(n541), .ZN(n2864) );
  OAI22_X1 U756 ( .A1(n43), .A2(n520), .B1(n521), .B2(n542), .ZN(n2865) );
  OAI22_X1 U757 ( .A1(n45), .A2(n520), .B1(n521), .B2(n543), .ZN(n2866) );
  OAI22_X1 U758 ( .A1(n47), .A2(n520), .B1(n521), .B2(n544), .ZN(n2867) );
  OAI22_X1 U759 ( .A1(n49), .A2(n520), .B1(n521), .B2(n545), .ZN(n2868) );
  OAI22_X1 U760 ( .A1(n51), .A2(n520), .B1(n521), .B2(n546), .ZN(n2869) );
  OAI22_X1 U761 ( .A1(n53), .A2(n520), .B1(n521), .B2(n547), .ZN(n2870) );
  OAI22_X1 U762 ( .A1(n55), .A2(n520), .B1(n521), .B2(n548), .ZN(n2871) );
  OAI22_X1 U763 ( .A1(n57), .A2(n520), .B1(n521), .B2(n549), .ZN(n2872) );
  OAI22_X1 U764 ( .A1(n59), .A2(n520), .B1(n521), .B2(n550), .ZN(n2873) );
  OAI22_X1 U765 ( .A1(n61), .A2(n520), .B1(n521), .B2(n551), .ZN(n2874) );
  OAI22_X1 U766 ( .A1(n63), .A2(n520), .B1(n521), .B2(n552), .ZN(n2875) );
  OAI22_X1 U767 ( .A1(n65), .A2(n520), .B1(n521), .B2(n553), .ZN(n2876) );
  OAI22_X1 U770 ( .A1(n2), .A2(n554), .B1(n555), .B2(n556), .ZN(n2877) );
  OAI22_X1 U771 ( .A1(n5), .A2(n554), .B1(n555), .B2(n557), .ZN(n2878) );
  OAI22_X1 U772 ( .A1(n7), .A2(n554), .B1(n555), .B2(n558), .ZN(n2879) );
  OAI22_X1 U773 ( .A1(n9), .A2(n554), .B1(n555), .B2(n559), .ZN(n2880) );
  OAI22_X1 U774 ( .A1(n11), .A2(n554), .B1(n555), .B2(n560), .ZN(n2881) );
  OAI22_X1 U775 ( .A1(n13), .A2(n554), .B1(n555), .B2(n561), .ZN(n2882) );
  OAI22_X1 U776 ( .A1(n15), .A2(n554), .B1(n555), .B2(n562), .ZN(n2883) );
  OAI22_X1 U777 ( .A1(n17), .A2(n554), .B1(n555), .B2(n563), .ZN(n2884) );
  OAI22_X1 U778 ( .A1(n19), .A2(n554), .B1(n555), .B2(n564), .ZN(n2885) );
  OAI22_X1 U779 ( .A1(n21), .A2(n554), .B1(n555), .B2(n565), .ZN(n2886) );
  OAI22_X1 U780 ( .A1(n23), .A2(n554), .B1(n555), .B2(n566), .ZN(n2887) );
  OAI22_X1 U781 ( .A1(n25), .A2(n554), .B1(n555), .B2(n567), .ZN(n2888) );
  OAI22_X1 U782 ( .A1(n27), .A2(n554), .B1(n555), .B2(n568), .ZN(n2889) );
  OAI22_X1 U783 ( .A1(n29), .A2(n554), .B1(n555), .B2(n569), .ZN(n2890) );
  OAI22_X1 U784 ( .A1(n31), .A2(n554), .B1(n555), .B2(n570), .ZN(n2891) );
  OAI22_X1 U785 ( .A1(n33), .A2(n554), .B1(n555), .B2(n571), .ZN(n2892) );
  OAI22_X1 U786 ( .A1(n35), .A2(n554), .B1(n555), .B2(n572), .ZN(n2893) );
  OAI22_X1 U787 ( .A1(n37), .A2(n554), .B1(n555), .B2(n573), .ZN(n2894) );
  OAI22_X1 U788 ( .A1(n39), .A2(n554), .B1(n555), .B2(n574), .ZN(n2895) );
  OAI22_X1 U789 ( .A1(n41), .A2(n554), .B1(n555), .B2(n575), .ZN(n2896) );
  OAI22_X1 U790 ( .A1(n43), .A2(n554), .B1(n555), .B2(n576), .ZN(n2897) );
  OAI22_X1 U791 ( .A1(n45), .A2(n554), .B1(n555), .B2(n577), .ZN(n2898) );
  OAI22_X1 U792 ( .A1(n47), .A2(n554), .B1(n555), .B2(n578), .ZN(n2899) );
  OAI22_X1 U793 ( .A1(n49), .A2(n554), .B1(n555), .B2(n579), .ZN(n2900) );
  OAI22_X1 U794 ( .A1(n51), .A2(n554), .B1(n555), .B2(n580), .ZN(n2901) );
  OAI22_X1 U795 ( .A1(n53), .A2(n554), .B1(n555), .B2(n581), .ZN(n2902) );
  OAI22_X1 U796 ( .A1(n55), .A2(n554), .B1(n555), .B2(n582), .ZN(n2903) );
  OAI22_X1 U797 ( .A1(n57), .A2(n554), .B1(n555), .B2(n583), .ZN(n2904) );
  OAI22_X1 U798 ( .A1(n59), .A2(n554), .B1(n555), .B2(n584), .ZN(n2905) );
  OAI22_X1 U799 ( .A1(n61), .A2(n554), .B1(n555), .B2(n585), .ZN(n2906) );
  OAI22_X1 U800 ( .A1(n63), .A2(n554), .B1(n555), .B2(n586), .ZN(n2907) );
  OAI22_X1 U801 ( .A1(n65), .A2(n554), .B1(n555), .B2(n587), .ZN(n2908) );
  AND3_X1 U804 ( .A1(n314), .A2(n588), .A3(ADD_WR[4]), .ZN(n349) );
  INV_X1 U805 ( .A(n589), .ZN(n2909) );
  AOI22_X1 U806 ( .A1(DATAIN[0]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][0] ), .ZN(n589) );
  INV_X1 U807 ( .A(n592), .ZN(n2910) );
  AOI22_X1 U808 ( .A1(DATAIN[1]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][1] ), .ZN(n592) );
  INV_X1 U809 ( .A(n593), .ZN(n2911) );
  AOI22_X1 U810 ( .A1(DATAIN[2]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][2] ), .ZN(n593) );
  INV_X1 U811 ( .A(n594), .ZN(n2912) );
  AOI22_X1 U812 ( .A1(DATAIN[3]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][3] ), .ZN(n594) );
  INV_X1 U813 ( .A(n595), .ZN(n2913) );
  AOI22_X1 U814 ( .A1(DATAIN[4]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][4] ), .ZN(n595) );
  INV_X1 U815 ( .A(n596), .ZN(n2914) );
  AOI22_X1 U816 ( .A1(DATAIN[5]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][5] ), .ZN(n596) );
  INV_X1 U817 ( .A(n597), .ZN(n2915) );
  AOI22_X1 U818 ( .A1(DATAIN[6]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][6] ), .ZN(n597) );
  INV_X1 U819 ( .A(n598), .ZN(n2916) );
  AOI22_X1 U820 ( .A1(DATAIN[7]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][7] ), .ZN(n598) );
  INV_X1 U821 ( .A(n599), .ZN(n2917) );
  AOI22_X1 U822 ( .A1(DATAIN[8]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][8] ), .ZN(n599) );
  INV_X1 U823 ( .A(n600), .ZN(n2918) );
  AOI22_X1 U824 ( .A1(DATAIN[9]), .A2(n590), .B1(n591), .B2(\REGISTERS[15][9] ), .ZN(n600) );
  INV_X1 U825 ( .A(n601), .ZN(n2919) );
  AOI22_X1 U826 ( .A1(DATAIN[10]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][10] ), .ZN(n601) );
  INV_X1 U827 ( .A(n602), .ZN(n2920) );
  AOI22_X1 U828 ( .A1(DATAIN[11]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][11] ), .ZN(n602) );
  INV_X1 U829 ( .A(n603), .ZN(n2921) );
  AOI22_X1 U830 ( .A1(DATAIN[12]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][12] ), .ZN(n603) );
  INV_X1 U831 ( .A(n604), .ZN(n2922) );
  AOI22_X1 U832 ( .A1(DATAIN[13]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][13] ), .ZN(n604) );
  INV_X1 U833 ( .A(n605), .ZN(n2923) );
  AOI22_X1 U834 ( .A1(DATAIN[14]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][14] ), .ZN(n605) );
  INV_X1 U835 ( .A(n606), .ZN(n2924) );
  AOI22_X1 U836 ( .A1(DATAIN[15]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][15] ), .ZN(n606) );
  INV_X1 U837 ( .A(n607), .ZN(n2925) );
  AOI22_X1 U838 ( .A1(DATAIN[16]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][16] ), .ZN(n607) );
  INV_X1 U839 ( .A(n608), .ZN(n2926) );
  AOI22_X1 U840 ( .A1(DATAIN[17]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][17] ), .ZN(n608) );
  INV_X1 U841 ( .A(n609), .ZN(n2927) );
  AOI22_X1 U842 ( .A1(DATAIN[18]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][18] ), .ZN(n609) );
  INV_X1 U843 ( .A(n610), .ZN(n2928) );
  AOI22_X1 U844 ( .A1(DATAIN[19]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][19] ), .ZN(n610) );
  INV_X1 U845 ( .A(n611), .ZN(n2929) );
  AOI22_X1 U846 ( .A1(DATAIN[20]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][20] ), .ZN(n611) );
  INV_X1 U847 ( .A(n612), .ZN(n2930) );
  AOI22_X1 U848 ( .A1(DATAIN[21]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][21] ), .ZN(n612) );
  INV_X1 U849 ( .A(n613), .ZN(n2931) );
  AOI22_X1 U850 ( .A1(DATAIN[22]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][22] ), .ZN(n613) );
  INV_X1 U851 ( .A(n614), .ZN(n2932) );
  AOI22_X1 U852 ( .A1(DATAIN[23]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][23] ), .ZN(n614) );
  INV_X1 U853 ( .A(n615), .ZN(n2933) );
  AOI22_X1 U854 ( .A1(DATAIN[24]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][24] ), .ZN(n615) );
  INV_X1 U855 ( .A(n616), .ZN(n2934) );
  AOI22_X1 U856 ( .A1(DATAIN[25]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][25] ), .ZN(n616) );
  INV_X1 U857 ( .A(n617), .ZN(n2935) );
  AOI22_X1 U858 ( .A1(DATAIN[26]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][26] ), .ZN(n617) );
  INV_X1 U859 ( .A(n618), .ZN(n2936) );
  AOI22_X1 U860 ( .A1(DATAIN[27]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][27] ), .ZN(n618) );
  INV_X1 U861 ( .A(n619), .ZN(n2937) );
  AOI22_X1 U862 ( .A1(DATAIN[28]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][28] ), .ZN(n619) );
  INV_X1 U863 ( .A(n620), .ZN(n2938) );
  AOI22_X1 U864 ( .A1(DATAIN[29]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][29] ), .ZN(n620) );
  INV_X1 U865 ( .A(n621), .ZN(n2939) );
  AOI22_X1 U866 ( .A1(DATAIN[30]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][30] ), .ZN(n621) );
  INV_X1 U867 ( .A(n622), .ZN(n2940) );
  AOI22_X1 U868 ( .A1(DATAIN[31]), .A2(n590), .B1(n591), .B2(
        \REGISTERS[15][31] ), .ZN(n622) );
  INV_X1 U871 ( .A(n624), .ZN(n2941) );
  AOI22_X1 U872 ( .A1(DATAIN[0]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][0] ), .ZN(n624) );
  INV_X1 U873 ( .A(n627), .ZN(n2942) );
  AOI22_X1 U874 ( .A1(DATAIN[1]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][1] ), .ZN(n627) );
  INV_X1 U875 ( .A(n628), .ZN(n2943) );
  AOI22_X1 U876 ( .A1(DATAIN[2]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][2] ), .ZN(n628) );
  INV_X1 U877 ( .A(n629), .ZN(n2944) );
  AOI22_X1 U878 ( .A1(DATAIN[3]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][3] ), .ZN(n629) );
  INV_X1 U879 ( .A(n630), .ZN(n2945) );
  AOI22_X1 U880 ( .A1(DATAIN[4]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][4] ), .ZN(n630) );
  INV_X1 U881 ( .A(n631), .ZN(n2946) );
  AOI22_X1 U882 ( .A1(DATAIN[5]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][5] ), .ZN(n631) );
  INV_X1 U883 ( .A(n632), .ZN(n2947) );
  AOI22_X1 U884 ( .A1(DATAIN[6]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][6] ), .ZN(n632) );
  INV_X1 U885 ( .A(n633), .ZN(n2948) );
  AOI22_X1 U886 ( .A1(DATAIN[7]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][7] ), .ZN(n633) );
  INV_X1 U887 ( .A(n634), .ZN(n2949) );
  AOI22_X1 U888 ( .A1(DATAIN[8]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][8] ), .ZN(n634) );
  INV_X1 U889 ( .A(n635), .ZN(n2950) );
  AOI22_X1 U890 ( .A1(DATAIN[9]), .A2(n625), .B1(n626), .B2(\REGISTERS[14][9] ), .ZN(n635) );
  INV_X1 U891 ( .A(n636), .ZN(n2951) );
  AOI22_X1 U892 ( .A1(DATAIN[10]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][10] ), .ZN(n636) );
  INV_X1 U893 ( .A(n637), .ZN(n2952) );
  AOI22_X1 U894 ( .A1(DATAIN[11]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][11] ), .ZN(n637) );
  INV_X1 U895 ( .A(n638), .ZN(n2953) );
  AOI22_X1 U896 ( .A1(DATAIN[12]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][12] ), .ZN(n638) );
  INV_X1 U897 ( .A(n639), .ZN(n2954) );
  AOI22_X1 U898 ( .A1(DATAIN[13]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][13] ), .ZN(n639) );
  INV_X1 U899 ( .A(n640), .ZN(n2955) );
  AOI22_X1 U900 ( .A1(DATAIN[14]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][14] ), .ZN(n640) );
  INV_X1 U901 ( .A(n641), .ZN(n2956) );
  AOI22_X1 U902 ( .A1(DATAIN[15]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][15] ), .ZN(n641) );
  INV_X1 U903 ( .A(n642), .ZN(n2957) );
  AOI22_X1 U904 ( .A1(DATAIN[16]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][16] ), .ZN(n642) );
  INV_X1 U905 ( .A(n643), .ZN(n2958) );
  AOI22_X1 U906 ( .A1(DATAIN[17]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][17] ), .ZN(n643) );
  INV_X1 U907 ( .A(n644), .ZN(n2959) );
  AOI22_X1 U908 ( .A1(DATAIN[18]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][18] ), .ZN(n644) );
  INV_X1 U909 ( .A(n645), .ZN(n2960) );
  AOI22_X1 U910 ( .A1(DATAIN[19]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][19] ), .ZN(n645) );
  INV_X1 U911 ( .A(n646), .ZN(n2961) );
  AOI22_X1 U912 ( .A1(DATAIN[20]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][20] ), .ZN(n646) );
  INV_X1 U913 ( .A(n647), .ZN(n2962) );
  AOI22_X1 U914 ( .A1(DATAIN[21]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][21] ), .ZN(n647) );
  INV_X1 U915 ( .A(n648), .ZN(n2963) );
  AOI22_X1 U916 ( .A1(DATAIN[22]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][22] ), .ZN(n648) );
  INV_X1 U917 ( .A(n649), .ZN(n2964) );
  AOI22_X1 U918 ( .A1(DATAIN[23]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][23] ), .ZN(n649) );
  INV_X1 U919 ( .A(n650), .ZN(n2965) );
  AOI22_X1 U920 ( .A1(DATAIN[24]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][24] ), .ZN(n650) );
  INV_X1 U921 ( .A(n651), .ZN(n2966) );
  AOI22_X1 U922 ( .A1(DATAIN[25]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][25] ), .ZN(n651) );
  INV_X1 U923 ( .A(n652), .ZN(n2967) );
  AOI22_X1 U924 ( .A1(DATAIN[26]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][26] ), .ZN(n652) );
  INV_X1 U925 ( .A(n653), .ZN(n2968) );
  AOI22_X1 U926 ( .A1(DATAIN[27]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][27] ), .ZN(n653) );
  INV_X1 U927 ( .A(n654), .ZN(n2969) );
  AOI22_X1 U928 ( .A1(DATAIN[28]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][28] ), .ZN(n654) );
  INV_X1 U929 ( .A(n655), .ZN(n2970) );
  AOI22_X1 U930 ( .A1(DATAIN[29]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][29] ), .ZN(n655) );
  INV_X1 U931 ( .A(n656), .ZN(n2971) );
  AOI22_X1 U932 ( .A1(DATAIN[30]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][30] ), .ZN(n656) );
  INV_X1 U933 ( .A(n657), .ZN(n2972) );
  AOI22_X1 U934 ( .A1(DATAIN[31]), .A2(n625), .B1(n626), .B2(
        \REGISTERS[14][31] ), .ZN(n657) );
  OAI22_X1 U937 ( .A1(n2), .A2(n658), .B1(n659), .B2(n660), .ZN(n2973) );
  OAI22_X1 U938 ( .A1(n5), .A2(n658), .B1(n659), .B2(n661), .ZN(n2974) );
  OAI22_X1 U939 ( .A1(n7), .A2(n658), .B1(n659), .B2(n662), .ZN(n2975) );
  OAI22_X1 U940 ( .A1(n9), .A2(n658), .B1(n659), .B2(n663), .ZN(n2976) );
  OAI22_X1 U941 ( .A1(n11), .A2(n658), .B1(n659), .B2(n664), .ZN(n2977) );
  OAI22_X1 U942 ( .A1(n13), .A2(n658), .B1(n659), .B2(n665), .ZN(n2978) );
  OAI22_X1 U943 ( .A1(n15), .A2(n658), .B1(n659), .B2(n666), .ZN(n2979) );
  OAI22_X1 U944 ( .A1(n17), .A2(n658), .B1(n659), .B2(n667), .ZN(n2980) );
  OAI22_X1 U945 ( .A1(n19), .A2(n658), .B1(n659), .B2(n668), .ZN(n2981) );
  OAI22_X1 U946 ( .A1(n21), .A2(n658), .B1(n659), .B2(n669), .ZN(n2982) );
  OAI22_X1 U947 ( .A1(n23), .A2(n658), .B1(n659), .B2(n670), .ZN(n2983) );
  OAI22_X1 U948 ( .A1(n25), .A2(n658), .B1(n659), .B2(n671), .ZN(n2984) );
  OAI22_X1 U949 ( .A1(n27), .A2(n658), .B1(n659), .B2(n672), .ZN(n2985) );
  OAI22_X1 U950 ( .A1(n29), .A2(n658), .B1(n659), .B2(n673), .ZN(n2986) );
  OAI22_X1 U951 ( .A1(n31), .A2(n658), .B1(n659), .B2(n674), .ZN(n2987) );
  OAI22_X1 U952 ( .A1(n33), .A2(n658), .B1(n659), .B2(n675), .ZN(n2988) );
  OAI22_X1 U953 ( .A1(n35), .A2(n658), .B1(n659), .B2(n676), .ZN(n2989) );
  OAI22_X1 U954 ( .A1(n37), .A2(n658), .B1(n659), .B2(n677), .ZN(n2990) );
  OAI22_X1 U955 ( .A1(n39), .A2(n658), .B1(n659), .B2(n678), .ZN(n2991) );
  OAI22_X1 U956 ( .A1(n41), .A2(n658), .B1(n659), .B2(n679), .ZN(n2992) );
  OAI22_X1 U957 ( .A1(n43), .A2(n658), .B1(n659), .B2(n680), .ZN(n2993) );
  OAI22_X1 U958 ( .A1(n45), .A2(n658), .B1(n659), .B2(n681), .ZN(n2994) );
  OAI22_X1 U959 ( .A1(n47), .A2(n658), .B1(n659), .B2(n682), .ZN(n2995) );
  OAI22_X1 U960 ( .A1(n49), .A2(n658), .B1(n659), .B2(n683), .ZN(n2996) );
  OAI22_X1 U961 ( .A1(n51), .A2(n658), .B1(n659), .B2(n684), .ZN(n2997) );
  OAI22_X1 U962 ( .A1(n53), .A2(n658), .B1(n659), .B2(n685), .ZN(n2998) );
  OAI22_X1 U963 ( .A1(n55), .A2(n658), .B1(n659), .B2(n686), .ZN(n2999) );
  OAI22_X1 U964 ( .A1(n57), .A2(n658), .B1(n659), .B2(n687), .ZN(n3000) );
  OAI22_X1 U965 ( .A1(n59), .A2(n658), .B1(n659), .B2(n688), .ZN(n3001) );
  OAI22_X1 U966 ( .A1(n61), .A2(n658), .B1(n659), .B2(n689), .ZN(n3002) );
  OAI22_X1 U967 ( .A1(n63), .A2(n658), .B1(n659), .B2(n690), .ZN(n3003) );
  OAI22_X1 U968 ( .A1(n65), .A2(n658), .B1(n659), .B2(n691), .ZN(n3004) );
  OAI22_X1 U971 ( .A1(n2), .A2(n692), .B1(n693), .B2(n694), .ZN(n3005) );
  OAI22_X1 U972 ( .A1(n5), .A2(n692), .B1(n693), .B2(n695), .ZN(n3006) );
  OAI22_X1 U973 ( .A1(n7), .A2(n692), .B1(n693), .B2(n696), .ZN(n3007) );
  OAI22_X1 U974 ( .A1(n9), .A2(n692), .B1(n693), .B2(n697), .ZN(n3008) );
  OAI22_X1 U975 ( .A1(n11), .A2(n692), .B1(n693), .B2(n698), .ZN(n3009) );
  OAI22_X1 U976 ( .A1(n13), .A2(n692), .B1(n693), .B2(n699), .ZN(n3010) );
  OAI22_X1 U977 ( .A1(n15), .A2(n692), .B1(n693), .B2(n700), .ZN(n3011) );
  OAI22_X1 U978 ( .A1(n17), .A2(n692), .B1(n693), .B2(n701), .ZN(n3012) );
  OAI22_X1 U979 ( .A1(n19), .A2(n692), .B1(n693), .B2(n702), .ZN(n3013) );
  OAI22_X1 U980 ( .A1(n21), .A2(n692), .B1(n693), .B2(n703), .ZN(n3014) );
  OAI22_X1 U981 ( .A1(n23), .A2(n692), .B1(n693), .B2(n704), .ZN(n3015) );
  OAI22_X1 U982 ( .A1(n25), .A2(n692), .B1(n693), .B2(n705), .ZN(n3016) );
  OAI22_X1 U983 ( .A1(n27), .A2(n692), .B1(n693), .B2(n706), .ZN(n3017) );
  OAI22_X1 U984 ( .A1(n29), .A2(n692), .B1(n693), .B2(n707), .ZN(n3018) );
  OAI22_X1 U985 ( .A1(n31), .A2(n692), .B1(n693), .B2(n708), .ZN(n3019) );
  OAI22_X1 U986 ( .A1(n33), .A2(n692), .B1(n693), .B2(n709), .ZN(n3020) );
  OAI22_X1 U987 ( .A1(n35), .A2(n692), .B1(n693), .B2(n710), .ZN(n3021) );
  OAI22_X1 U988 ( .A1(n37), .A2(n692), .B1(n693), .B2(n711), .ZN(n3022) );
  OAI22_X1 U989 ( .A1(n39), .A2(n692), .B1(n693), .B2(n712), .ZN(n3023) );
  OAI22_X1 U990 ( .A1(n41), .A2(n692), .B1(n693), .B2(n713), .ZN(n3024) );
  OAI22_X1 U991 ( .A1(n43), .A2(n692), .B1(n693), .B2(n714), .ZN(n3025) );
  OAI22_X1 U992 ( .A1(n45), .A2(n692), .B1(n693), .B2(n715), .ZN(n3026) );
  OAI22_X1 U993 ( .A1(n47), .A2(n692), .B1(n693), .B2(n716), .ZN(n3027) );
  OAI22_X1 U994 ( .A1(n49), .A2(n692), .B1(n693), .B2(n717), .ZN(n3028) );
  OAI22_X1 U995 ( .A1(n51), .A2(n692), .B1(n693), .B2(n718), .ZN(n3029) );
  OAI22_X1 U996 ( .A1(n53), .A2(n692), .B1(n693), .B2(n719), .ZN(n3030) );
  OAI22_X1 U997 ( .A1(n55), .A2(n692), .B1(n693), .B2(n720), .ZN(n3031) );
  OAI22_X1 U998 ( .A1(n57), .A2(n692), .B1(n693), .B2(n721), .ZN(n3032) );
  OAI22_X1 U999 ( .A1(n59), .A2(n692), .B1(n693), .B2(n722), .ZN(n3033) );
  OAI22_X1 U1000 ( .A1(n61), .A2(n692), .B1(n693), .B2(n723), .ZN(n3034) );
  OAI22_X1 U1001 ( .A1(n63), .A2(n692), .B1(n693), .B2(n724), .ZN(n3035) );
  OAI22_X1 U1002 ( .A1(n65), .A2(n692), .B1(n693), .B2(n725), .ZN(n3036) );
  INV_X1 U1005 ( .A(n726), .ZN(n3037) );
  AOI22_X1 U1006 ( .A1(DATAIN[0]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][0] ), .ZN(n726) );
  INV_X1 U1007 ( .A(n729), .ZN(n3038) );
  AOI22_X1 U1008 ( .A1(DATAIN[1]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][1] ), .ZN(n729) );
  INV_X1 U1009 ( .A(n730), .ZN(n3039) );
  AOI22_X1 U1010 ( .A1(DATAIN[2]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][2] ), .ZN(n730) );
  INV_X1 U1011 ( .A(n731), .ZN(n3040) );
  AOI22_X1 U1012 ( .A1(DATAIN[3]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][3] ), .ZN(n731) );
  INV_X1 U1013 ( .A(n732), .ZN(n3041) );
  AOI22_X1 U1014 ( .A1(DATAIN[4]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][4] ), .ZN(n732) );
  INV_X1 U1015 ( .A(n733), .ZN(n3042) );
  AOI22_X1 U1016 ( .A1(DATAIN[5]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][5] ), .ZN(n733) );
  INV_X1 U1017 ( .A(n734), .ZN(n3043) );
  AOI22_X1 U1018 ( .A1(DATAIN[6]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][6] ), .ZN(n734) );
  INV_X1 U1019 ( .A(n735), .ZN(n3044) );
  AOI22_X1 U1020 ( .A1(DATAIN[7]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][7] ), .ZN(n735) );
  INV_X1 U1021 ( .A(n736), .ZN(n3045) );
  AOI22_X1 U1022 ( .A1(DATAIN[8]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][8] ), .ZN(n736) );
  INV_X1 U1023 ( .A(n737), .ZN(n3046) );
  AOI22_X1 U1024 ( .A1(DATAIN[9]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][9] ), .ZN(n737) );
  INV_X1 U1025 ( .A(n738), .ZN(n3047) );
  AOI22_X1 U1026 ( .A1(DATAIN[10]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][10] ), .ZN(n738) );
  INV_X1 U1027 ( .A(n739), .ZN(n3048) );
  AOI22_X1 U1028 ( .A1(DATAIN[11]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][11] ), .ZN(n739) );
  INV_X1 U1029 ( .A(n740), .ZN(n3049) );
  AOI22_X1 U1030 ( .A1(DATAIN[12]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][12] ), .ZN(n740) );
  INV_X1 U1031 ( .A(n741), .ZN(n3050) );
  AOI22_X1 U1032 ( .A1(DATAIN[13]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][13] ), .ZN(n741) );
  INV_X1 U1033 ( .A(n742), .ZN(n3051) );
  AOI22_X1 U1034 ( .A1(DATAIN[14]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][14] ), .ZN(n742) );
  INV_X1 U1035 ( .A(n743), .ZN(n3052) );
  AOI22_X1 U1036 ( .A1(DATAIN[15]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][15] ), .ZN(n743) );
  INV_X1 U1037 ( .A(n744), .ZN(n3053) );
  AOI22_X1 U1038 ( .A1(DATAIN[16]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][16] ), .ZN(n744) );
  INV_X1 U1039 ( .A(n745), .ZN(n3054) );
  AOI22_X1 U1040 ( .A1(DATAIN[17]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][17] ), .ZN(n745) );
  INV_X1 U1041 ( .A(n746), .ZN(n3055) );
  AOI22_X1 U1042 ( .A1(DATAIN[18]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][18] ), .ZN(n746) );
  INV_X1 U1043 ( .A(n747), .ZN(n3056) );
  AOI22_X1 U1044 ( .A1(DATAIN[19]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][19] ), .ZN(n747) );
  INV_X1 U1045 ( .A(n748), .ZN(n3057) );
  AOI22_X1 U1046 ( .A1(DATAIN[20]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][20] ), .ZN(n748) );
  INV_X1 U1047 ( .A(n749), .ZN(n3058) );
  AOI22_X1 U1048 ( .A1(DATAIN[21]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][21] ), .ZN(n749) );
  INV_X1 U1049 ( .A(n750), .ZN(n3059) );
  AOI22_X1 U1050 ( .A1(DATAIN[22]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][22] ), .ZN(n750) );
  INV_X1 U1051 ( .A(n751), .ZN(n3060) );
  AOI22_X1 U1052 ( .A1(DATAIN[23]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][23] ), .ZN(n751) );
  INV_X1 U1053 ( .A(n752), .ZN(n3061) );
  AOI22_X1 U1054 ( .A1(DATAIN[24]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][24] ), .ZN(n752) );
  INV_X1 U1055 ( .A(n753), .ZN(n3062) );
  AOI22_X1 U1056 ( .A1(DATAIN[25]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][25] ), .ZN(n753) );
  INV_X1 U1057 ( .A(n754), .ZN(n3063) );
  AOI22_X1 U1058 ( .A1(DATAIN[26]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][26] ), .ZN(n754) );
  INV_X1 U1059 ( .A(n755), .ZN(n3064) );
  AOI22_X1 U1060 ( .A1(DATAIN[27]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][27] ), .ZN(n755) );
  INV_X1 U1061 ( .A(n756), .ZN(n3065) );
  AOI22_X1 U1062 ( .A1(DATAIN[28]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][28] ), .ZN(n756) );
  INV_X1 U1063 ( .A(n757), .ZN(n3066) );
  AOI22_X1 U1064 ( .A1(DATAIN[29]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][29] ), .ZN(n757) );
  INV_X1 U1065 ( .A(n758), .ZN(n3067) );
  AOI22_X1 U1066 ( .A1(DATAIN[30]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][30] ), .ZN(n758) );
  INV_X1 U1067 ( .A(n759), .ZN(n3068) );
  AOI22_X1 U1068 ( .A1(DATAIN[31]), .A2(n727), .B1(n728), .B2(
        \REGISTERS[11][31] ), .ZN(n759) );
  INV_X1 U1071 ( .A(n760), .ZN(n3069) );
  AOI22_X1 U1072 ( .A1(DATAIN[0]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][0] ), .ZN(n760) );
  INV_X1 U1073 ( .A(n763), .ZN(n3070) );
  AOI22_X1 U1074 ( .A1(DATAIN[1]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][1] ), .ZN(n763) );
  INV_X1 U1075 ( .A(n764), .ZN(n3071) );
  AOI22_X1 U1076 ( .A1(DATAIN[2]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][2] ), .ZN(n764) );
  INV_X1 U1077 ( .A(n765), .ZN(n3072) );
  AOI22_X1 U1078 ( .A1(DATAIN[3]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][3] ), .ZN(n765) );
  INV_X1 U1079 ( .A(n766), .ZN(n3073) );
  AOI22_X1 U1080 ( .A1(DATAIN[4]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][4] ), .ZN(n766) );
  INV_X1 U1081 ( .A(n767), .ZN(n3074) );
  AOI22_X1 U1082 ( .A1(DATAIN[5]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][5] ), .ZN(n767) );
  INV_X1 U1083 ( .A(n768), .ZN(n3075) );
  AOI22_X1 U1084 ( .A1(DATAIN[6]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][6] ), .ZN(n768) );
  INV_X1 U1085 ( .A(n769), .ZN(n3076) );
  AOI22_X1 U1086 ( .A1(DATAIN[7]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][7] ), .ZN(n769) );
  INV_X1 U1087 ( .A(n770), .ZN(n3077) );
  AOI22_X1 U1088 ( .A1(DATAIN[8]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][8] ), .ZN(n770) );
  INV_X1 U1089 ( .A(n771), .ZN(n3078) );
  AOI22_X1 U1090 ( .A1(DATAIN[9]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][9] ), .ZN(n771) );
  INV_X1 U1091 ( .A(n772), .ZN(n3079) );
  AOI22_X1 U1092 ( .A1(DATAIN[10]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][10] ), .ZN(n772) );
  INV_X1 U1093 ( .A(n773), .ZN(n3080) );
  AOI22_X1 U1094 ( .A1(DATAIN[11]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][11] ), .ZN(n773) );
  INV_X1 U1095 ( .A(n774), .ZN(n3081) );
  AOI22_X1 U1096 ( .A1(DATAIN[12]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][12] ), .ZN(n774) );
  INV_X1 U1097 ( .A(n775), .ZN(n3082) );
  AOI22_X1 U1098 ( .A1(DATAIN[13]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][13] ), .ZN(n775) );
  INV_X1 U1099 ( .A(n776), .ZN(n3083) );
  AOI22_X1 U1100 ( .A1(DATAIN[14]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][14] ), .ZN(n776) );
  INV_X1 U1101 ( .A(n777), .ZN(n3084) );
  AOI22_X1 U1102 ( .A1(DATAIN[15]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][15] ), .ZN(n777) );
  INV_X1 U1103 ( .A(n778), .ZN(n3085) );
  AOI22_X1 U1104 ( .A1(DATAIN[16]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][16] ), .ZN(n778) );
  INV_X1 U1105 ( .A(n779), .ZN(n3086) );
  AOI22_X1 U1106 ( .A1(DATAIN[17]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][17] ), .ZN(n779) );
  INV_X1 U1107 ( .A(n780), .ZN(n3087) );
  AOI22_X1 U1108 ( .A1(DATAIN[18]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][18] ), .ZN(n780) );
  INV_X1 U1109 ( .A(n781), .ZN(n3088) );
  AOI22_X1 U1110 ( .A1(DATAIN[19]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][19] ), .ZN(n781) );
  INV_X1 U1111 ( .A(n782), .ZN(n3089) );
  AOI22_X1 U1112 ( .A1(DATAIN[20]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][20] ), .ZN(n782) );
  INV_X1 U1113 ( .A(n783), .ZN(n3090) );
  AOI22_X1 U1114 ( .A1(DATAIN[21]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][21] ), .ZN(n783) );
  INV_X1 U1115 ( .A(n784), .ZN(n3091) );
  AOI22_X1 U1116 ( .A1(DATAIN[22]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][22] ), .ZN(n784) );
  INV_X1 U1117 ( .A(n785), .ZN(n3092) );
  AOI22_X1 U1118 ( .A1(DATAIN[23]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][23] ), .ZN(n785) );
  INV_X1 U1119 ( .A(n786), .ZN(n3093) );
  AOI22_X1 U1120 ( .A1(DATAIN[24]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][24] ), .ZN(n786) );
  INV_X1 U1121 ( .A(n787), .ZN(n3094) );
  AOI22_X1 U1122 ( .A1(DATAIN[25]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][25] ), .ZN(n787) );
  INV_X1 U1123 ( .A(n788), .ZN(n3095) );
  AOI22_X1 U1124 ( .A1(DATAIN[26]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][26] ), .ZN(n788) );
  INV_X1 U1125 ( .A(n789), .ZN(n3096) );
  AOI22_X1 U1126 ( .A1(DATAIN[27]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][27] ), .ZN(n789) );
  INV_X1 U1127 ( .A(n790), .ZN(n3097) );
  AOI22_X1 U1128 ( .A1(DATAIN[28]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][28] ), .ZN(n790) );
  INV_X1 U1129 ( .A(n791), .ZN(n3098) );
  AOI22_X1 U1130 ( .A1(DATAIN[29]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][29] ), .ZN(n791) );
  INV_X1 U1131 ( .A(n792), .ZN(n3099) );
  AOI22_X1 U1132 ( .A1(DATAIN[30]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][30] ), .ZN(n792) );
  INV_X1 U1133 ( .A(n793), .ZN(n3100) );
  AOI22_X1 U1134 ( .A1(DATAIN[31]), .A2(n761), .B1(n762), .B2(
        \REGISTERS[10][31] ), .ZN(n793) );
  OAI22_X1 U1137 ( .A1(n2), .A2(n794), .B1(n795), .B2(n796), .ZN(n3101) );
  OAI22_X1 U1138 ( .A1(n5), .A2(n794), .B1(n795), .B2(n797), .ZN(n3102) );
  OAI22_X1 U1139 ( .A1(n7), .A2(n794), .B1(n795), .B2(n798), .ZN(n3103) );
  OAI22_X1 U1140 ( .A1(n9), .A2(n794), .B1(n795), .B2(n799), .ZN(n3104) );
  OAI22_X1 U1141 ( .A1(n11), .A2(n794), .B1(n795), .B2(n800), .ZN(n3105) );
  OAI22_X1 U1142 ( .A1(n13), .A2(n794), .B1(n795), .B2(n801), .ZN(n3106) );
  OAI22_X1 U1143 ( .A1(n15), .A2(n794), .B1(n795), .B2(n802), .ZN(n3107) );
  OAI22_X1 U1144 ( .A1(n17), .A2(n794), .B1(n795), .B2(n803), .ZN(n3108) );
  OAI22_X1 U1145 ( .A1(n19), .A2(n794), .B1(n795), .B2(n804), .ZN(n3109) );
  OAI22_X1 U1146 ( .A1(n21), .A2(n794), .B1(n795), .B2(n805), .ZN(n3110) );
  OAI22_X1 U1147 ( .A1(n23), .A2(n794), .B1(n795), .B2(n806), .ZN(n3111) );
  OAI22_X1 U1148 ( .A1(n25), .A2(n794), .B1(n795), .B2(n807), .ZN(n3112) );
  OAI22_X1 U1149 ( .A1(n27), .A2(n794), .B1(n795), .B2(n808), .ZN(n3113) );
  OAI22_X1 U1150 ( .A1(n29), .A2(n794), .B1(n795), .B2(n809), .ZN(n3114) );
  OAI22_X1 U1151 ( .A1(n31), .A2(n794), .B1(n795), .B2(n810), .ZN(n3115) );
  OAI22_X1 U1152 ( .A1(n33), .A2(n794), .B1(n795), .B2(n811), .ZN(n3116) );
  OAI22_X1 U1153 ( .A1(n35), .A2(n794), .B1(n795), .B2(n812), .ZN(n3117) );
  OAI22_X1 U1154 ( .A1(n37), .A2(n794), .B1(n795), .B2(n813), .ZN(n3118) );
  OAI22_X1 U1155 ( .A1(n39), .A2(n794), .B1(n795), .B2(n814), .ZN(n3119) );
  OAI22_X1 U1156 ( .A1(n41), .A2(n794), .B1(n795), .B2(n815), .ZN(n3120) );
  OAI22_X1 U1157 ( .A1(n43), .A2(n794), .B1(n795), .B2(n816), .ZN(n3121) );
  OAI22_X1 U1158 ( .A1(n45), .A2(n794), .B1(n795), .B2(n817), .ZN(n3122) );
  OAI22_X1 U1159 ( .A1(n47), .A2(n794), .B1(n795), .B2(n818), .ZN(n3123) );
  OAI22_X1 U1160 ( .A1(n49), .A2(n794), .B1(n795), .B2(n819), .ZN(n3124) );
  OAI22_X1 U1161 ( .A1(n51), .A2(n794), .B1(n795), .B2(n820), .ZN(n3125) );
  OAI22_X1 U1162 ( .A1(n53), .A2(n794), .B1(n795), .B2(n821), .ZN(n3126) );
  OAI22_X1 U1163 ( .A1(n55), .A2(n794), .B1(n795), .B2(n822), .ZN(n3127) );
  OAI22_X1 U1164 ( .A1(n57), .A2(n794), .B1(n795), .B2(n823), .ZN(n3128) );
  OAI22_X1 U1165 ( .A1(n59), .A2(n794), .B1(n795), .B2(n824), .ZN(n3129) );
  OAI22_X1 U1166 ( .A1(n61), .A2(n794), .B1(n795), .B2(n825), .ZN(n3130) );
  OAI22_X1 U1167 ( .A1(n63), .A2(n794), .B1(n795), .B2(n826), .ZN(n3131) );
  OAI22_X1 U1168 ( .A1(n65), .A2(n794), .B1(n795), .B2(n827), .ZN(n3132) );
  OAI22_X1 U1171 ( .A1(n2), .A2(n828), .B1(n829), .B2(n830), .ZN(n3133) );
  OAI22_X1 U1172 ( .A1(n5), .A2(n828), .B1(n829), .B2(n831), .ZN(n3134) );
  OAI22_X1 U1173 ( .A1(n7), .A2(n828), .B1(n829), .B2(n832), .ZN(n3135) );
  OAI22_X1 U1174 ( .A1(n9), .A2(n828), .B1(n829), .B2(n833), .ZN(n3136) );
  OAI22_X1 U1175 ( .A1(n11), .A2(n828), .B1(n829), .B2(n834), .ZN(n3137) );
  OAI22_X1 U1176 ( .A1(n13), .A2(n828), .B1(n829), .B2(n835), .ZN(n3138) );
  OAI22_X1 U1177 ( .A1(n15), .A2(n828), .B1(n829), .B2(n836), .ZN(n3139) );
  OAI22_X1 U1178 ( .A1(n17), .A2(n828), .B1(n829), .B2(n837), .ZN(n3140) );
  OAI22_X1 U1179 ( .A1(n19), .A2(n828), .B1(n829), .B2(n838), .ZN(n3141) );
  OAI22_X1 U1180 ( .A1(n21), .A2(n828), .B1(n829), .B2(n839), .ZN(n3142) );
  OAI22_X1 U1181 ( .A1(n23), .A2(n828), .B1(n829), .B2(n840), .ZN(n3143) );
  OAI22_X1 U1182 ( .A1(n25), .A2(n828), .B1(n829), .B2(n841), .ZN(n3144) );
  OAI22_X1 U1183 ( .A1(n27), .A2(n828), .B1(n829), .B2(n842), .ZN(n3145) );
  OAI22_X1 U1184 ( .A1(n29), .A2(n828), .B1(n829), .B2(n843), .ZN(n3146) );
  OAI22_X1 U1185 ( .A1(n31), .A2(n828), .B1(n829), .B2(n844), .ZN(n3147) );
  OAI22_X1 U1186 ( .A1(n33), .A2(n828), .B1(n829), .B2(n845), .ZN(n3148) );
  OAI22_X1 U1187 ( .A1(n35), .A2(n828), .B1(n829), .B2(n846), .ZN(n3149) );
  OAI22_X1 U1188 ( .A1(n37), .A2(n828), .B1(n829), .B2(n847), .ZN(n3150) );
  OAI22_X1 U1189 ( .A1(n39), .A2(n828), .B1(n829), .B2(n848), .ZN(n3151) );
  OAI22_X1 U1190 ( .A1(n41), .A2(n828), .B1(n829), .B2(n849), .ZN(n3152) );
  OAI22_X1 U1191 ( .A1(n43), .A2(n828), .B1(n829), .B2(n850), .ZN(n3153) );
  OAI22_X1 U1192 ( .A1(n45), .A2(n828), .B1(n829), .B2(n851), .ZN(n3154) );
  OAI22_X1 U1193 ( .A1(n47), .A2(n828), .B1(n829), .B2(n852), .ZN(n3155) );
  OAI22_X1 U1194 ( .A1(n49), .A2(n828), .B1(n829), .B2(n853), .ZN(n3156) );
  OAI22_X1 U1195 ( .A1(n51), .A2(n828), .B1(n829), .B2(n854), .ZN(n3157) );
  OAI22_X1 U1196 ( .A1(n53), .A2(n828), .B1(n829), .B2(n855), .ZN(n3158) );
  OAI22_X1 U1197 ( .A1(n55), .A2(n828), .B1(n829), .B2(n856), .ZN(n3159) );
  OAI22_X1 U1198 ( .A1(n57), .A2(n828), .B1(n829), .B2(n857), .ZN(n3160) );
  OAI22_X1 U1199 ( .A1(n59), .A2(n828), .B1(n829), .B2(n858), .ZN(n3161) );
  OAI22_X1 U1200 ( .A1(n61), .A2(n828), .B1(n829), .B2(n859), .ZN(n3162) );
  OAI22_X1 U1201 ( .A1(n63), .A2(n828), .B1(n829), .B2(n860), .ZN(n3163) );
  OAI22_X1 U1202 ( .A1(n65), .A2(n828), .B1(n829), .B2(n861), .ZN(n3164) );
  AND3_X1 U1205 ( .A1(n314), .A2(n862), .A3(ADD_WR[3]), .ZN(n623) );
  INV_X1 U1206 ( .A(n863), .ZN(n3165) );
  AOI22_X1 U1207 ( .A1(DATAIN[0]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][0] ), .ZN(n863) );
  INV_X1 U1208 ( .A(n866), .ZN(n3166) );
  AOI22_X1 U1209 ( .A1(DATAIN[1]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][1] ), .ZN(n866) );
  INV_X1 U1210 ( .A(n867), .ZN(n3167) );
  AOI22_X1 U1211 ( .A1(DATAIN[2]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][2] ), .ZN(n867) );
  INV_X1 U1212 ( .A(n868), .ZN(n3168) );
  AOI22_X1 U1213 ( .A1(DATAIN[3]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][3] ), .ZN(n868) );
  INV_X1 U1214 ( .A(n869), .ZN(n3169) );
  AOI22_X1 U1215 ( .A1(DATAIN[4]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][4] ), .ZN(n869) );
  INV_X1 U1216 ( .A(n870), .ZN(n3170) );
  AOI22_X1 U1217 ( .A1(DATAIN[5]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][5] ), .ZN(n870) );
  INV_X1 U1218 ( .A(n871), .ZN(n3171) );
  AOI22_X1 U1219 ( .A1(DATAIN[6]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][6] ), .ZN(n871) );
  INV_X1 U1220 ( .A(n872), .ZN(n3172) );
  AOI22_X1 U1221 ( .A1(DATAIN[7]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][7] ), .ZN(n872) );
  INV_X1 U1222 ( .A(n873), .ZN(n3173) );
  AOI22_X1 U1223 ( .A1(DATAIN[8]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][8] ), .ZN(n873) );
  INV_X1 U1224 ( .A(n874), .ZN(n3174) );
  AOI22_X1 U1225 ( .A1(DATAIN[9]), .A2(n864), .B1(n865), .B2(\REGISTERS[7][9] ), .ZN(n874) );
  INV_X1 U1226 ( .A(n875), .ZN(n3175) );
  AOI22_X1 U1227 ( .A1(DATAIN[10]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][10] ), .ZN(n875) );
  INV_X1 U1228 ( .A(n876), .ZN(n3176) );
  AOI22_X1 U1229 ( .A1(DATAIN[11]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][11] ), .ZN(n876) );
  INV_X1 U1230 ( .A(n877), .ZN(n3177) );
  AOI22_X1 U1231 ( .A1(DATAIN[12]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][12] ), .ZN(n877) );
  INV_X1 U1232 ( .A(n878), .ZN(n3178) );
  AOI22_X1 U1233 ( .A1(DATAIN[13]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][13] ), .ZN(n878) );
  INV_X1 U1234 ( .A(n879), .ZN(n3179) );
  AOI22_X1 U1235 ( .A1(DATAIN[14]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][14] ), .ZN(n879) );
  INV_X1 U1236 ( .A(n880), .ZN(n3180) );
  AOI22_X1 U1237 ( .A1(DATAIN[15]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][15] ), .ZN(n880) );
  INV_X1 U1238 ( .A(n881), .ZN(n3181) );
  AOI22_X1 U1239 ( .A1(DATAIN[16]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][16] ), .ZN(n881) );
  INV_X1 U1240 ( .A(n882), .ZN(n3182) );
  AOI22_X1 U1241 ( .A1(DATAIN[17]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][17] ), .ZN(n882) );
  INV_X1 U1242 ( .A(n883), .ZN(n3183) );
  AOI22_X1 U1243 ( .A1(DATAIN[18]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][18] ), .ZN(n883) );
  INV_X1 U1244 ( .A(n884), .ZN(n3184) );
  AOI22_X1 U1245 ( .A1(DATAIN[19]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][19] ), .ZN(n884) );
  INV_X1 U1246 ( .A(n885), .ZN(n3185) );
  AOI22_X1 U1247 ( .A1(DATAIN[20]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][20] ), .ZN(n885) );
  INV_X1 U1248 ( .A(n886), .ZN(n3186) );
  AOI22_X1 U1249 ( .A1(DATAIN[21]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][21] ), .ZN(n886) );
  INV_X1 U1250 ( .A(n887), .ZN(n3187) );
  AOI22_X1 U1251 ( .A1(DATAIN[22]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][22] ), .ZN(n887) );
  INV_X1 U1252 ( .A(n888), .ZN(n3188) );
  AOI22_X1 U1253 ( .A1(DATAIN[23]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][23] ), .ZN(n888) );
  INV_X1 U1254 ( .A(n889), .ZN(n3189) );
  AOI22_X1 U1255 ( .A1(DATAIN[24]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][24] ), .ZN(n889) );
  INV_X1 U1256 ( .A(n890), .ZN(n3190) );
  AOI22_X1 U1257 ( .A1(DATAIN[25]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][25] ), .ZN(n890) );
  INV_X1 U1258 ( .A(n891), .ZN(n3191) );
  AOI22_X1 U1259 ( .A1(DATAIN[26]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][26] ), .ZN(n891) );
  INV_X1 U1260 ( .A(n892), .ZN(n3192) );
  AOI22_X1 U1261 ( .A1(DATAIN[27]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][27] ), .ZN(n892) );
  INV_X1 U1262 ( .A(n893), .ZN(n3193) );
  AOI22_X1 U1263 ( .A1(DATAIN[28]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][28] ), .ZN(n893) );
  INV_X1 U1264 ( .A(n894), .ZN(n3194) );
  AOI22_X1 U1265 ( .A1(DATAIN[29]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][29] ), .ZN(n894) );
  INV_X1 U1266 ( .A(n895), .ZN(n3195) );
  AOI22_X1 U1267 ( .A1(DATAIN[30]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][30] ), .ZN(n895) );
  INV_X1 U1268 ( .A(n896), .ZN(n3196) );
  AOI22_X1 U1269 ( .A1(DATAIN[31]), .A2(n864), .B1(n865), .B2(
        \REGISTERS[7][31] ), .ZN(n896) );
  NOR3_X1 U1272 ( .A1(n898), .A2(n899), .A3(n900), .ZN(n67) );
  INV_X1 U1273 ( .A(n901), .ZN(n3197) );
  AOI22_X1 U1274 ( .A1(DATAIN[0]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][0] ), .ZN(n901) );
  INV_X1 U1275 ( .A(n904), .ZN(n3198) );
  AOI22_X1 U1276 ( .A1(DATAIN[1]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][1] ), .ZN(n904) );
  INV_X1 U1277 ( .A(n905), .ZN(n3199) );
  AOI22_X1 U1278 ( .A1(DATAIN[2]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][2] ), .ZN(n905) );
  INV_X1 U1279 ( .A(n906), .ZN(n3200) );
  AOI22_X1 U1280 ( .A1(DATAIN[3]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][3] ), .ZN(n906) );
  INV_X1 U1281 ( .A(n907), .ZN(n3201) );
  AOI22_X1 U1282 ( .A1(DATAIN[4]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][4] ), .ZN(n907) );
  INV_X1 U1283 ( .A(n908), .ZN(n3202) );
  AOI22_X1 U1284 ( .A1(DATAIN[5]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][5] ), .ZN(n908) );
  INV_X1 U1285 ( .A(n909), .ZN(n3203) );
  AOI22_X1 U1286 ( .A1(DATAIN[6]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][6] ), .ZN(n909) );
  INV_X1 U1287 ( .A(n910), .ZN(n3204) );
  AOI22_X1 U1288 ( .A1(DATAIN[7]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][7] ), .ZN(n910) );
  INV_X1 U1289 ( .A(n911), .ZN(n3205) );
  AOI22_X1 U1290 ( .A1(DATAIN[8]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][8] ), .ZN(n911) );
  INV_X1 U1291 ( .A(n912), .ZN(n3206) );
  AOI22_X1 U1292 ( .A1(DATAIN[9]), .A2(n902), .B1(n903), .B2(\REGISTERS[6][9] ), .ZN(n912) );
  INV_X1 U1293 ( .A(n913), .ZN(n3207) );
  AOI22_X1 U1294 ( .A1(DATAIN[10]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][10] ), .ZN(n913) );
  INV_X1 U1295 ( .A(n914), .ZN(n3208) );
  AOI22_X1 U1296 ( .A1(DATAIN[11]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][11] ), .ZN(n914) );
  INV_X1 U1297 ( .A(n915), .ZN(n3209) );
  AOI22_X1 U1298 ( .A1(DATAIN[12]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][12] ), .ZN(n915) );
  INV_X1 U1299 ( .A(n916), .ZN(n3210) );
  AOI22_X1 U1300 ( .A1(DATAIN[13]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][13] ), .ZN(n916) );
  INV_X1 U1301 ( .A(n917), .ZN(n3211) );
  AOI22_X1 U1302 ( .A1(DATAIN[14]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][14] ), .ZN(n917) );
  INV_X1 U1303 ( .A(n918), .ZN(n3212) );
  AOI22_X1 U1304 ( .A1(DATAIN[15]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][15] ), .ZN(n918) );
  INV_X1 U1305 ( .A(n919), .ZN(n3213) );
  AOI22_X1 U1306 ( .A1(DATAIN[16]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][16] ), .ZN(n919) );
  INV_X1 U1307 ( .A(n920), .ZN(n3214) );
  AOI22_X1 U1308 ( .A1(DATAIN[17]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][17] ), .ZN(n920) );
  INV_X1 U1309 ( .A(n921), .ZN(n3215) );
  AOI22_X1 U1310 ( .A1(DATAIN[18]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][18] ), .ZN(n921) );
  INV_X1 U1311 ( .A(n922), .ZN(n3216) );
  AOI22_X1 U1312 ( .A1(DATAIN[19]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][19] ), .ZN(n922) );
  INV_X1 U1313 ( .A(n923), .ZN(n3217) );
  AOI22_X1 U1314 ( .A1(DATAIN[20]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][20] ), .ZN(n923) );
  INV_X1 U1315 ( .A(n924), .ZN(n3218) );
  AOI22_X1 U1316 ( .A1(DATAIN[21]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][21] ), .ZN(n924) );
  INV_X1 U1317 ( .A(n925), .ZN(n3219) );
  AOI22_X1 U1318 ( .A1(DATAIN[22]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][22] ), .ZN(n925) );
  INV_X1 U1319 ( .A(n926), .ZN(n3220) );
  AOI22_X1 U1320 ( .A1(DATAIN[23]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][23] ), .ZN(n926) );
  INV_X1 U1321 ( .A(n927), .ZN(n3221) );
  AOI22_X1 U1322 ( .A1(DATAIN[24]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][24] ), .ZN(n927) );
  INV_X1 U1323 ( .A(n928), .ZN(n3222) );
  AOI22_X1 U1324 ( .A1(DATAIN[25]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][25] ), .ZN(n928) );
  INV_X1 U1325 ( .A(n929), .ZN(n3223) );
  AOI22_X1 U1326 ( .A1(DATAIN[26]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][26] ), .ZN(n929) );
  INV_X1 U1327 ( .A(n930), .ZN(n3224) );
  AOI22_X1 U1328 ( .A1(DATAIN[27]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][27] ), .ZN(n930) );
  INV_X1 U1329 ( .A(n931), .ZN(n3225) );
  AOI22_X1 U1330 ( .A1(DATAIN[28]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][28] ), .ZN(n931) );
  INV_X1 U1331 ( .A(n932), .ZN(n3226) );
  AOI22_X1 U1332 ( .A1(DATAIN[29]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][29] ), .ZN(n932) );
  INV_X1 U1333 ( .A(n933), .ZN(n3227) );
  AOI22_X1 U1334 ( .A1(DATAIN[30]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][30] ), .ZN(n933) );
  INV_X1 U1335 ( .A(n934), .ZN(n3228) );
  AOI22_X1 U1336 ( .A1(DATAIN[31]), .A2(n902), .B1(n903), .B2(
        \REGISTERS[6][31] ), .ZN(n934) );
  NOR3_X1 U1339 ( .A1(n898), .A2(ADD_WR[0]), .A3(n900), .ZN(n103) );
  OAI22_X1 U1340 ( .A1(n2), .A2(n935), .B1(n936), .B2(n937), .ZN(n3229) );
  OAI22_X1 U1341 ( .A1(n5), .A2(n935), .B1(n936), .B2(n938), .ZN(n3230) );
  OAI22_X1 U1342 ( .A1(n7), .A2(n935), .B1(n936), .B2(n939), .ZN(n3231) );
  OAI22_X1 U1343 ( .A1(n9), .A2(n935), .B1(n936), .B2(n940), .ZN(n3232) );
  OAI22_X1 U1344 ( .A1(n11), .A2(n935), .B1(n936), .B2(n941), .ZN(n3233) );
  OAI22_X1 U1345 ( .A1(n13), .A2(n935), .B1(n936), .B2(n942), .ZN(n3234) );
  OAI22_X1 U1346 ( .A1(n15), .A2(n935), .B1(n936), .B2(n943), .ZN(n3235) );
  OAI22_X1 U1347 ( .A1(n17), .A2(n935), .B1(n936), .B2(n944), .ZN(n3236) );
  OAI22_X1 U1348 ( .A1(n19), .A2(n935), .B1(n936), .B2(n945), .ZN(n3237) );
  OAI22_X1 U1349 ( .A1(n21), .A2(n935), .B1(n936), .B2(n946), .ZN(n3238) );
  OAI22_X1 U1350 ( .A1(n23), .A2(n935), .B1(n936), .B2(n947), .ZN(n3239) );
  OAI22_X1 U1351 ( .A1(n25), .A2(n935), .B1(n936), .B2(n948), .ZN(n3240) );
  OAI22_X1 U1352 ( .A1(n27), .A2(n935), .B1(n936), .B2(n949), .ZN(n3241) );
  OAI22_X1 U1353 ( .A1(n29), .A2(n935), .B1(n936), .B2(n950), .ZN(n3242) );
  OAI22_X1 U1354 ( .A1(n31), .A2(n935), .B1(n936), .B2(n951), .ZN(n3243) );
  OAI22_X1 U1355 ( .A1(n33), .A2(n935), .B1(n936), .B2(n952), .ZN(n3244) );
  OAI22_X1 U1356 ( .A1(n35), .A2(n935), .B1(n936), .B2(n953), .ZN(n3245) );
  OAI22_X1 U1357 ( .A1(n37), .A2(n935), .B1(n936), .B2(n954), .ZN(n3246) );
  OAI22_X1 U1358 ( .A1(n39), .A2(n935), .B1(n936), .B2(n955), .ZN(n3247) );
  OAI22_X1 U1359 ( .A1(n41), .A2(n935), .B1(n936), .B2(n956), .ZN(n3248) );
  OAI22_X1 U1360 ( .A1(n43), .A2(n935), .B1(n936), .B2(n957), .ZN(n3249) );
  OAI22_X1 U1361 ( .A1(n45), .A2(n935), .B1(n936), .B2(n958), .ZN(n3250) );
  OAI22_X1 U1362 ( .A1(n47), .A2(n935), .B1(n936), .B2(n959), .ZN(n3251) );
  OAI22_X1 U1363 ( .A1(n49), .A2(n935), .B1(n936), .B2(n960), .ZN(n3252) );
  OAI22_X1 U1364 ( .A1(n51), .A2(n935), .B1(n936), .B2(n961), .ZN(n3253) );
  OAI22_X1 U1365 ( .A1(n53), .A2(n935), .B1(n936), .B2(n962), .ZN(n3254) );
  OAI22_X1 U1366 ( .A1(n55), .A2(n935), .B1(n936), .B2(n963), .ZN(n3255) );
  OAI22_X1 U1367 ( .A1(n57), .A2(n935), .B1(n936), .B2(n964), .ZN(n3256) );
  OAI22_X1 U1368 ( .A1(n59), .A2(n935), .B1(n936), .B2(n965), .ZN(n3257) );
  OAI22_X1 U1369 ( .A1(n61), .A2(n935), .B1(n936), .B2(n966), .ZN(n3258) );
  OAI22_X1 U1370 ( .A1(n63), .A2(n935), .B1(n936), .B2(n967), .ZN(n3259) );
  OAI22_X1 U1371 ( .A1(n65), .A2(n935), .B1(n936), .B2(n968), .ZN(n3260) );
  NOR3_X1 U1374 ( .A1(n899), .A2(ADD_WR[1]), .A3(n900), .ZN(n138) );
  OAI22_X1 U1375 ( .A1(n2), .A2(n969), .B1(n970), .B2(n971), .ZN(n3261) );
  OAI22_X1 U1376 ( .A1(n5), .A2(n969), .B1(n970), .B2(n972), .ZN(n3262) );
  OAI22_X1 U1377 ( .A1(n7), .A2(n969), .B1(n970), .B2(n973), .ZN(n3263) );
  OAI22_X1 U1378 ( .A1(n9), .A2(n969), .B1(n970), .B2(n974), .ZN(n3264) );
  OAI22_X1 U1379 ( .A1(n11), .A2(n969), .B1(n970), .B2(n975), .ZN(n3265) );
  OAI22_X1 U1380 ( .A1(n13), .A2(n969), .B1(n970), .B2(n976), .ZN(n3266) );
  OAI22_X1 U1381 ( .A1(n15), .A2(n969), .B1(n970), .B2(n977), .ZN(n3267) );
  OAI22_X1 U1382 ( .A1(n17), .A2(n969), .B1(n970), .B2(n978), .ZN(n3268) );
  OAI22_X1 U1383 ( .A1(n19), .A2(n969), .B1(n970), .B2(n979), .ZN(n3269) );
  OAI22_X1 U1384 ( .A1(n21), .A2(n969), .B1(n970), .B2(n980), .ZN(n3270) );
  OAI22_X1 U1385 ( .A1(n23), .A2(n969), .B1(n970), .B2(n981), .ZN(n3271) );
  OAI22_X1 U1386 ( .A1(n25), .A2(n969), .B1(n970), .B2(n982), .ZN(n3272) );
  OAI22_X1 U1387 ( .A1(n27), .A2(n969), .B1(n970), .B2(n983), .ZN(n3273) );
  OAI22_X1 U1388 ( .A1(n29), .A2(n969), .B1(n970), .B2(n984), .ZN(n3274) );
  OAI22_X1 U1389 ( .A1(n31), .A2(n969), .B1(n970), .B2(n985), .ZN(n3275) );
  OAI22_X1 U1390 ( .A1(n33), .A2(n969), .B1(n970), .B2(n986), .ZN(n3276) );
  OAI22_X1 U1391 ( .A1(n35), .A2(n969), .B1(n970), .B2(n987), .ZN(n3277) );
  OAI22_X1 U1392 ( .A1(n37), .A2(n969), .B1(n970), .B2(n988), .ZN(n3278) );
  OAI22_X1 U1393 ( .A1(n39), .A2(n969), .B1(n970), .B2(n989), .ZN(n3279) );
  OAI22_X1 U1394 ( .A1(n41), .A2(n969), .B1(n970), .B2(n990), .ZN(n3280) );
  OAI22_X1 U1395 ( .A1(n43), .A2(n969), .B1(n970), .B2(n991), .ZN(n3281) );
  OAI22_X1 U1396 ( .A1(n45), .A2(n969), .B1(n970), .B2(n992), .ZN(n3282) );
  OAI22_X1 U1397 ( .A1(n47), .A2(n969), .B1(n970), .B2(n993), .ZN(n3283) );
  OAI22_X1 U1398 ( .A1(n49), .A2(n969), .B1(n970), .B2(n994), .ZN(n3284) );
  OAI22_X1 U1399 ( .A1(n51), .A2(n969), .B1(n970), .B2(n995), .ZN(n3285) );
  OAI22_X1 U1400 ( .A1(n53), .A2(n969), .B1(n970), .B2(n996), .ZN(n3286) );
  OAI22_X1 U1401 ( .A1(n55), .A2(n969), .B1(n970), .B2(n997), .ZN(n3287) );
  OAI22_X1 U1402 ( .A1(n57), .A2(n969), .B1(n970), .B2(n998), .ZN(n3288) );
  OAI22_X1 U1403 ( .A1(n59), .A2(n969), .B1(n970), .B2(n999), .ZN(n3289) );
  OAI22_X1 U1404 ( .A1(n61), .A2(n969), .B1(n970), .B2(n1000), .ZN(n3290) );
  OAI22_X1 U1405 ( .A1(n63), .A2(n969), .B1(n970), .B2(n1001), .ZN(n3291) );
  OAI22_X1 U1406 ( .A1(n65), .A2(n969), .B1(n970), .B2(n1002), .ZN(n3292) );
  NOR3_X1 U1409 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n900), .ZN(n173) );
  INV_X1 U1410 ( .A(ADD_WR[2]), .ZN(n900) );
  INV_X1 U1411 ( .A(n1003), .ZN(n3293) );
  AOI22_X1 U1412 ( .A1(DATAIN[0]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][0] ), .ZN(n1003) );
  INV_X1 U1413 ( .A(n1006), .ZN(n3294) );
  AOI22_X1 U1414 ( .A1(DATAIN[1]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][1] ), .ZN(n1006) );
  INV_X1 U1415 ( .A(n1007), .ZN(n3295) );
  AOI22_X1 U1416 ( .A1(DATAIN[2]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][2] ), .ZN(n1007) );
  INV_X1 U1417 ( .A(n1008), .ZN(n3296) );
  AOI22_X1 U1418 ( .A1(DATAIN[3]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][3] ), .ZN(n1008) );
  INV_X1 U1419 ( .A(n1009), .ZN(n3297) );
  AOI22_X1 U1420 ( .A1(DATAIN[4]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][4] ), .ZN(n1009) );
  INV_X1 U1421 ( .A(n1010), .ZN(n3298) );
  AOI22_X1 U1422 ( .A1(DATAIN[5]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][5] ), .ZN(n1010) );
  INV_X1 U1423 ( .A(n1011), .ZN(n3299) );
  AOI22_X1 U1424 ( .A1(DATAIN[6]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][6] ), .ZN(n1011) );
  INV_X1 U1425 ( .A(n1012), .ZN(n3300) );
  AOI22_X1 U1426 ( .A1(DATAIN[7]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][7] ), .ZN(n1012) );
  INV_X1 U1427 ( .A(n1013), .ZN(n3301) );
  AOI22_X1 U1428 ( .A1(DATAIN[8]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][8] ), .ZN(n1013) );
  INV_X1 U1429 ( .A(n1014), .ZN(n3302) );
  AOI22_X1 U1430 ( .A1(DATAIN[9]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][9] ), .ZN(n1014) );
  INV_X1 U1431 ( .A(n1015), .ZN(n3303) );
  AOI22_X1 U1432 ( .A1(DATAIN[10]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][10] ), .ZN(n1015) );
  INV_X1 U1433 ( .A(n1016), .ZN(n3304) );
  AOI22_X1 U1434 ( .A1(DATAIN[11]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][11] ), .ZN(n1016) );
  INV_X1 U1435 ( .A(n1017), .ZN(n3305) );
  AOI22_X1 U1436 ( .A1(DATAIN[12]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][12] ), .ZN(n1017) );
  INV_X1 U1437 ( .A(n1018), .ZN(n3306) );
  AOI22_X1 U1438 ( .A1(DATAIN[13]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][13] ), .ZN(n1018) );
  INV_X1 U1439 ( .A(n1019), .ZN(n3307) );
  AOI22_X1 U1440 ( .A1(DATAIN[14]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][14] ), .ZN(n1019) );
  INV_X1 U1441 ( .A(n1020), .ZN(n3308) );
  AOI22_X1 U1442 ( .A1(DATAIN[15]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][15] ), .ZN(n1020) );
  INV_X1 U1443 ( .A(n1021), .ZN(n3309) );
  AOI22_X1 U1444 ( .A1(DATAIN[16]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][16] ), .ZN(n1021) );
  INV_X1 U1445 ( .A(n1022), .ZN(n3310) );
  AOI22_X1 U1446 ( .A1(DATAIN[17]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][17] ), .ZN(n1022) );
  INV_X1 U1447 ( .A(n1023), .ZN(n3311) );
  AOI22_X1 U1448 ( .A1(DATAIN[18]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][18] ), .ZN(n1023) );
  INV_X1 U1449 ( .A(n1024), .ZN(n3312) );
  AOI22_X1 U1450 ( .A1(DATAIN[19]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][19] ), .ZN(n1024) );
  INV_X1 U1451 ( .A(n1025), .ZN(n3313) );
  AOI22_X1 U1452 ( .A1(DATAIN[20]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][20] ), .ZN(n1025) );
  INV_X1 U1453 ( .A(n1026), .ZN(n3314) );
  AOI22_X1 U1454 ( .A1(DATAIN[21]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][21] ), .ZN(n1026) );
  INV_X1 U1455 ( .A(n1027), .ZN(n3315) );
  AOI22_X1 U1456 ( .A1(DATAIN[22]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][22] ), .ZN(n1027) );
  INV_X1 U1457 ( .A(n1028), .ZN(n3316) );
  AOI22_X1 U1458 ( .A1(DATAIN[23]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][23] ), .ZN(n1028) );
  INV_X1 U1459 ( .A(n1029), .ZN(n3317) );
  AOI22_X1 U1460 ( .A1(DATAIN[24]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][24] ), .ZN(n1029) );
  INV_X1 U1461 ( .A(n1030), .ZN(n3318) );
  AOI22_X1 U1462 ( .A1(DATAIN[25]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][25] ), .ZN(n1030) );
  INV_X1 U1463 ( .A(n1031), .ZN(n3319) );
  AOI22_X1 U1464 ( .A1(DATAIN[26]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][26] ), .ZN(n1031) );
  INV_X1 U1465 ( .A(n1032), .ZN(n3320) );
  AOI22_X1 U1466 ( .A1(DATAIN[27]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][27] ), .ZN(n1032) );
  INV_X1 U1467 ( .A(n1033), .ZN(n3321) );
  AOI22_X1 U1468 ( .A1(DATAIN[28]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][28] ), .ZN(n1033) );
  INV_X1 U1469 ( .A(n1034), .ZN(n3322) );
  AOI22_X1 U1470 ( .A1(DATAIN[29]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][29] ), .ZN(n1034) );
  INV_X1 U1471 ( .A(n1035), .ZN(n3323) );
  AOI22_X1 U1472 ( .A1(DATAIN[30]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][30] ), .ZN(n1035) );
  INV_X1 U1473 ( .A(n1036), .ZN(n3324) );
  AOI22_X1 U1474 ( .A1(DATAIN[31]), .A2(n1004), .B1(n1005), .B2(
        \REGISTERS[3][31] ), .ZN(n1036) );
  NOR3_X1 U1477 ( .A1(n899), .A2(ADD_WR[2]), .A3(n898), .ZN(n208) );
  INV_X1 U1478 ( .A(n1037), .ZN(n3325) );
  AOI22_X1 U1479 ( .A1(DATAIN[0]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][0] ), .ZN(n1037) );
  INV_X1 U1480 ( .A(n1040), .ZN(n3326) );
  AOI22_X1 U1481 ( .A1(DATAIN[1]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][1] ), .ZN(n1040) );
  INV_X1 U1482 ( .A(n1041), .ZN(n3327) );
  AOI22_X1 U1483 ( .A1(DATAIN[2]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][2] ), .ZN(n1041) );
  INV_X1 U1484 ( .A(n1042), .ZN(n3328) );
  AOI22_X1 U1485 ( .A1(DATAIN[3]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][3] ), .ZN(n1042) );
  INV_X1 U1486 ( .A(n1043), .ZN(n3329) );
  AOI22_X1 U1487 ( .A1(DATAIN[4]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][4] ), .ZN(n1043) );
  INV_X1 U1488 ( .A(n1044), .ZN(n3330) );
  AOI22_X1 U1489 ( .A1(DATAIN[5]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][5] ), .ZN(n1044) );
  INV_X1 U1490 ( .A(n1045), .ZN(n3331) );
  AOI22_X1 U1491 ( .A1(DATAIN[6]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][6] ), .ZN(n1045) );
  INV_X1 U1492 ( .A(n1046), .ZN(n3332) );
  AOI22_X1 U1493 ( .A1(DATAIN[7]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][7] ), .ZN(n1046) );
  INV_X1 U1494 ( .A(n1047), .ZN(n3333) );
  AOI22_X1 U1495 ( .A1(DATAIN[8]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][8] ), .ZN(n1047) );
  INV_X1 U1496 ( .A(n1048), .ZN(n3334) );
  AOI22_X1 U1497 ( .A1(DATAIN[9]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][9] ), .ZN(n1048) );
  INV_X1 U1498 ( .A(n1049), .ZN(n3335) );
  AOI22_X1 U1499 ( .A1(DATAIN[10]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][10] ), .ZN(n1049) );
  INV_X1 U1500 ( .A(n1050), .ZN(n3336) );
  AOI22_X1 U1501 ( .A1(DATAIN[11]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][11] ), .ZN(n1050) );
  INV_X1 U1502 ( .A(n1051), .ZN(n3337) );
  AOI22_X1 U1503 ( .A1(DATAIN[12]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][12] ), .ZN(n1051) );
  INV_X1 U1504 ( .A(n1052), .ZN(n3338) );
  AOI22_X1 U1505 ( .A1(DATAIN[13]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][13] ), .ZN(n1052) );
  INV_X1 U1506 ( .A(n1053), .ZN(n3339) );
  AOI22_X1 U1507 ( .A1(DATAIN[14]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][14] ), .ZN(n1053) );
  INV_X1 U1508 ( .A(n1054), .ZN(n3340) );
  AOI22_X1 U1509 ( .A1(DATAIN[15]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][15] ), .ZN(n1054) );
  INV_X1 U1510 ( .A(n1055), .ZN(n3341) );
  AOI22_X1 U1511 ( .A1(DATAIN[16]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][16] ), .ZN(n1055) );
  INV_X1 U1512 ( .A(n1056), .ZN(n3342) );
  AOI22_X1 U1513 ( .A1(DATAIN[17]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][17] ), .ZN(n1056) );
  INV_X1 U1514 ( .A(n1057), .ZN(n3343) );
  AOI22_X1 U1515 ( .A1(DATAIN[18]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][18] ), .ZN(n1057) );
  INV_X1 U1516 ( .A(n1058), .ZN(n3344) );
  AOI22_X1 U1517 ( .A1(DATAIN[19]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][19] ), .ZN(n1058) );
  INV_X1 U1518 ( .A(n1059), .ZN(n3345) );
  AOI22_X1 U1519 ( .A1(DATAIN[20]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][20] ), .ZN(n1059) );
  INV_X1 U1520 ( .A(n1060), .ZN(n3346) );
  AOI22_X1 U1521 ( .A1(DATAIN[21]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][21] ), .ZN(n1060) );
  INV_X1 U1522 ( .A(n1061), .ZN(n3347) );
  AOI22_X1 U1523 ( .A1(DATAIN[22]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][22] ), .ZN(n1061) );
  INV_X1 U1524 ( .A(n1062), .ZN(n3348) );
  AOI22_X1 U1525 ( .A1(DATAIN[23]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][23] ), .ZN(n1062) );
  INV_X1 U1526 ( .A(n1063), .ZN(n3349) );
  AOI22_X1 U1527 ( .A1(DATAIN[24]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][24] ), .ZN(n1063) );
  INV_X1 U1528 ( .A(n1064), .ZN(n3350) );
  AOI22_X1 U1529 ( .A1(DATAIN[25]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][25] ), .ZN(n1064) );
  INV_X1 U1530 ( .A(n1065), .ZN(n3351) );
  AOI22_X1 U1531 ( .A1(DATAIN[26]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][26] ), .ZN(n1065) );
  INV_X1 U1532 ( .A(n1066), .ZN(n3352) );
  AOI22_X1 U1533 ( .A1(DATAIN[27]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][27] ), .ZN(n1066) );
  INV_X1 U1534 ( .A(n1067), .ZN(n3353) );
  AOI22_X1 U1535 ( .A1(DATAIN[28]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][28] ), .ZN(n1067) );
  INV_X1 U1536 ( .A(n1068), .ZN(n3354) );
  AOI22_X1 U1537 ( .A1(DATAIN[29]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][29] ), .ZN(n1068) );
  INV_X1 U1538 ( .A(n1069), .ZN(n3355) );
  AOI22_X1 U1539 ( .A1(DATAIN[30]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][30] ), .ZN(n1069) );
  INV_X1 U1540 ( .A(n1070), .ZN(n3356) );
  AOI22_X1 U1541 ( .A1(DATAIN[31]), .A2(n1038), .B1(n1039), .B2(
        \REGISTERS[2][31] ), .ZN(n1070) );
  NOR3_X1 U1544 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n898), .ZN(n243) );
  INV_X1 U1545 ( .A(ADD_WR[1]), .ZN(n898) );
  OAI22_X1 U1546 ( .A1(n2), .A2(n1071), .B1(n1072), .B2(n1073), .ZN(n3357) );
  OAI22_X1 U1547 ( .A1(n5), .A2(n1071), .B1(n1072), .B2(n1074), .ZN(n3358) );
  OAI22_X1 U1548 ( .A1(n7), .A2(n1071), .B1(n1072), .B2(n1075), .ZN(n3359) );
  OAI22_X1 U1549 ( .A1(n9), .A2(n1071), .B1(n1072), .B2(n1076), .ZN(n3360) );
  OAI22_X1 U1550 ( .A1(n11), .A2(n1071), .B1(n1072), .B2(n1077), .ZN(n3361) );
  OAI22_X1 U1551 ( .A1(n13), .A2(n1071), .B1(n1072), .B2(n1078), .ZN(n3362) );
  OAI22_X1 U1552 ( .A1(n15), .A2(n1071), .B1(n1072), .B2(n1079), .ZN(n3363) );
  OAI22_X1 U1553 ( .A1(n17), .A2(n1071), .B1(n1072), .B2(n1080), .ZN(n3364) );
  OAI22_X1 U1554 ( .A1(n19), .A2(n1071), .B1(n1072), .B2(n1081), .ZN(n3365) );
  OAI22_X1 U1555 ( .A1(n21), .A2(n1071), .B1(n1072), .B2(n1082), .ZN(n3366) );
  OAI22_X1 U1556 ( .A1(n23), .A2(n1071), .B1(n1072), .B2(n1083), .ZN(n3367) );
  OAI22_X1 U1557 ( .A1(n25), .A2(n1071), .B1(n1072), .B2(n1084), .ZN(n3368) );
  OAI22_X1 U1558 ( .A1(n27), .A2(n1071), .B1(n1072), .B2(n1085), .ZN(n3369) );
  OAI22_X1 U1559 ( .A1(n29), .A2(n1071), .B1(n1072), .B2(n1086), .ZN(n3370) );
  OAI22_X1 U1560 ( .A1(n31), .A2(n1071), .B1(n1072), .B2(n1087), .ZN(n3371) );
  OAI22_X1 U1561 ( .A1(n33), .A2(n1071), .B1(n1072), .B2(n1088), .ZN(n3372) );
  OAI22_X1 U1562 ( .A1(n35), .A2(n1071), .B1(n1072), .B2(n1089), .ZN(n3373) );
  OAI22_X1 U1563 ( .A1(n37), .A2(n1071), .B1(n1072), .B2(n1090), .ZN(n3374) );
  OAI22_X1 U1564 ( .A1(n39), .A2(n1071), .B1(n1072), .B2(n1091), .ZN(n3375) );
  OAI22_X1 U1565 ( .A1(n41), .A2(n1071), .B1(n1072), .B2(n1092), .ZN(n3376) );
  OAI22_X1 U1566 ( .A1(n43), .A2(n1071), .B1(n1072), .B2(n1093), .ZN(n3377) );
  OAI22_X1 U1567 ( .A1(n45), .A2(n1071), .B1(n1072), .B2(n1094), .ZN(n3378) );
  OAI22_X1 U1568 ( .A1(n47), .A2(n1071), .B1(n1072), .B2(n1095), .ZN(n3379) );
  OAI22_X1 U1569 ( .A1(n49), .A2(n1071), .B1(n1072), .B2(n1096), .ZN(n3380) );
  OAI22_X1 U1570 ( .A1(n51), .A2(n1071), .B1(n1072), .B2(n1097), .ZN(n3381) );
  OAI22_X1 U1571 ( .A1(n53), .A2(n1071), .B1(n1072), .B2(n1098), .ZN(n3382) );
  OAI22_X1 U1572 ( .A1(n55), .A2(n1071), .B1(n1072), .B2(n1099), .ZN(n3383) );
  OAI22_X1 U1573 ( .A1(n57), .A2(n1071), .B1(n1072), .B2(n1100), .ZN(n3384) );
  OAI22_X1 U1574 ( .A1(n59), .A2(n1071), .B1(n1072), .B2(n1101), .ZN(n3385) );
  OAI22_X1 U1575 ( .A1(n61), .A2(n1071), .B1(n1072), .B2(n1102), .ZN(n3386) );
  OAI22_X1 U1576 ( .A1(n63), .A2(n1071), .B1(n1072), .B2(n1103), .ZN(n3387) );
  OAI22_X1 U1577 ( .A1(n65), .A2(n1071), .B1(n1072), .B2(n1104), .ZN(n3388) );
  NOR3_X1 U1580 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n899), .ZN(n278) );
  INV_X1 U1581 ( .A(ADD_WR[0]), .ZN(n899) );
  OAI22_X1 U1582 ( .A1(n2), .A2(n1105), .B1(n1106), .B2(n1107), .ZN(n3389) );
  INV_X1 U1583 ( .A(DATAIN[0]), .ZN(n2) );
  OAI22_X1 U1584 ( .A1(n5), .A2(n1105), .B1(n1106), .B2(n1108), .ZN(n3390) );
  INV_X1 U1585 ( .A(DATAIN[1]), .ZN(n5) );
  OAI22_X1 U1586 ( .A1(n7), .A2(n1105), .B1(n1106), .B2(n1109), .ZN(n3391) );
  INV_X1 U1587 ( .A(DATAIN[2]), .ZN(n7) );
  OAI22_X1 U1588 ( .A1(n9), .A2(n1105), .B1(n1106), .B2(n1110), .ZN(n3392) );
  INV_X1 U1589 ( .A(DATAIN[3]), .ZN(n9) );
  OAI22_X1 U1590 ( .A1(n11), .A2(n1105), .B1(n1106), .B2(n1111), .ZN(n3393) );
  INV_X1 U1591 ( .A(DATAIN[4]), .ZN(n11) );
  OAI22_X1 U1592 ( .A1(n13), .A2(n1105), .B1(n1106), .B2(n1112), .ZN(n3394) );
  INV_X1 U1593 ( .A(DATAIN[5]), .ZN(n13) );
  OAI22_X1 U1594 ( .A1(n15), .A2(n1105), .B1(n1106), .B2(n1113), .ZN(n3395) );
  INV_X1 U1595 ( .A(DATAIN[6]), .ZN(n15) );
  OAI22_X1 U1596 ( .A1(n17), .A2(n1105), .B1(n1106), .B2(n1114), .ZN(n3396) );
  INV_X1 U1597 ( .A(DATAIN[7]), .ZN(n17) );
  OAI22_X1 U1598 ( .A1(n19), .A2(n1105), .B1(n1106), .B2(n1115), .ZN(n3397) );
  INV_X1 U1599 ( .A(DATAIN[8]), .ZN(n19) );
  OAI22_X1 U1600 ( .A1(n21), .A2(n1105), .B1(n1106), .B2(n1116), .ZN(n3398) );
  INV_X1 U1601 ( .A(DATAIN[9]), .ZN(n21) );
  OAI22_X1 U1602 ( .A1(n23), .A2(n1105), .B1(n1106), .B2(n1117), .ZN(n3399) );
  INV_X1 U1603 ( .A(DATAIN[10]), .ZN(n23) );
  OAI22_X1 U1604 ( .A1(n25), .A2(n1105), .B1(n1106), .B2(n1118), .ZN(n3400) );
  INV_X1 U1605 ( .A(DATAIN[11]), .ZN(n25) );
  OAI22_X1 U1606 ( .A1(n27), .A2(n1105), .B1(n1106), .B2(n1119), .ZN(n3401) );
  INV_X1 U1607 ( .A(DATAIN[12]), .ZN(n27) );
  OAI22_X1 U1608 ( .A1(n29), .A2(n1105), .B1(n1106), .B2(n1120), .ZN(n3402) );
  INV_X1 U1609 ( .A(DATAIN[13]), .ZN(n29) );
  OAI22_X1 U1610 ( .A1(n31), .A2(n1105), .B1(n1106), .B2(n1121), .ZN(n3403) );
  INV_X1 U1611 ( .A(DATAIN[14]), .ZN(n31) );
  OAI22_X1 U1612 ( .A1(n33), .A2(n1105), .B1(n1106), .B2(n1122), .ZN(n3404) );
  INV_X1 U1613 ( .A(DATAIN[15]), .ZN(n33) );
  OAI22_X1 U1614 ( .A1(n35), .A2(n1105), .B1(n1106), .B2(n1123), .ZN(n3405) );
  INV_X1 U1615 ( .A(DATAIN[16]), .ZN(n35) );
  OAI22_X1 U1616 ( .A1(n37), .A2(n1105), .B1(n1106), .B2(n1124), .ZN(n3406) );
  INV_X1 U1617 ( .A(DATAIN[17]), .ZN(n37) );
  OAI22_X1 U1618 ( .A1(n39), .A2(n1105), .B1(n1106), .B2(n1125), .ZN(n3407) );
  INV_X1 U1619 ( .A(DATAIN[18]), .ZN(n39) );
  OAI22_X1 U1620 ( .A1(n41), .A2(n1105), .B1(n1106), .B2(n1126), .ZN(n3408) );
  INV_X1 U1621 ( .A(DATAIN[19]), .ZN(n41) );
  OAI22_X1 U1622 ( .A1(n43), .A2(n1105), .B1(n1106), .B2(n1127), .ZN(n3409) );
  INV_X1 U1623 ( .A(DATAIN[20]), .ZN(n43) );
  OAI22_X1 U1624 ( .A1(n45), .A2(n1105), .B1(n1106), .B2(n1128), .ZN(n3410) );
  INV_X1 U1625 ( .A(DATAIN[21]), .ZN(n45) );
  OAI22_X1 U1626 ( .A1(n47), .A2(n1105), .B1(n1106), .B2(n1129), .ZN(n3411) );
  INV_X1 U1627 ( .A(DATAIN[22]), .ZN(n47) );
  OAI22_X1 U1628 ( .A1(n49), .A2(n1105), .B1(n1106), .B2(n1130), .ZN(n3412) );
  INV_X1 U1629 ( .A(DATAIN[23]), .ZN(n49) );
  OAI22_X1 U1630 ( .A1(n51), .A2(n1105), .B1(n1106), .B2(n1131), .ZN(n3413) );
  INV_X1 U1631 ( .A(DATAIN[24]), .ZN(n51) );
  OAI22_X1 U1632 ( .A1(n53), .A2(n1105), .B1(n1106), .B2(n1132), .ZN(n3414) );
  INV_X1 U1633 ( .A(DATAIN[25]), .ZN(n53) );
  OAI22_X1 U1634 ( .A1(n55), .A2(n1105), .B1(n1106), .B2(n1133), .ZN(n3415) );
  INV_X1 U1635 ( .A(DATAIN[26]), .ZN(n55) );
  OAI22_X1 U1636 ( .A1(n57), .A2(n1105), .B1(n1106), .B2(n1134), .ZN(n3416) );
  INV_X1 U1637 ( .A(DATAIN[27]), .ZN(n57) );
  OAI22_X1 U1638 ( .A1(n59), .A2(n1105), .B1(n1106), .B2(n1135), .ZN(n3417) );
  INV_X1 U1639 ( .A(DATAIN[28]), .ZN(n59) );
  OAI22_X1 U1640 ( .A1(n61), .A2(n1105), .B1(n1106), .B2(n1136), .ZN(n3418) );
  INV_X1 U1641 ( .A(DATAIN[29]), .ZN(n61) );
  OAI22_X1 U1642 ( .A1(n63), .A2(n1105), .B1(n1106), .B2(n1137), .ZN(n3419) );
  INV_X1 U1643 ( .A(DATAIN[30]), .ZN(n63) );
  OAI22_X1 U1644 ( .A1(n65), .A2(n1105), .B1(n1106), .B2(n1138), .ZN(n3420) );
  NOR3_X1 U1647 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n313) );
  AND3_X1 U1648 ( .A1(n588), .A2(n862), .A3(n314), .ZN(n897) );
  AND3_X1 U1649 ( .A1(WR), .A2(ENABLE), .A3(wr_signal), .ZN(n314) );
  INV_X1 U1650 ( .A(ADD_WR[4]), .ZN(n862) );
  INV_X1 U1651 ( .A(ADD_WR[3]), .ZN(n588) );
  INV_X1 U1652 ( .A(DATAIN[31]), .ZN(n65) );
  AOI21_X1 U1653 ( .B1(n1139), .B2(n1140), .A(N352), .ZN(N351) );
  NOR4_X1 U1654 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1140)
         );
  OAI221_X1 U1655 ( .B1(n553), .B2(n1145), .C1(n587), .C2(n1146), .A(n1147), 
        .ZN(n1144) );
  AOI22_X1 U1656 ( .A1(n1148), .A2(\REGISTERS[19][31] ), .B1(n1149), .B2(
        \REGISTERS[18][31] ), .ZN(n1147) );
  OAI221_X1 U1657 ( .B1(n417), .B2(n1150), .C1(n451), .C2(n1151), .A(n1152), 
        .ZN(n1143) );
  AOI22_X1 U1658 ( .A1(n1153), .A2(\REGISTERS[23][31] ), .B1(n1154), .B2(
        \REGISTERS[22][31] ), .ZN(n1152) );
  OAI221_X1 U1659 ( .B1(n277), .B2(n1155), .C1(n312), .C2(n1156), .A(n1157), 
        .ZN(n1142) );
  AOI22_X1 U1660 ( .A1(n1158), .A2(\REGISTERS[27][31] ), .B1(n1159), .B2(
        \REGISTERS[26][31] ), .ZN(n1157) );
  OAI221_X1 U1661 ( .B1(n66), .B2(n1160), .C1(n102), .C2(n1161), .A(n1162), 
        .ZN(n1141) );
  AOI22_X1 U1662 ( .A1(n1163), .A2(\REGISTERS[29][31] ), .B1(n1164), .B2(
        \REGISTERS[28][31] ), .ZN(n1162) );
  NOR4_X1 U1663 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1139)
         );
  OAI221_X1 U1664 ( .B1(n1104), .B2(n1169), .C1(n1138), .C2(n1170), .A(n1171), 
        .ZN(n1168) );
  AOI22_X1 U1665 ( .A1(n1172), .A2(\REGISTERS[3][31] ), .B1(n1173), .B2(
        \REGISTERS[2][31] ), .ZN(n1171) );
  OAI221_X1 U1666 ( .B1(n968), .B2(n1174), .C1(n1002), .C2(n1175), .A(n1176), 
        .ZN(n1167) );
  AOI22_X1 U1667 ( .A1(n1177), .A2(\REGISTERS[7][31] ), .B1(n1178), .B2(
        \REGISTERS[6][31] ), .ZN(n1176) );
  OAI221_X1 U1668 ( .B1(n827), .B2(n1179), .C1(n861), .C2(n1180), .A(n1181), 
        .ZN(n1166) );
  AOI22_X1 U1669 ( .A1(n1182), .A2(\REGISTERS[11][31] ), .B1(n1183), .B2(
        \REGISTERS[10][31] ), .ZN(n1181) );
  OAI221_X1 U1670 ( .B1(n691), .B2(n1184), .C1(n725), .C2(n1185), .A(n1186), 
        .ZN(n1165) );
  AOI22_X1 U1671 ( .A1(n1187), .A2(\REGISTERS[15][31] ), .B1(n1188), .B2(
        \REGISTERS[14][31] ), .ZN(n1186) );
  AOI21_X1 U1672 ( .B1(n1189), .B2(n1190), .A(N352), .ZN(N350) );
  NOR4_X1 U1673 ( .A1(n1191), .A2(n1192), .A3(n1193), .A4(n1194), .ZN(n1190)
         );
  OAI221_X1 U1674 ( .B1(n552), .B2(n1145), .C1(n586), .C2(n1146), .A(n1195), 
        .ZN(n1194) );
  AOI22_X1 U1675 ( .A1(n1148), .A2(\REGISTERS[19][30] ), .B1(n1149), .B2(
        \REGISTERS[18][30] ), .ZN(n1195) );
  OAI221_X1 U1676 ( .B1(n416), .B2(n1150), .C1(n450), .C2(n1151), .A(n1196), 
        .ZN(n1193) );
  AOI22_X1 U1677 ( .A1(n1153), .A2(\REGISTERS[23][30] ), .B1(n1154), .B2(
        \REGISTERS[22][30] ), .ZN(n1196) );
  OAI221_X1 U1678 ( .B1(n276), .B2(n1155), .C1(n311), .C2(n1156), .A(n1197), 
        .ZN(n1192) );
  AOI22_X1 U1679 ( .A1(n1158), .A2(\REGISTERS[27][30] ), .B1(n1159), .B2(
        \REGISTERS[26][30] ), .ZN(n1197) );
  OAI221_X1 U1680 ( .B1(n64), .B2(n1160), .C1(n101), .C2(n1161), .A(n1198), 
        .ZN(n1191) );
  AOI22_X1 U1681 ( .A1(n1163), .A2(\REGISTERS[29][30] ), .B1(n1164), .B2(
        \REGISTERS[28][30] ), .ZN(n1198) );
  NOR4_X1 U1682 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n1189)
         );
  OAI221_X1 U1683 ( .B1(n1103), .B2(n1169), .C1(n1137), .C2(n1170), .A(n1203), 
        .ZN(n1202) );
  AOI22_X1 U1684 ( .A1(n1172), .A2(\REGISTERS[3][30] ), .B1(n1173), .B2(
        \REGISTERS[2][30] ), .ZN(n1203) );
  OAI221_X1 U1685 ( .B1(n967), .B2(n1174), .C1(n1001), .C2(n1175), .A(n1204), 
        .ZN(n1201) );
  AOI22_X1 U1686 ( .A1(n1177), .A2(\REGISTERS[7][30] ), .B1(n1178), .B2(
        \REGISTERS[6][30] ), .ZN(n1204) );
  OAI221_X1 U1687 ( .B1(n826), .B2(n1179), .C1(n860), .C2(n1180), .A(n1205), 
        .ZN(n1200) );
  AOI22_X1 U1688 ( .A1(n1182), .A2(\REGISTERS[11][30] ), .B1(n1183), .B2(
        \REGISTERS[10][30] ), .ZN(n1205) );
  OAI221_X1 U1689 ( .B1(n690), .B2(n1184), .C1(n724), .C2(n1185), .A(n1206), 
        .ZN(n1199) );
  AOI22_X1 U1690 ( .A1(n1187), .A2(\REGISTERS[15][30] ), .B1(n1188), .B2(
        \REGISTERS[14][30] ), .ZN(n1206) );
  AOI21_X1 U1691 ( .B1(n1207), .B2(n1208), .A(N352), .ZN(N349) );
  NOR4_X1 U1692 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1208)
         );
  OAI221_X1 U1693 ( .B1(n551), .B2(n1145), .C1(n585), .C2(n1146), .A(n1213), 
        .ZN(n1212) );
  AOI22_X1 U1694 ( .A1(n1148), .A2(\REGISTERS[19][29] ), .B1(n1149), .B2(
        \REGISTERS[18][29] ), .ZN(n1213) );
  OAI221_X1 U1695 ( .B1(n415), .B2(n1150), .C1(n449), .C2(n1151), .A(n1214), 
        .ZN(n1211) );
  AOI22_X1 U1696 ( .A1(n1153), .A2(\REGISTERS[23][29] ), .B1(n1154), .B2(
        \REGISTERS[22][29] ), .ZN(n1214) );
  OAI221_X1 U1697 ( .B1(n275), .B2(n1155), .C1(n310), .C2(n1156), .A(n1215), 
        .ZN(n1210) );
  AOI22_X1 U1698 ( .A1(n1158), .A2(\REGISTERS[27][29] ), .B1(n1159), .B2(
        \REGISTERS[26][29] ), .ZN(n1215) );
  OAI221_X1 U1699 ( .B1(n62), .B2(n1160), .C1(n100), .C2(n1161), .A(n1216), 
        .ZN(n1209) );
  AOI22_X1 U1700 ( .A1(n1163), .A2(\REGISTERS[29][29] ), .B1(n1164), .B2(
        \REGISTERS[28][29] ), .ZN(n1216) );
  NOR4_X1 U1701 ( .A1(n1217), .A2(n1218), .A3(n1219), .A4(n1220), .ZN(n1207)
         );
  OAI221_X1 U1702 ( .B1(n1102), .B2(n1169), .C1(n1136), .C2(n1170), .A(n1221), 
        .ZN(n1220) );
  AOI22_X1 U1703 ( .A1(n1172), .A2(\REGISTERS[3][29] ), .B1(n1173), .B2(
        \REGISTERS[2][29] ), .ZN(n1221) );
  OAI221_X1 U1704 ( .B1(n966), .B2(n1174), .C1(n1000), .C2(n1175), .A(n1222), 
        .ZN(n1219) );
  AOI22_X1 U1705 ( .A1(n1177), .A2(\REGISTERS[7][29] ), .B1(n1178), .B2(
        \REGISTERS[6][29] ), .ZN(n1222) );
  OAI221_X1 U1706 ( .B1(n825), .B2(n1179), .C1(n859), .C2(n1180), .A(n1223), 
        .ZN(n1218) );
  AOI22_X1 U1707 ( .A1(n1182), .A2(\REGISTERS[11][29] ), .B1(n1183), .B2(
        \REGISTERS[10][29] ), .ZN(n1223) );
  OAI221_X1 U1708 ( .B1(n689), .B2(n1184), .C1(n723), .C2(n1185), .A(n1224), 
        .ZN(n1217) );
  AOI22_X1 U1709 ( .A1(n1187), .A2(\REGISTERS[15][29] ), .B1(n1188), .B2(
        \REGISTERS[14][29] ), .ZN(n1224) );
  AOI21_X1 U1710 ( .B1(n1225), .B2(n1226), .A(N352), .ZN(N348) );
  NOR4_X1 U1711 ( .A1(n1227), .A2(n1228), .A3(n1229), .A4(n1230), .ZN(n1226)
         );
  OAI221_X1 U1712 ( .B1(n550), .B2(n1145), .C1(n584), .C2(n1146), .A(n1231), 
        .ZN(n1230) );
  AOI22_X1 U1713 ( .A1(n1148), .A2(\REGISTERS[19][28] ), .B1(n1149), .B2(
        \REGISTERS[18][28] ), .ZN(n1231) );
  OAI221_X1 U1714 ( .B1(n414), .B2(n1150), .C1(n448), .C2(n1151), .A(n1232), 
        .ZN(n1229) );
  AOI22_X1 U1715 ( .A1(n1153), .A2(\REGISTERS[23][28] ), .B1(n1154), .B2(
        \REGISTERS[22][28] ), .ZN(n1232) );
  OAI221_X1 U1716 ( .B1(n274), .B2(n1155), .C1(n309), .C2(n1156), .A(n1233), 
        .ZN(n1228) );
  AOI22_X1 U1717 ( .A1(n1158), .A2(\REGISTERS[27][28] ), .B1(n1159), .B2(
        \REGISTERS[26][28] ), .ZN(n1233) );
  OAI221_X1 U1718 ( .B1(n60), .B2(n1160), .C1(n99), .C2(n1161), .A(n1234), 
        .ZN(n1227) );
  AOI22_X1 U1719 ( .A1(n1163), .A2(\REGISTERS[29][28] ), .B1(n1164), .B2(
        \REGISTERS[28][28] ), .ZN(n1234) );
  NOR4_X1 U1720 ( .A1(n1235), .A2(n1236), .A3(n1237), .A4(n1238), .ZN(n1225)
         );
  OAI221_X1 U1721 ( .B1(n1101), .B2(n1169), .C1(n1135), .C2(n1170), .A(n1239), 
        .ZN(n1238) );
  AOI22_X1 U1722 ( .A1(n1172), .A2(\REGISTERS[3][28] ), .B1(n1173), .B2(
        \REGISTERS[2][28] ), .ZN(n1239) );
  OAI221_X1 U1723 ( .B1(n965), .B2(n1174), .C1(n999), .C2(n1175), .A(n1240), 
        .ZN(n1237) );
  AOI22_X1 U1724 ( .A1(n1177), .A2(\REGISTERS[7][28] ), .B1(n1178), .B2(
        \REGISTERS[6][28] ), .ZN(n1240) );
  OAI221_X1 U1725 ( .B1(n824), .B2(n1179), .C1(n858), .C2(n1180), .A(n1241), 
        .ZN(n1236) );
  AOI22_X1 U1726 ( .A1(n1182), .A2(\REGISTERS[11][28] ), .B1(n1183), .B2(
        \REGISTERS[10][28] ), .ZN(n1241) );
  OAI221_X1 U1727 ( .B1(n688), .B2(n1184), .C1(n722), .C2(n1185), .A(n1242), 
        .ZN(n1235) );
  AOI22_X1 U1728 ( .A1(n1187), .A2(\REGISTERS[15][28] ), .B1(n1188), .B2(
        \REGISTERS[14][28] ), .ZN(n1242) );
  AOI21_X1 U1729 ( .B1(n1243), .B2(n1244), .A(N352), .ZN(N347) );
  NOR4_X1 U1730 ( .A1(n1245), .A2(n1246), .A3(n1247), .A4(n1248), .ZN(n1244)
         );
  OAI221_X1 U1731 ( .B1(n549), .B2(n1145), .C1(n583), .C2(n1146), .A(n1249), 
        .ZN(n1248) );
  AOI22_X1 U1732 ( .A1(n1148), .A2(\REGISTERS[19][27] ), .B1(n1149), .B2(
        \REGISTERS[18][27] ), .ZN(n1249) );
  OAI221_X1 U1733 ( .B1(n413), .B2(n1150), .C1(n447), .C2(n1151), .A(n1250), 
        .ZN(n1247) );
  AOI22_X1 U1734 ( .A1(n1153), .A2(\REGISTERS[23][27] ), .B1(n1154), .B2(
        \REGISTERS[22][27] ), .ZN(n1250) );
  OAI221_X1 U1735 ( .B1(n273), .B2(n1155), .C1(n308), .C2(n1156), .A(n1251), 
        .ZN(n1246) );
  AOI22_X1 U1736 ( .A1(n1158), .A2(\REGISTERS[27][27] ), .B1(n1159), .B2(
        \REGISTERS[26][27] ), .ZN(n1251) );
  OAI221_X1 U1737 ( .B1(n58), .B2(n1160), .C1(n98), .C2(n1161), .A(n1252), 
        .ZN(n1245) );
  AOI22_X1 U1738 ( .A1(n1163), .A2(\REGISTERS[29][27] ), .B1(n1164), .B2(
        \REGISTERS[28][27] ), .ZN(n1252) );
  NOR4_X1 U1739 ( .A1(n1253), .A2(n1254), .A3(n1255), .A4(n1256), .ZN(n1243)
         );
  OAI221_X1 U1740 ( .B1(n1100), .B2(n1169), .C1(n1134), .C2(n1170), .A(n1257), 
        .ZN(n1256) );
  AOI22_X1 U1741 ( .A1(n1172), .A2(\REGISTERS[3][27] ), .B1(n1173), .B2(
        \REGISTERS[2][27] ), .ZN(n1257) );
  OAI221_X1 U1742 ( .B1(n964), .B2(n1174), .C1(n998), .C2(n1175), .A(n1258), 
        .ZN(n1255) );
  AOI22_X1 U1743 ( .A1(n1177), .A2(\REGISTERS[7][27] ), .B1(n1178), .B2(
        \REGISTERS[6][27] ), .ZN(n1258) );
  OAI221_X1 U1744 ( .B1(n823), .B2(n1179), .C1(n857), .C2(n1180), .A(n1259), 
        .ZN(n1254) );
  AOI22_X1 U1745 ( .A1(n1182), .A2(\REGISTERS[11][27] ), .B1(n1183), .B2(
        \REGISTERS[10][27] ), .ZN(n1259) );
  OAI221_X1 U1746 ( .B1(n687), .B2(n1184), .C1(n721), .C2(n1185), .A(n1260), 
        .ZN(n1253) );
  AOI22_X1 U1747 ( .A1(n1187), .A2(\REGISTERS[15][27] ), .B1(n1188), .B2(
        \REGISTERS[14][27] ), .ZN(n1260) );
  AOI21_X1 U1748 ( .B1(n1261), .B2(n1262), .A(N352), .ZN(N346) );
  NOR4_X1 U1749 ( .A1(n1263), .A2(n1264), .A3(n1265), .A4(n1266), .ZN(n1262)
         );
  OAI221_X1 U1750 ( .B1(n548), .B2(n1145), .C1(n582), .C2(n1146), .A(n1267), 
        .ZN(n1266) );
  AOI22_X1 U1751 ( .A1(n1148), .A2(\REGISTERS[19][26] ), .B1(n1149), .B2(
        \REGISTERS[18][26] ), .ZN(n1267) );
  OAI221_X1 U1752 ( .B1(n412), .B2(n1150), .C1(n446), .C2(n1151), .A(n1268), 
        .ZN(n1265) );
  AOI22_X1 U1753 ( .A1(n1153), .A2(\REGISTERS[23][26] ), .B1(n1154), .B2(
        \REGISTERS[22][26] ), .ZN(n1268) );
  OAI221_X1 U1754 ( .B1(n272), .B2(n1155), .C1(n307), .C2(n1156), .A(n1269), 
        .ZN(n1264) );
  AOI22_X1 U1755 ( .A1(n1158), .A2(\REGISTERS[27][26] ), .B1(n1159), .B2(
        \REGISTERS[26][26] ), .ZN(n1269) );
  OAI221_X1 U1756 ( .B1(n56), .B2(n1160), .C1(n97), .C2(n1161), .A(n1270), 
        .ZN(n1263) );
  AOI22_X1 U1757 ( .A1(n1163), .A2(\REGISTERS[29][26] ), .B1(n1164), .B2(
        \REGISTERS[28][26] ), .ZN(n1270) );
  NOR4_X1 U1758 ( .A1(n1271), .A2(n1272), .A3(n1273), .A4(n1274), .ZN(n1261)
         );
  OAI221_X1 U1759 ( .B1(n1099), .B2(n1169), .C1(n1133), .C2(n1170), .A(n1275), 
        .ZN(n1274) );
  AOI22_X1 U1760 ( .A1(n1172), .A2(\REGISTERS[3][26] ), .B1(n1173), .B2(
        \REGISTERS[2][26] ), .ZN(n1275) );
  OAI221_X1 U1761 ( .B1(n963), .B2(n1174), .C1(n997), .C2(n1175), .A(n1276), 
        .ZN(n1273) );
  AOI22_X1 U1762 ( .A1(n1177), .A2(\REGISTERS[7][26] ), .B1(n1178), .B2(
        \REGISTERS[6][26] ), .ZN(n1276) );
  OAI221_X1 U1763 ( .B1(n822), .B2(n1179), .C1(n856), .C2(n1180), .A(n1277), 
        .ZN(n1272) );
  AOI22_X1 U1764 ( .A1(n1182), .A2(\REGISTERS[11][26] ), .B1(n1183), .B2(
        \REGISTERS[10][26] ), .ZN(n1277) );
  OAI221_X1 U1765 ( .B1(n686), .B2(n1184), .C1(n720), .C2(n1185), .A(n1278), 
        .ZN(n1271) );
  AOI22_X1 U1766 ( .A1(n1187), .A2(\REGISTERS[15][26] ), .B1(n1188), .B2(
        \REGISTERS[14][26] ), .ZN(n1278) );
  AOI21_X1 U1767 ( .B1(n1279), .B2(n1280), .A(N352), .ZN(N345) );
  NOR4_X1 U1768 ( .A1(n1281), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1280)
         );
  OAI221_X1 U1769 ( .B1(n547), .B2(n1145), .C1(n581), .C2(n1146), .A(n1285), 
        .ZN(n1284) );
  AOI22_X1 U1770 ( .A1(n1148), .A2(\REGISTERS[19][25] ), .B1(n1149), .B2(
        \REGISTERS[18][25] ), .ZN(n1285) );
  OAI221_X1 U1771 ( .B1(n411), .B2(n1150), .C1(n445), .C2(n1151), .A(n1286), 
        .ZN(n1283) );
  AOI22_X1 U1772 ( .A1(n1153), .A2(\REGISTERS[23][25] ), .B1(n1154), .B2(
        \REGISTERS[22][25] ), .ZN(n1286) );
  OAI221_X1 U1773 ( .B1(n271), .B2(n1155), .C1(n306), .C2(n1156), .A(n1287), 
        .ZN(n1282) );
  AOI22_X1 U1774 ( .A1(n1158), .A2(\REGISTERS[27][25] ), .B1(n1159), .B2(
        \REGISTERS[26][25] ), .ZN(n1287) );
  OAI221_X1 U1775 ( .B1(n54), .B2(n1160), .C1(n96), .C2(n1161), .A(n1288), 
        .ZN(n1281) );
  AOI22_X1 U1776 ( .A1(n1163), .A2(\REGISTERS[29][25] ), .B1(n1164), .B2(
        \REGISTERS[28][25] ), .ZN(n1288) );
  NOR4_X1 U1777 ( .A1(n1289), .A2(n1290), .A3(n1291), .A4(n1292), .ZN(n1279)
         );
  OAI221_X1 U1778 ( .B1(n1098), .B2(n1169), .C1(n1132), .C2(n1170), .A(n1293), 
        .ZN(n1292) );
  AOI22_X1 U1779 ( .A1(n1172), .A2(\REGISTERS[3][25] ), .B1(n1173), .B2(
        \REGISTERS[2][25] ), .ZN(n1293) );
  OAI221_X1 U1780 ( .B1(n962), .B2(n1174), .C1(n996), .C2(n1175), .A(n1294), 
        .ZN(n1291) );
  AOI22_X1 U1781 ( .A1(n1177), .A2(\REGISTERS[7][25] ), .B1(n1178), .B2(
        \REGISTERS[6][25] ), .ZN(n1294) );
  OAI221_X1 U1782 ( .B1(n821), .B2(n1179), .C1(n855), .C2(n1180), .A(n1295), 
        .ZN(n1290) );
  AOI22_X1 U1783 ( .A1(n1182), .A2(\REGISTERS[11][25] ), .B1(n1183), .B2(
        \REGISTERS[10][25] ), .ZN(n1295) );
  OAI221_X1 U1784 ( .B1(n685), .B2(n1184), .C1(n719), .C2(n1185), .A(n1296), 
        .ZN(n1289) );
  AOI22_X1 U1785 ( .A1(n1187), .A2(\REGISTERS[15][25] ), .B1(n1188), .B2(
        \REGISTERS[14][25] ), .ZN(n1296) );
  AOI21_X1 U1786 ( .B1(n1297), .B2(n1298), .A(N352), .ZN(N344) );
  NOR4_X1 U1787 ( .A1(n1299), .A2(n1300), .A3(n1301), .A4(n1302), .ZN(n1298)
         );
  OAI221_X1 U1788 ( .B1(n546), .B2(n1145), .C1(n580), .C2(n1146), .A(n1303), 
        .ZN(n1302) );
  AOI22_X1 U1789 ( .A1(n1148), .A2(\REGISTERS[19][24] ), .B1(n1149), .B2(
        \REGISTERS[18][24] ), .ZN(n1303) );
  OAI221_X1 U1790 ( .B1(n410), .B2(n1150), .C1(n444), .C2(n1151), .A(n1304), 
        .ZN(n1301) );
  AOI22_X1 U1791 ( .A1(n1153), .A2(\REGISTERS[23][24] ), .B1(n1154), .B2(
        \REGISTERS[22][24] ), .ZN(n1304) );
  OAI221_X1 U1792 ( .B1(n270), .B2(n1155), .C1(n305), .C2(n1156), .A(n1305), 
        .ZN(n1300) );
  AOI22_X1 U1793 ( .A1(n1158), .A2(\REGISTERS[27][24] ), .B1(n1159), .B2(
        \REGISTERS[26][24] ), .ZN(n1305) );
  OAI221_X1 U1794 ( .B1(n52), .B2(n1160), .C1(n95), .C2(n1161), .A(n1306), 
        .ZN(n1299) );
  AOI22_X1 U1795 ( .A1(n1163), .A2(\REGISTERS[29][24] ), .B1(n1164), .B2(
        \REGISTERS[28][24] ), .ZN(n1306) );
  NOR4_X1 U1796 ( .A1(n1307), .A2(n1308), .A3(n1309), .A4(n1310), .ZN(n1297)
         );
  OAI221_X1 U1797 ( .B1(n1097), .B2(n1169), .C1(n1131), .C2(n1170), .A(n1311), 
        .ZN(n1310) );
  AOI22_X1 U1798 ( .A1(n1172), .A2(\REGISTERS[3][24] ), .B1(n1173), .B2(
        \REGISTERS[2][24] ), .ZN(n1311) );
  OAI221_X1 U1799 ( .B1(n961), .B2(n1174), .C1(n995), .C2(n1175), .A(n1312), 
        .ZN(n1309) );
  AOI22_X1 U1800 ( .A1(n1177), .A2(\REGISTERS[7][24] ), .B1(n1178), .B2(
        \REGISTERS[6][24] ), .ZN(n1312) );
  OAI221_X1 U1801 ( .B1(n820), .B2(n1179), .C1(n854), .C2(n1180), .A(n1313), 
        .ZN(n1308) );
  AOI22_X1 U1802 ( .A1(n1182), .A2(\REGISTERS[11][24] ), .B1(n1183), .B2(
        \REGISTERS[10][24] ), .ZN(n1313) );
  OAI221_X1 U1803 ( .B1(n684), .B2(n1184), .C1(n718), .C2(n1185), .A(n1314), 
        .ZN(n1307) );
  AOI22_X1 U1804 ( .A1(n1187), .A2(\REGISTERS[15][24] ), .B1(n1188), .B2(
        \REGISTERS[14][24] ), .ZN(n1314) );
  AOI21_X1 U1805 ( .B1(n1315), .B2(n1316), .A(N352), .ZN(N343) );
  NOR4_X1 U1806 ( .A1(n1317), .A2(n1318), .A3(n1319), .A4(n1320), .ZN(n1316)
         );
  OAI221_X1 U1807 ( .B1(n545), .B2(n1145), .C1(n579), .C2(n1146), .A(n1321), 
        .ZN(n1320) );
  AOI22_X1 U1808 ( .A1(n1148), .A2(\REGISTERS[19][23] ), .B1(n1149), .B2(
        \REGISTERS[18][23] ), .ZN(n1321) );
  OAI221_X1 U1809 ( .B1(n409), .B2(n1150), .C1(n443), .C2(n1151), .A(n1322), 
        .ZN(n1319) );
  AOI22_X1 U1810 ( .A1(n1153), .A2(\REGISTERS[23][23] ), .B1(n1154), .B2(
        \REGISTERS[22][23] ), .ZN(n1322) );
  OAI221_X1 U1811 ( .B1(n269), .B2(n1155), .C1(n304), .C2(n1156), .A(n1323), 
        .ZN(n1318) );
  AOI22_X1 U1812 ( .A1(n1158), .A2(\REGISTERS[27][23] ), .B1(n1159), .B2(
        \REGISTERS[26][23] ), .ZN(n1323) );
  OAI221_X1 U1813 ( .B1(n50), .B2(n1160), .C1(n94), .C2(n1161), .A(n1324), 
        .ZN(n1317) );
  AOI22_X1 U1814 ( .A1(n1163), .A2(\REGISTERS[29][23] ), .B1(n1164), .B2(
        \REGISTERS[28][23] ), .ZN(n1324) );
  NOR4_X1 U1815 ( .A1(n1325), .A2(n1326), .A3(n1327), .A4(n1328), .ZN(n1315)
         );
  OAI221_X1 U1816 ( .B1(n1096), .B2(n1169), .C1(n1130), .C2(n1170), .A(n1329), 
        .ZN(n1328) );
  AOI22_X1 U1817 ( .A1(n1172), .A2(\REGISTERS[3][23] ), .B1(n1173), .B2(
        \REGISTERS[2][23] ), .ZN(n1329) );
  OAI221_X1 U1818 ( .B1(n960), .B2(n1174), .C1(n994), .C2(n1175), .A(n1330), 
        .ZN(n1327) );
  AOI22_X1 U1819 ( .A1(n1177), .A2(\REGISTERS[7][23] ), .B1(n1178), .B2(
        \REGISTERS[6][23] ), .ZN(n1330) );
  OAI221_X1 U1820 ( .B1(n819), .B2(n1179), .C1(n853), .C2(n1180), .A(n1331), 
        .ZN(n1326) );
  AOI22_X1 U1821 ( .A1(n1182), .A2(\REGISTERS[11][23] ), .B1(n1183), .B2(
        \REGISTERS[10][23] ), .ZN(n1331) );
  OAI221_X1 U1822 ( .B1(n683), .B2(n1184), .C1(n717), .C2(n1185), .A(n1332), 
        .ZN(n1325) );
  AOI22_X1 U1823 ( .A1(n1187), .A2(\REGISTERS[15][23] ), .B1(n1188), .B2(
        \REGISTERS[14][23] ), .ZN(n1332) );
  AOI21_X1 U1824 ( .B1(n1333), .B2(n1334), .A(N352), .ZN(N342) );
  NOR4_X1 U1825 ( .A1(n1335), .A2(n1336), .A3(n1337), .A4(n1338), .ZN(n1334)
         );
  OAI221_X1 U1826 ( .B1(n544), .B2(n1145), .C1(n578), .C2(n1146), .A(n1339), 
        .ZN(n1338) );
  AOI22_X1 U1827 ( .A1(n1148), .A2(\REGISTERS[19][22] ), .B1(n1149), .B2(
        \REGISTERS[18][22] ), .ZN(n1339) );
  OAI221_X1 U1828 ( .B1(n408), .B2(n1150), .C1(n442), .C2(n1151), .A(n1340), 
        .ZN(n1337) );
  AOI22_X1 U1829 ( .A1(n1153), .A2(\REGISTERS[23][22] ), .B1(n1154), .B2(
        \REGISTERS[22][22] ), .ZN(n1340) );
  OAI221_X1 U1830 ( .B1(n268), .B2(n1155), .C1(n303), .C2(n1156), .A(n1341), 
        .ZN(n1336) );
  AOI22_X1 U1831 ( .A1(n1158), .A2(\REGISTERS[27][22] ), .B1(n1159), .B2(
        \REGISTERS[26][22] ), .ZN(n1341) );
  OAI221_X1 U1832 ( .B1(n48), .B2(n1160), .C1(n93), .C2(n1161), .A(n1342), 
        .ZN(n1335) );
  AOI22_X1 U1833 ( .A1(n1163), .A2(\REGISTERS[29][22] ), .B1(n1164), .B2(
        \REGISTERS[28][22] ), .ZN(n1342) );
  NOR4_X1 U1834 ( .A1(n1343), .A2(n1344), .A3(n1345), .A4(n1346), .ZN(n1333)
         );
  OAI221_X1 U1835 ( .B1(n1095), .B2(n1169), .C1(n1129), .C2(n1170), .A(n1347), 
        .ZN(n1346) );
  AOI22_X1 U1836 ( .A1(n1172), .A2(\REGISTERS[3][22] ), .B1(n1173), .B2(
        \REGISTERS[2][22] ), .ZN(n1347) );
  OAI221_X1 U1837 ( .B1(n959), .B2(n1174), .C1(n993), .C2(n1175), .A(n1348), 
        .ZN(n1345) );
  AOI22_X1 U1838 ( .A1(n1177), .A2(\REGISTERS[7][22] ), .B1(n1178), .B2(
        \REGISTERS[6][22] ), .ZN(n1348) );
  OAI221_X1 U1839 ( .B1(n818), .B2(n1179), .C1(n852), .C2(n1180), .A(n1349), 
        .ZN(n1344) );
  AOI22_X1 U1840 ( .A1(n1182), .A2(\REGISTERS[11][22] ), .B1(n1183), .B2(
        \REGISTERS[10][22] ), .ZN(n1349) );
  OAI221_X1 U1841 ( .B1(n682), .B2(n1184), .C1(n716), .C2(n1185), .A(n1350), 
        .ZN(n1343) );
  AOI22_X1 U1842 ( .A1(n1187), .A2(\REGISTERS[15][22] ), .B1(n1188), .B2(
        \REGISTERS[14][22] ), .ZN(n1350) );
  AOI21_X1 U1843 ( .B1(n1351), .B2(n1352), .A(N352), .ZN(N341) );
  NOR4_X1 U1844 ( .A1(n1353), .A2(n1354), .A3(n1355), .A4(n1356), .ZN(n1352)
         );
  OAI221_X1 U1845 ( .B1(n543), .B2(n1145), .C1(n577), .C2(n1146), .A(n1357), 
        .ZN(n1356) );
  AOI22_X1 U1846 ( .A1(n1148), .A2(\REGISTERS[19][21] ), .B1(n1149), .B2(
        \REGISTERS[18][21] ), .ZN(n1357) );
  OAI221_X1 U1847 ( .B1(n407), .B2(n1150), .C1(n441), .C2(n1151), .A(n1358), 
        .ZN(n1355) );
  AOI22_X1 U1848 ( .A1(n1153), .A2(\REGISTERS[23][21] ), .B1(n1154), .B2(
        \REGISTERS[22][21] ), .ZN(n1358) );
  OAI221_X1 U1849 ( .B1(n267), .B2(n1155), .C1(n302), .C2(n1156), .A(n1359), 
        .ZN(n1354) );
  AOI22_X1 U1850 ( .A1(n1158), .A2(\REGISTERS[27][21] ), .B1(n1159), .B2(
        \REGISTERS[26][21] ), .ZN(n1359) );
  OAI221_X1 U1851 ( .B1(n46), .B2(n1160), .C1(n92), .C2(n1161), .A(n1360), 
        .ZN(n1353) );
  AOI22_X1 U1852 ( .A1(n1163), .A2(\REGISTERS[29][21] ), .B1(n1164), .B2(
        \REGISTERS[28][21] ), .ZN(n1360) );
  NOR4_X1 U1853 ( .A1(n1361), .A2(n1362), .A3(n1363), .A4(n1364), .ZN(n1351)
         );
  OAI221_X1 U1854 ( .B1(n1094), .B2(n1169), .C1(n1128), .C2(n1170), .A(n1365), 
        .ZN(n1364) );
  AOI22_X1 U1855 ( .A1(n1172), .A2(\REGISTERS[3][21] ), .B1(n1173), .B2(
        \REGISTERS[2][21] ), .ZN(n1365) );
  OAI221_X1 U1856 ( .B1(n958), .B2(n1174), .C1(n992), .C2(n1175), .A(n1366), 
        .ZN(n1363) );
  AOI22_X1 U1857 ( .A1(n1177), .A2(\REGISTERS[7][21] ), .B1(n1178), .B2(
        \REGISTERS[6][21] ), .ZN(n1366) );
  OAI221_X1 U1858 ( .B1(n817), .B2(n1179), .C1(n851), .C2(n1180), .A(n1367), 
        .ZN(n1362) );
  AOI22_X1 U1859 ( .A1(n1182), .A2(\REGISTERS[11][21] ), .B1(n1183), .B2(
        \REGISTERS[10][21] ), .ZN(n1367) );
  OAI221_X1 U1860 ( .B1(n681), .B2(n1184), .C1(n715), .C2(n1185), .A(n1368), 
        .ZN(n1361) );
  AOI22_X1 U1861 ( .A1(n1187), .A2(\REGISTERS[15][21] ), .B1(n1188), .B2(
        \REGISTERS[14][21] ), .ZN(n1368) );
  AOI21_X1 U1862 ( .B1(n1369), .B2(n1370), .A(N352), .ZN(N340) );
  NOR4_X1 U1863 ( .A1(n1371), .A2(n1372), .A3(n1373), .A4(n1374), .ZN(n1370)
         );
  OAI221_X1 U1864 ( .B1(n542), .B2(n1145), .C1(n576), .C2(n1146), .A(n1375), 
        .ZN(n1374) );
  AOI22_X1 U1865 ( .A1(n1148), .A2(\REGISTERS[19][20] ), .B1(n1149), .B2(
        \REGISTERS[18][20] ), .ZN(n1375) );
  OAI221_X1 U1866 ( .B1(n406), .B2(n1150), .C1(n440), .C2(n1151), .A(n1376), 
        .ZN(n1373) );
  AOI22_X1 U1867 ( .A1(n1153), .A2(\REGISTERS[23][20] ), .B1(n1154), .B2(
        \REGISTERS[22][20] ), .ZN(n1376) );
  OAI221_X1 U1868 ( .B1(n266), .B2(n1155), .C1(n301), .C2(n1156), .A(n1377), 
        .ZN(n1372) );
  AOI22_X1 U1869 ( .A1(n1158), .A2(\REGISTERS[27][20] ), .B1(n1159), .B2(
        \REGISTERS[26][20] ), .ZN(n1377) );
  OAI221_X1 U1870 ( .B1(n44), .B2(n1160), .C1(n91), .C2(n1161), .A(n1378), 
        .ZN(n1371) );
  AOI22_X1 U1871 ( .A1(n1163), .A2(\REGISTERS[29][20] ), .B1(n1164), .B2(
        \REGISTERS[28][20] ), .ZN(n1378) );
  NOR4_X1 U1872 ( .A1(n1379), .A2(n1380), .A3(n1381), .A4(n1382), .ZN(n1369)
         );
  OAI221_X1 U1873 ( .B1(n1093), .B2(n1169), .C1(n1127), .C2(n1170), .A(n1383), 
        .ZN(n1382) );
  AOI22_X1 U1874 ( .A1(n1172), .A2(\REGISTERS[3][20] ), .B1(n1173), .B2(
        \REGISTERS[2][20] ), .ZN(n1383) );
  OAI221_X1 U1875 ( .B1(n957), .B2(n1174), .C1(n991), .C2(n1175), .A(n1384), 
        .ZN(n1381) );
  AOI22_X1 U1876 ( .A1(n1177), .A2(\REGISTERS[7][20] ), .B1(n1178), .B2(
        \REGISTERS[6][20] ), .ZN(n1384) );
  OAI221_X1 U1877 ( .B1(n816), .B2(n1179), .C1(n850), .C2(n1180), .A(n1385), 
        .ZN(n1380) );
  AOI22_X1 U1878 ( .A1(n1182), .A2(\REGISTERS[11][20] ), .B1(n1183), .B2(
        \REGISTERS[10][20] ), .ZN(n1385) );
  OAI221_X1 U1879 ( .B1(n680), .B2(n1184), .C1(n714), .C2(n1185), .A(n1386), 
        .ZN(n1379) );
  AOI22_X1 U1880 ( .A1(n1187), .A2(\REGISTERS[15][20] ), .B1(n1188), .B2(
        \REGISTERS[14][20] ), .ZN(n1386) );
  AOI21_X1 U1881 ( .B1(n1387), .B2(n1388), .A(N352), .ZN(N339) );
  NOR4_X1 U1882 ( .A1(n1389), .A2(n1390), .A3(n1391), .A4(n1392), .ZN(n1388)
         );
  OAI221_X1 U1883 ( .B1(n541), .B2(n1145), .C1(n575), .C2(n1146), .A(n1393), 
        .ZN(n1392) );
  AOI22_X1 U1884 ( .A1(n1148), .A2(\REGISTERS[19][19] ), .B1(n1149), .B2(
        \REGISTERS[18][19] ), .ZN(n1393) );
  OAI221_X1 U1885 ( .B1(n405), .B2(n1150), .C1(n439), .C2(n1151), .A(n1394), 
        .ZN(n1391) );
  AOI22_X1 U1886 ( .A1(n1153), .A2(\REGISTERS[23][19] ), .B1(n1154), .B2(
        \REGISTERS[22][19] ), .ZN(n1394) );
  OAI221_X1 U1887 ( .B1(n265), .B2(n1155), .C1(n300), .C2(n1156), .A(n1395), 
        .ZN(n1390) );
  AOI22_X1 U1888 ( .A1(n1158), .A2(\REGISTERS[27][19] ), .B1(n1159), .B2(
        \REGISTERS[26][19] ), .ZN(n1395) );
  OAI221_X1 U1889 ( .B1(n42), .B2(n1160), .C1(n90), .C2(n1161), .A(n1396), 
        .ZN(n1389) );
  AOI22_X1 U1890 ( .A1(n1163), .A2(\REGISTERS[29][19] ), .B1(n1164), .B2(
        \REGISTERS[28][19] ), .ZN(n1396) );
  NOR4_X1 U1891 ( .A1(n1397), .A2(n1398), .A3(n1399), .A4(n1400), .ZN(n1387)
         );
  OAI221_X1 U1892 ( .B1(n1092), .B2(n1169), .C1(n1126), .C2(n1170), .A(n1401), 
        .ZN(n1400) );
  AOI22_X1 U1893 ( .A1(n1172), .A2(\REGISTERS[3][19] ), .B1(n1173), .B2(
        \REGISTERS[2][19] ), .ZN(n1401) );
  OAI221_X1 U1894 ( .B1(n956), .B2(n1174), .C1(n990), .C2(n1175), .A(n1402), 
        .ZN(n1399) );
  AOI22_X1 U1895 ( .A1(n1177), .A2(\REGISTERS[7][19] ), .B1(n1178), .B2(
        \REGISTERS[6][19] ), .ZN(n1402) );
  OAI221_X1 U1896 ( .B1(n815), .B2(n1179), .C1(n849), .C2(n1180), .A(n1403), 
        .ZN(n1398) );
  AOI22_X1 U1897 ( .A1(n1182), .A2(\REGISTERS[11][19] ), .B1(n1183), .B2(
        \REGISTERS[10][19] ), .ZN(n1403) );
  OAI221_X1 U1898 ( .B1(n679), .B2(n1184), .C1(n713), .C2(n1185), .A(n1404), 
        .ZN(n1397) );
  AOI22_X1 U1899 ( .A1(n1187), .A2(\REGISTERS[15][19] ), .B1(n1188), .B2(
        \REGISTERS[14][19] ), .ZN(n1404) );
  AOI21_X1 U1900 ( .B1(n1405), .B2(n1406), .A(N352), .ZN(N338) );
  NOR4_X1 U1901 ( .A1(n1407), .A2(n1408), .A3(n1409), .A4(n1410), .ZN(n1406)
         );
  OAI221_X1 U1902 ( .B1(n540), .B2(n1145), .C1(n574), .C2(n1146), .A(n1411), 
        .ZN(n1410) );
  AOI22_X1 U1903 ( .A1(n1148), .A2(\REGISTERS[19][18] ), .B1(n1149), .B2(
        \REGISTERS[18][18] ), .ZN(n1411) );
  OAI221_X1 U1904 ( .B1(n404), .B2(n1150), .C1(n438), .C2(n1151), .A(n1412), 
        .ZN(n1409) );
  AOI22_X1 U1905 ( .A1(n1153), .A2(\REGISTERS[23][18] ), .B1(n1154), .B2(
        \REGISTERS[22][18] ), .ZN(n1412) );
  OAI221_X1 U1906 ( .B1(n264), .B2(n1155), .C1(n299), .C2(n1156), .A(n1413), 
        .ZN(n1408) );
  AOI22_X1 U1907 ( .A1(n1158), .A2(\REGISTERS[27][18] ), .B1(n1159), .B2(
        \REGISTERS[26][18] ), .ZN(n1413) );
  OAI221_X1 U1908 ( .B1(n40), .B2(n1160), .C1(n89), .C2(n1161), .A(n1414), 
        .ZN(n1407) );
  AOI22_X1 U1909 ( .A1(n1163), .A2(\REGISTERS[29][18] ), .B1(n1164), .B2(
        \REGISTERS[28][18] ), .ZN(n1414) );
  NOR4_X1 U1910 ( .A1(n1415), .A2(n1416), .A3(n1417), .A4(n1418), .ZN(n1405)
         );
  OAI221_X1 U1911 ( .B1(n1091), .B2(n1169), .C1(n1125), .C2(n1170), .A(n1419), 
        .ZN(n1418) );
  AOI22_X1 U1912 ( .A1(n1172), .A2(\REGISTERS[3][18] ), .B1(n1173), .B2(
        \REGISTERS[2][18] ), .ZN(n1419) );
  OAI221_X1 U1913 ( .B1(n955), .B2(n1174), .C1(n989), .C2(n1175), .A(n1420), 
        .ZN(n1417) );
  AOI22_X1 U1914 ( .A1(n1177), .A2(\REGISTERS[7][18] ), .B1(n1178), .B2(
        \REGISTERS[6][18] ), .ZN(n1420) );
  OAI221_X1 U1915 ( .B1(n814), .B2(n1179), .C1(n848), .C2(n1180), .A(n1421), 
        .ZN(n1416) );
  AOI22_X1 U1916 ( .A1(n1182), .A2(\REGISTERS[11][18] ), .B1(n1183), .B2(
        \REGISTERS[10][18] ), .ZN(n1421) );
  OAI221_X1 U1917 ( .B1(n678), .B2(n1184), .C1(n712), .C2(n1185), .A(n1422), 
        .ZN(n1415) );
  AOI22_X1 U1918 ( .A1(n1187), .A2(\REGISTERS[15][18] ), .B1(n1188), .B2(
        \REGISTERS[14][18] ), .ZN(n1422) );
  AOI21_X1 U1919 ( .B1(n1423), .B2(n1424), .A(N352), .ZN(N337) );
  NOR4_X1 U1920 ( .A1(n1425), .A2(n1426), .A3(n1427), .A4(n1428), .ZN(n1424)
         );
  OAI221_X1 U1921 ( .B1(n539), .B2(n1145), .C1(n573), .C2(n1146), .A(n1429), 
        .ZN(n1428) );
  AOI22_X1 U1922 ( .A1(n1148), .A2(\REGISTERS[19][17] ), .B1(n1149), .B2(
        \REGISTERS[18][17] ), .ZN(n1429) );
  OAI221_X1 U1923 ( .B1(n403), .B2(n1150), .C1(n437), .C2(n1151), .A(n1430), 
        .ZN(n1427) );
  AOI22_X1 U1924 ( .A1(n1153), .A2(\REGISTERS[23][17] ), .B1(n1154), .B2(
        \REGISTERS[22][17] ), .ZN(n1430) );
  OAI221_X1 U1925 ( .B1(n263), .B2(n1155), .C1(n298), .C2(n1156), .A(n1431), 
        .ZN(n1426) );
  AOI22_X1 U1926 ( .A1(n1158), .A2(\REGISTERS[27][17] ), .B1(n1159), .B2(
        \REGISTERS[26][17] ), .ZN(n1431) );
  OAI221_X1 U1927 ( .B1(n38), .B2(n1160), .C1(n88), .C2(n1161), .A(n1432), 
        .ZN(n1425) );
  AOI22_X1 U1928 ( .A1(n1163), .A2(\REGISTERS[29][17] ), .B1(n1164), .B2(
        \REGISTERS[28][17] ), .ZN(n1432) );
  NOR4_X1 U1929 ( .A1(n1433), .A2(n1434), .A3(n1435), .A4(n1436), .ZN(n1423)
         );
  OAI221_X1 U1930 ( .B1(n1090), .B2(n1169), .C1(n1124), .C2(n1170), .A(n1437), 
        .ZN(n1436) );
  AOI22_X1 U1931 ( .A1(n1172), .A2(\REGISTERS[3][17] ), .B1(n1173), .B2(
        \REGISTERS[2][17] ), .ZN(n1437) );
  OAI221_X1 U1932 ( .B1(n954), .B2(n1174), .C1(n988), .C2(n1175), .A(n1438), 
        .ZN(n1435) );
  AOI22_X1 U1933 ( .A1(n1177), .A2(\REGISTERS[7][17] ), .B1(n1178), .B2(
        \REGISTERS[6][17] ), .ZN(n1438) );
  OAI221_X1 U1934 ( .B1(n813), .B2(n1179), .C1(n847), .C2(n1180), .A(n1439), 
        .ZN(n1434) );
  AOI22_X1 U1935 ( .A1(n1182), .A2(\REGISTERS[11][17] ), .B1(n1183), .B2(
        \REGISTERS[10][17] ), .ZN(n1439) );
  OAI221_X1 U1936 ( .B1(n677), .B2(n1184), .C1(n711), .C2(n1185), .A(n1440), 
        .ZN(n1433) );
  AOI22_X1 U1937 ( .A1(n1187), .A2(\REGISTERS[15][17] ), .B1(n1188), .B2(
        \REGISTERS[14][17] ), .ZN(n1440) );
  AOI21_X1 U1938 ( .B1(n1441), .B2(n1442), .A(N352), .ZN(N336) );
  NOR4_X1 U1939 ( .A1(n1443), .A2(n1444), .A3(n1445), .A4(n1446), .ZN(n1442)
         );
  OAI221_X1 U1940 ( .B1(n538), .B2(n1145), .C1(n572), .C2(n1146), .A(n1447), 
        .ZN(n1446) );
  AOI22_X1 U1941 ( .A1(n1148), .A2(\REGISTERS[19][16] ), .B1(n1149), .B2(
        \REGISTERS[18][16] ), .ZN(n1447) );
  OAI221_X1 U1942 ( .B1(n402), .B2(n1150), .C1(n436), .C2(n1151), .A(n1448), 
        .ZN(n1445) );
  AOI22_X1 U1943 ( .A1(n1153), .A2(\REGISTERS[23][16] ), .B1(n1154), .B2(
        \REGISTERS[22][16] ), .ZN(n1448) );
  OAI221_X1 U1944 ( .B1(n262), .B2(n1155), .C1(n297), .C2(n1156), .A(n1449), 
        .ZN(n1444) );
  AOI22_X1 U1945 ( .A1(n1158), .A2(\REGISTERS[27][16] ), .B1(n1159), .B2(
        \REGISTERS[26][16] ), .ZN(n1449) );
  OAI221_X1 U1946 ( .B1(n36), .B2(n1160), .C1(n87), .C2(n1161), .A(n1450), 
        .ZN(n1443) );
  AOI22_X1 U1947 ( .A1(n1163), .A2(\REGISTERS[29][16] ), .B1(n1164), .B2(
        \REGISTERS[28][16] ), .ZN(n1450) );
  NOR4_X1 U1948 ( .A1(n1451), .A2(n1452), .A3(n1453), .A4(n1454), .ZN(n1441)
         );
  OAI221_X1 U1949 ( .B1(n1089), .B2(n1169), .C1(n1123), .C2(n1170), .A(n1455), 
        .ZN(n1454) );
  AOI22_X1 U1950 ( .A1(n1172), .A2(\REGISTERS[3][16] ), .B1(n1173), .B2(
        \REGISTERS[2][16] ), .ZN(n1455) );
  OAI221_X1 U1951 ( .B1(n953), .B2(n1174), .C1(n987), .C2(n1175), .A(n1456), 
        .ZN(n1453) );
  AOI22_X1 U1952 ( .A1(n1177), .A2(\REGISTERS[7][16] ), .B1(n1178), .B2(
        \REGISTERS[6][16] ), .ZN(n1456) );
  OAI221_X1 U1953 ( .B1(n812), .B2(n1179), .C1(n846), .C2(n1180), .A(n1457), 
        .ZN(n1452) );
  AOI22_X1 U1954 ( .A1(n1182), .A2(\REGISTERS[11][16] ), .B1(n1183), .B2(
        \REGISTERS[10][16] ), .ZN(n1457) );
  OAI221_X1 U1955 ( .B1(n676), .B2(n1184), .C1(n710), .C2(n1185), .A(n1458), 
        .ZN(n1451) );
  AOI22_X1 U1956 ( .A1(n1187), .A2(\REGISTERS[15][16] ), .B1(n1188), .B2(
        \REGISTERS[14][16] ), .ZN(n1458) );
  AOI21_X1 U1957 ( .B1(n1459), .B2(n1460), .A(N352), .ZN(N335) );
  NOR4_X1 U1958 ( .A1(n1461), .A2(n1462), .A3(n1463), .A4(n1464), .ZN(n1460)
         );
  OAI221_X1 U1959 ( .B1(n537), .B2(n1145), .C1(n571), .C2(n1146), .A(n1465), 
        .ZN(n1464) );
  AOI22_X1 U1960 ( .A1(n1148), .A2(\REGISTERS[19][15] ), .B1(n1149), .B2(
        \REGISTERS[18][15] ), .ZN(n1465) );
  OAI221_X1 U1961 ( .B1(n401), .B2(n1150), .C1(n435), .C2(n1151), .A(n1466), 
        .ZN(n1463) );
  AOI22_X1 U1962 ( .A1(n1153), .A2(\REGISTERS[23][15] ), .B1(n1154), .B2(
        \REGISTERS[22][15] ), .ZN(n1466) );
  OAI221_X1 U1963 ( .B1(n261), .B2(n1155), .C1(n296), .C2(n1156), .A(n1467), 
        .ZN(n1462) );
  AOI22_X1 U1964 ( .A1(n1158), .A2(\REGISTERS[27][15] ), .B1(n1159), .B2(
        \REGISTERS[26][15] ), .ZN(n1467) );
  OAI221_X1 U1965 ( .B1(n34), .B2(n1160), .C1(n86), .C2(n1161), .A(n1468), 
        .ZN(n1461) );
  AOI22_X1 U1966 ( .A1(n1163), .A2(\REGISTERS[29][15] ), .B1(n1164), .B2(
        \REGISTERS[28][15] ), .ZN(n1468) );
  NOR4_X1 U1967 ( .A1(n1469), .A2(n1470), .A3(n1471), .A4(n1472), .ZN(n1459)
         );
  OAI221_X1 U1968 ( .B1(n1088), .B2(n1169), .C1(n1122), .C2(n1170), .A(n1473), 
        .ZN(n1472) );
  AOI22_X1 U1969 ( .A1(n1172), .A2(\REGISTERS[3][15] ), .B1(n1173), .B2(
        \REGISTERS[2][15] ), .ZN(n1473) );
  OAI221_X1 U1970 ( .B1(n952), .B2(n1174), .C1(n986), .C2(n1175), .A(n1474), 
        .ZN(n1471) );
  AOI22_X1 U1971 ( .A1(n1177), .A2(\REGISTERS[7][15] ), .B1(n1178), .B2(
        \REGISTERS[6][15] ), .ZN(n1474) );
  OAI221_X1 U1972 ( .B1(n811), .B2(n1179), .C1(n845), .C2(n1180), .A(n1475), 
        .ZN(n1470) );
  AOI22_X1 U1973 ( .A1(n1182), .A2(\REGISTERS[11][15] ), .B1(n1183), .B2(
        \REGISTERS[10][15] ), .ZN(n1475) );
  OAI221_X1 U1974 ( .B1(n675), .B2(n1184), .C1(n709), .C2(n1185), .A(n1476), 
        .ZN(n1469) );
  AOI22_X1 U1975 ( .A1(n1187), .A2(\REGISTERS[15][15] ), .B1(n1188), .B2(
        \REGISTERS[14][15] ), .ZN(n1476) );
  AOI21_X1 U1976 ( .B1(n1477), .B2(n1478), .A(N352), .ZN(N334) );
  NOR4_X1 U1977 ( .A1(n1479), .A2(n1480), .A3(n1481), .A4(n1482), .ZN(n1478)
         );
  OAI221_X1 U1978 ( .B1(n536), .B2(n1145), .C1(n570), .C2(n1146), .A(n1483), 
        .ZN(n1482) );
  AOI22_X1 U1979 ( .A1(n1148), .A2(\REGISTERS[19][14] ), .B1(n1149), .B2(
        \REGISTERS[18][14] ), .ZN(n1483) );
  OAI221_X1 U1980 ( .B1(n400), .B2(n1150), .C1(n434), .C2(n1151), .A(n1484), 
        .ZN(n1481) );
  AOI22_X1 U1981 ( .A1(n1153), .A2(\REGISTERS[23][14] ), .B1(n1154), .B2(
        \REGISTERS[22][14] ), .ZN(n1484) );
  OAI221_X1 U1982 ( .B1(n260), .B2(n1155), .C1(n295), .C2(n1156), .A(n1485), 
        .ZN(n1480) );
  AOI22_X1 U1983 ( .A1(n1158), .A2(\REGISTERS[27][14] ), .B1(n1159), .B2(
        \REGISTERS[26][14] ), .ZN(n1485) );
  OAI221_X1 U1984 ( .B1(n32), .B2(n1160), .C1(n85), .C2(n1161), .A(n1486), 
        .ZN(n1479) );
  AOI22_X1 U1985 ( .A1(n1163), .A2(\REGISTERS[29][14] ), .B1(n1164), .B2(
        \REGISTERS[28][14] ), .ZN(n1486) );
  NOR4_X1 U1986 ( .A1(n1487), .A2(n1488), .A3(n1489), .A4(n1490), .ZN(n1477)
         );
  OAI221_X1 U1987 ( .B1(n1087), .B2(n1169), .C1(n1121), .C2(n1170), .A(n1491), 
        .ZN(n1490) );
  AOI22_X1 U1988 ( .A1(n1172), .A2(\REGISTERS[3][14] ), .B1(n1173), .B2(
        \REGISTERS[2][14] ), .ZN(n1491) );
  OAI221_X1 U1989 ( .B1(n951), .B2(n1174), .C1(n985), .C2(n1175), .A(n1492), 
        .ZN(n1489) );
  AOI22_X1 U1990 ( .A1(n1177), .A2(\REGISTERS[7][14] ), .B1(n1178), .B2(
        \REGISTERS[6][14] ), .ZN(n1492) );
  OAI221_X1 U1991 ( .B1(n810), .B2(n1179), .C1(n844), .C2(n1180), .A(n1493), 
        .ZN(n1488) );
  AOI22_X1 U1992 ( .A1(n1182), .A2(\REGISTERS[11][14] ), .B1(n1183), .B2(
        \REGISTERS[10][14] ), .ZN(n1493) );
  OAI221_X1 U1993 ( .B1(n674), .B2(n1184), .C1(n708), .C2(n1185), .A(n1494), 
        .ZN(n1487) );
  AOI22_X1 U1994 ( .A1(n1187), .A2(\REGISTERS[15][14] ), .B1(n1188), .B2(
        \REGISTERS[14][14] ), .ZN(n1494) );
  AOI21_X1 U1995 ( .B1(n1495), .B2(n1496), .A(N352), .ZN(N333) );
  NOR4_X1 U1996 ( .A1(n1497), .A2(n1498), .A3(n1499), .A4(n1500), .ZN(n1496)
         );
  OAI221_X1 U1997 ( .B1(n535), .B2(n1145), .C1(n569), .C2(n1146), .A(n1501), 
        .ZN(n1500) );
  AOI22_X1 U1998 ( .A1(n1148), .A2(\REGISTERS[19][13] ), .B1(n1149), .B2(
        \REGISTERS[18][13] ), .ZN(n1501) );
  OAI221_X1 U1999 ( .B1(n399), .B2(n1150), .C1(n433), .C2(n1151), .A(n1502), 
        .ZN(n1499) );
  AOI22_X1 U2000 ( .A1(n1153), .A2(\REGISTERS[23][13] ), .B1(n1154), .B2(
        \REGISTERS[22][13] ), .ZN(n1502) );
  OAI221_X1 U2001 ( .B1(n259), .B2(n1155), .C1(n294), .C2(n1156), .A(n1503), 
        .ZN(n1498) );
  AOI22_X1 U2002 ( .A1(n1158), .A2(\REGISTERS[27][13] ), .B1(n1159), .B2(
        \REGISTERS[26][13] ), .ZN(n1503) );
  OAI221_X1 U2003 ( .B1(n30), .B2(n1160), .C1(n84), .C2(n1161), .A(n1504), 
        .ZN(n1497) );
  AOI22_X1 U2004 ( .A1(n1163), .A2(\REGISTERS[29][13] ), .B1(n1164), .B2(
        \REGISTERS[28][13] ), .ZN(n1504) );
  NOR4_X1 U2005 ( .A1(n1505), .A2(n1506), .A3(n1507), .A4(n1508), .ZN(n1495)
         );
  OAI221_X1 U2006 ( .B1(n1086), .B2(n1169), .C1(n1120), .C2(n1170), .A(n1509), 
        .ZN(n1508) );
  AOI22_X1 U2007 ( .A1(n1172), .A2(\REGISTERS[3][13] ), .B1(n1173), .B2(
        \REGISTERS[2][13] ), .ZN(n1509) );
  OAI221_X1 U2008 ( .B1(n950), .B2(n1174), .C1(n984), .C2(n1175), .A(n1510), 
        .ZN(n1507) );
  AOI22_X1 U2009 ( .A1(n1177), .A2(\REGISTERS[7][13] ), .B1(n1178), .B2(
        \REGISTERS[6][13] ), .ZN(n1510) );
  OAI221_X1 U2010 ( .B1(n809), .B2(n1179), .C1(n843), .C2(n1180), .A(n1511), 
        .ZN(n1506) );
  AOI22_X1 U2011 ( .A1(n1182), .A2(\REGISTERS[11][13] ), .B1(n1183), .B2(
        \REGISTERS[10][13] ), .ZN(n1511) );
  OAI221_X1 U2012 ( .B1(n673), .B2(n1184), .C1(n707), .C2(n1185), .A(n1512), 
        .ZN(n1505) );
  AOI22_X1 U2013 ( .A1(n1187), .A2(\REGISTERS[15][13] ), .B1(n1188), .B2(
        \REGISTERS[14][13] ), .ZN(n1512) );
  AOI21_X1 U2014 ( .B1(n1513), .B2(n1514), .A(N352), .ZN(N332) );
  NOR4_X1 U2015 ( .A1(n1515), .A2(n1516), .A3(n1517), .A4(n1518), .ZN(n1514)
         );
  OAI221_X1 U2016 ( .B1(n534), .B2(n1145), .C1(n568), .C2(n1146), .A(n1519), 
        .ZN(n1518) );
  AOI22_X1 U2017 ( .A1(n1148), .A2(\REGISTERS[19][12] ), .B1(n1149), .B2(
        \REGISTERS[18][12] ), .ZN(n1519) );
  OAI221_X1 U2018 ( .B1(n398), .B2(n1150), .C1(n432), .C2(n1151), .A(n1520), 
        .ZN(n1517) );
  AOI22_X1 U2019 ( .A1(n1153), .A2(\REGISTERS[23][12] ), .B1(n1154), .B2(
        \REGISTERS[22][12] ), .ZN(n1520) );
  OAI221_X1 U2020 ( .B1(n258), .B2(n1155), .C1(n293), .C2(n1156), .A(n1521), 
        .ZN(n1516) );
  AOI22_X1 U2021 ( .A1(n1158), .A2(\REGISTERS[27][12] ), .B1(n1159), .B2(
        \REGISTERS[26][12] ), .ZN(n1521) );
  OAI221_X1 U2022 ( .B1(n28), .B2(n1160), .C1(n83), .C2(n1161), .A(n1522), 
        .ZN(n1515) );
  AOI22_X1 U2023 ( .A1(n1163), .A2(\REGISTERS[29][12] ), .B1(n1164), .B2(
        \REGISTERS[28][12] ), .ZN(n1522) );
  NOR4_X1 U2024 ( .A1(n1523), .A2(n1524), .A3(n1525), .A4(n1526), .ZN(n1513)
         );
  OAI221_X1 U2025 ( .B1(n1085), .B2(n1169), .C1(n1119), .C2(n1170), .A(n1527), 
        .ZN(n1526) );
  AOI22_X1 U2026 ( .A1(n1172), .A2(\REGISTERS[3][12] ), .B1(n1173), .B2(
        \REGISTERS[2][12] ), .ZN(n1527) );
  OAI221_X1 U2027 ( .B1(n949), .B2(n1174), .C1(n983), .C2(n1175), .A(n1528), 
        .ZN(n1525) );
  AOI22_X1 U2028 ( .A1(n1177), .A2(\REGISTERS[7][12] ), .B1(n1178), .B2(
        \REGISTERS[6][12] ), .ZN(n1528) );
  OAI221_X1 U2029 ( .B1(n808), .B2(n1179), .C1(n842), .C2(n1180), .A(n1529), 
        .ZN(n1524) );
  AOI22_X1 U2030 ( .A1(n1182), .A2(\REGISTERS[11][12] ), .B1(n1183), .B2(
        \REGISTERS[10][12] ), .ZN(n1529) );
  OAI221_X1 U2031 ( .B1(n672), .B2(n1184), .C1(n706), .C2(n1185), .A(n1530), 
        .ZN(n1523) );
  AOI22_X1 U2032 ( .A1(n1187), .A2(\REGISTERS[15][12] ), .B1(n1188), .B2(
        \REGISTERS[14][12] ), .ZN(n1530) );
  AOI21_X1 U2033 ( .B1(n1531), .B2(n1532), .A(N352), .ZN(N331) );
  NOR4_X1 U2034 ( .A1(n1533), .A2(n1534), .A3(n1535), .A4(n1536), .ZN(n1532)
         );
  OAI221_X1 U2035 ( .B1(n533), .B2(n1145), .C1(n567), .C2(n1146), .A(n1537), 
        .ZN(n1536) );
  AOI22_X1 U2036 ( .A1(n1148), .A2(\REGISTERS[19][11] ), .B1(n1149), .B2(
        \REGISTERS[18][11] ), .ZN(n1537) );
  OAI221_X1 U2037 ( .B1(n397), .B2(n1150), .C1(n431), .C2(n1151), .A(n1538), 
        .ZN(n1535) );
  AOI22_X1 U2038 ( .A1(n1153), .A2(\REGISTERS[23][11] ), .B1(n1154), .B2(
        \REGISTERS[22][11] ), .ZN(n1538) );
  OAI221_X1 U2039 ( .B1(n257), .B2(n1155), .C1(n292), .C2(n1156), .A(n1539), 
        .ZN(n1534) );
  AOI22_X1 U2040 ( .A1(n1158), .A2(\REGISTERS[27][11] ), .B1(n1159), .B2(
        \REGISTERS[26][11] ), .ZN(n1539) );
  OAI221_X1 U2041 ( .B1(n26), .B2(n1160), .C1(n82), .C2(n1161), .A(n1540), 
        .ZN(n1533) );
  AOI22_X1 U2042 ( .A1(n1163), .A2(\REGISTERS[29][11] ), .B1(n1164), .B2(
        \REGISTERS[28][11] ), .ZN(n1540) );
  NOR4_X1 U2043 ( .A1(n1541), .A2(n1542), .A3(n1543), .A4(n1544), .ZN(n1531)
         );
  OAI221_X1 U2044 ( .B1(n1084), .B2(n1169), .C1(n1118), .C2(n1170), .A(n1545), 
        .ZN(n1544) );
  AOI22_X1 U2045 ( .A1(n1172), .A2(\REGISTERS[3][11] ), .B1(n1173), .B2(
        \REGISTERS[2][11] ), .ZN(n1545) );
  OAI221_X1 U2046 ( .B1(n948), .B2(n1174), .C1(n982), .C2(n1175), .A(n1546), 
        .ZN(n1543) );
  AOI22_X1 U2047 ( .A1(n1177), .A2(\REGISTERS[7][11] ), .B1(n1178), .B2(
        \REGISTERS[6][11] ), .ZN(n1546) );
  OAI221_X1 U2048 ( .B1(n807), .B2(n1179), .C1(n841), .C2(n1180), .A(n1547), 
        .ZN(n1542) );
  AOI22_X1 U2049 ( .A1(n1182), .A2(\REGISTERS[11][11] ), .B1(n1183), .B2(
        \REGISTERS[10][11] ), .ZN(n1547) );
  OAI221_X1 U2050 ( .B1(n671), .B2(n1184), .C1(n705), .C2(n1185), .A(n1548), 
        .ZN(n1541) );
  AOI22_X1 U2051 ( .A1(n1187), .A2(\REGISTERS[15][11] ), .B1(n1188), .B2(
        \REGISTERS[14][11] ), .ZN(n1548) );
  AOI21_X1 U2052 ( .B1(n1549), .B2(n1550), .A(N352), .ZN(N330) );
  NOR4_X1 U2053 ( .A1(n1551), .A2(n1552), .A3(n1553), .A4(n1554), .ZN(n1550)
         );
  OAI221_X1 U2054 ( .B1(n532), .B2(n1145), .C1(n566), .C2(n1146), .A(n1555), 
        .ZN(n1554) );
  AOI22_X1 U2055 ( .A1(n1148), .A2(\REGISTERS[19][10] ), .B1(n1149), .B2(
        \REGISTERS[18][10] ), .ZN(n1555) );
  OAI221_X1 U2056 ( .B1(n396), .B2(n1150), .C1(n430), .C2(n1151), .A(n1556), 
        .ZN(n1553) );
  AOI22_X1 U2057 ( .A1(n1153), .A2(\REGISTERS[23][10] ), .B1(n1154), .B2(
        \REGISTERS[22][10] ), .ZN(n1556) );
  OAI221_X1 U2058 ( .B1(n256), .B2(n1155), .C1(n291), .C2(n1156), .A(n1557), 
        .ZN(n1552) );
  AOI22_X1 U2059 ( .A1(n1158), .A2(\REGISTERS[27][10] ), .B1(n1159), .B2(
        \REGISTERS[26][10] ), .ZN(n1557) );
  OAI221_X1 U2060 ( .B1(n24), .B2(n1160), .C1(n81), .C2(n1161), .A(n1558), 
        .ZN(n1551) );
  AOI22_X1 U2061 ( .A1(n1163), .A2(\REGISTERS[29][10] ), .B1(n1164), .B2(
        \REGISTERS[28][10] ), .ZN(n1558) );
  NOR4_X1 U2062 ( .A1(n1559), .A2(n1560), .A3(n1561), .A4(n1562), .ZN(n1549)
         );
  OAI221_X1 U2063 ( .B1(n1083), .B2(n1169), .C1(n1117), .C2(n1170), .A(n1563), 
        .ZN(n1562) );
  AOI22_X1 U2064 ( .A1(n1172), .A2(\REGISTERS[3][10] ), .B1(n1173), .B2(
        \REGISTERS[2][10] ), .ZN(n1563) );
  OAI221_X1 U2065 ( .B1(n947), .B2(n1174), .C1(n981), .C2(n1175), .A(n1564), 
        .ZN(n1561) );
  AOI22_X1 U2066 ( .A1(n1177), .A2(\REGISTERS[7][10] ), .B1(n1178), .B2(
        \REGISTERS[6][10] ), .ZN(n1564) );
  OAI221_X1 U2067 ( .B1(n806), .B2(n1179), .C1(n840), .C2(n1180), .A(n1565), 
        .ZN(n1560) );
  AOI22_X1 U2068 ( .A1(n1182), .A2(\REGISTERS[11][10] ), .B1(n1183), .B2(
        \REGISTERS[10][10] ), .ZN(n1565) );
  OAI221_X1 U2069 ( .B1(n670), .B2(n1184), .C1(n704), .C2(n1185), .A(n1566), 
        .ZN(n1559) );
  AOI22_X1 U2070 ( .A1(n1187), .A2(\REGISTERS[15][10] ), .B1(n1188), .B2(
        \REGISTERS[14][10] ), .ZN(n1566) );
  AOI21_X1 U2071 ( .B1(n1567), .B2(n1568), .A(N352), .ZN(N329) );
  NOR4_X1 U2072 ( .A1(n1569), .A2(n1570), .A3(n1571), .A4(n1572), .ZN(n1568)
         );
  OAI221_X1 U2073 ( .B1(n531), .B2(n1145), .C1(n565), .C2(n1146), .A(n1573), 
        .ZN(n1572) );
  AOI22_X1 U2074 ( .A1(n1148), .A2(\REGISTERS[19][9] ), .B1(n1149), .B2(
        \REGISTERS[18][9] ), .ZN(n1573) );
  OAI221_X1 U2075 ( .B1(n395), .B2(n1150), .C1(n429), .C2(n1151), .A(n1574), 
        .ZN(n1571) );
  AOI22_X1 U2076 ( .A1(n1153), .A2(\REGISTERS[23][9] ), .B1(n1154), .B2(
        \REGISTERS[22][9] ), .ZN(n1574) );
  OAI221_X1 U2077 ( .B1(n255), .B2(n1155), .C1(n290), .C2(n1156), .A(n1575), 
        .ZN(n1570) );
  AOI22_X1 U2078 ( .A1(n1158), .A2(\REGISTERS[27][9] ), .B1(n1159), .B2(
        \REGISTERS[26][9] ), .ZN(n1575) );
  OAI221_X1 U2079 ( .B1(n22), .B2(n1160), .C1(n80), .C2(n1161), .A(n1576), 
        .ZN(n1569) );
  AOI22_X1 U2080 ( .A1(n1163), .A2(\REGISTERS[29][9] ), .B1(n1164), .B2(
        \REGISTERS[28][9] ), .ZN(n1576) );
  NOR4_X1 U2081 ( .A1(n1577), .A2(n1578), .A3(n1579), .A4(n1580), .ZN(n1567)
         );
  OAI221_X1 U2082 ( .B1(n1082), .B2(n1169), .C1(n1116), .C2(n1170), .A(n1581), 
        .ZN(n1580) );
  AOI22_X1 U2083 ( .A1(n1172), .A2(\REGISTERS[3][9] ), .B1(n1173), .B2(
        \REGISTERS[2][9] ), .ZN(n1581) );
  OAI221_X1 U2084 ( .B1(n946), .B2(n1174), .C1(n980), .C2(n1175), .A(n1582), 
        .ZN(n1579) );
  AOI22_X1 U2085 ( .A1(n1177), .A2(\REGISTERS[7][9] ), .B1(n1178), .B2(
        \REGISTERS[6][9] ), .ZN(n1582) );
  OAI221_X1 U2086 ( .B1(n805), .B2(n1179), .C1(n839), .C2(n1180), .A(n1583), 
        .ZN(n1578) );
  AOI22_X1 U2087 ( .A1(n1182), .A2(\REGISTERS[11][9] ), .B1(n1183), .B2(
        \REGISTERS[10][9] ), .ZN(n1583) );
  OAI221_X1 U2088 ( .B1(n669), .B2(n1184), .C1(n703), .C2(n1185), .A(n1584), 
        .ZN(n1577) );
  AOI22_X1 U2089 ( .A1(n1187), .A2(\REGISTERS[15][9] ), .B1(n1188), .B2(
        \REGISTERS[14][9] ), .ZN(n1584) );
  AOI21_X1 U2090 ( .B1(n1585), .B2(n1586), .A(N352), .ZN(N328) );
  NOR4_X1 U2091 ( .A1(n1587), .A2(n1588), .A3(n1589), .A4(n1590), .ZN(n1586)
         );
  OAI221_X1 U2092 ( .B1(n530), .B2(n1145), .C1(n564), .C2(n1146), .A(n1591), 
        .ZN(n1590) );
  AOI22_X1 U2093 ( .A1(n1148), .A2(\REGISTERS[19][8] ), .B1(n1149), .B2(
        \REGISTERS[18][8] ), .ZN(n1591) );
  OAI221_X1 U2094 ( .B1(n394), .B2(n1150), .C1(n428), .C2(n1151), .A(n1592), 
        .ZN(n1589) );
  AOI22_X1 U2095 ( .A1(n1153), .A2(\REGISTERS[23][8] ), .B1(n1154), .B2(
        \REGISTERS[22][8] ), .ZN(n1592) );
  OAI221_X1 U2096 ( .B1(n254), .B2(n1155), .C1(n289), .C2(n1156), .A(n1593), 
        .ZN(n1588) );
  AOI22_X1 U2097 ( .A1(n1158), .A2(\REGISTERS[27][8] ), .B1(n1159), .B2(
        \REGISTERS[26][8] ), .ZN(n1593) );
  OAI221_X1 U2098 ( .B1(n20), .B2(n1160), .C1(n79), .C2(n1161), .A(n1594), 
        .ZN(n1587) );
  AOI22_X1 U2099 ( .A1(n1163), .A2(\REGISTERS[29][8] ), .B1(n1164), .B2(
        \REGISTERS[28][8] ), .ZN(n1594) );
  NOR4_X1 U2100 ( .A1(n1595), .A2(n1596), .A3(n1597), .A4(n1598), .ZN(n1585)
         );
  OAI221_X1 U2101 ( .B1(n1081), .B2(n1169), .C1(n1115), .C2(n1170), .A(n1599), 
        .ZN(n1598) );
  AOI22_X1 U2102 ( .A1(n1172), .A2(\REGISTERS[3][8] ), .B1(n1173), .B2(
        \REGISTERS[2][8] ), .ZN(n1599) );
  OAI221_X1 U2103 ( .B1(n945), .B2(n1174), .C1(n979), .C2(n1175), .A(n1600), 
        .ZN(n1597) );
  AOI22_X1 U2104 ( .A1(n1177), .A2(\REGISTERS[7][8] ), .B1(n1178), .B2(
        \REGISTERS[6][8] ), .ZN(n1600) );
  OAI221_X1 U2105 ( .B1(n804), .B2(n1179), .C1(n838), .C2(n1180), .A(n1601), 
        .ZN(n1596) );
  AOI22_X1 U2106 ( .A1(n1182), .A2(\REGISTERS[11][8] ), .B1(n1183), .B2(
        \REGISTERS[10][8] ), .ZN(n1601) );
  OAI221_X1 U2107 ( .B1(n668), .B2(n1184), .C1(n702), .C2(n1185), .A(n1602), 
        .ZN(n1595) );
  AOI22_X1 U2108 ( .A1(n1187), .A2(\REGISTERS[15][8] ), .B1(n1188), .B2(
        \REGISTERS[14][8] ), .ZN(n1602) );
  AOI21_X1 U2109 ( .B1(n1603), .B2(n1604), .A(N352), .ZN(N327) );
  NOR4_X1 U2110 ( .A1(n1605), .A2(n1606), .A3(n1607), .A4(n1608), .ZN(n1604)
         );
  OAI221_X1 U2111 ( .B1(n529), .B2(n1145), .C1(n563), .C2(n1146), .A(n1609), 
        .ZN(n1608) );
  AOI22_X1 U2112 ( .A1(n1148), .A2(\REGISTERS[19][7] ), .B1(n1149), .B2(
        \REGISTERS[18][7] ), .ZN(n1609) );
  OAI221_X1 U2113 ( .B1(n393), .B2(n1150), .C1(n427), .C2(n1151), .A(n1610), 
        .ZN(n1607) );
  AOI22_X1 U2114 ( .A1(n1153), .A2(\REGISTERS[23][7] ), .B1(n1154), .B2(
        \REGISTERS[22][7] ), .ZN(n1610) );
  OAI221_X1 U2115 ( .B1(n253), .B2(n1155), .C1(n288), .C2(n1156), .A(n1611), 
        .ZN(n1606) );
  AOI22_X1 U2116 ( .A1(n1158), .A2(\REGISTERS[27][7] ), .B1(n1159), .B2(
        \REGISTERS[26][7] ), .ZN(n1611) );
  OAI221_X1 U2117 ( .B1(n18), .B2(n1160), .C1(n78), .C2(n1161), .A(n1612), 
        .ZN(n1605) );
  AOI22_X1 U2118 ( .A1(n1163), .A2(\REGISTERS[29][7] ), .B1(n1164), .B2(
        \REGISTERS[28][7] ), .ZN(n1612) );
  NOR4_X1 U2119 ( .A1(n1613), .A2(n1614), .A3(n1615), .A4(n1616), .ZN(n1603)
         );
  OAI221_X1 U2120 ( .B1(n1080), .B2(n1169), .C1(n1114), .C2(n1170), .A(n1617), 
        .ZN(n1616) );
  AOI22_X1 U2121 ( .A1(n1172), .A2(\REGISTERS[3][7] ), .B1(n1173), .B2(
        \REGISTERS[2][7] ), .ZN(n1617) );
  OAI221_X1 U2122 ( .B1(n944), .B2(n1174), .C1(n978), .C2(n1175), .A(n1618), 
        .ZN(n1615) );
  AOI22_X1 U2123 ( .A1(n1177), .A2(\REGISTERS[7][7] ), .B1(n1178), .B2(
        \REGISTERS[6][7] ), .ZN(n1618) );
  OAI221_X1 U2124 ( .B1(n803), .B2(n1179), .C1(n837), .C2(n1180), .A(n1619), 
        .ZN(n1614) );
  AOI22_X1 U2125 ( .A1(n1182), .A2(\REGISTERS[11][7] ), .B1(n1183), .B2(
        \REGISTERS[10][7] ), .ZN(n1619) );
  OAI221_X1 U2126 ( .B1(n667), .B2(n1184), .C1(n701), .C2(n1185), .A(n1620), 
        .ZN(n1613) );
  AOI22_X1 U2127 ( .A1(n1187), .A2(\REGISTERS[15][7] ), .B1(n1188), .B2(
        \REGISTERS[14][7] ), .ZN(n1620) );
  AOI21_X1 U2128 ( .B1(n1621), .B2(n1622), .A(N352), .ZN(N326) );
  NOR4_X1 U2129 ( .A1(n1623), .A2(n1624), .A3(n1625), .A4(n1626), .ZN(n1622)
         );
  OAI221_X1 U2130 ( .B1(n528), .B2(n1145), .C1(n562), .C2(n1146), .A(n1627), 
        .ZN(n1626) );
  AOI22_X1 U2131 ( .A1(n1148), .A2(\REGISTERS[19][6] ), .B1(n1149), .B2(
        \REGISTERS[18][6] ), .ZN(n1627) );
  OAI221_X1 U2132 ( .B1(n392), .B2(n1150), .C1(n426), .C2(n1151), .A(n1628), 
        .ZN(n1625) );
  AOI22_X1 U2133 ( .A1(n1153), .A2(\REGISTERS[23][6] ), .B1(n1154), .B2(
        \REGISTERS[22][6] ), .ZN(n1628) );
  OAI221_X1 U2134 ( .B1(n252), .B2(n1155), .C1(n287), .C2(n1156), .A(n1629), 
        .ZN(n1624) );
  AOI22_X1 U2135 ( .A1(n1158), .A2(\REGISTERS[27][6] ), .B1(n1159), .B2(
        \REGISTERS[26][6] ), .ZN(n1629) );
  OAI221_X1 U2136 ( .B1(n16), .B2(n1160), .C1(n77), .C2(n1161), .A(n1630), 
        .ZN(n1623) );
  AOI22_X1 U2137 ( .A1(n1163), .A2(\REGISTERS[29][6] ), .B1(n1164), .B2(
        \REGISTERS[28][6] ), .ZN(n1630) );
  NOR4_X1 U2138 ( .A1(n1631), .A2(n1632), .A3(n1633), .A4(n1634), .ZN(n1621)
         );
  OAI221_X1 U2139 ( .B1(n1079), .B2(n1169), .C1(n1113), .C2(n1170), .A(n1635), 
        .ZN(n1634) );
  AOI22_X1 U2140 ( .A1(n1172), .A2(\REGISTERS[3][6] ), .B1(n1173), .B2(
        \REGISTERS[2][6] ), .ZN(n1635) );
  OAI221_X1 U2141 ( .B1(n943), .B2(n1174), .C1(n977), .C2(n1175), .A(n1636), 
        .ZN(n1633) );
  AOI22_X1 U2142 ( .A1(n1177), .A2(\REGISTERS[7][6] ), .B1(n1178), .B2(
        \REGISTERS[6][6] ), .ZN(n1636) );
  OAI221_X1 U2143 ( .B1(n802), .B2(n1179), .C1(n836), .C2(n1180), .A(n1637), 
        .ZN(n1632) );
  AOI22_X1 U2144 ( .A1(n1182), .A2(\REGISTERS[11][6] ), .B1(n1183), .B2(
        \REGISTERS[10][6] ), .ZN(n1637) );
  OAI221_X1 U2145 ( .B1(n666), .B2(n1184), .C1(n700), .C2(n1185), .A(n1638), 
        .ZN(n1631) );
  AOI22_X1 U2146 ( .A1(n1187), .A2(\REGISTERS[15][6] ), .B1(n1188), .B2(
        \REGISTERS[14][6] ), .ZN(n1638) );
  AOI21_X1 U2147 ( .B1(n1639), .B2(n1640), .A(N352), .ZN(N325) );
  NOR4_X1 U2148 ( .A1(n1641), .A2(n1642), .A3(n1643), .A4(n1644), .ZN(n1640)
         );
  OAI221_X1 U2149 ( .B1(n527), .B2(n1145), .C1(n561), .C2(n1146), .A(n1645), 
        .ZN(n1644) );
  AOI22_X1 U2150 ( .A1(n1148), .A2(\REGISTERS[19][5] ), .B1(n1149), .B2(
        \REGISTERS[18][5] ), .ZN(n1645) );
  OAI221_X1 U2151 ( .B1(n391), .B2(n1150), .C1(n425), .C2(n1151), .A(n1646), 
        .ZN(n1643) );
  AOI22_X1 U2152 ( .A1(n1153), .A2(\REGISTERS[23][5] ), .B1(n1154), .B2(
        \REGISTERS[22][5] ), .ZN(n1646) );
  OAI221_X1 U2153 ( .B1(n251), .B2(n1155), .C1(n286), .C2(n1156), .A(n1647), 
        .ZN(n1642) );
  AOI22_X1 U2154 ( .A1(n1158), .A2(\REGISTERS[27][5] ), .B1(n1159), .B2(
        \REGISTERS[26][5] ), .ZN(n1647) );
  OAI221_X1 U2155 ( .B1(n14), .B2(n1160), .C1(n76), .C2(n1161), .A(n1648), 
        .ZN(n1641) );
  AOI22_X1 U2156 ( .A1(n1163), .A2(\REGISTERS[29][5] ), .B1(n1164), .B2(
        \REGISTERS[28][5] ), .ZN(n1648) );
  NOR4_X1 U2157 ( .A1(n1649), .A2(n1650), .A3(n1651), .A4(n1652), .ZN(n1639)
         );
  OAI221_X1 U2158 ( .B1(n1078), .B2(n1169), .C1(n1112), .C2(n1170), .A(n1653), 
        .ZN(n1652) );
  AOI22_X1 U2159 ( .A1(n1172), .A2(\REGISTERS[3][5] ), .B1(n1173), .B2(
        \REGISTERS[2][5] ), .ZN(n1653) );
  OAI221_X1 U2160 ( .B1(n942), .B2(n1174), .C1(n976), .C2(n1175), .A(n1654), 
        .ZN(n1651) );
  AOI22_X1 U2161 ( .A1(n1177), .A2(\REGISTERS[7][5] ), .B1(n1178), .B2(
        \REGISTERS[6][5] ), .ZN(n1654) );
  OAI221_X1 U2162 ( .B1(n801), .B2(n1179), .C1(n835), .C2(n1180), .A(n1655), 
        .ZN(n1650) );
  AOI22_X1 U2163 ( .A1(n1182), .A2(\REGISTERS[11][5] ), .B1(n1183), .B2(
        \REGISTERS[10][5] ), .ZN(n1655) );
  OAI221_X1 U2164 ( .B1(n665), .B2(n1184), .C1(n699), .C2(n1185), .A(n1656), 
        .ZN(n1649) );
  AOI22_X1 U2165 ( .A1(n1187), .A2(\REGISTERS[15][5] ), .B1(n1188), .B2(
        \REGISTERS[14][5] ), .ZN(n1656) );
  AOI21_X1 U2166 ( .B1(n1657), .B2(n1658), .A(N352), .ZN(N324) );
  NOR4_X1 U2167 ( .A1(n1659), .A2(n1660), .A3(n1661), .A4(n1662), .ZN(n1658)
         );
  OAI221_X1 U2168 ( .B1(n526), .B2(n1145), .C1(n560), .C2(n1146), .A(n1663), 
        .ZN(n1662) );
  AOI22_X1 U2169 ( .A1(n1148), .A2(\REGISTERS[19][4] ), .B1(n1149), .B2(
        \REGISTERS[18][4] ), .ZN(n1663) );
  OAI221_X1 U2170 ( .B1(n390), .B2(n1150), .C1(n424), .C2(n1151), .A(n1664), 
        .ZN(n1661) );
  AOI22_X1 U2171 ( .A1(n1153), .A2(\REGISTERS[23][4] ), .B1(n1154), .B2(
        \REGISTERS[22][4] ), .ZN(n1664) );
  OAI221_X1 U2172 ( .B1(n250), .B2(n1155), .C1(n285), .C2(n1156), .A(n1665), 
        .ZN(n1660) );
  AOI22_X1 U2173 ( .A1(n1158), .A2(\REGISTERS[27][4] ), .B1(n1159), .B2(
        \REGISTERS[26][4] ), .ZN(n1665) );
  OAI221_X1 U2174 ( .B1(n12), .B2(n1160), .C1(n75), .C2(n1161), .A(n1666), 
        .ZN(n1659) );
  AOI22_X1 U2175 ( .A1(n1163), .A2(\REGISTERS[29][4] ), .B1(n1164), .B2(
        \REGISTERS[28][4] ), .ZN(n1666) );
  NOR4_X1 U2176 ( .A1(n1667), .A2(n1668), .A3(n1669), .A4(n1670), .ZN(n1657)
         );
  OAI221_X1 U2177 ( .B1(n1077), .B2(n1169), .C1(n1111), .C2(n1170), .A(n1671), 
        .ZN(n1670) );
  AOI22_X1 U2178 ( .A1(n1172), .A2(\REGISTERS[3][4] ), .B1(n1173), .B2(
        \REGISTERS[2][4] ), .ZN(n1671) );
  OAI221_X1 U2179 ( .B1(n941), .B2(n1174), .C1(n975), .C2(n1175), .A(n1672), 
        .ZN(n1669) );
  AOI22_X1 U2180 ( .A1(n1177), .A2(\REGISTERS[7][4] ), .B1(n1178), .B2(
        \REGISTERS[6][4] ), .ZN(n1672) );
  OAI221_X1 U2181 ( .B1(n800), .B2(n1179), .C1(n834), .C2(n1180), .A(n1673), 
        .ZN(n1668) );
  AOI22_X1 U2182 ( .A1(n1182), .A2(\REGISTERS[11][4] ), .B1(n1183), .B2(
        \REGISTERS[10][4] ), .ZN(n1673) );
  OAI221_X1 U2183 ( .B1(n664), .B2(n1184), .C1(n698), .C2(n1185), .A(n1674), 
        .ZN(n1667) );
  AOI22_X1 U2184 ( .A1(n1187), .A2(\REGISTERS[15][4] ), .B1(n1188), .B2(
        \REGISTERS[14][4] ), .ZN(n1674) );
  AOI21_X1 U2185 ( .B1(n1675), .B2(n1676), .A(N352), .ZN(N323) );
  NOR4_X1 U2186 ( .A1(n1677), .A2(n1678), .A3(n1679), .A4(n1680), .ZN(n1676)
         );
  OAI221_X1 U2187 ( .B1(n525), .B2(n1145), .C1(n559), .C2(n1146), .A(n1681), 
        .ZN(n1680) );
  AOI22_X1 U2188 ( .A1(n1148), .A2(\REGISTERS[19][3] ), .B1(n1149), .B2(
        \REGISTERS[18][3] ), .ZN(n1681) );
  OAI221_X1 U2189 ( .B1(n389), .B2(n1150), .C1(n423), .C2(n1151), .A(n1682), 
        .ZN(n1679) );
  AOI22_X1 U2190 ( .A1(n1153), .A2(\REGISTERS[23][3] ), .B1(n1154), .B2(
        \REGISTERS[22][3] ), .ZN(n1682) );
  OAI221_X1 U2191 ( .B1(n249), .B2(n1155), .C1(n284), .C2(n1156), .A(n1683), 
        .ZN(n1678) );
  AOI22_X1 U2192 ( .A1(n1158), .A2(\REGISTERS[27][3] ), .B1(n1159), .B2(
        \REGISTERS[26][3] ), .ZN(n1683) );
  OAI221_X1 U2193 ( .B1(n10), .B2(n1160), .C1(n74), .C2(n1161), .A(n1684), 
        .ZN(n1677) );
  AOI22_X1 U2194 ( .A1(n1163), .A2(\REGISTERS[29][3] ), .B1(n1164), .B2(
        \REGISTERS[28][3] ), .ZN(n1684) );
  NOR4_X1 U2195 ( .A1(n1685), .A2(n1686), .A3(n1687), .A4(n1688), .ZN(n1675)
         );
  OAI221_X1 U2196 ( .B1(n1076), .B2(n1169), .C1(n1110), .C2(n1170), .A(n1689), 
        .ZN(n1688) );
  AOI22_X1 U2197 ( .A1(n1172), .A2(\REGISTERS[3][3] ), .B1(n1173), .B2(
        \REGISTERS[2][3] ), .ZN(n1689) );
  OAI221_X1 U2198 ( .B1(n940), .B2(n1174), .C1(n974), .C2(n1175), .A(n1690), 
        .ZN(n1687) );
  AOI22_X1 U2199 ( .A1(n1177), .A2(\REGISTERS[7][3] ), .B1(n1178), .B2(
        \REGISTERS[6][3] ), .ZN(n1690) );
  OAI221_X1 U2200 ( .B1(n799), .B2(n1179), .C1(n833), .C2(n1180), .A(n1691), 
        .ZN(n1686) );
  AOI22_X1 U2201 ( .A1(n1182), .A2(\REGISTERS[11][3] ), .B1(n1183), .B2(
        \REGISTERS[10][3] ), .ZN(n1691) );
  OAI221_X1 U2202 ( .B1(n663), .B2(n1184), .C1(n697), .C2(n1185), .A(n1692), 
        .ZN(n1685) );
  AOI22_X1 U2203 ( .A1(n1187), .A2(\REGISTERS[15][3] ), .B1(n1188), .B2(
        \REGISTERS[14][3] ), .ZN(n1692) );
  AOI21_X1 U2204 ( .B1(n1693), .B2(n1694), .A(N352), .ZN(N322) );
  NOR4_X1 U2205 ( .A1(n1695), .A2(n1696), .A3(n1697), .A4(n1698), .ZN(n1694)
         );
  OAI221_X1 U2206 ( .B1(n524), .B2(n1145), .C1(n558), .C2(n1146), .A(n1699), 
        .ZN(n1698) );
  AOI22_X1 U2207 ( .A1(n1148), .A2(\REGISTERS[19][2] ), .B1(n1149), .B2(
        \REGISTERS[18][2] ), .ZN(n1699) );
  OAI221_X1 U2208 ( .B1(n388), .B2(n1150), .C1(n422), .C2(n1151), .A(n1700), 
        .ZN(n1697) );
  AOI22_X1 U2209 ( .A1(n1153), .A2(\REGISTERS[23][2] ), .B1(n1154), .B2(
        \REGISTERS[22][2] ), .ZN(n1700) );
  OAI221_X1 U2210 ( .B1(n248), .B2(n1155), .C1(n283), .C2(n1156), .A(n1701), 
        .ZN(n1696) );
  AOI22_X1 U2211 ( .A1(n1158), .A2(\REGISTERS[27][2] ), .B1(n1159), .B2(
        \REGISTERS[26][2] ), .ZN(n1701) );
  OAI221_X1 U2212 ( .B1(n8), .B2(n1160), .C1(n73), .C2(n1161), .A(n1702), .ZN(
        n1695) );
  AOI22_X1 U2213 ( .A1(n1163), .A2(\REGISTERS[29][2] ), .B1(n1164), .B2(
        \REGISTERS[28][2] ), .ZN(n1702) );
  NOR4_X1 U2214 ( .A1(n1703), .A2(n1704), .A3(n1705), .A4(n1706), .ZN(n1693)
         );
  OAI221_X1 U2215 ( .B1(n1075), .B2(n1169), .C1(n1109), .C2(n1170), .A(n1707), 
        .ZN(n1706) );
  AOI22_X1 U2216 ( .A1(n1172), .A2(\REGISTERS[3][2] ), .B1(n1173), .B2(
        \REGISTERS[2][2] ), .ZN(n1707) );
  OAI221_X1 U2217 ( .B1(n939), .B2(n1174), .C1(n973), .C2(n1175), .A(n1708), 
        .ZN(n1705) );
  AOI22_X1 U2218 ( .A1(n1177), .A2(\REGISTERS[7][2] ), .B1(n1178), .B2(
        \REGISTERS[6][2] ), .ZN(n1708) );
  OAI221_X1 U2219 ( .B1(n798), .B2(n1179), .C1(n832), .C2(n1180), .A(n1709), 
        .ZN(n1704) );
  AOI22_X1 U2220 ( .A1(n1182), .A2(\REGISTERS[11][2] ), .B1(n1183), .B2(
        \REGISTERS[10][2] ), .ZN(n1709) );
  OAI221_X1 U2221 ( .B1(n662), .B2(n1184), .C1(n696), .C2(n1185), .A(n1710), 
        .ZN(n1703) );
  AOI22_X1 U2222 ( .A1(n1187), .A2(\REGISTERS[15][2] ), .B1(n1188), .B2(
        \REGISTERS[14][2] ), .ZN(n1710) );
  AOI21_X1 U2223 ( .B1(n1711), .B2(n1712), .A(N352), .ZN(N321) );
  NOR4_X1 U2224 ( .A1(n1713), .A2(n1714), .A3(n1715), .A4(n1716), .ZN(n1712)
         );
  OAI221_X1 U2225 ( .B1(n523), .B2(n1145), .C1(n557), .C2(n1146), .A(n1717), 
        .ZN(n1716) );
  AOI22_X1 U2226 ( .A1(n1148), .A2(\REGISTERS[19][1] ), .B1(n1149), .B2(
        \REGISTERS[18][1] ), .ZN(n1717) );
  OAI221_X1 U2227 ( .B1(n387), .B2(n1150), .C1(n421), .C2(n1151), .A(n1718), 
        .ZN(n1715) );
  AOI22_X1 U2228 ( .A1(n1153), .A2(\REGISTERS[23][1] ), .B1(n1154), .B2(
        \REGISTERS[22][1] ), .ZN(n1718) );
  OAI221_X1 U2229 ( .B1(n247), .B2(n1155), .C1(n282), .C2(n1156), .A(n1719), 
        .ZN(n1714) );
  AOI22_X1 U2230 ( .A1(n1158), .A2(\REGISTERS[27][1] ), .B1(n1159), .B2(
        \REGISTERS[26][1] ), .ZN(n1719) );
  OAI221_X1 U2231 ( .B1(n6), .B2(n1160), .C1(n72), .C2(n1161), .A(n1720), .ZN(
        n1713) );
  AOI22_X1 U2232 ( .A1(n1163), .A2(\REGISTERS[29][1] ), .B1(n1164), .B2(
        \REGISTERS[28][1] ), .ZN(n1720) );
  NOR4_X1 U2233 ( .A1(n1721), .A2(n1722), .A3(n1723), .A4(n1724), .ZN(n1711)
         );
  OAI221_X1 U2234 ( .B1(n1074), .B2(n1169), .C1(n1108), .C2(n1170), .A(n1725), 
        .ZN(n1724) );
  AOI22_X1 U2235 ( .A1(n1172), .A2(\REGISTERS[3][1] ), .B1(n1173), .B2(
        \REGISTERS[2][1] ), .ZN(n1725) );
  OAI221_X1 U2236 ( .B1(n938), .B2(n1174), .C1(n972), .C2(n1175), .A(n1726), 
        .ZN(n1723) );
  AOI22_X1 U2237 ( .A1(n1177), .A2(\REGISTERS[7][1] ), .B1(n1178), .B2(
        \REGISTERS[6][1] ), .ZN(n1726) );
  OAI221_X1 U2238 ( .B1(n797), .B2(n1179), .C1(n831), .C2(n1180), .A(n1727), 
        .ZN(n1722) );
  AOI22_X1 U2239 ( .A1(n1182), .A2(\REGISTERS[11][1] ), .B1(n1183), .B2(
        \REGISTERS[10][1] ), .ZN(n1727) );
  OAI221_X1 U2240 ( .B1(n661), .B2(n1184), .C1(n695), .C2(n1185), .A(n1728), 
        .ZN(n1721) );
  AOI22_X1 U2241 ( .A1(n1187), .A2(\REGISTERS[15][1] ), .B1(n1188), .B2(
        \REGISTERS[14][1] ), .ZN(n1728) );
  AOI21_X1 U2242 ( .B1(n1729), .B2(n1730), .A(N352), .ZN(N320) );
  NOR4_X1 U2243 ( .A1(n1731), .A2(n1732), .A3(n1733), .A4(n1734), .ZN(n1730)
         );
  OAI221_X1 U2244 ( .B1(n522), .B2(n1145), .C1(n556), .C2(n1146), .A(n1735), 
        .ZN(n1734) );
  AOI22_X1 U2245 ( .A1(n1148), .A2(\REGISTERS[19][0] ), .B1(n1149), .B2(
        \REGISTERS[18][0] ), .ZN(n1735) );
  OAI221_X1 U2250 ( .B1(n386), .B2(n1150), .C1(n420), .C2(n1151), .A(n1740), 
        .ZN(n1733) );
  AOI22_X1 U2251 ( .A1(n1153), .A2(\REGISTERS[23][0] ), .B1(n1154), .B2(
        \REGISTERS[22][0] ), .ZN(n1740) );
  AND2_X1 U2255 ( .A1(n1743), .A2(n1744), .ZN(n1736) );
  AND2_X1 U2257 ( .A1(n1743), .A2(ADD_RD2[0]), .ZN(n1738) );
  AND2_X1 U2258 ( .A1(ADD_RD2[4]), .A2(n1745), .ZN(n1743) );
  OAI221_X1 U2259 ( .B1(n246), .B2(n1155), .C1(n281), .C2(n1156), .A(n1746), 
        .ZN(n1732) );
  AOI22_X1 U2260 ( .A1(n1158), .A2(\REGISTERS[27][0] ), .B1(n1159), .B2(
        \REGISTERS[26][0] ), .ZN(n1746) );
  OAI221_X1 U2265 ( .B1(n4), .B2(n1160), .C1(n71), .C2(n1161), .A(n1749), .ZN(
        n1731) );
  AOI22_X1 U2266 ( .A1(n1163), .A2(\REGISTERS[29][0] ), .B1(n1164), .B2(
        \REGISTERS[28][0] ), .ZN(n1749) );
  AND2_X1 U2270 ( .A1(n1750), .A2(n1744), .ZN(n1747) );
  AND2_X1 U2272 ( .A1(ADD_RD2[0]), .A2(n1750), .ZN(n1748) );
  AND2_X1 U2273 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n1750) );
  NOR4_X1 U2274 ( .A1(n1751), .A2(n1752), .A3(n1753), .A4(n1754), .ZN(n1729)
         );
  OAI221_X1 U2275 ( .B1(n1073), .B2(n1169), .C1(n1107), .C2(n1170), .A(n1755), 
        .ZN(n1754) );
  AOI22_X1 U2276 ( .A1(n1172), .A2(\REGISTERS[3][0] ), .B1(n1173), .B2(
        \REGISTERS[2][0] ), .ZN(n1755) );
  OAI221_X1 U2281 ( .B1(n937), .B2(n1174), .C1(n971), .C2(n1175), .A(n1758), 
        .ZN(n1753) );
  AOI22_X1 U2282 ( .A1(n1177), .A2(\REGISTERS[7][0] ), .B1(n1178), .B2(
        \REGISTERS[6][0] ), .ZN(n1758) );
  AND2_X1 U2286 ( .A1(n1759), .A2(n1744), .ZN(n1756) );
  AND2_X1 U2288 ( .A1(n1759), .A2(ADD_RD2[0]), .ZN(n1757) );
  NOR2_X1 U2289 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .ZN(n1759) );
  OAI221_X1 U2290 ( .B1(n796), .B2(n1179), .C1(n830), .C2(n1180), .A(n1760), 
        .ZN(n1752) );
  AOI22_X1 U2291 ( .A1(n1182), .A2(\REGISTERS[11][0] ), .B1(n1183), .B2(
        \REGISTERS[10][0] ), .ZN(n1760) );
  NOR2_X1 U2294 ( .A1(n1763), .A2(ADD_RD2[2]), .ZN(n1737) );
  OAI221_X1 U2298 ( .B1(n660), .B2(n1184), .C1(n694), .C2(n1185), .A(n1764), 
        .ZN(n1751) );
  AOI22_X1 U2299 ( .A1(n1187), .A2(\REGISTERS[15][0] ), .B1(n1188), .B2(
        \REGISTERS[14][0] ), .ZN(n1764) );
  NOR2_X1 U2302 ( .A1(n1765), .A2(n1763), .ZN(n1741) );
  INV_X1 U2303 ( .A(ADD_RD2[1]), .ZN(n1763) );
  AND2_X1 U2305 ( .A1(n1766), .A2(n1744), .ZN(n1761) );
  INV_X1 U2306 ( .A(ADD_RD2[0]), .ZN(n1744) );
  INV_X1 U2309 ( .A(ADD_RD2[2]), .ZN(n1765) );
  AND2_X1 U2310 ( .A1(n1766), .A2(ADD_RD2[0]), .ZN(n1762) );
  NOR2_X1 U2311 ( .A1(n1745), .A2(ADD_RD2[4]), .ZN(n1766) );
  INV_X1 U2312 ( .A(ADD_RD2[3]), .ZN(n1745) );
  NAND2_X1 U2313 ( .A1(n1767), .A2(RESET), .ZN(N319) );
  NAND2_X1 U2314 ( .A1(RD2), .A2(ENABLE), .ZN(n1767) );
  AOI21_X1 U2315 ( .B1(n1768), .B2(n1769), .A(N352), .ZN(N318) );
  NOR4_X1 U2316 ( .A1(n1770), .A2(n1771), .A3(n1772), .A4(n1773), .ZN(n1769)
         );
  OAI221_X1 U2317 ( .B1(n553), .B2(n1774), .C1(n587), .C2(n1775), .A(n1776), 
        .ZN(n1773) );
  AOI22_X1 U2318 ( .A1(n1777), .A2(\REGISTERS[19][31] ), .B1(n1778), .B2(
        \REGISTERS[18][31] ), .ZN(n1776) );
  OAI221_X1 U2319 ( .B1(n417), .B2(n1779), .C1(n451), .C2(n1780), .A(n1781), 
        .ZN(n1772) );
  AOI22_X1 U2320 ( .A1(n1782), .A2(\REGISTERS[23][31] ), .B1(n1783), .B2(
        \REGISTERS[22][31] ), .ZN(n1781) );
  OAI221_X1 U2321 ( .B1(n277), .B2(n1784), .C1(n312), .C2(n1785), .A(n1786), 
        .ZN(n1771) );
  AOI22_X1 U2322 ( .A1(n1787), .A2(\REGISTERS[27][31] ), .B1(n1788), .B2(
        \REGISTERS[26][31] ), .ZN(n1786) );
  OAI221_X1 U2323 ( .B1(n66), .B2(n1789), .C1(n102), .C2(n1790), .A(n1791), 
        .ZN(n1770) );
  AOI22_X1 U2324 ( .A1(n1792), .A2(\REGISTERS[29][31] ), .B1(n1793), .B2(
        \REGISTERS[28][31] ), .ZN(n1791) );
  NOR4_X1 U2325 ( .A1(n1794), .A2(n1795), .A3(n1796), .A4(n1797), .ZN(n1768)
         );
  OAI221_X1 U2326 ( .B1(n1104), .B2(n1798), .C1(n1138), .C2(n1799), .A(n1800), 
        .ZN(n1797) );
  AOI22_X1 U2327 ( .A1(n1801), .A2(\REGISTERS[3][31] ), .B1(n1802), .B2(
        \REGISTERS[2][31] ), .ZN(n1800) );
  OAI221_X1 U2328 ( .B1(n968), .B2(n1803), .C1(n1002), .C2(n1804), .A(n1805), 
        .ZN(n1796) );
  AOI22_X1 U2329 ( .A1(n1806), .A2(\REGISTERS[7][31] ), .B1(n1807), .B2(
        \REGISTERS[6][31] ), .ZN(n1805) );
  OAI221_X1 U2330 ( .B1(n827), .B2(n1808), .C1(n861), .C2(n1809), .A(n1810), 
        .ZN(n1795) );
  AOI22_X1 U2331 ( .A1(n1811), .A2(\REGISTERS[11][31] ), .B1(n1812), .B2(
        \REGISTERS[10][31] ), .ZN(n1810) );
  OAI221_X1 U2332 ( .B1(n691), .B2(n1813), .C1(n725), .C2(n1814), .A(n1815), 
        .ZN(n1794) );
  AOI22_X1 U2333 ( .A1(n1816), .A2(\REGISTERS[15][31] ), .B1(n1817), .B2(
        \REGISTERS[14][31] ), .ZN(n1815) );
  AOI21_X1 U2334 ( .B1(n1818), .B2(n1819), .A(N352), .ZN(N317) );
  NOR4_X1 U2335 ( .A1(n1820), .A2(n1821), .A3(n1822), .A4(n1823), .ZN(n1819)
         );
  OAI221_X1 U2336 ( .B1(n552), .B2(n1774), .C1(n586), .C2(n1775), .A(n1824), 
        .ZN(n1823) );
  AOI22_X1 U2337 ( .A1(n1777), .A2(\REGISTERS[19][30] ), .B1(n1778), .B2(
        \REGISTERS[18][30] ), .ZN(n1824) );
  OAI221_X1 U2338 ( .B1(n416), .B2(n1779), .C1(n450), .C2(n1780), .A(n1825), 
        .ZN(n1822) );
  AOI22_X1 U2339 ( .A1(n1782), .A2(\REGISTERS[23][30] ), .B1(n1783), .B2(
        \REGISTERS[22][30] ), .ZN(n1825) );
  OAI221_X1 U2340 ( .B1(n276), .B2(n1784), .C1(n311), .C2(n1785), .A(n1826), 
        .ZN(n1821) );
  AOI22_X1 U2341 ( .A1(n1787), .A2(\REGISTERS[27][30] ), .B1(n1788), .B2(
        \REGISTERS[26][30] ), .ZN(n1826) );
  OAI221_X1 U2342 ( .B1(n64), .B2(n1789), .C1(n101), .C2(n1790), .A(n1827), 
        .ZN(n1820) );
  AOI22_X1 U2343 ( .A1(n1792), .A2(\REGISTERS[29][30] ), .B1(n1793), .B2(
        \REGISTERS[28][30] ), .ZN(n1827) );
  NOR4_X1 U2344 ( .A1(n1828), .A2(n1829), .A3(n1830), .A4(n1831), .ZN(n1818)
         );
  OAI221_X1 U2345 ( .B1(n1103), .B2(n1798), .C1(n1137), .C2(n1799), .A(n1832), 
        .ZN(n1831) );
  AOI22_X1 U2346 ( .A1(n1801), .A2(\REGISTERS[3][30] ), .B1(n1802), .B2(
        \REGISTERS[2][30] ), .ZN(n1832) );
  OAI221_X1 U2347 ( .B1(n967), .B2(n1803), .C1(n1001), .C2(n1804), .A(n1833), 
        .ZN(n1830) );
  AOI22_X1 U2348 ( .A1(n1806), .A2(\REGISTERS[7][30] ), .B1(n1807), .B2(
        \REGISTERS[6][30] ), .ZN(n1833) );
  OAI221_X1 U2349 ( .B1(n826), .B2(n1808), .C1(n860), .C2(n1809), .A(n1834), 
        .ZN(n1829) );
  AOI22_X1 U2350 ( .A1(n1811), .A2(\REGISTERS[11][30] ), .B1(n1812), .B2(
        \REGISTERS[10][30] ), .ZN(n1834) );
  OAI221_X1 U2351 ( .B1(n690), .B2(n1813), .C1(n724), .C2(n1814), .A(n1835), 
        .ZN(n1828) );
  AOI22_X1 U2352 ( .A1(n1816), .A2(\REGISTERS[15][30] ), .B1(n1817), .B2(
        \REGISTERS[14][30] ), .ZN(n1835) );
  AOI21_X1 U2353 ( .B1(n1836), .B2(n1837), .A(N352), .ZN(N316) );
  NOR4_X1 U2354 ( .A1(n1838), .A2(n1839), .A3(n1840), .A4(n1841), .ZN(n1837)
         );
  OAI221_X1 U2355 ( .B1(n551), .B2(n1774), .C1(n585), .C2(n1775), .A(n1842), 
        .ZN(n1841) );
  AOI22_X1 U2356 ( .A1(n1777), .A2(\REGISTERS[19][29] ), .B1(n1778), .B2(
        \REGISTERS[18][29] ), .ZN(n1842) );
  OAI221_X1 U2357 ( .B1(n415), .B2(n1779), .C1(n449), .C2(n1780), .A(n1843), 
        .ZN(n1840) );
  AOI22_X1 U2358 ( .A1(n1782), .A2(\REGISTERS[23][29] ), .B1(n1783), .B2(
        \REGISTERS[22][29] ), .ZN(n1843) );
  OAI221_X1 U2359 ( .B1(n275), .B2(n1784), .C1(n310), .C2(n1785), .A(n1844), 
        .ZN(n1839) );
  AOI22_X1 U2360 ( .A1(n1787), .A2(\REGISTERS[27][29] ), .B1(n1788), .B2(
        \REGISTERS[26][29] ), .ZN(n1844) );
  OAI221_X1 U2361 ( .B1(n62), .B2(n1789), .C1(n100), .C2(n1790), .A(n1845), 
        .ZN(n1838) );
  AOI22_X1 U2362 ( .A1(n1792), .A2(\REGISTERS[29][29] ), .B1(n1793), .B2(
        \REGISTERS[28][29] ), .ZN(n1845) );
  NOR4_X1 U2363 ( .A1(n1846), .A2(n1847), .A3(n1848), .A4(n1849), .ZN(n1836)
         );
  OAI221_X1 U2364 ( .B1(n1102), .B2(n1798), .C1(n1136), .C2(n1799), .A(n1850), 
        .ZN(n1849) );
  AOI22_X1 U2365 ( .A1(n1801), .A2(\REGISTERS[3][29] ), .B1(n1802), .B2(
        \REGISTERS[2][29] ), .ZN(n1850) );
  OAI221_X1 U2366 ( .B1(n966), .B2(n1803), .C1(n1000), .C2(n1804), .A(n1851), 
        .ZN(n1848) );
  AOI22_X1 U2367 ( .A1(n1806), .A2(\REGISTERS[7][29] ), .B1(n1807), .B2(
        \REGISTERS[6][29] ), .ZN(n1851) );
  OAI221_X1 U2368 ( .B1(n825), .B2(n1808), .C1(n859), .C2(n1809), .A(n1852), 
        .ZN(n1847) );
  AOI22_X1 U2369 ( .A1(n1811), .A2(\REGISTERS[11][29] ), .B1(n1812), .B2(
        \REGISTERS[10][29] ), .ZN(n1852) );
  OAI221_X1 U2370 ( .B1(n689), .B2(n1813), .C1(n723), .C2(n1814), .A(n1853), 
        .ZN(n1846) );
  AOI22_X1 U2371 ( .A1(n1816), .A2(\REGISTERS[15][29] ), .B1(n1817), .B2(
        \REGISTERS[14][29] ), .ZN(n1853) );
  AOI21_X1 U2372 ( .B1(n1854), .B2(n1855), .A(N352), .ZN(N315) );
  NOR4_X1 U2373 ( .A1(n1856), .A2(n1857), .A3(n1858), .A4(n1859), .ZN(n1855)
         );
  OAI221_X1 U2374 ( .B1(n550), .B2(n1774), .C1(n584), .C2(n1775), .A(n1860), 
        .ZN(n1859) );
  AOI22_X1 U2375 ( .A1(n1777), .A2(\REGISTERS[19][28] ), .B1(n1778), .B2(
        \REGISTERS[18][28] ), .ZN(n1860) );
  OAI221_X1 U2376 ( .B1(n414), .B2(n1779), .C1(n448), .C2(n1780), .A(n1861), 
        .ZN(n1858) );
  AOI22_X1 U2377 ( .A1(n1782), .A2(\REGISTERS[23][28] ), .B1(n1783), .B2(
        \REGISTERS[22][28] ), .ZN(n1861) );
  OAI221_X1 U2378 ( .B1(n274), .B2(n1784), .C1(n309), .C2(n1785), .A(n1862), 
        .ZN(n1857) );
  AOI22_X1 U2379 ( .A1(n1787), .A2(\REGISTERS[27][28] ), .B1(n1788), .B2(
        \REGISTERS[26][28] ), .ZN(n1862) );
  OAI221_X1 U2380 ( .B1(n60), .B2(n1789), .C1(n99), .C2(n1790), .A(n1863), 
        .ZN(n1856) );
  AOI22_X1 U2381 ( .A1(n1792), .A2(\REGISTERS[29][28] ), .B1(n1793), .B2(
        \REGISTERS[28][28] ), .ZN(n1863) );
  NOR4_X1 U2382 ( .A1(n1864), .A2(n1865), .A3(n1866), .A4(n1867), .ZN(n1854)
         );
  OAI221_X1 U2383 ( .B1(n1101), .B2(n1798), .C1(n1135), .C2(n1799), .A(n1868), 
        .ZN(n1867) );
  AOI22_X1 U2384 ( .A1(n1801), .A2(\REGISTERS[3][28] ), .B1(n1802), .B2(
        \REGISTERS[2][28] ), .ZN(n1868) );
  OAI221_X1 U2385 ( .B1(n965), .B2(n1803), .C1(n999), .C2(n1804), .A(n1869), 
        .ZN(n1866) );
  AOI22_X1 U2386 ( .A1(n1806), .A2(\REGISTERS[7][28] ), .B1(n1807), .B2(
        \REGISTERS[6][28] ), .ZN(n1869) );
  OAI221_X1 U2387 ( .B1(n824), .B2(n1808), .C1(n858), .C2(n1809), .A(n1870), 
        .ZN(n1865) );
  AOI22_X1 U2388 ( .A1(n1811), .A2(\REGISTERS[11][28] ), .B1(n1812), .B2(
        \REGISTERS[10][28] ), .ZN(n1870) );
  OAI221_X1 U2389 ( .B1(n688), .B2(n1813), .C1(n722), .C2(n1814), .A(n1871), 
        .ZN(n1864) );
  AOI22_X1 U2390 ( .A1(n1816), .A2(\REGISTERS[15][28] ), .B1(n1817), .B2(
        \REGISTERS[14][28] ), .ZN(n1871) );
  AOI21_X1 U2391 ( .B1(n1872), .B2(n1873), .A(N352), .ZN(N314) );
  NOR4_X1 U2392 ( .A1(n1874), .A2(n1875), .A3(n1876), .A4(n1877), .ZN(n1873)
         );
  OAI221_X1 U2393 ( .B1(n549), .B2(n1774), .C1(n583), .C2(n1775), .A(n1878), 
        .ZN(n1877) );
  AOI22_X1 U2394 ( .A1(n1777), .A2(\REGISTERS[19][27] ), .B1(n1778), .B2(
        \REGISTERS[18][27] ), .ZN(n1878) );
  OAI221_X1 U2395 ( .B1(n413), .B2(n1779), .C1(n447), .C2(n1780), .A(n1879), 
        .ZN(n1876) );
  AOI22_X1 U2396 ( .A1(n1782), .A2(\REGISTERS[23][27] ), .B1(n1783), .B2(
        \REGISTERS[22][27] ), .ZN(n1879) );
  OAI221_X1 U2397 ( .B1(n273), .B2(n1784), .C1(n308), .C2(n1785), .A(n1880), 
        .ZN(n1875) );
  AOI22_X1 U2398 ( .A1(n1787), .A2(\REGISTERS[27][27] ), .B1(n1788), .B2(
        \REGISTERS[26][27] ), .ZN(n1880) );
  OAI221_X1 U2399 ( .B1(n58), .B2(n1789), .C1(n98), .C2(n1790), .A(n1881), 
        .ZN(n1874) );
  AOI22_X1 U2400 ( .A1(n1792), .A2(\REGISTERS[29][27] ), .B1(n1793), .B2(
        \REGISTERS[28][27] ), .ZN(n1881) );
  NOR4_X1 U2401 ( .A1(n1882), .A2(n1883), .A3(n1884), .A4(n1885), .ZN(n1872)
         );
  OAI221_X1 U2402 ( .B1(n1100), .B2(n1798), .C1(n1134), .C2(n1799), .A(n1886), 
        .ZN(n1885) );
  AOI22_X1 U2403 ( .A1(n1801), .A2(\REGISTERS[3][27] ), .B1(n1802), .B2(
        \REGISTERS[2][27] ), .ZN(n1886) );
  OAI221_X1 U2404 ( .B1(n964), .B2(n1803), .C1(n998), .C2(n1804), .A(n1887), 
        .ZN(n1884) );
  AOI22_X1 U2405 ( .A1(n1806), .A2(\REGISTERS[7][27] ), .B1(n1807), .B2(
        \REGISTERS[6][27] ), .ZN(n1887) );
  OAI221_X1 U2406 ( .B1(n823), .B2(n1808), .C1(n857), .C2(n1809), .A(n1888), 
        .ZN(n1883) );
  AOI22_X1 U2407 ( .A1(n1811), .A2(\REGISTERS[11][27] ), .B1(n1812), .B2(
        \REGISTERS[10][27] ), .ZN(n1888) );
  OAI221_X1 U2408 ( .B1(n687), .B2(n1813), .C1(n721), .C2(n1814), .A(n1889), 
        .ZN(n1882) );
  AOI22_X1 U2409 ( .A1(n1816), .A2(\REGISTERS[15][27] ), .B1(n1817), .B2(
        \REGISTERS[14][27] ), .ZN(n1889) );
  AOI21_X1 U2410 ( .B1(n1890), .B2(n1891), .A(N352), .ZN(N313) );
  NOR4_X1 U2411 ( .A1(n1892), .A2(n1893), .A3(n1894), .A4(n1895), .ZN(n1891)
         );
  OAI221_X1 U2412 ( .B1(n548), .B2(n1774), .C1(n582), .C2(n1775), .A(n1896), 
        .ZN(n1895) );
  AOI22_X1 U2413 ( .A1(n1777), .A2(\REGISTERS[19][26] ), .B1(n1778), .B2(
        \REGISTERS[18][26] ), .ZN(n1896) );
  OAI221_X1 U2414 ( .B1(n412), .B2(n1779), .C1(n446), .C2(n1780), .A(n1897), 
        .ZN(n1894) );
  AOI22_X1 U2415 ( .A1(n1782), .A2(\REGISTERS[23][26] ), .B1(n1783), .B2(
        \REGISTERS[22][26] ), .ZN(n1897) );
  OAI221_X1 U2416 ( .B1(n272), .B2(n1784), .C1(n307), .C2(n1785), .A(n1898), 
        .ZN(n1893) );
  AOI22_X1 U2417 ( .A1(n1787), .A2(\REGISTERS[27][26] ), .B1(n1788), .B2(
        \REGISTERS[26][26] ), .ZN(n1898) );
  OAI221_X1 U2418 ( .B1(n56), .B2(n1789), .C1(n97), .C2(n1790), .A(n1899), 
        .ZN(n1892) );
  AOI22_X1 U2419 ( .A1(n1792), .A2(\REGISTERS[29][26] ), .B1(n1793), .B2(
        \REGISTERS[28][26] ), .ZN(n1899) );
  NOR4_X1 U2420 ( .A1(n1900), .A2(n1901), .A3(n1902), .A4(n1903), .ZN(n1890)
         );
  OAI221_X1 U2421 ( .B1(n1099), .B2(n1798), .C1(n1133), .C2(n1799), .A(n1904), 
        .ZN(n1903) );
  AOI22_X1 U2422 ( .A1(n1801), .A2(\REGISTERS[3][26] ), .B1(n1802), .B2(
        \REGISTERS[2][26] ), .ZN(n1904) );
  OAI221_X1 U2423 ( .B1(n963), .B2(n1803), .C1(n997), .C2(n1804), .A(n1905), 
        .ZN(n1902) );
  AOI22_X1 U2424 ( .A1(n1806), .A2(\REGISTERS[7][26] ), .B1(n1807), .B2(
        \REGISTERS[6][26] ), .ZN(n1905) );
  OAI221_X1 U2425 ( .B1(n822), .B2(n1808), .C1(n856), .C2(n1809), .A(n1906), 
        .ZN(n1901) );
  AOI22_X1 U2426 ( .A1(n1811), .A2(\REGISTERS[11][26] ), .B1(n1812), .B2(
        \REGISTERS[10][26] ), .ZN(n1906) );
  OAI221_X1 U2427 ( .B1(n686), .B2(n1813), .C1(n720), .C2(n1814), .A(n1907), 
        .ZN(n1900) );
  AOI22_X1 U2428 ( .A1(n1816), .A2(\REGISTERS[15][26] ), .B1(n1817), .B2(
        \REGISTERS[14][26] ), .ZN(n1907) );
  AOI21_X1 U2429 ( .B1(n1908), .B2(n1909), .A(N352), .ZN(N312) );
  NOR4_X1 U2430 ( .A1(n1910), .A2(n1911), .A3(n1912), .A4(n1913), .ZN(n1909)
         );
  OAI221_X1 U2431 ( .B1(n547), .B2(n1774), .C1(n581), .C2(n1775), .A(n1914), 
        .ZN(n1913) );
  AOI22_X1 U2432 ( .A1(n1777), .A2(\REGISTERS[19][25] ), .B1(n1778), .B2(
        \REGISTERS[18][25] ), .ZN(n1914) );
  OAI221_X1 U2433 ( .B1(n411), .B2(n1779), .C1(n445), .C2(n1780), .A(n1915), 
        .ZN(n1912) );
  AOI22_X1 U2434 ( .A1(n1782), .A2(\REGISTERS[23][25] ), .B1(n1783), .B2(
        \REGISTERS[22][25] ), .ZN(n1915) );
  OAI221_X1 U2435 ( .B1(n271), .B2(n1784), .C1(n306), .C2(n1785), .A(n1916), 
        .ZN(n1911) );
  AOI22_X1 U2436 ( .A1(n1787), .A2(\REGISTERS[27][25] ), .B1(n1788), .B2(
        \REGISTERS[26][25] ), .ZN(n1916) );
  OAI221_X1 U2437 ( .B1(n54), .B2(n1789), .C1(n96), .C2(n1790), .A(n1917), 
        .ZN(n1910) );
  AOI22_X1 U2438 ( .A1(n1792), .A2(\REGISTERS[29][25] ), .B1(n1793), .B2(
        \REGISTERS[28][25] ), .ZN(n1917) );
  NOR4_X1 U2439 ( .A1(n1918), .A2(n1919), .A3(n1920), .A4(n1921), .ZN(n1908)
         );
  OAI221_X1 U2440 ( .B1(n1098), .B2(n1798), .C1(n1132), .C2(n1799), .A(n1922), 
        .ZN(n1921) );
  AOI22_X1 U2441 ( .A1(n1801), .A2(\REGISTERS[3][25] ), .B1(n1802), .B2(
        \REGISTERS[2][25] ), .ZN(n1922) );
  OAI221_X1 U2442 ( .B1(n962), .B2(n1803), .C1(n996), .C2(n1804), .A(n1923), 
        .ZN(n1920) );
  AOI22_X1 U2443 ( .A1(n1806), .A2(\REGISTERS[7][25] ), .B1(n1807), .B2(
        \REGISTERS[6][25] ), .ZN(n1923) );
  OAI221_X1 U2444 ( .B1(n821), .B2(n1808), .C1(n855), .C2(n1809), .A(n1924), 
        .ZN(n1919) );
  AOI22_X1 U2445 ( .A1(n1811), .A2(\REGISTERS[11][25] ), .B1(n1812), .B2(
        \REGISTERS[10][25] ), .ZN(n1924) );
  OAI221_X1 U2446 ( .B1(n685), .B2(n1813), .C1(n719), .C2(n1814), .A(n1925), 
        .ZN(n1918) );
  AOI22_X1 U2447 ( .A1(n1816), .A2(\REGISTERS[15][25] ), .B1(n1817), .B2(
        \REGISTERS[14][25] ), .ZN(n1925) );
  AOI21_X1 U2448 ( .B1(n1926), .B2(n1927), .A(N352), .ZN(N311) );
  NOR4_X1 U2449 ( .A1(n1928), .A2(n1929), .A3(n1930), .A4(n1931), .ZN(n1927)
         );
  OAI221_X1 U2450 ( .B1(n546), .B2(n1774), .C1(n580), .C2(n1775), .A(n1932), 
        .ZN(n1931) );
  AOI22_X1 U2451 ( .A1(n1777), .A2(\REGISTERS[19][24] ), .B1(n1778), .B2(
        \REGISTERS[18][24] ), .ZN(n1932) );
  OAI221_X1 U2452 ( .B1(n410), .B2(n1779), .C1(n444), .C2(n1780), .A(n1933), 
        .ZN(n1930) );
  AOI22_X1 U2453 ( .A1(n1782), .A2(\REGISTERS[23][24] ), .B1(n1783), .B2(
        \REGISTERS[22][24] ), .ZN(n1933) );
  OAI221_X1 U2454 ( .B1(n270), .B2(n1784), .C1(n305), .C2(n1785), .A(n1934), 
        .ZN(n1929) );
  AOI22_X1 U2455 ( .A1(n1787), .A2(\REGISTERS[27][24] ), .B1(n1788), .B2(
        \REGISTERS[26][24] ), .ZN(n1934) );
  OAI221_X1 U2456 ( .B1(n52), .B2(n1789), .C1(n95), .C2(n1790), .A(n1935), 
        .ZN(n1928) );
  AOI22_X1 U2457 ( .A1(n1792), .A2(\REGISTERS[29][24] ), .B1(n1793), .B2(
        \REGISTERS[28][24] ), .ZN(n1935) );
  NOR4_X1 U2458 ( .A1(n1936), .A2(n1937), .A3(n1938), .A4(n1939), .ZN(n1926)
         );
  OAI221_X1 U2459 ( .B1(n1097), .B2(n1798), .C1(n1131), .C2(n1799), .A(n1940), 
        .ZN(n1939) );
  AOI22_X1 U2460 ( .A1(n1801), .A2(\REGISTERS[3][24] ), .B1(n1802), .B2(
        \REGISTERS[2][24] ), .ZN(n1940) );
  OAI221_X1 U2461 ( .B1(n961), .B2(n1803), .C1(n995), .C2(n1804), .A(n1941), 
        .ZN(n1938) );
  AOI22_X1 U2462 ( .A1(n1806), .A2(\REGISTERS[7][24] ), .B1(n1807), .B2(
        \REGISTERS[6][24] ), .ZN(n1941) );
  OAI221_X1 U2463 ( .B1(n820), .B2(n1808), .C1(n854), .C2(n1809), .A(n1942), 
        .ZN(n1937) );
  AOI22_X1 U2464 ( .A1(n1811), .A2(\REGISTERS[11][24] ), .B1(n1812), .B2(
        \REGISTERS[10][24] ), .ZN(n1942) );
  OAI221_X1 U2465 ( .B1(n684), .B2(n1813), .C1(n718), .C2(n1814), .A(n1943), 
        .ZN(n1936) );
  AOI22_X1 U2466 ( .A1(n1816), .A2(\REGISTERS[15][24] ), .B1(n1817), .B2(
        \REGISTERS[14][24] ), .ZN(n1943) );
  AOI21_X1 U2467 ( .B1(n1944), .B2(n1945), .A(N352), .ZN(N310) );
  NOR4_X1 U2468 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(n1945)
         );
  OAI221_X1 U2469 ( .B1(n545), .B2(n1774), .C1(n579), .C2(n1775), .A(n1950), 
        .ZN(n1949) );
  AOI22_X1 U2470 ( .A1(n1777), .A2(\REGISTERS[19][23] ), .B1(n1778), .B2(
        \REGISTERS[18][23] ), .ZN(n1950) );
  OAI221_X1 U2471 ( .B1(n409), .B2(n1779), .C1(n443), .C2(n1780), .A(n1951), 
        .ZN(n1948) );
  AOI22_X1 U2472 ( .A1(n1782), .A2(\REGISTERS[23][23] ), .B1(n1783), .B2(
        \REGISTERS[22][23] ), .ZN(n1951) );
  OAI221_X1 U2473 ( .B1(n269), .B2(n1784), .C1(n304), .C2(n1785), .A(n1952), 
        .ZN(n1947) );
  AOI22_X1 U2474 ( .A1(n1787), .A2(\REGISTERS[27][23] ), .B1(n1788), .B2(
        \REGISTERS[26][23] ), .ZN(n1952) );
  OAI221_X1 U2475 ( .B1(n50), .B2(n1789), .C1(n94), .C2(n1790), .A(n1953), 
        .ZN(n1946) );
  AOI22_X1 U2476 ( .A1(n1792), .A2(\REGISTERS[29][23] ), .B1(n1793), .B2(
        \REGISTERS[28][23] ), .ZN(n1953) );
  NOR4_X1 U2477 ( .A1(n1954), .A2(n1955), .A3(n1956), .A4(n1957), .ZN(n1944)
         );
  OAI221_X1 U2478 ( .B1(n1096), .B2(n1798), .C1(n1130), .C2(n1799), .A(n1958), 
        .ZN(n1957) );
  AOI22_X1 U2479 ( .A1(n1801), .A2(\REGISTERS[3][23] ), .B1(n1802), .B2(
        \REGISTERS[2][23] ), .ZN(n1958) );
  OAI221_X1 U2480 ( .B1(n960), .B2(n1803), .C1(n994), .C2(n1804), .A(n1959), 
        .ZN(n1956) );
  AOI22_X1 U2481 ( .A1(n1806), .A2(\REGISTERS[7][23] ), .B1(n1807), .B2(
        \REGISTERS[6][23] ), .ZN(n1959) );
  OAI221_X1 U2482 ( .B1(n819), .B2(n1808), .C1(n853), .C2(n1809), .A(n1960), 
        .ZN(n1955) );
  AOI22_X1 U2483 ( .A1(n1811), .A2(\REGISTERS[11][23] ), .B1(n1812), .B2(
        \REGISTERS[10][23] ), .ZN(n1960) );
  OAI221_X1 U2484 ( .B1(n683), .B2(n1813), .C1(n717), .C2(n1814), .A(n1961), 
        .ZN(n1954) );
  AOI22_X1 U2485 ( .A1(n1816), .A2(\REGISTERS[15][23] ), .B1(n1817), .B2(
        \REGISTERS[14][23] ), .ZN(n1961) );
  AOI21_X1 U2486 ( .B1(n1962), .B2(n1963), .A(N352), .ZN(N309) );
  NOR4_X1 U2487 ( .A1(n1964), .A2(n1965), .A3(n1966), .A4(n1967), .ZN(n1963)
         );
  OAI221_X1 U2488 ( .B1(n544), .B2(n1774), .C1(n578), .C2(n1775), .A(n1968), 
        .ZN(n1967) );
  AOI22_X1 U2489 ( .A1(n1777), .A2(\REGISTERS[19][22] ), .B1(n1778), .B2(
        \REGISTERS[18][22] ), .ZN(n1968) );
  OAI221_X1 U2490 ( .B1(n408), .B2(n1779), .C1(n442), .C2(n1780), .A(n1969), 
        .ZN(n1966) );
  AOI22_X1 U2491 ( .A1(n1782), .A2(\REGISTERS[23][22] ), .B1(n1783), .B2(
        \REGISTERS[22][22] ), .ZN(n1969) );
  OAI221_X1 U2492 ( .B1(n268), .B2(n1784), .C1(n303), .C2(n1785), .A(n1970), 
        .ZN(n1965) );
  AOI22_X1 U2493 ( .A1(n1787), .A2(\REGISTERS[27][22] ), .B1(n1788), .B2(
        \REGISTERS[26][22] ), .ZN(n1970) );
  OAI221_X1 U2494 ( .B1(n48), .B2(n1789), .C1(n93), .C2(n1790), .A(n1971), 
        .ZN(n1964) );
  AOI22_X1 U2495 ( .A1(n1792), .A2(\REGISTERS[29][22] ), .B1(n1793), .B2(
        \REGISTERS[28][22] ), .ZN(n1971) );
  NOR4_X1 U2496 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .ZN(n1962)
         );
  OAI221_X1 U2497 ( .B1(n1095), .B2(n1798), .C1(n1129), .C2(n1799), .A(n1976), 
        .ZN(n1975) );
  AOI22_X1 U2498 ( .A1(n1801), .A2(\REGISTERS[3][22] ), .B1(n1802), .B2(
        \REGISTERS[2][22] ), .ZN(n1976) );
  OAI221_X1 U2499 ( .B1(n959), .B2(n1803), .C1(n993), .C2(n1804), .A(n1977), 
        .ZN(n1974) );
  AOI22_X1 U2500 ( .A1(n1806), .A2(\REGISTERS[7][22] ), .B1(n1807), .B2(
        \REGISTERS[6][22] ), .ZN(n1977) );
  OAI221_X1 U2501 ( .B1(n818), .B2(n1808), .C1(n852), .C2(n1809), .A(n1978), 
        .ZN(n1973) );
  AOI22_X1 U2502 ( .A1(n1811), .A2(\REGISTERS[11][22] ), .B1(n1812), .B2(
        \REGISTERS[10][22] ), .ZN(n1978) );
  OAI221_X1 U2503 ( .B1(n682), .B2(n1813), .C1(n716), .C2(n1814), .A(n1979), 
        .ZN(n1972) );
  AOI22_X1 U2504 ( .A1(n1816), .A2(\REGISTERS[15][22] ), .B1(n1817), .B2(
        \REGISTERS[14][22] ), .ZN(n1979) );
  AOI21_X1 U2505 ( .B1(n1980), .B2(n1981), .A(N352), .ZN(N308) );
  NOR4_X1 U2506 ( .A1(n1982), .A2(n1983), .A3(n1984), .A4(n1985), .ZN(n1981)
         );
  OAI221_X1 U2507 ( .B1(n543), .B2(n1774), .C1(n577), .C2(n1775), .A(n1986), 
        .ZN(n1985) );
  AOI22_X1 U2508 ( .A1(n1777), .A2(\REGISTERS[19][21] ), .B1(n1778), .B2(
        \REGISTERS[18][21] ), .ZN(n1986) );
  OAI221_X1 U2509 ( .B1(n407), .B2(n1779), .C1(n441), .C2(n1780), .A(n1987), 
        .ZN(n1984) );
  AOI22_X1 U2510 ( .A1(n1782), .A2(\REGISTERS[23][21] ), .B1(n1783), .B2(
        \REGISTERS[22][21] ), .ZN(n1987) );
  OAI221_X1 U2511 ( .B1(n267), .B2(n1784), .C1(n302), .C2(n1785), .A(n1988), 
        .ZN(n1983) );
  AOI22_X1 U2512 ( .A1(n1787), .A2(\REGISTERS[27][21] ), .B1(n1788), .B2(
        \REGISTERS[26][21] ), .ZN(n1988) );
  OAI221_X1 U2513 ( .B1(n46), .B2(n1789), .C1(n92), .C2(n1790), .A(n1989), 
        .ZN(n1982) );
  AOI22_X1 U2514 ( .A1(n1792), .A2(\REGISTERS[29][21] ), .B1(n1793), .B2(
        \REGISTERS[28][21] ), .ZN(n1989) );
  NOR4_X1 U2515 ( .A1(n1990), .A2(n1991), .A3(n1992), .A4(n1993), .ZN(n1980)
         );
  OAI221_X1 U2516 ( .B1(n1094), .B2(n1798), .C1(n1128), .C2(n1799), .A(n1994), 
        .ZN(n1993) );
  AOI22_X1 U2517 ( .A1(n1801), .A2(\REGISTERS[3][21] ), .B1(n1802), .B2(
        \REGISTERS[2][21] ), .ZN(n1994) );
  OAI221_X1 U2518 ( .B1(n958), .B2(n1803), .C1(n992), .C2(n1804), .A(n1995), 
        .ZN(n1992) );
  AOI22_X1 U2519 ( .A1(n1806), .A2(\REGISTERS[7][21] ), .B1(n1807), .B2(
        \REGISTERS[6][21] ), .ZN(n1995) );
  OAI221_X1 U2520 ( .B1(n817), .B2(n1808), .C1(n851), .C2(n1809), .A(n1996), 
        .ZN(n1991) );
  AOI22_X1 U2521 ( .A1(n1811), .A2(\REGISTERS[11][21] ), .B1(n1812), .B2(
        \REGISTERS[10][21] ), .ZN(n1996) );
  OAI221_X1 U2522 ( .B1(n681), .B2(n1813), .C1(n715), .C2(n1814), .A(n1997), 
        .ZN(n1990) );
  AOI22_X1 U2523 ( .A1(n1816), .A2(\REGISTERS[15][21] ), .B1(n1817), .B2(
        \REGISTERS[14][21] ), .ZN(n1997) );
  AOI21_X1 U2524 ( .B1(n1998), .B2(n1999), .A(N352), .ZN(N307) );
  NOR4_X1 U2525 ( .A1(n2000), .A2(n2001), .A3(n2002), .A4(n2003), .ZN(n1999)
         );
  OAI221_X1 U2526 ( .B1(n542), .B2(n1774), .C1(n576), .C2(n1775), .A(n2004), 
        .ZN(n2003) );
  AOI22_X1 U2527 ( .A1(n1777), .A2(\REGISTERS[19][20] ), .B1(n1778), .B2(
        \REGISTERS[18][20] ), .ZN(n2004) );
  OAI221_X1 U2528 ( .B1(n406), .B2(n1779), .C1(n440), .C2(n1780), .A(n2005), 
        .ZN(n2002) );
  AOI22_X1 U2529 ( .A1(n1782), .A2(\REGISTERS[23][20] ), .B1(n1783), .B2(
        \REGISTERS[22][20] ), .ZN(n2005) );
  OAI221_X1 U2530 ( .B1(n266), .B2(n1784), .C1(n301), .C2(n1785), .A(n2006), 
        .ZN(n2001) );
  AOI22_X1 U2531 ( .A1(n1787), .A2(\REGISTERS[27][20] ), .B1(n1788), .B2(
        \REGISTERS[26][20] ), .ZN(n2006) );
  OAI221_X1 U2532 ( .B1(n44), .B2(n1789), .C1(n91), .C2(n1790), .A(n2007), 
        .ZN(n2000) );
  AOI22_X1 U2533 ( .A1(n1792), .A2(\REGISTERS[29][20] ), .B1(n1793), .B2(
        \REGISTERS[28][20] ), .ZN(n2007) );
  NOR4_X1 U2534 ( .A1(n2008), .A2(n2009), .A3(n2010), .A4(n2011), .ZN(n1998)
         );
  OAI221_X1 U2535 ( .B1(n1093), .B2(n1798), .C1(n1127), .C2(n1799), .A(n2012), 
        .ZN(n2011) );
  AOI22_X1 U2536 ( .A1(n1801), .A2(\REGISTERS[3][20] ), .B1(n1802), .B2(
        \REGISTERS[2][20] ), .ZN(n2012) );
  OAI221_X1 U2537 ( .B1(n957), .B2(n1803), .C1(n991), .C2(n1804), .A(n2013), 
        .ZN(n2010) );
  AOI22_X1 U2538 ( .A1(n1806), .A2(\REGISTERS[7][20] ), .B1(n1807), .B2(
        \REGISTERS[6][20] ), .ZN(n2013) );
  OAI221_X1 U2539 ( .B1(n816), .B2(n1808), .C1(n850), .C2(n1809), .A(n2014), 
        .ZN(n2009) );
  AOI22_X1 U2540 ( .A1(n1811), .A2(\REGISTERS[11][20] ), .B1(n1812), .B2(
        \REGISTERS[10][20] ), .ZN(n2014) );
  OAI221_X1 U2541 ( .B1(n680), .B2(n1813), .C1(n714), .C2(n1814), .A(n2015), 
        .ZN(n2008) );
  AOI22_X1 U2542 ( .A1(n1816), .A2(\REGISTERS[15][20] ), .B1(n1817), .B2(
        \REGISTERS[14][20] ), .ZN(n2015) );
  AOI21_X1 U2543 ( .B1(n2016), .B2(n2017), .A(N352), .ZN(N306) );
  NOR4_X1 U2544 ( .A1(n2018), .A2(n2019), .A3(n2020), .A4(n2021), .ZN(n2017)
         );
  OAI221_X1 U2545 ( .B1(n541), .B2(n1774), .C1(n575), .C2(n1775), .A(n2022), 
        .ZN(n2021) );
  AOI22_X1 U2546 ( .A1(n1777), .A2(\REGISTERS[19][19] ), .B1(n1778), .B2(
        \REGISTERS[18][19] ), .ZN(n2022) );
  OAI221_X1 U2547 ( .B1(n405), .B2(n1779), .C1(n439), .C2(n1780), .A(n2023), 
        .ZN(n2020) );
  AOI22_X1 U2548 ( .A1(n1782), .A2(\REGISTERS[23][19] ), .B1(n1783), .B2(
        \REGISTERS[22][19] ), .ZN(n2023) );
  OAI221_X1 U2549 ( .B1(n265), .B2(n1784), .C1(n300), .C2(n1785), .A(n2024), 
        .ZN(n2019) );
  AOI22_X1 U2550 ( .A1(n1787), .A2(\REGISTERS[27][19] ), .B1(n1788), .B2(
        \REGISTERS[26][19] ), .ZN(n2024) );
  OAI221_X1 U2551 ( .B1(n42), .B2(n1789), .C1(n90), .C2(n1790), .A(n2025), 
        .ZN(n2018) );
  AOI22_X1 U2552 ( .A1(n1792), .A2(\REGISTERS[29][19] ), .B1(n1793), .B2(
        \REGISTERS[28][19] ), .ZN(n2025) );
  NOR4_X1 U2553 ( .A1(n2026), .A2(n2027), .A3(n2028), .A4(n2029), .ZN(n2016)
         );
  OAI221_X1 U2554 ( .B1(n1092), .B2(n1798), .C1(n1126), .C2(n1799), .A(n2030), 
        .ZN(n2029) );
  AOI22_X1 U2555 ( .A1(n1801), .A2(\REGISTERS[3][19] ), .B1(n1802), .B2(
        \REGISTERS[2][19] ), .ZN(n2030) );
  OAI221_X1 U2556 ( .B1(n956), .B2(n1803), .C1(n990), .C2(n1804), .A(n2031), 
        .ZN(n2028) );
  AOI22_X1 U2557 ( .A1(n1806), .A2(\REGISTERS[7][19] ), .B1(n1807), .B2(
        \REGISTERS[6][19] ), .ZN(n2031) );
  OAI221_X1 U2558 ( .B1(n815), .B2(n1808), .C1(n849), .C2(n1809), .A(n2032), 
        .ZN(n2027) );
  AOI22_X1 U2559 ( .A1(n1811), .A2(\REGISTERS[11][19] ), .B1(n1812), .B2(
        \REGISTERS[10][19] ), .ZN(n2032) );
  OAI221_X1 U2560 ( .B1(n679), .B2(n1813), .C1(n713), .C2(n1814), .A(n2033), 
        .ZN(n2026) );
  AOI22_X1 U2561 ( .A1(n1816), .A2(\REGISTERS[15][19] ), .B1(n1817), .B2(
        \REGISTERS[14][19] ), .ZN(n2033) );
  AOI21_X1 U2562 ( .B1(n2034), .B2(n2035), .A(N352), .ZN(N305) );
  NOR4_X1 U2563 ( .A1(n2036), .A2(n2037), .A3(n2038), .A4(n2039), .ZN(n2035)
         );
  OAI221_X1 U2564 ( .B1(n540), .B2(n1774), .C1(n574), .C2(n1775), .A(n2040), 
        .ZN(n2039) );
  AOI22_X1 U2565 ( .A1(n1777), .A2(\REGISTERS[19][18] ), .B1(n1778), .B2(
        \REGISTERS[18][18] ), .ZN(n2040) );
  OAI221_X1 U2566 ( .B1(n404), .B2(n1779), .C1(n438), .C2(n1780), .A(n2041), 
        .ZN(n2038) );
  AOI22_X1 U2567 ( .A1(n1782), .A2(\REGISTERS[23][18] ), .B1(n1783), .B2(
        \REGISTERS[22][18] ), .ZN(n2041) );
  OAI221_X1 U2568 ( .B1(n264), .B2(n1784), .C1(n299), .C2(n1785), .A(n2042), 
        .ZN(n2037) );
  AOI22_X1 U2569 ( .A1(n1787), .A2(\REGISTERS[27][18] ), .B1(n1788), .B2(
        \REGISTERS[26][18] ), .ZN(n2042) );
  OAI221_X1 U2570 ( .B1(n40), .B2(n1789), .C1(n89), .C2(n1790), .A(n2043), 
        .ZN(n2036) );
  AOI22_X1 U2571 ( .A1(n1792), .A2(\REGISTERS[29][18] ), .B1(n1793), .B2(
        \REGISTERS[28][18] ), .ZN(n2043) );
  NOR4_X1 U2572 ( .A1(n2044), .A2(n2045), .A3(n2046), .A4(n2047), .ZN(n2034)
         );
  OAI221_X1 U2573 ( .B1(n1091), .B2(n1798), .C1(n1125), .C2(n1799), .A(n2048), 
        .ZN(n2047) );
  AOI22_X1 U2574 ( .A1(n1801), .A2(\REGISTERS[3][18] ), .B1(n1802), .B2(
        \REGISTERS[2][18] ), .ZN(n2048) );
  OAI221_X1 U2575 ( .B1(n955), .B2(n1803), .C1(n989), .C2(n1804), .A(n2049), 
        .ZN(n2046) );
  AOI22_X1 U2576 ( .A1(n1806), .A2(\REGISTERS[7][18] ), .B1(n1807), .B2(
        \REGISTERS[6][18] ), .ZN(n2049) );
  OAI221_X1 U2577 ( .B1(n814), .B2(n1808), .C1(n848), .C2(n1809), .A(n2050), 
        .ZN(n2045) );
  AOI22_X1 U2578 ( .A1(n1811), .A2(\REGISTERS[11][18] ), .B1(n1812), .B2(
        \REGISTERS[10][18] ), .ZN(n2050) );
  OAI221_X1 U2579 ( .B1(n678), .B2(n1813), .C1(n712), .C2(n1814), .A(n2051), 
        .ZN(n2044) );
  AOI22_X1 U2580 ( .A1(n1816), .A2(\REGISTERS[15][18] ), .B1(n1817), .B2(
        \REGISTERS[14][18] ), .ZN(n2051) );
  AOI21_X1 U2581 ( .B1(n2052), .B2(n2053), .A(N352), .ZN(N304) );
  NOR4_X1 U2582 ( .A1(n2054), .A2(n2055), .A3(n2056), .A4(n2057), .ZN(n2053)
         );
  OAI221_X1 U2583 ( .B1(n539), .B2(n1774), .C1(n573), .C2(n1775), .A(n2058), 
        .ZN(n2057) );
  AOI22_X1 U2584 ( .A1(n1777), .A2(\REGISTERS[19][17] ), .B1(n1778), .B2(
        \REGISTERS[18][17] ), .ZN(n2058) );
  OAI221_X1 U2585 ( .B1(n403), .B2(n1779), .C1(n437), .C2(n1780), .A(n2059), 
        .ZN(n2056) );
  AOI22_X1 U2586 ( .A1(n1782), .A2(\REGISTERS[23][17] ), .B1(n1783), .B2(
        \REGISTERS[22][17] ), .ZN(n2059) );
  OAI221_X1 U2587 ( .B1(n263), .B2(n1784), .C1(n298), .C2(n1785), .A(n2060), 
        .ZN(n2055) );
  AOI22_X1 U2588 ( .A1(n1787), .A2(\REGISTERS[27][17] ), .B1(n1788), .B2(
        \REGISTERS[26][17] ), .ZN(n2060) );
  OAI221_X1 U2589 ( .B1(n38), .B2(n1789), .C1(n88), .C2(n1790), .A(n2061), 
        .ZN(n2054) );
  AOI22_X1 U2590 ( .A1(n1792), .A2(\REGISTERS[29][17] ), .B1(n1793), .B2(
        \REGISTERS[28][17] ), .ZN(n2061) );
  NOR4_X1 U2591 ( .A1(n2062), .A2(n2063), .A3(n2064), .A4(n2065), .ZN(n2052)
         );
  OAI221_X1 U2592 ( .B1(n1090), .B2(n1798), .C1(n1124), .C2(n1799), .A(n2066), 
        .ZN(n2065) );
  AOI22_X1 U2593 ( .A1(n1801), .A2(\REGISTERS[3][17] ), .B1(n1802), .B2(
        \REGISTERS[2][17] ), .ZN(n2066) );
  OAI221_X1 U2594 ( .B1(n954), .B2(n1803), .C1(n988), .C2(n1804), .A(n2067), 
        .ZN(n2064) );
  AOI22_X1 U2595 ( .A1(n1806), .A2(\REGISTERS[7][17] ), .B1(n1807), .B2(
        \REGISTERS[6][17] ), .ZN(n2067) );
  OAI221_X1 U2596 ( .B1(n813), .B2(n1808), .C1(n847), .C2(n1809), .A(n2068), 
        .ZN(n2063) );
  AOI22_X1 U2597 ( .A1(n1811), .A2(\REGISTERS[11][17] ), .B1(n1812), .B2(
        \REGISTERS[10][17] ), .ZN(n2068) );
  OAI221_X1 U2598 ( .B1(n677), .B2(n1813), .C1(n711), .C2(n1814), .A(n2069), 
        .ZN(n2062) );
  AOI22_X1 U2599 ( .A1(n1816), .A2(\REGISTERS[15][17] ), .B1(n1817), .B2(
        \REGISTERS[14][17] ), .ZN(n2069) );
  AOI21_X1 U2600 ( .B1(n2070), .B2(n2071), .A(N352), .ZN(N303) );
  NOR4_X1 U2601 ( .A1(n2072), .A2(n2073), .A3(n2074), .A4(n2075), .ZN(n2071)
         );
  OAI221_X1 U2602 ( .B1(n538), .B2(n1774), .C1(n572), .C2(n1775), .A(n2076), 
        .ZN(n2075) );
  AOI22_X1 U2603 ( .A1(n1777), .A2(\REGISTERS[19][16] ), .B1(n1778), .B2(
        \REGISTERS[18][16] ), .ZN(n2076) );
  OAI221_X1 U2604 ( .B1(n402), .B2(n1779), .C1(n436), .C2(n1780), .A(n2077), 
        .ZN(n2074) );
  AOI22_X1 U2605 ( .A1(n1782), .A2(\REGISTERS[23][16] ), .B1(n1783), .B2(
        \REGISTERS[22][16] ), .ZN(n2077) );
  OAI221_X1 U2606 ( .B1(n262), .B2(n1784), .C1(n297), .C2(n1785), .A(n2078), 
        .ZN(n2073) );
  AOI22_X1 U2607 ( .A1(n1787), .A2(\REGISTERS[27][16] ), .B1(n1788), .B2(
        \REGISTERS[26][16] ), .ZN(n2078) );
  OAI221_X1 U2608 ( .B1(n36), .B2(n1789), .C1(n87), .C2(n1790), .A(n2079), 
        .ZN(n2072) );
  AOI22_X1 U2609 ( .A1(n1792), .A2(\REGISTERS[29][16] ), .B1(n1793), .B2(
        \REGISTERS[28][16] ), .ZN(n2079) );
  NOR4_X1 U2610 ( .A1(n2080), .A2(n2081), .A3(n2082), .A4(n2083), .ZN(n2070)
         );
  OAI221_X1 U2611 ( .B1(n1089), .B2(n1798), .C1(n1123), .C2(n1799), .A(n2084), 
        .ZN(n2083) );
  AOI22_X1 U2612 ( .A1(n1801), .A2(\REGISTERS[3][16] ), .B1(n1802), .B2(
        \REGISTERS[2][16] ), .ZN(n2084) );
  OAI221_X1 U2613 ( .B1(n953), .B2(n1803), .C1(n987), .C2(n1804), .A(n2085), 
        .ZN(n2082) );
  AOI22_X1 U2614 ( .A1(n1806), .A2(\REGISTERS[7][16] ), .B1(n1807), .B2(
        \REGISTERS[6][16] ), .ZN(n2085) );
  OAI221_X1 U2615 ( .B1(n812), .B2(n1808), .C1(n846), .C2(n1809), .A(n2086), 
        .ZN(n2081) );
  AOI22_X1 U2616 ( .A1(n1811), .A2(\REGISTERS[11][16] ), .B1(n1812), .B2(
        \REGISTERS[10][16] ), .ZN(n2086) );
  OAI221_X1 U2617 ( .B1(n676), .B2(n1813), .C1(n710), .C2(n1814), .A(n2087), 
        .ZN(n2080) );
  AOI22_X1 U2618 ( .A1(n1816), .A2(\REGISTERS[15][16] ), .B1(n1817), .B2(
        \REGISTERS[14][16] ), .ZN(n2087) );
  AOI21_X1 U2619 ( .B1(n2088), .B2(n2089), .A(N352), .ZN(N302) );
  NOR4_X1 U2620 ( .A1(n2090), .A2(n2091), .A3(n2092), .A4(n2093), .ZN(n2089)
         );
  OAI221_X1 U2621 ( .B1(n537), .B2(n1774), .C1(n571), .C2(n1775), .A(n2094), 
        .ZN(n2093) );
  AOI22_X1 U2622 ( .A1(n1777), .A2(\REGISTERS[19][15] ), .B1(n1778), .B2(
        \REGISTERS[18][15] ), .ZN(n2094) );
  OAI221_X1 U2623 ( .B1(n401), .B2(n1779), .C1(n435), .C2(n1780), .A(n2095), 
        .ZN(n2092) );
  AOI22_X1 U2624 ( .A1(n1782), .A2(\REGISTERS[23][15] ), .B1(n1783), .B2(
        \REGISTERS[22][15] ), .ZN(n2095) );
  OAI221_X1 U2625 ( .B1(n261), .B2(n1784), .C1(n296), .C2(n1785), .A(n2096), 
        .ZN(n2091) );
  AOI22_X1 U2626 ( .A1(n1787), .A2(\REGISTERS[27][15] ), .B1(n1788), .B2(
        \REGISTERS[26][15] ), .ZN(n2096) );
  OAI221_X1 U2627 ( .B1(n34), .B2(n1789), .C1(n86), .C2(n1790), .A(n2097), 
        .ZN(n2090) );
  AOI22_X1 U2628 ( .A1(n1792), .A2(\REGISTERS[29][15] ), .B1(n1793), .B2(
        \REGISTERS[28][15] ), .ZN(n2097) );
  NOR4_X1 U2629 ( .A1(n2098), .A2(n2099), .A3(n2100), .A4(n2101), .ZN(n2088)
         );
  OAI221_X1 U2630 ( .B1(n1088), .B2(n1798), .C1(n1122), .C2(n1799), .A(n2102), 
        .ZN(n2101) );
  AOI22_X1 U2631 ( .A1(n1801), .A2(\REGISTERS[3][15] ), .B1(n1802), .B2(
        \REGISTERS[2][15] ), .ZN(n2102) );
  OAI221_X1 U2632 ( .B1(n952), .B2(n1803), .C1(n986), .C2(n1804), .A(n2103), 
        .ZN(n2100) );
  AOI22_X1 U2633 ( .A1(n1806), .A2(\REGISTERS[7][15] ), .B1(n1807), .B2(
        \REGISTERS[6][15] ), .ZN(n2103) );
  OAI221_X1 U2634 ( .B1(n811), .B2(n1808), .C1(n845), .C2(n1809), .A(n2104), 
        .ZN(n2099) );
  AOI22_X1 U2635 ( .A1(n1811), .A2(\REGISTERS[11][15] ), .B1(n1812), .B2(
        \REGISTERS[10][15] ), .ZN(n2104) );
  OAI221_X1 U2636 ( .B1(n675), .B2(n1813), .C1(n709), .C2(n1814), .A(n2105), 
        .ZN(n2098) );
  AOI22_X1 U2637 ( .A1(n1816), .A2(\REGISTERS[15][15] ), .B1(n1817), .B2(
        \REGISTERS[14][15] ), .ZN(n2105) );
  AOI21_X1 U2638 ( .B1(n2106), .B2(n2107), .A(N352), .ZN(N301) );
  NOR4_X1 U2639 ( .A1(n2108), .A2(n2109), .A3(n2110), .A4(n2111), .ZN(n2107)
         );
  OAI221_X1 U2640 ( .B1(n536), .B2(n1774), .C1(n570), .C2(n1775), .A(n2112), 
        .ZN(n2111) );
  AOI22_X1 U2641 ( .A1(n1777), .A2(\REGISTERS[19][14] ), .B1(n1778), .B2(
        \REGISTERS[18][14] ), .ZN(n2112) );
  OAI221_X1 U2642 ( .B1(n400), .B2(n1779), .C1(n434), .C2(n1780), .A(n2113), 
        .ZN(n2110) );
  AOI22_X1 U2643 ( .A1(n1782), .A2(\REGISTERS[23][14] ), .B1(n1783), .B2(
        \REGISTERS[22][14] ), .ZN(n2113) );
  OAI221_X1 U2644 ( .B1(n260), .B2(n1784), .C1(n295), .C2(n1785), .A(n2114), 
        .ZN(n2109) );
  AOI22_X1 U2645 ( .A1(n1787), .A2(\REGISTERS[27][14] ), .B1(n1788), .B2(
        \REGISTERS[26][14] ), .ZN(n2114) );
  OAI221_X1 U2646 ( .B1(n32), .B2(n1789), .C1(n85), .C2(n1790), .A(n2115), 
        .ZN(n2108) );
  AOI22_X1 U2647 ( .A1(n1792), .A2(\REGISTERS[29][14] ), .B1(n1793), .B2(
        \REGISTERS[28][14] ), .ZN(n2115) );
  NOR4_X1 U2648 ( .A1(n2116), .A2(n2117), .A3(n2118), .A4(n2119), .ZN(n2106)
         );
  OAI221_X1 U2649 ( .B1(n1087), .B2(n1798), .C1(n1121), .C2(n1799), .A(n2120), 
        .ZN(n2119) );
  AOI22_X1 U2650 ( .A1(n1801), .A2(\REGISTERS[3][14] ), .B1(n1802), .B2(
        \REGISTERS[2][14] ), .ZN(n2120) );
  OAI221_X1 U2651 ( .B1(n951), .B2(n1803), .C1(n985), .C2(n1804), .A(n2121), 
        .ZN(n2118) );
  AOI22_X1 U2652 ( .A1(n1806), .A2(\REGISTERS[7][14] ), .B1(n1807), .B2(
        \REGISTERS[6][14] ), .ZN(n2121) );
  OAI221_X1 U2653 ( .B1(n810), .B2(n1808), .C1(n844), .C2(n1809), .A(n2122), 
        .ZN(n2117) );
  AOI22_X1 U2654 ( .A1(n1811), .A2(\REGISTERS[11][14] ), .B1(n1812), .B2(
        \REGISTERS[10][14] ), .ZN(n2122) );
  OAI221_X1 U2655 ( .B1(n674), .B2(n1813), .C1(n708), .C2(n1814), .A(n2123), 
        .ZN(n2116) );
  AOI22_X1 U2656 ( .A1(n1816), .A2(\REGISTERS[15][14] ), .B1(n1817), .B2(
        \REGISTERS[14][14] ), .ZN(n2123) );
  AOI21_X1 U2657 ( .B1(n2124), .B2(n2125), .A(N352), .ZN(N300) );
  NOR4_X1 U2658 ( .A1(n2126), .A2(n2127), .A3(n2128), .A4(n2129), .ZN(n2125)
         );
  OAI221_X1 U2659 ( .B1(n535), .B2(n1774), .C1(n569), .C2(n1775), .A(n2130), 
        .ZN(n2129) );
  AOI22_X1 U2660 ( .A1(n1777), .A2(\REGISTERS[19][13] ), .B1(n1778), .B2(
        \REGISTERS[18][13] ), .ZN(n2130) );
  OAI221_X1 U2661 ( .B1(n399), .B2(n1779), .C1(n433), .C2(n1780), .A(n2131), 
        .ZN(n2128) );
  AOI22_X1 U2662 ( .A1(n1782), .A2(\REGISTERS[23][13] ), .B1(n1783), .B2(
        \REGISTERS[22][13] ), .ZN(n2131) );
  OAI221_X1 U2663 ( .B1(n259), .B2(n1784), .C1(n294), .C2(n1785), .A(n2132), 
        .ZN(n2127) );
  AOI22_X1 U2664 ( .A1(n1787), .A2(\REGISTERS[27][13] ), .B1(n1788), .B2(
        \REGISTERS[26][13] ), .ZN(n2132) );
  OAI221_X1 U2665 ( .B1(n30), .B2(n1789), .C1(n84), .C2(n1790), .A(n2133), 
        .ZN(n2126) );
  AOI22_X1 U2666 ( .A1(n1792), .A2(\REGISTERS[29][13] ), .B1(n1793), .B2(
        \REGISTERS[28][13] ), .ZN(n2133) );
  NOR4_X1 U2667 ( .A1(n2134), .A2(n2135), .A3(n2136), .A4(n2137), .ZN(n2124)
         );
  OAI221_X1 U2668 ( .B1(n1086), .B2(n1798), .C1(n1120), .C2(n1799), .A(n2138), 
        .ZN(n2137) );
  AOI22_X1 U2669 ( .A1(n1801), .A2(\REGISTERS[3][13] ), .B1(n1802), .B2(
        \REGISTERS[2][13] ), .ZN(n2138) );
  OAI221_X1 U2670 ( .B1(n950), .B2(n1803), .C1(n984), .C2(n1804), .A(n2139), 
        .ZN(n2136) );
  AOI22_X1 U2671 ( .A1(n1806), .A2(\REGISTERS[7][13] ), .B1(n1807), .B2(
        \REGISTERS[6][13] ), .ZN(n2139) );
  OAI221_X1 U2672 ( .B1(n809), .B2(n1808), .C1(n843), .C2(n1809), .A(n2140), 
        .ZN(n2135) );
  AOI22_X1 U2673 ( .A1(n1811), .A2(\REGISTERS[11][13] ), .B1(n1812), .B2(
        \REGISTERS[10][13] ), .ZN(n2140) );
  OAI221_X1 U2674 ( .B1(n673), .B2(n1813), .C1(n707), .C2(n1814), .A(n2141), 
        .ZN(n2134) );
  AOI22_X1 U2675 ( .A1(n1816), .A2(\REGISTERS[15][13] ), .B1(n1817), .B2(
        \REGISTERS[14][13] ), .ZN(n2141) );
  AOI21_X1 U2676 ( .B1(n2142), .B2(n2143), .A(N352), .ZN(N299) );
  NOR4_X1 U2677 ( .A1(n2144), .A2(n2145), .A3(n2146), .A4(n2147), .ZN(n2143)
         );
  OAI221_X1 U2678 ( .B1(n534), .B2(n1774), .C1(n568), .C2(n1775), .A(n2148), 
        .ZN(n2147) );
  AOI22_X1 U2679 ( .A1(n1777), .A2(\REGISTERS[19][12] ), .B1(n1778), .B2(
        \REGISTERS[18][12] ), .ZN(n2148) );
  OAI221_X1 U2680 ( .B1(n398), .B2(n1779), .C1(n432), .C2(n1780), .A(n2149), 
        .ZN(n2146) );
  AOI22_X1 U2681 ( .A1(n1782), .A2(\REGISTERS[23][12] ), .B1(n1783), .B2(
        \REGISTERS[22][12] ), .ZN(n2149) );
  OAI221_X1 U2682 ( .B1(n258), .B2(n1784), .C1(n293), .C2(n1785), .A(n2150), 
        .ZN(n2145) );
  AOI22_X1 U2683 ( .A1(n1787), .A2(\REGISTERS[27][12] ), .B1(n1788), .B2(
        \REGISTERS[26][12] ), .ZN(n2150) );
  OAI221_X1 U2684 ( .B1(n28), .B2(n1789), .C1(n83), .C2(n1790), .A(n2151), 
        .ZN(n2144) );
  AOI22_X1 U2685 ( .A1(n1792), .A2(\REGISTERS[29][12] ), .B1(n1793), .B2(
        \REGISTERS[28][12] ), .ZN(n2151) );
  NOR4_X1 U2686 ( .A1(n2152), .A2(n2153), .A3(n2154), .A4(n2155), .ZN(n2142)
         );
  OAI221_X1 U2687 ( .B1(n1085), .B2(n1798), .C1(n1119), .C2(n1799), .A(n2156), 
        .ZN(n2155) );
  AOI22_X1 U2688 ( .A1(n1801), .A2(\REGISTERS[3][12] ), .B1(n1802), .B2(
        \REGISTERS[2][12] ), .ZN(n2156) );
  OAI221_X1 U2689 ( .B1(n949), .B2(n1803), .C1(n983), .C2(n1804), .A(n2157), 
        .ZN(n2154) );
  AOI22_X1 U2690 ( .A1(n1806), .A2(\REGISTERS[7][12] ), .B1(n1807), .B2(
        \REGISTERS[6][12] ), .ZN(n2157) );
  OAI221_X1 U2691 ( .B1(n808), .B2(n1808), .C1(n842), .C2(n1809), .A(n2158), 
        .ZN(n2153) );
  AOI22_X1 U2692 ( .A1(n1811), .A2(\REGISTERS[11][12] ), .B1(n1812), .B2(
        \REGISTERS[10][12] ), .ZN(n2158) );
  OAI221_X1 U2693 ( .B1(n672), .B2(n1813), .C1(n706), .C2(n1814), .A(n2159), 
        .ZN(n2152) );
  AOI22_X1 U2694 ( .A1(n1816), .A2(\REGISTERS[15][12] ), .B1(n1817), .B2(
        \REGISTERS[14][12] ), .ZN(n2159) );
  AOI21_X1 U2695 ( .B1(n2160), .B2(n2161), .A(N352), .ZN(N298) );
  NOR4_X1 U2696 ( .A1(n2162), .A2(n2163), .A3(n2164), .A4(n2165), .ZN(n2161)
         );
  OAI221_X1 U2697 ( .B1(n533), .B2(n1774), .C1(n567), .C2(n1775), .A(n2166), 
        .ZN(n2165) );
  AOI22_X1 U2698 ( .A1(n1777), .A2(\REGISTERS[19][11] ), .B1(n1778), .B2(
        \REGISTERS[18][11] ), .ZN(n2166) );
  OAI221_X1 U2699 ( .B1(n397), .B2(n1779), .C1(n431), .C2(n1780), .A(n2167), 
        .ZN(n2164) );
  AOI22_X1 U2700 ( .A1(n1782), .A2(\REGISTERS[23][11] ), .B1(n1783), .B2(
        \REGISTERS[22][11] ), .ZN(n2167) );
  OAI221_X1 U2701 ( .B1(n257), .B2(n1784), .C1(n292), .C2(n1785), .A(n2168), 
        .ZN(n2163) );
  AOI22_X1 U2702 ( .A1(n1787), .A2(\REGISTERS[27][11] ), .B1(n1788), .B2(
        \REGISTERS[26][11] ), .ZN(n2168) );
  OAI221_X1 U2703 ( .B1(n26), .B2(n1789), .C1(n82), .C2(n1790), .A(n2169), 
        .ZN(n2162) );
  AOI22_X1 U2704 ( .A1(n1792), .A2(\REGISTERS[29][11] ), .B1(n1793), .B2(
        \REGISTERS[28][11] ), .ZN(n2169) );
  NOR4_X1 U2705 ( .A1(n2170), .A2(n2171), .A3(n2172), .A4(n2173), .ZN(n2160)
         );
  OAI221_X1 U2706 ( .B1(n1084), .B2(n1798), .C1(n1118), .C2(n1799), .A(n2174), 
        .ZN(n2173) );
  AOI22_X1 U2707 ( .A1(n1801), .A2(\REGISTERS[3][11] ), .B1(n1802), .B2(
        \REGISTERS[2][11] ), .ZN(n2174) );
  OAI221_X1 U2708 ( .B1(n948), .B2(n1803), .C1(n982), .C2(n1804), .A(n2175), 
        .ZN(n2172) );
  AOI22_X1 U2709 ( .A1(n1806), .A2(\REGISTERS[7][11] ), .B1(n1807), .B2(
        \REGISTERS[6][11] ), .ZN(n2175) );
  OAI221_X1 U2710 ( .B1(n807), .B2(n1808), .C1(n841), .C2(n1809), .A(n2176), 
        .ZN(n2171) );
  AOI22_X1 U2711 ( .A1(n1811), .A2(\REGISTERS[11][11] ), .B1(n1812), .B2(
        \REGISTERS[10][11] ), .ZN(n2176) );
  OAI221_X1 U2712 ( .B1(n671), .B2(n1813), .C1(n705), .C2(n1814), .A(n2177), 
        .ZN(n2170) );
  AOI22_X1 U2713 ( .A1(n1816), .A2(\REGISTERS[15][11] ), .B1(n1817), .B2(
        \REGISTERS[14][11] ), .ZN(n2177) );
  AOI21_X1 U2714 ( .B1(n2178), .B2(n2179), .A(N352), .ZN(N297) );
  NOR4_X1 U2715 ( .A1(n2180), .A2(n2181), .A3(n2182), .A4(n2183), .ZN(n2179)
         );
  OAI221_X1 U2716 ( .B1(n532), .B2(n1774), .C1(n566), .C2(n1775), .A(n2184), 
        .ZN(n2183) );
  AOI22_X1 U2717 ( .A1(n1777), .A2(\REGISTERS[19][10] ), .B1(n1778), .B2(
        \REGISTERS[18][10] ), .ZN(n2184) );
  OAI221_X1 U2718 ( .B1(n396), .B2(n1779), .C1(n430), .C2(n1780), .A(n2185), 
        .ZN(n2182) );
  AOI22_X1 U2719 ( .A1(n1782), .A2(\REGISTERS[23][10] ), .B1(n1783), .B2(
        \REGISTERS[22][10] ), .ZN(n2185) );
  OAI221_X1 U2720 ( .B1(n256), .B2(n1784), .C1(n291), .C2(n1785), .A(n2186), 
        .ZN(n2181) );
  AOI22_X1 U2721 ( .A1(n1787), .A2(\REGISTERS[27][10] ), .B1(n1788), .B2(
        \REGISTERS[26][10] ), .ZN(n2186) );
  OAI221_X1 U2722 ( .B1(n24), .B2(n1789), .C1(n81), .C2(n1790), .A(n2187), 
        .ZN(n2180) );
  AOI22_X1 U2723 ( .A1(n1792), .A2(\REGISTERS[29][10] ), .B1(n1793), .B2(
        \REGISTERS[28][10] ), .ZN(n2187) );
  NOR4_X1 U2724 ( .A1(n2188), .A2(n2189), .A3(n2190), .A4(n2191), .ZN(n2178)
         );
  OAI221_X1 U2725 ( .B1(n1083), .B2(n1798), .C1(n1117), .C2(n1799), .A(n2192), 
        .ZN(n2191) );
  AOI22_X1 U2726 ( .A1(n1801), .A2(\REGISTERS[3][10] ), .B1(n1802), .B2(
        \REGISTERS[2][10] ), .ZN(n2192) );
  OAI221_X1 U2727 ( .B1(n947), .B2(n1803), .C1(n981), .C2(n1804), .A(n2193), 
        .ZN(n2190) );
  AOI22_X1 U2728 ( .A1(n1806), .A2(\REGISTERS[7][10] ), .B1(n1807), .B2(
        \REGISTERS[6][10] ), .ZN(n2193) );
  OAI221_X1 U2729 ( .B1(n806), .B2(n1808), .C1(n840), .C2(n1809), .A(n2194), 
        .ZN(n2189) );
  AOI22_X1 U2730 ( .A1(n1811), .A2(\REGISTERS[11][10] ), .B1(n1812), .B2(
        \REGISTERS[10][10] ), .ZN(n2194) );
  OAI221_X1 U2731 ( .B1(n670), .B2(n1813), .C1(n704), .C2(n1814), .A(n2195), 
        .ZN(n2188) );
  AOI22_X1 U2732 ( .A1(n1816), .A2(\REGISTERS[15][10] ), .B1(n1817), .B2(
        \REGISTERS[14][10] ), .ZN(n2195) );
  AOI21_X1 U2733 ( .B1(n2196), .B2(n2197), .A(N352), .ZN(N296) );
  NOR4_X1 U2734 ( .A1(n2198), .A2(n2199), .A3(n2200), .A4(n2201), .ZN(n2197)
         );
  OAI221_X1 U2735 ( .B1(n531), .B2(n1774), .C1(n565), .C2(n1775), .A(n2202), 
        .ZN(n2201) );
  AOI22_X1 U2736 ( .A1(n1777), .A2(\REGISTERS[19][9] ), .B1(n1778), .B2(
        \REGISTERS[18][9] ), .ZN(n2202) );
  OAI221_X1 U2737 ( .B1(n395), .B2(n1779), .C1(n429), .C2(n1780), .A(n2203), 
        .ZN(n2200) );
  AOI22_X1 U2738 ( .A1(n1782), .A2(\REGISTERS[23][9] ), .B1(n1783), .B2(
        \REGISTERS[22][9] ), .ZN(n2203) );
  OAI221_X1 U2739 ( .B1(n255), .B2(n1784), .C1(n290), .C2(n1785), .A(n2204), 
        .ZN(n2199) );
  AOI22_X1 U2740 ( .A1(n1787), .A2(\REGISTERS[27][9] ), .B1(n1788), .B2(
        \REGISTERS[26][9] ), .ZN(n2204) );
  OAI221_X1 U2741 ( .B1(n22), .B2(n1789), .C1(n80), .C2(n1790), .A(n2205), 
        .ZN(n2198) );
  AOI22_X1 U2742 ( .A1(n1792), .A2(\REGISTERS[29][9] ), .B1(n1793), .B2(
        \REGISTERS[28][9] ), .ZN(n2205) );
  NOR4_X1 U2743 ( .A1(n2206), .A2(n2207), .A3(n2208), .A4(n2209), .ZN(n2196)
         );
  OAI221_X1 U2744 ( .B1(n1082), .B2(n1798), .C1(n1116), .C2(n1799), .A(n2210), 
        .ZN(n2209) );
  AOI22_X1 U2745 ( .A1(n1801), .A2(\REGISTERS[3][9] ), .B1(n1802), .B2(
        \REGISTERS[2][9] ), .ZN(n2210) );
  OAI221_X1 U2746 ( .B1(n946), .B2(n1803), .C1(n980), .C2(n1804), .A(n2211), 
        .ZN(n2208) );
  AOI22_X1 U2747 ( .A1(n1806), .A2(\REGISTERS[7][9] ), .B1(n1807), .B2(
        \REGISTERS[6][9] ), .ZN(n2211) );
  OAI221_X1 U2748 ( .B1(n805), .B2(n1808), .C1(n839), .C2(n1809), .A(n2212), 
        .ZN(n2207) );
  AOI22_X1 U2749 ( .A1(n1811), .A2(\REGISTERS[11][9] ), .B1(n1812), .B2(
        \REGISTERS[10][9] ), .ZN(n2212) );
  OAI221_X1 U2750 ( .B1(n669), .B2(n1813), .C1(n703), .C2(n1814), .A(n2213), 
        .ZN(n2206) );
  AOI22_X1 U2751 ( .A1(n1816), .A2(\REGISTERS[15][9] ), .B1(n1817), .B2(
        \REGISTERS[14][9] ), .ZN(n2213) );
  AOI21_X1 U2752 ( .B1(n2214), .B2(n2215), .A(N352), .ZN(N295) );
  NOR4_X1 U2753 ( .A1(n2216), .A2(n2217), .A3(n2218), .A4(n2219), .ZN(n2215)
         );
  OAI221_X1 U2754 ( .B1(n530), .B2(n1774), .C1(n564), .C2(n1775), .A(n2220), 
        .ZN(n2219) );
  AOI22_X1 U2755 ( .A1(n1777), .A2(\REGISTERS[19][8] ), .B1(n1778), .B2(
        \REGISTERS[18][8] ), .ZN(n2220) );
  OAI221_X1 U2756 ( .B1(n394), .B2(n1779), .C1(n428), .C2(n1780), .A(n2221), 
        .ZN(n2218) );
  AOI22_X1 U2757 ( .A1(n1782), .A2(\REGISTERS[23][8] ), .B1(n1783), .B2(
        \REGISTERS[22][8] ), .ZN(n2221) );
  OAI221_X1 U2758 ( .B1(n254), .B2(n1784), .C1(n289), .C2(n1785), .A(n2222), 
        .ZN(n2217) );
  AOI22_X1 U2759 ( .A1(n1787), .A2(\REGISTERS[27][8] ), .B1(n1788), .B2(
        \REGISTERS[26][8] ), .ZN(n2222) );
  OAI221_X1 U2760 ( .B1(n20), .B2(n1789), .C1(n79), .C2(n1790), .A(n2223), 
        .ZN(n2216) );
  AOI22_X1 U2761 ( .A1(n1792), .A2(\REGISTERS[29][8] ), .B1(n1793), .B2(
        \REGISTERS[28][8] ), .ZN(n2223) );
  NOR4_X1 U2762 ( .A1(n2224), .A2(n2225), .A3(n2226), .A4(n2227), .ZN(n2214)
         );
  OAI221_X1 U2763 ( .B1(n1081), .B2(n1798), .C1(n1115), .C2(n1799), .A(n2228), 
        .ZN(n2227) );
  AOI22_X1 U2764 ( .A1(n1801), .A2(\REGISTERS[3][8] ), .B1(n1802), .B2(
        \REGISTERS[2][8] ), .ZN(n2228) );
  OAI221_X1 U2765 ( .B1(n945), .B2(n1803), .C1(n979), .C2(n1804), .A(n2229), 
        .ZN(n2226) );
  AOI22_X1 U2766 ( .A1(n1806), .A2(\REGISTERS[7][8] ), .B1(n1807), .B2(
        \REGISTERS[6][8] ), .ZN(n2229) );
  OAI221_X1 U2767 ( .B1(n804), .B2(n1808), .C1(n838), .C2(n1809), .A(n2230), 
        .ZN(n2225) );
  AOI22_X1 U2768 ( .A1(n1811), .A2(\REGISTERS[11][8] ), .B1(n1812), .B2(
        \REGISTERS[10][8] ), .ZN(n2230) );
  OAI221_X1 U2769 ( .B1(n668), .B2(n1813), .C1(n702), .C2(n1814), .A(n2231), 
        .ZN(n2224) );
  AOI22_X1 U2770 ( .A1(n1816), .A2(\REGISTERS[15][8] ), .B1(n1817), .B2(
        \REGISTERS[14][8] ), .ZN(n2231) );
  AOI21_X1 U2771 ( .B1(n2232), .B2(n2233), .A(N352), .ZN(N294) );
  NOR4_X1 U2772 ( .A1(n2234), .A2(n2235), .A3(n2236), .A4(n2237), .ZN(n2233)
         );
  OAI221_X1 U2773 ( .B1(n529), .B2(n1774), .C1(n563), .C2(n1775), .A(n2238), 
        .ZN(n2237) );
  AOI22_X1 U2774 ( .A1(n1777), .A2(\REGISTERS[19][7] ), .B1(n1778), .B2(
        \REGISTERS[18][7] ), .ZN(n2238) );
  OAI221_X1 U2775 ( .B1(n393), .B2(n1779), .C1(n427), .C2(n1780), .A(n2239), 
        .ZN(n2236) );
  AOI22_X1 U2776 ( .A1(n1782), .A2(\REGISTERS[23][7] ), .B1(n1783), .B2(
        \REGISTERS[22][7] ), .ZN(n2239) );
  OAI221_X1 U2777 ( .B1(n253), .B2(n1784), .C1(n288), .C2(n1785), .A(n2240), 
        .ZN(n2235) );
  AOI22_X1 U2778 ( .A1(n1787), .A2(\REGISTERS[27][7] ), .B1(n1788), .B2(
        \REGISTERS[26][7] ), .ZN(n2240) );
  OAI221_X1 U2779 ( .B1(n18), .B2(n1789), .C1(n78), .C2(n1790), .A(n2241), 
        .ZN(n2234) );
  AOI22_X1 U2780 ( .A1(n1792), .A2(\REGISTERS[29][7] ), .B1(n1793), .B2(
        \REGISTERS[28][7] ), .ZN(n2241) );
  NOR4_X1 U2781 ( .A1(n2242), .A2(n2243), .A3(n2244), .A4(n2245), .ZN(n2232)
         );
  OAI221_X1 U2782 ( .B1(n1080), .B2(n1798), .C1(n1114), .C2(n1799), .A(n2246), 
        .ZN(n2245) );
  AOI22_X1 U2783 ( .A1(n1801), .A2(\REGISTERS[3][7] ), .B1(n1802), .B2(
        \REGISTERS[2][7] ), .ZN(n2246) );
  OAI221_X1 U2784 ( .B1(n944), .B2(n1803), .C1(n978), .C2(n1804), .A(n2247), 
        .ZN(n2244) );
  AOI22_X1 U2785 ( .A1(n1806), .A2(\REGISTERS[7][7] ), .B1(n1807), .B2(
        \REGISTERS[6][7] ), .ZN(n2247) );
  OAI221_X1 U2786 ( .B1(n803), .B2(n1808), .C1(n837), .C2(n1809), .A(n2248), 
        .ZN(n2243) );
  AOI22_X1 U2787 ( .A1(n1811), .A2(\REGISTERS[11][7] ), .B1(n1812), .B2(
        \REGISTERS[10][7] ), .ZN(n2248) );
  OAI221_X1 U2788 ( .B1(n667), .B2(n1813), .C1(n701), .C2(n1814), .A(n2249), 
        .ZN(n2242) );
  AOI22_X1 U2789 ( .A1(n1816), .A2(\REGISTERS[15][7] ), .B1(n1817), .B2(
        \REGISTERS[14][7] ), .ZN(n2249) );
  AOI21_X1 U2790 ( .B1(n2250), .B2(n2251), .A(N352), .ZN(N293) );
  NOR4_X1 U2791 ( .A1(n2252), .A2(n2253), .A3(n2254), .A4(n2255), .ZN(n2251)
         );
  OAI221_X1 U2792 ( .B1(n528), .B2(n1774), .C1(n562), .C2(n1775), .A(n2256), 
        .ZN(n2255) );
  AOI22_X1 U2793 ( .A1(n1777), .A2(\REGISTERS[19][6] ), .B1(n1778), .B2(
        \REGISTERS[18][6] ), .ZN(n2256) );
  OAI221_X1 U2794 ( .B1(n392), .B2(n1779), .C1(n426), .C2(n1780), .A(n2257), 
        .ZN(n2254) );
  AOI22_X1 U2795 ( .A1(n1782), .A2(\REGISTERS[23][6] ), .B1(n1783), .B2(
        \REGISTERS[22][6] ), .ZN(n2257) );
  OAI221_X1 U2796 ( .B1(n252), .B2(n1784), .C1(n287), .C2(n1785), .A(n2258), 
        .ZN(n2253) );
  AOI22_X1 U2797 ( .A1(n1787), .A2(\REGISTERS[27][6] ), .B1(n1788), .B2(
        \REGISTERS[26][6] ), .ZN(n2258) );
  OAI221_X1 U2798 ( .B1(n16), .B2(n1789), .C1(n77), .C2(n1790), .A(n2259), 
        .ZN(n2252) );
  AOI22_X1 U2799 ( .A1(n1792), .A2(\REGISTERS[29][6] ), .B1(n1793), .B2(
        \REGISTERS[28][6] ), .ZN(n2259) );
  NOR4_X1 U2800 ( .A1(n2260), .A2(n2261), .A3(n2262), .A4(n2263), .ZN(n2250)
         );
  OAI221_X1 U2801 ( .B1(n1079), .B2(n1798), .C1(n1113), .C2(n1799), .A(n2264), 
        .ZN(n2263) );
  AOI22_X1 U2802 ( .A1(n1801), .A2(\REGISTERS[3][6] ), .B1(n1802), .B2(
        \REGISTERS[2][6] ), .ZN(n2264) );
  OAI221_X1 U2803 ( .B1(n943), .B2(n1803), .C1(n977), .C2(n1804), .A(n2265), 
        .ZN(n2262) );
  AOI22_X1 U2804 ( .A1(n1806), .A2(\REGISTERS[7][6] ), .B1(n1807), .B2(
        \REGISTERS[6][6] ), .ZN(n2265) );
  OAI221_X1 U2805 ( .B1(n802), .B2(n1808), .C1(n836), .C2(n1809), .A(n2266), 
        .ZN(n2261) );
  AOI22_X1 U2806 ( .A1(n1811), .A2(\REGISTERS[11][6] ), .B1(n1812), .B2(
        \REGISTERS[10][6] ), .ZN(n2266) );
  OAI221_X1 U2807 ( .B1(n666), .B2(n1813), .C1(n700), .C2(n1814), .A(n2267), 
        .ZN(n2260) );
  AOI22_X1 U2808 ( .A1(n1816), .A2(\REGISTERS[15][6] ), .B1(n1817), .B2(
        \REGISTERS[14][6] ), .ZN(n2267) );
  AOI21_X1 U2809 ( .B1(n2268), .B2(n2269), .A(N352), .ZN(N292) );
  NOR4_X1 U2810 ( .A1(n2270), .A2(n2271), .A3(n2272), .A4(n2273), .ZN(n2269)
         );
  OAI221_X1 U2811 ( .B1(n527), .B2(n1774), .C1(n561), .C2(n1775), .A(n2274), 
        .ZN(n2273) );
  AOI22_X1 U2812 ( .A1(n1777), .A2(\REGISTERS[19][5] ), .B1(n1778), .B2(
        \REGISTERS[18][5] ), .ZN(n2274) );
  OAI221_X1 U2813 ( .B1(n391), .B2(n1779), .C1(n425), .C2(n1780), .A(n2275), 
        .ZN(n2272) );
  AOI22_X1 U2814 ( .A1(n1782), .A2(\REGISTERS[23][5] ), .B1(n1783), .B2(
        \REGISTERS[22][5] ), .ZN(n2275) );
  OAI221_X1 U2815 ( .B1(n251), .B2(n1784), .C1(n286), .C2(n1785), .A(n2276), 
        .ZN(n2271) );
  AOI22_X1 U2816 ( .A1(n1787), .A2(\REGISTERS[27][5] ), .B1(n1788), .B2(
        \REGISTERS[26][5] ), .ZN(n2276) );
  OAI221_X1 U2817 ( .B1(n14), .B2(n1789), .C1(n76), .C2(n1790), .A(n2277), 
        .ZN(n2270) );
  AOI22_X1 U2818 ( .A1(n1792), .A2(\REGISTERS[29][5] ), .B1(n1793), .B2(
        \REGISTERS[28][5] ), .ZN(n2277) );
  NOR4_X1 U2819 ( .A1(n2278), .A2(n2279), .A3(n2280), .A4(n2281), .ZN(n2268)
         );
  OAI221_X1 U2820 ( .B1(n1078), .B2(n1798), .C1(n1112), .C2(n1799), .A(n2282), 
        .ZN(n2281) );
  AOI22_X1 U2821 ( .A1(n1801), .A2(\REGISTERS[3][5] ), .B1(n1802), .B2(
        \REGISTERS[2][5] ), .ZN(n2282) );
  OAI221_X1 U2822 ( .B1(n942), .B2(n1803), .C1(n976), .C2(n1804), .A(n2283), 
        .ZN(n2280) );
  AOI22_X1 U2823 ( .A1(n1806), .A2(\REGISTERS[7][5] ), .B1(n1807), .B2(
        \REGISTERS[6][5] ), .ZN(n2283) );
  OAI221_X1 U2824 ( .B1(n801), .B2(n1808), .C1(n835), .C2(n1809), .A(n2284), 
        .ZN(n2279) );
  AOI22_X1 U2825 ( .A1(n1811), .A2(\REGISTERS[11][5] ), .B1(n1812), .B2(
        \REGISTERS[10][5] ), .ZN(n2284) );
  OAI221_X1 U2826 ( .B1(n665), .B2(n1813), .C1(n699), .C2(n1814), .A(n2285), 
        .ZN(n2278) );
  AOI22_X1 U2827 ( .A1(n1816), .A2(\REGISTERS[15][5] ), .B1(n1817), .B2(
        \REGISTERS[14][5] ), .ZN(n2285) );
  AOI21_X1 U2828 ( .B1(n2286), .B2(n2287), .A(N352), .ZN(N291) );
  NOR4_X1 U2829 ( .A1(n2288), .A2(n2289), .A3(n2290), .A4(n2291), .ZN(n2287)
         );
  OAI221_X1 U2830 ( .B1(n526), .B2(n1774), .C1(n560), .C2(n1775), .A(n2292), 
        .ZN(n2291) );
  AOI22_X1 U2831 ( .A1(n1777), .A2(\REGISTERS[19][4] ), .B1(n1778), .B2(
        \REGISTERS[18][4] ), .ZN(n2292) );
  OAI221_X1 U2832 ( .B1(n390), .B2(n1779), .C1(n424), .C2(n1780), .A(n2293), 
        .ZN(n2290) );
  AOI22_X1 U2833 ( .A1(n1782), .A2(\REGISTERS[23][4] ), .B1(n1783), .B2(
        \REGISTERS[22][4] ), .ZN(n2293) );
  OAI221_X1 U2834 ( .B1(n250), .B2(n1784), .C1(n285), .C2(n1785), .A(n2294), 
        .ZN(n2289) );
  AOI22_X1 U2835 ( .A1(n1787), .A2(\REGISTERS[27][4] ), .B1(n1788), .B2(
        \REGISTERS[26][4] ), .ZN(n2294) );
  OAI221_X1 U2836 ( .B1(n12), .B2(n1789), .C1(n75), .C2(n1790), .A(n2295), 
        .ZN(n2288) );
  AOI22_X1 U2837 ( .A1(n1792), .A2(\REGISTERS[29][4] ), .B1(n1793), .B2(
        \REGISTERS[28][4] ), .ZN(n2295) );
  NOR4_X1 U2838 ( .A1(n2296), .A2(n2297), .A3(n2298), .A4(n2299), .ZN(n2286)
         );
  OAI221_X1 U2839 ( .B1(n1077), .B2(n1798), .C1(n1111), .C2(n1799), .A(n2300), 
        .ZN(n2299) );
  AOI22_X1 U2840 ( .A1(n1801), .A2(\REGISTERS[3][4] ), .B1(n1802), .B2(
        \REGISTERS[2][4] ), .ZN(n2300) );
  OAI221_X1 U2841 ( .B1(n941), .B2(n1803), .C1(n975), .C2(n1804), .A(n2301), 
        .ZN(n2298) );
  AOI22_X1 U2842 ( .A1(n1806), .A2(\REGISTERS[7][4] ), .B1(n1807), .B2(
        \REGISTERS[6][4] ), .ZN(n2301) );
  OAI221_X1 U2843 ( .B1(n800), .B2(n1808), .C1(n834), .C2(n1809), .A(n2302), 
        .ZN(n2297) );
  AOI22_X1 U2844 ( .A1(n1811), .A2(\REGISTERS[11][4] ), .B1(n1812), .B2(
        \REGISTERS[10][4] ), .ZN(n2302) );
  OAI221_X1 U2845 ( .B1(n664), .B2(n1813), .C1(n698), .C2(n1814), .A(n2303), 
        .ZN(n2296) );
  AOI22_X1 U2846 ( .A1(n1816), .A2(\REGISTERS[15][4] ), .B1(n1817), .B2(
        \REGISTERS[14][4] ), .ZN(n2303) );
  AOI21_X1 U2847 ( .B1(n2304), .B2(n2305), .A(N352), .ZN(N290) );
  NOR4_X1 U2848 ( .A1(n2306), .A2(n2307), .A3(n2308), .A4(n2309), .ZN(n2305)
         );
  OAI221_X1 U2849 ( .B1(n525), .B2(n1774), .C1(n559), .C2(n1775), .A(n2310), 
        .ZN(n2309) );
  AOI22_X1 U2850 ( .A1(n1777), .A2(\REGISTERS[19][3] ), .B1(n1778), .B2(
        \REGISTERS[18][3] ), .ZN(n2310) );
  OAI221_X1 U2851 ( .B1(n389), .B2(n1779), .C1(n423), .C2(n1780), .A(n2311), 
        .ZN(n2308) );
  AOI22_X1 U2852 ( .A1(n1782), .A2(\REGISTERS[23][3] ), .B1(n1783), .B2(
        \REGISTERS[22][3] ), .ZN(n2311) );
  OAI221_X1 U2853 ( .B1(n249), .B2(n1784), .C1(n284), .C2(n1785), .A(n2312), 
        .ZN(n2307) );
  AOI22_X1 U2854 ( .A1(n1787), .A2(\REGISTERS[27][3] ), .B1(n1788), .B2(
        \REGISTERS[26][3] ), .ZN(n2312) );
  OAI221_X1 U2855 ( .B1(n10), .B2(n1789), .C1(n74), .C2(n1790), .A(n2313), 
        .ZN(n2306) );
  AOI22_X1 U2856 ( .A1(n1792), .A2(\REGISTERS[29][3] ), .B1(n1793), .B2(
        \REGISTERS[28][3] ), .ZN(n2313) );
  NOR4_X1 U2857 ( .A1(n2314), .A2(n2315), .A3(n2316), .A4(n2317), .ZN(n2304)
         );
  OAI221_X1 U2858 ( .B1(n1076), .B2(n1798), .C1(n1110), .C2(n1799), .A(n2318), 
        .ZN(n2317) );
  AOI22_X1 U2859 ( .A1(n1801), .A2(\REGISTERS[3][3] ), .B1(n1802), .B2(
        \REGISTERS[2][3] ), .ZN(n2318) );
  OAI221_X1 U2860 ( .B1(n940), .B2(n1803), .C1(n974), .C2(n1804), .A(n2319), 
        .ZN(n2316) );
  AOI22_X1 U2861 ( .A1(n1806), .A2(\REGISTERS[7][3] ), .B1(n1807), .B2(
        \REGISTERS[6][3] ), .ZN(n2319) );
  OAI221_X1 U2862 ( .B1(n799), .B2(n1808), .C1(n833), .C2(n1809), .A(n2320), 
        .ZN(n2315) );
  AOI22_X1 U2863 ( .A1(n1811), .A2(\REGISTERS[11][3] ), .B1(n1812), .B2(
        \REGISTERS[10][3] ), .ZN(n2320) );
  OAI221_X1 U2864 ( .B1(n663), .B2(n1813), .C1(n697), .C2(n1814), .A(n2321), 
        .ZN(n2314) );
  AOI22_X1 U2865 ( .A1(n1816), .A2(\REGISTERS[15][3] ), .B1(n1817), .B2(
        \REGISTERS[14][3] ), .ZN(n2321) );
  AOI21_X1 U2866 ( .B1(n2322), .B2(n2323), .A(N352), .ZN(N289) );
  NOR4_X1 U2867 ( .A1(n2324), .A2(n2325), .A3(n2326), .A4(n2327), .ZN(n2323)
         );
  OAI221_X1 U2868 ( .B1(n524), .B2(n1774), .C1(n558), .C2(n1775), .A(n2328), 
        .ZN(n2327) );
  AOI22_X1 U2869 ( .A1(n1777), .A2(\REGISTERS[19][2] ), .B1(n1778), .B2(
        \REGISTERS[18][2] ), .ZN(n2328) );
  OAI221_X1 U2870 ( .B1(n388), .B2(n1779), .C1(n422), .C2(n1780), .A(n2329), 
        .ZN(n2326) );
  AOI22_X1 U2871 ( .A1(n1782), .A2(\REGISTERS[23][2] ), .B1(n1783), .B2(
        \REGISTERS[22][2] ), .ZN(n2329) );
  OAI221_X1 U2872 ( .B1(n248), .B2(n1784), .C1(n283), .C2(n1785), .A(n2330), 
        .ZN(n2325) );
  AOI22_X1 U2873 ( .A1(n1787), .A2(\REGISTERS[27][2] ), .B1(n1788), .B2(
        \REGISTERS[26][2] ), .ZN(n2330) );
  OAI221_X1 U2874 ( .B1(n8), .B2(n1789), .C1(n73), .C2(n1790), .A(n2331), .ZN(
        n2324) );
  AOI22_X1 U2875 ( .A1(n1792), .A2(\REGISTERS[29][2] ), .B1(n1793), .B2(
        \REGISTERS[28][2] ), .ZN(n2331) );
  NOR4_X1 U2876 ( .A1(n2332), .A2(n2333), .A3(n2334), .A4(n2335), .ZN(n2322)
         );
  OAI221_X1 U2877 ( .B1(n1075), .B2(n1798), .C1(n1109), .C2(n1799), .A(n2336), 
        .ZN(n2335) );
  AOI22_X1 U2878 ( .A1(n1801), .A2(\REGISTERS[3][2] ), .B1(n1802), .B2(
        \REGISTERS[2][2] ), .ZN(n2336) );
  OAI221_X1 U2879 ( .B1(n939), .B2(n1803), .C1(n973), .C2(n1804), .A(n2337), 
        .ZN(n2334) );
  AOI22_X1 U2880 ( .A1(n1806), .A2(\REGISTERS[7][2] ), .B1(n1807), .B2(
        \REGISTERS[6][2] ), .ZN(n2337) );
  OAI221_X1 U2881 ( .B1(n798), .B2(n1808), .C1(n832), .C2(n1809), .A(n2338), 
        .ZN(n2333) );
  AOI22_X1 U2882 ( .A1(n1811), .A2(\REGISTERS[11][2] ), .B1(n1812), .B2(
        \REGISTERS[10][2] ), .ZN(n2338) );
  OAI221_X1 U2883 ( .B1(n662), .B2(n1813), .C1(n696), .C2(n1814), .A(n2339), 
        .ZN(n2332) );
  AOI22_X1 U2884 ( .A1(n1816), .A2(\REGISTERS[15][2] ), .B1(n1817), .B2(
        \REGISTERS[14][2] ), .ZN(n2339) );
  AOI21_X1 U2885 ( .B1(n2340), .B2(n2341), .A(N352), .ZN(N288) );
  NOR4_X1 U2886 ( .A1(n2342), .A2(n2343), .A3(n2344), .A4(n2345), .ZN(n2341)
         );
  OAI221_X1 U2887 ( .B1(n523), .B2(n1774), .C1(n557), .C2(n1775), .A(n2346), 
        .ZN(n2345) );
  AOI22_X1 U2888 ( .A1(n1777), .A2(\REGISTERS[19][1] ), .B1(n1778), .B2(
        \REGISTERS[18][1] ), .ZN(n2346) );
  OAI221_X1 U2889 ( .B1(n387), .B2(n1779), .C1(n421), .C2(n1780), .A(n2347), 
        .ZN(n2344) );
  AOI22_X1 U2890 ( .A1(n1782), .A2(\REGISTERS[23][1] ), .B1(n1783), .B2(
        \REGISTERS[22][1] ), .ZN(n2347) );
  OAI221_X1 U2891 ( .B1(n247), .B2(n1784), .C1(n282), .C2(n1785), .A(n2348), 
        .ZN(n2343) );
  AOI22_X1 U2892 ( .A1(n1787), .A2(\REGISTERS[27][1] ), .B1(n1788), .B2(
        \REGISTERS[26][1] ), .ZN(n2348) );
  OAI221_X1 U2893 ( .B1(n6), .B2(n1789), .C1(n72), .C2(n1790), .A(n2349), .ZN(
        n2342) );
  AOI22_X1 U2894 ( .A1(n1792), .A2(\REGISTERS[29][1] ), .B1(n1793), .B2(
        \REGISTERS[28][1] ), .ZN(n2349) );
  NOR4_X1 U2895 ( .A1(n2350), .A2(n2351), .A3(n2352), .A4(n2353), .ZN(n2340)
         );
  OAI221_X1 U2896 ( .B1(n1074), .B2(n1798), .C1(n1108), .C2(n1799), .A(n2354), 
        .ZN(n2353) );
  AOI22_X1 U2897 ( .A1(n1801), .A2(\REGISTERS[3][1] ), .B1(n1802), .B2(
        \REGISTERS[2][1] ), .ZN(n2354) );
  OAI221_X1 U2898 ( .B1(n938), .B2(n1803), .C1(n972), .C2(n1804), .A(n2355), 
        .ZN(n2352) );
  AOI22_X1 U2899 ( .A1(n1806), .A2(\REGISTERS[7][1] ), .B1(n1807), .B2(
        \REGISTERS[6][1] ), .ZN(n2355) );
  OAI221_X1 U2900 ( .B1(n797), .B2(n1808), .C1(n831), .C2(n1809), .A(n2356), 
        .ZN(n2351) );
  AOI22_X1 U2901 ( .A1(n1811), .A2(\REGISTERS[11][1] ), .B1(n1812), .B2(
        \REGISTERS[10][1] ), .ZN(n2356) );
  OAI221_X1 U2902 ( .B1(n661), .B2(n1813), .C1(n695), .C2(n1814), .A(n2357), 
        .ZN(n2350) );
  AOI22_X1 U2903 ( .A1(n1816), .A2(\REGISTERS[15][1] ), .B1(n1817), .B2(
        \REGISTERS[14][1] ), .ZN(n2357) );
  AOI21_X1 U2904 ( .B1(n2358), .B2(n2359), .A(N352), .ZN(N287) );
  NOR4_X1 U2906 ( .A1(n2360), .A2(n2361), .A3(n2362), .A4(n2363), .ZN(n2359)
         );
  OAI221_X1 U2907 ( .B1(n522), .B2(n1774), .C1(n556), .C2(n1775), .A(n2364), 
        .ZN(n2363) );
  AOI22_X1 U2908 ( .A1(n1777), .A2(\REGISTERS[19][0] ), .B1(n1778), .B2(
        \REGISTERS[18][0] ), .ZN(n2364) );
  OAI221_X1 U2913 ( .B1(n386), .B2(n1779), .C1(n420), .C2(n1780), .A(n2369), 
        .ZN(n2362) );
  AOI22_X1 U2914 ( .A1(n1782), .A2(\REGISTERS[23][0] ), .B1(n1783), .B2(
        \REGISTERS[22][0] ), .ZN(n2369) );
  AND2_X1 U2918 ( .A1(n2372), .A2(n2373), .ZN(n2365) );
  AND2_X1 U2920 ( .A1(n2372), .A2(ADD_RD1[0]), .ZN(n2367) );
  AND2_X1 U2921 ( .A1(ADD_RD1[4]), .A2(n2374), .ZN(n2372) );
  OAI221_X1 U2922 ( .B1(n246), .B2(n1784), .C1(n281), .C2(n1785), .A(n2375), 
        .ZN(n2361) );
  AOI22_X1 U2923 ( .A1(n1787), .A2(\REGISTERS[27][0] ), .B1(n1788), .B2(
        \REGISTERS[26][0] ), .ZN(n2375) );
  OAI221_X1 U2928 ( .B1(n4), .B2(n1789), .C1(n71), .C2(n1790), .A(n2378), .ZN(
        n2360) );
  AOI22_X1 U2929 ( .A1(n1792), .A2(\REGISTERS[29][0] ), .B1(n1793), .B2(
        \REGISTERS[28][0] ), .ZN(n2378) );
  AND2_X1 U2933 ( .A1(n2379), .A2(n2373), .ZN(n2376) );
  AND2_X1 U2935 ( .A1(ADD_RD1[0]), .A2(n2379), .ZN(n2377) );
  AND2_X1 U2936 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n2379) );
  NOR4_X1 U2937 ( .A1(n2380), .A2(n2381), .A3(n2382), .A4(n2383), .ZN(n2358)
         );
  OAI221_X1 U2938 ( .B1(n1073), .B2(n1798), .C1(n1107), .C2(n1799), .A(n2384), 
        .ZN(n2383) );
  AOI22_X1 U2939 ( .A1(n1801), .A2(\REGISTERS[3][0] ), .B1(n1802), .B2(
        \REGISTERS[2][0] ), .ZN(n2384) );
  OAI221_X1 U2944 ( .B1(n937), .B2(n1803), .C1(n971), .C2(n1804), .A(n2387), 
        .ZN(n2382) );
  AOI22_X1 U2945 ( .A1(n1806), .A2(\REGISTERS[7][0] ), .B1(n1807), .B2(
        \REGISTERS[6][0] ), .ZN(n2387) );
  AND2_X1 U2949 ( .A1(n2388), .A2(n2373), .ZN(n2385) );
  AND2_X1 U2951 ( .A1(n2388), .A2(ADD_RD1[0]), .ZN(n2386) );
  NOR2_X1 U2952 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .ZN(n2388) );
  OAI221_X1 U2953 ( .B1(n796), .B2(n1808), .C1(n830), .C2(n1809), .A(n2389), 
        .ZN(n2381) );
  AOI22_X1 U2954 ( .A1(n1811), .A2(\REGISTERS[11][0] ), .B1(n1812), .B2(
        \REGISTERS[10][0] ), .ZN(n2389) );
  NOR2_X1 U2957 ( .A1(n2392), .A2(ADD_RD1[2]), .ZN(n2366) );
  OAI221_X1 U2961 ( .B1(n660), .B2(n1813), .C1(n694), .C2(n1814), .A(n2393), 
        .ZN(n2380) );
  AOI22_X1 U2962 ( .A1(n1816), .A2(\REGISTERS[15][0] ), .B1(n1817), .B2(
        \REGISTERS[14][0] ), .ZN(n2393) );
  NOR2_X1 U2965 ( .A1(n2394), .A2(n2392), .ZN(n2370) );
  INV_X1 U2966 ( .A(ADD_RD1[1]), .ZN(n2392) );
  AND2_X1 U2968 ( .A1(n2395), .A2(n2373), .ZN(n2390) );
  INV_X1 U2969 ( .A(ADD_RD1[0]), .ZN(n2373) );
  INV_X1 U2972 ( .A(ADD_RD1[2]), .ZN(n2394) );
  AND2_X1 U2973 ( .A1(n2395), .A2(ADD_RD1[0]), .ZN(n2391) );
  NOR2_X1 U2974 ( .A1(n2374), .A2(ADD_RD1[4]), .ZN(n2395) );
  INV_X1 U2975 ( .A(ADD_RD1[3]), .ZN(n2374) );
  NAND2_X1 U2976 ( .A1(n2396), .A2(RESET), .ZN(N286) );
  NAND2_X1 U2977 ( .A1(RD1), .A2(ENABLE), .ZN(n2396) );
  AND2_X2 U35 ( .A1(n2390), .A2(n2370), .ZN(n1817) );
  AND2_X2 U36 ( .A1(n2390), .A2(n2366), .ZN(n1812) );
  AND2_X2 U69 ( .A1(n2385), .A2(n2370), .ZN(n1807) );
  AND2_X2 U70 ( .A1(n2385), .A2(n2366), .ZN(n1802) );
  AND2_X2 U135 ( .A1(n2371), .A2(n2376), .ZN(n1793) );
  AND2_X2 U136 ( .A1(n2366), .A2(n2376), .ZN(n1788) );
  AND2_X2 U201 ( .A1(n2365), .A2(n2370), .ZN(n1783) );
  AND2_X2 U202 ( .A1(n2365), .A2(n2366), .ZN(n1778) );
  AND2_X2 U267 ( .A1(n1761), .A2(n1741), .ZN(n1188) );
  AND2_X2 U268 ( .A1(n1761), .A2(n1737), .ZN(n1183) );
  AND2_X2 U333 ( .A1(n1756), .A2(n1741), .ZN(n1178) );
  AND2_X2 U334 ( .A1(n1756), .A2(n1737), .ZN(n1173) );
  AND2_X2 U367 ( .A1(n1742), .A2(n1747), .ZN(n1164) );
  AND2_X2 U368 ( .A1(n1737), .A2(n1747), .ZN(n1159) );
  AND2_X2 U401 ( .A1(n1736), .A2(n1741), .ZN(n1154) );
  AND2_X2 U402 ( .A1(n1736), .A2(n1737), .ZN(n1149) );
  NAND2_X2 U468 ( .A1(n2385), .A2(n2368), .ZN(n1799) );
  NAND2_X2 U469 ( .A1(n2376), .A2(n2370), .ZN(n1790) );
  NAND2_X2 U534 ( .A1(n2368), .A2(n2376), .ZN(n1785) );
  NAND2_X2 U535 ( .A1(n2365), .A2(n2371), .ZN(n1780) );
  NOR2_X2 U568 ( .A1(n2394), .A2(ADD_RD1[1]), .ZN(n2371) );
  NAND2_X2 U569 ( .A1(n2365), .A2(n2368), .ZN(n1775) );
  NOR2_X2 U602 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n2368) );
  NAND2_X2 U603 ( .A1(n1761), .A2(n1742), .ZN(n1185) );
  NOR2_X2 U668 ( .A1(n1765), .A2(ADD_RD2[1]), .ZN(n1742) );
  NAND2_X2 U669 ( .A1(n1761), .A2(n1739), .ZN(n1180) );
  NAND2_X2 U734 ( .A1(n1756), .A2(n1742), .ZN(n1175) );
  NAND2_X2 U735 ( .A1(n1756), .A2(n1739), .ZN(n1170) );
  NAND2_X2 U768 ( .A1(n1747), .A2(n1741), .ZN(n1161) );
  NAND2_X2 U769 ( .A1(n1739), .A2(n1747), .ZN(n1156) );
  NOR2_X2 U802 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n1739) );
  NAND2_X2 U803 ( .A1(n1736), .A2(n1742), .ZN(n1151) );
  NAND2_X2 U869 ( .A1(n1736), .A2(n1739), .ZN(n1146) );
  NAND2_X2 U870 ( .A1(n2390), .A2(n2368), .ZN(n1809) );
  NAND2_X2 U935 ( .A1(n2385), .A2(n2371), .ZN(n1804) );
  NAND2_X2 U936 ( .A1(n2390), .A2(n2371), .ZN(n1814) );
  NAND2_X2 U969 ( .A1(n1738), .A2(n1739), .ZN(n1145) );
  NAND2_X2 U970 ( .A1(n1739), .A2(n1748), .ZN(n1155) );
  NAND2_X2 U1003 ( .A1(n1738), .A2(n1742), .ZN(n1150) );
  NAND2_X2 U1004 ( .A1(n1757), .A2(n1739), .ZN(n1169) );
  NAND2_X2 U1069 ( .A1(n1741), .A2(n1748), .ZN(n1160) );
  NAND2_X2 U1070 ( .A1(n1762), .A2(n1739), .ZN(n1179) );
  NAND2_X2 U1135 ( .A1(n1757), .A2(n1742), .ZN(n1174) );
  NAND2_X2 U1136 ( .A1(n2367), .A2(n2368), .ZN(n1774) );
  NAND2_X2 U1169 ( .A1(n1762), .A2(n1742), .ZN(n1184) );
  NAND2_X2 U1170 ( .A1(n2368), .A2(n2377), .ZN(n1784) );
  NAND2_X2 U1203 ( .A1(n2367), .A2(n2371), .ZN(n1779) );
  NAND2_X2 U1204 ( .A1(n2386), .A2(n2368), .ZN(n1798) );
  NAND2_X2 U1270 ( .A1(n2370), .A2(n2377), .ZN(n1789) );
  NAND2_X2 U1271 ( .A1(n2391), .A2(n2368), .ZN(n1808) );
  NAND2_X2 U1337 ( .A1(n2386), .A2(n2371), .ZN(n1803) );
  NAND2_X2 U1338 ( .A1(n2391), .A2(n2371), .ZN(n1813) );
  AND2_X2 U1372 ( .A1(n1738), .A2(n1741), .ZN(n1153) );
  AND2_X2 U1373 ( .A1(n1738), .A2(n1737), .ZN(n1148) );
  AND2_X2 U1407 ( .A1(n1742), .A2(n1748), .ZN(n1163) );
  AND2_X2 U1408 ( .A1(n1737), .A2(n1748), .ZN(n1158) );
  AND2_X2 U1475 ( .A1(n1757), .A2(n1741), .ZN(n1177) );
  AND2_X2 U1476 ( .A1(n1757), .A2(n1737), .ZN(n1172) );
  AND2_X2 U1542 ( .A1(n1762), .A2(n1741), .ZN(n1187) );
  AND2_X2 U1543 ( .A1(n1762), .A2(n1737), .ZN(n1182) );
  AND2_X2 U1578 ( .A1(n2367), .A2(n2370), .ZN(n1782) );
  AND2_X2 U1579 ( .A1(n2367), .A2(n2366), .ZN(n1777) );
  AND2_X2 U1645 ( .A1(n2371), .A2(n2377), .ZN(n1792) );
  AND2_X2 U1646 ( .A1(n2366), .A2(n2377), .ZN(n1787) );
  AND2_X2 U2246 ( .A1(n2386), .A2(n2370), .ZN(n1806) );
  AND2_X2 U2247 ( .A1(n2386), .A2(n2366), .ZN(n1801) );
  AND2_X2 U2248 ( .A1(n2391), .A2(n2370), .ZN(n1816) );
  AND2_X2 U2249 ( .A1(n2391), .A2(n2366), .ZN(n1811) );
  INV_X2 U2252 ( .A(n106), .ZN(n105) );
  NAND2_X2 U2253 ( .A1(n138), .A2(n68), .ZN(n106) );
  INV_X2 U2254 ( .A(n176), .ZN(n175) );
  NAND2_X2 U2256 ( .A1(n208), .A2(n68), .ZN(n176) );
  INV_X2 U2261 ( .A(n141), .ZN(n140) );
  NAND2_X2 U2262 ( .A1(n173), .A2(n68), .ZN(n141) );
  INV_X2 U2263 ( .A(n317), .ZN(n316) );
  NAND2_X2 U2264 ( .A1(n349), .A2(n67), .ZN(n317) );
  INV_X2 U2267 ( .A(n211), .ZN(n210) );
  NAND2_X2 U2268 ( .A1(n243), .A2(n68), .ZN(n211) );
  INV_X2 U2269 ( .A(n454), .ZN(n453) );
  NAND2_X2 U2271 ( .A1(n349), .A2(n208), .ZN(n454) );
  INV_X2 U2277 ( .A(n352), .ZN(n351) );
  NAND2_X2 U2278 ( .A1(n349), .A2(n103), .ZN(n352) );
  INV_X2 U2279 ( .A(n591), .ZN(n590) );
  NAND2_X2 U2280 ( .A1(n623), .A2(n67), .ZN(n591) );
  INV_X2 U2283 ( .A(n488), .ZN(n487) );
  NAND2_X2 U2284 ( .A1(n349), .A2(n243), .ZN(n488) );
  INV_X2 U2285 ( .A(n728), .ZN(n727) );
  NAND2_X2 U2287 ( .A1(n623), .A2(n208), .ZN(n728) );
  INV_X2 U2292 ( .A(n626), .ZN(n625) );
  NAND2_X2 U2293 ( .A1(n623), .A2(n103), .ZN(n626) );
  INV_X2 U2295 ( .A(n865), .ZN(n864) );
  NAND2_X2 U2296 ( .A1(n897), .A2(n67), .ZN(n865) );
  INV_X2 U2297 ( .A(n762), .ZN(n761) );
  NAND2_X2 U2300 ( .A1(n623), .A2(n243), .ZN(n762) );
  INV_X2 U2301 ( .A(n1005), .ZN(n1004) );
  NAND2_X2 U2304 ( .A1(n897), .A2(n208), .ZN(n1005) );
  INV_X2 U2307 ( .A(n903), .ZN(n902) );
  NAND2_X2 U2308 ( .A1(n897), .A2(n103), .ZN(n903) );
  INV_X2 U2905 ( .A(n69), .ZN(n70) );
  NAND2_X2 U2909 ( .A1(n103), .A2(n68), .ZN(n69) );
  INV_X2 U2910 ( .A(n1039), .ZN(n1038) );
  NAND2_X2 U2911 ( .A1(n897), .A2(n243), .ZN(n1039) );
  INV_X2 U2912 ( .A(n279), .ZN(n280) );
  NAND2_X2 U2915 ( .A1(n313), .A2(n68), .ZN(n279) );
  INV_X2 U2916 ( .A(n244), .ZN(n245) );
  NAND2_X2 U2917 ( .A1(n278), .A2(n68), .ZN(n244) );
  INV_X2 U2919 ( .A(n418), .ZN(n419) );
  NAND2_X2 U2924 ( .A1(n349), .A2(n173), .ZN(n418) );
  INV_X2 U2925 ( .A(n384), .ZN(n385) );
  NAND2_X2 U2926 ( .A1(n349), .A2(n138), .ZN(n384) );
  INV_X2 U2927 ( .A(n554), .ZN(n555) );
  NAND2_X2 U2930 ( .A1(n349), .A2(n313), .ZN(n554) );
  INV_X2 U2931 ( .A(n520), .ZN(n521) );
  NAND2_X2 U2932 ( .A1(n349), .A2(n278), .ZN(n520) );
  INV_X2 U2934 ( .A(n692), .ZN(n693) );
  NAND2_X2 U2940 ( .A1(n623), .A2(n173), .ZN(n692) );
  INV_X2 U2941 ( .A(n658), .ZN(n659) );
  NAND2_X2 U2942 ( .A1(n623), .A2(n138), .ZN(n658) );
  INV_X2 U2943 ( .A(n828), .ZN(n829) );
  NAND2_X2 U2946 ( .A1(n623), .A2(n313), .ZN(n828) );
  INV_X2 U2947 ( .A(n794), .ZN(n795) );
  NAND2_X2 U2948 ( .A1(n623), .A2(n278), .ZN(n794) );
  INV_X2 U2950 ( .A(n969), .ZN(n970) );
  NAND2_X2 U2955 ( .A1(n897), .A2(n173), .ZN(n969) );
  INV_X2 U2956 ( .A(n935), .ZN(n936) );
  NAND2_X2 U2958 ( .A1(n897), .A2(n138), .ZN(n935) );
  INV_X2 U2959 ( .A(n1105), .ZN(n1106) );
  NAND2_X2 U2960 ( .A1(n897), .A2(n313), .ZN(n1105) );
  INV_X2 U2963 ( .A(n1071), .ZN(n1072) );
  NAND2_X2 U2964 ( .A1(n897), .A2(n278), .ZN(n1071) );
  INV_X2 U2967 ( .A(n1), .ZN(n3) );
  NAND2_X2 U2970 ( .A1(n67), .A2(n68), .ZN(n1) );
  INV_X4 U2971 ( .A(RESET), .ZN(N352) );
endmodule


module FF_0 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n1, n2, n3, n4;

  DFF_X1 Q_reg ( .D(n4), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n1), .A2(n2), .ZN(n4) );
  INV_X1 U4 ( .A(RESET), .ZN(n2) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n3), .ZN(n1) );
  INV_X1 U6 ( .A(EN), .ZN(n3) );
endmodule


module regFFD_NBIT32_10 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_9 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_8 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_7 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT5_0 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  DFFR_X1 \Q_reg[4]  ( .D(n15), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n10) );
  DFFR_X1 \Q_reg[3]  ( .D(n14), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n9) );
  DFFR_X1 \Q_reg[2]  ( .D(n13), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n8) );
  DFFR_X1 \Q_reg[1]  ( .D(n12), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n7) );
  DFFR_X1 \Q_reg[0]  ( .D(n11), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n6) );
  OAI21_X1 U2 ( .B1(n6), .B2(ENABLE), .A(n1), .ZN(n11) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n7), .B2(ENABLE), .A(n2), .ZN(n12) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n2) );
  OAI21_X1 U6 ( .B1(n8), .B2(ENABLE), .A(n3), .ZN(n13) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n3) );
  OAI21_X1 U8 ( .B1(n9), .B2(ENABLE), .A(n4), .ZN(n14) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n4) );
  OAI21_X1 U10 ( .B1(n10), .B2(ENABLE), .A(n5), .ZN(n15) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n5) );
endmodule


module FF_7 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n5, n6, n7, n8;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n8), .A2(n7), .ZN(n5) );
  INV_X1 U4 ( .A(RESET), .ZN(n7) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n6), .ZN(n8) );
  INV_X1 U6 ( .A(EN), .ZN(n6) );
endmodule


module regFFD_NBIT6_0 ( CK, RESET, ENABLE, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  DFFR_X1 \Q_reg[5]  ( .D(n18), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n12) );
  DFFR_X1 \Q_reg[4]  ( .D(n17), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n11) );
  DFFR_X1 \Q_reg[3]  ( .D(n16), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n10) );
  DFFR_X1 \Q_reg[2]  ( .D(n15), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n9) );
  DFFR_X1 \Q_reg[1]  ( .D(n14), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n8) );
  DFFR_X1 \Q_reg[0]  ( .D(n13), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n7) );
  OAI21_X1 U2 ( .B1(n7), .B2(ENABLE), .A(n1), .ZN(n13) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(n8), .B2(ENABLE), .A(n2), .ZN(n14) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n2) );
  OAI21_X1 U6 ( .B1(n9), .B2(ENABLE), .A(n3), .ZN(n15) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n3) );
  OAI21_X1 U8 ( .B1(n10), .B2(ENABLE), .A(n4), .ZN(n16) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n4) );
  OAI21_X1 U10 ( .B1(n11), .B2(ENABLE), .A(n5), .ZN(n17) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n5) );
  OAI21_X1 U12 ( .B1(n12), .B2(ENABLE), .A(n6), .ZN(n18) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n6) );
endmodule


module regFFD_NBIT32_6 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module IV_224 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_672 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_671 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_670 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_224 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_224 UIV ( .A(S), .Y(SB) );
  ND2_672 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_671 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_670 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_223 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_669 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_668 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_667 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_223 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_223 UIV ( .A(S), .Y(SB) );
  ND2_669 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_668 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_667 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_222 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_666 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_665 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_664 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_222 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_222 UIV ( .A(S), .Y(SB) );
  ND2_666 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_665 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_664 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_221 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_663 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_662 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_661 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_221 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_221 UIV ( .A(S), .Y(SB) );
  ND2_663 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_662 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_661 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_220 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_660 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_659 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_658 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_220 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_220 UIV ( .A(S), .Y(SB) );
  ND2_660 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_659 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_658 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_219 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_657 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_656 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_655 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_219 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_219 UIV ( .A(S), .Y(SB) );
  ND2_657 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_656 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_655 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_218 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_654 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_653 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_652 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_218 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_218 UIV ( .A(S), .Y(SB) );
  ND2_654 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_653 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_652 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_217 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_651 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_650 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_649 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_217 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_217 UIV ( .A(S), .Y(SB) );
  ND2_651 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_650 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_649 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_216 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_648 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_647 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_646 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_216 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_216 UIV ( .A(S), .Y(SB) );
  ND2_648 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_647 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_646 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_215 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_645 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_644 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_643 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_215 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_215 UIV ( .A(S), .Y(SB) );
  ND2_645 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_644 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_643 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_214 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_642 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_641 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_640 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_214 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_214 UIV ( .A(S), .Y(SB) );
  ND2_642 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_641 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_640 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_213 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_639 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_638 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_637 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_213 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_213 UIV ( .A(S), .Y(SB) );
  ND2_639 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_638 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_637 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_212 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_636 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_635 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_634 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_212 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_212 UIV ( .A(S), .Y(SB) );
  ND2_636 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_635 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_634 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_211 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_633 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_632 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_631 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_211 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_211 UIV ( .A(S), .Y(SB) );
  ND2_633 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_632 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_631 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_210 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_630 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_629 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_628 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_210 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_210 UIV ( .A(S), .Y(SB) );
  ND2_630 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_629 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_628 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_209 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_627 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_626 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_625 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_209 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_209 UIV ( .A(S), .Y(SB) );
  ND2_627 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_626 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_625 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_208 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_624 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_623 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_622 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_208 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_208 UIV ( .A(S), .Y(SB) );
  ND2_624 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_623 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_622 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_207 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_621 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_620 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_619 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_207 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_207 UIV ( .A(S), .Y(SB) );
  ND2_621 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_620 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_619 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_206 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_618 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_617 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_616 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_206 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_206 UIV ( .A(S), .Y(SB) );
  ND2_618 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_617 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_616 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_205 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_615 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_614 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_613 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_205 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_205 UIV ( .A(S), .Y(SB) );
  ND2_615 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_614 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_613 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_204 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_612 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_611 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_610 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_204 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_204 UIV ( .A(S), .Y(SB) );
  ND2_612 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_611 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_610 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_203 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_609 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_608 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_607 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_203 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_203 UIV ( .A(S), .Y(SB) );
  ND2_609 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_608 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_607 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_202 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_606 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_605 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_604 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_202 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_202 UIV ( .A(S), .Y(SB) );
  ND2_606 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_605 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_604 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_201 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_603 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_602 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_601 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_201 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_201 UIV ( .A(S), .Y(SB) );
  ND2_603 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_602 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_601 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_200 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_600 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_599 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_598 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_200 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_200 UIV ( .A(S), .Y(SB) );
  ND2_600 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_599 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_598 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_199 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_597 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_596 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_595 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_199 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_199 UIV ( .A(S), .Y(SB) );
  ND2_597 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_596 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_595 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_198 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_594 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_593 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_592 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_198 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_198 UIV ( .A(S), .Y(SB) );
  ND2_594 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_593 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_592 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_197 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_591 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_590 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_589 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_197 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_197 UIV ( .A(S), .Y(SB) );
  ND2_591 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_590 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_589 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_196 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_588 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_587 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_586 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_196 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_196 UIV ( .A(S), .Y(SB) );
  ND2_588 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_587 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_586 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_195 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_585 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_584 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_583 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_195 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_195 UIV ( .A(S), .Y(SB) );
  ND2_585 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_584 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_583 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_194 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_582 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_581 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_580 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_194 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_194 UIV ( .A(S), .Y(SB) );
  ND2_582 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_581 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_580 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_193 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_579 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_578 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_577 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_193 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_193 UIV ( .A(S), .Y(SB) );
  ND2_579 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_578 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_577 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_6 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_224 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_223 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_222 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_221 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_220 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_219 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_218 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_217 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_216 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_215 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_214 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_213 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_212 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_211 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_210 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_209 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_208 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_207 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_206 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_205 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_204 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_203 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_202 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_201 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_200 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_199 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_198 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_197 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_196 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_195 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_194 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_193 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_192 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_576 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_575 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_574 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1, n1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
  INV_X1 U2 ( .A(N1), .ZN(n1) );
  INV_X8 U3 ( .A(n1), .ZN(Y) );
endmodule


module MUX21_192 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_192 UIV ( .A(S), .Y(SB) );
  ND2_576 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_575 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_574 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_191 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_573 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_572 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_571 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1, n1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
  INV_X1 U2 ( .A(N1), .ZN(n1) );
  INV_X8 U3 ( .A(n1), .ZN(Y) );
endmodule


module MUX21_191 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_191 UIV ( .A(S), .Y(SB) );
  ND2_573 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_572 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_571 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_190 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_570 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_569 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_568 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1, n1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
  INV_X1 U2 ( .A(N1), .ZN(n1) );
  INV_X8 U3 ( .A(n1), .ZN(Y) );
endmodule


module MUX21_190 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_190 UIV ( .A(S), .Y(SB) );
  ND2_570 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_569 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_568 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_189 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_567 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_566 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_565 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1, n1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
  INV_X1 U2 ( .A(N1), .ZN(n1) );
  INV_X8 U3 ( .A(n1), .ZN(Y) );
endmodule


module MUX21_189 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_189 UIV ( .A(S), .Y(SB) );
  ND2_567 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_566 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_565 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_188 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_564 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_563 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_562 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_188 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_188 UIV ( .A(S), .Y(SB) );
  ND2_564 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_563 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_562 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_187 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_561 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_560 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_559 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_187 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_187 UIV ( .A(S), .Y(SB) );
  ND2_561 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_560 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_559 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_186 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_558 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_557 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_556 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_186 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_186 UIV ( .A(S), .Y(SB) );
  ND2_558 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_557 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_556 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_185 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_555 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_554 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_553 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_185 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_185 UIV ( .A(S), .Y(SB) );
  ND2_555 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_554 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_553 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_184 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_552 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_551 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_550 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_184 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_184 UIV ( .A(S), .Y(SB) );
  ND2_552 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_551 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_550 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_183 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_549 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_548 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_547 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_183 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_183 UIV ( .A(S), .Y(SB) );
  ND2_549 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_548 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_547 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_182 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_546 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_545 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_544 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_182 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_182 UIV ( .A(S), .Y(SB) );
  ND2_546 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_545 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_544 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_181 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_543 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_542 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_541 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_181 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_181 UIV ( .A(S), .Y(SB) );
  ND2_543 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_542 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_541 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_180 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_540 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_539 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_538 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_180 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_180 UIV ( .A(S), .Y(SB) );
  ND2_540 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_539 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_538 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_179 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_537 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_536 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_535 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_179 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_179 UIV ( .A(S), .Y(SB) );
  ND2_537 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_536 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_535 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_178 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_534 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_533 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_532 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_178 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_178 UIV ( .A(S), .Y(SB) );
  ND2_534 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_533 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_532 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_177 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_531 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_530 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_529 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_177 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_177 UIV ( .A(S), .Y(SB) );
  ND2_531 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_530 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_529 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_176 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_528 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_527 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_526 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_176 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_176 UIV ( .A(S), .Y(SB) );
  ND2_528 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_527 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_526 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_175 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_525 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_524 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_523 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_175 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_175 UIV ( .A(S), .Y(SB) );
  ND2_525 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_524 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_523 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_174 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_522 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_521 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_520 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_174 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_174 UIV ( .A(S), .Y(SB) );
  ND2_522 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_521 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_520 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_173 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_519 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_518 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_517 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_173 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_173 UIV ( .A(S), .Y(SB) );
  ND2_519 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_518 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_517 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_172 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_516 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_515 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_514 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_172 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_172 UIV ( .A(S), .Y(SB) );
  ND2_516 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_515 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_514 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_171 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_513 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_512 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_511 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_171 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_171 UIV ( .A(S), .Y(SB) );
  ND2_513 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_512 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_511 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_170 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_510 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_509 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_508 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_170 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_170 UIV ( .A(S), .Y(SB) );
  ND2_510 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_509 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_508 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_507 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_506 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_505 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_169 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_169 UIV ( .A(S), .Y(SB) );
  ND2_507 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_506 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_505 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_504 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_503 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_502 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_168 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_168 UIV ( .A(S), .Y(SB) );
  ND2_504 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_503 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_502 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_501 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_500 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_499 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_167 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_167 UIV ( .A(S), .Y(SB) );
  ND2_501 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_500 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_499 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_498 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_497 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_496 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_166 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_166 UIV ( .A(S), .Y(SB) );
  ND2_498 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_497 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_496 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_495 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_494 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_493 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_165 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_165 UIV ( .A(S), .Y(SB) );
  ND2_495 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_494 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_493 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_492 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_491 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_490 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_164 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_164 UIV ( .A(S), .Y(SB) );
  ND2_492 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_491 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_490 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_489 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_488 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_487 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_163 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_163 UIV ( .A(S), .Y(SB) );
  ND2_489 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_488 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_487 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_486 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_485 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_484 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_162 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_162 UIV ( .A(S), .Y(SB) );
  ND2_486 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_485 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_484 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_483 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_482 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_481 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_161 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_161 UIV ( .A(S), .Y(SB) );
  ND2_483 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_482 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_481 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_5 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_192 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_191 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_190 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_189 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_188 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_187 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_186 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_185 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_184 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_183 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_182 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_181 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_180 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_179 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_178 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_177 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_176 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_175 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_174 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_173 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_172 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_171 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_170 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_169 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_168 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_167 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_166 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_165 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_164 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_163 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_162 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_161 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module logic_N32 ( .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , 
        \FUNC[1] , \FUNC[0] }), DATA1, DATA2, OUT_ALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUT_ALU;
  input \FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n25, n141, n142, n143, n144
;
  wire   [5:0] FUNC;

  OAI22_X1 U2 ( .A1(n1), .A2(n2), .B1(n3), .B2(n4), .ZN(OUT_ALU[9]) );
  AOI21_X1 U3 ( .B1(n5), .B2(n2), .A(n143), .ZN(n3) );
  INV_X1 U4 ( .A(DATA2[9]), .ZN(n2) );
  AOI221_X1 U5 ( .B1(n5), .B2(n4), .C1(n141), .C2(DATA1[9]), .A(n143), .ZN(n1)
         );
  INV_X1 U6 ( .A(DATA1[9]), .ZN(n4) );
  OAI22_X1 U7 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .ZN(OUT_ALU[8]) );
  AOI21_X1 U8 ( .B1(n5), .B2(n9), .A(n143), .ZN(n10) );
  INV_X1 U9 ( .A(DATA2[8]), .ZN(n9) );
  AOI221_X1 U10 ( .B1(n5), .B2(n11), .C1(DATA1[8]), .C2(n141), .A(n143), .ZN(
        n8) );
  INV_X1 U11 ( .A(DATA1[8]), .ZN(n11) );
  OAI22_X1 U12 ( .A1(n12), .A2(n13), .B1(n14), .B2(n15), .ZN(OUT_ALU[7]) );
  AOI21_X1 U13 ( .B1(n5), .B2(n13), .A(n143), .ZN(n14) );
  INV_X1 U14 ( .A(DATA2[7]), .ZN(n13) );
  AOI221_X1 U15 ( .B1(n5), .B2(n15), .C1(DATA1[7]), .C2(n141), .A(n143), .ZN(
        n12) );
  INV_X1 U16 ( .A(DATA1[7]), .ZN(n15) );
  OAI22_X1 U17 ( .A1(n16), .A2(n17), .B1(n18), .B2(n19), .ZN(OUT_ALU[6]) );
  AOI21_X1 U18 ( .B1(n5), .B2(n17), .A(n143), .ZN(n18) );
  INV_X1 U19 ( .A(DATA2[6]), .ZN(n17) );
  AOI221_X1 U20 ( .B1(n5), .B2(n19), .C1(DATA1[6]), .C2(n141), .A(n143), .ZN(
        n16) );
  INV_X1 U21 ( .A(DATA1[6]), .ZN(n19) );
  OAI22_X1 U22 ( .A1(n20), .A2(n21), .B1(n22), .B2(n23), .ZN(OUT_ALU[5]) );
  AOI21_X1 U23 ( .B1(n5), .B2(n21), .A(n143), .ZN(n22) );
  INV_X1 U24 ( .A(DATA2[5]), .ZN(n21) );
  AOI221_X1 U25 ( .B1(n5), .B2(n23), .C1(DATA1[5]), .C2(n141), .A(n143), .ZN(
        n20) );
  INV_X1 U26 ( .A(DATA1[5]), .ZN(n23) );
  OAI22_X1 U27 ( .A1(n24), .A2(n144), .B1(n26), .B2(n27), .ZN(OUT_ALU[4]) );
  AOI21_X1 U28 ( .B1(n5), .B2(n144), .A(n143), .ZN(n26) );
  AOI221_X1 U30 ( .B1(n5), .B2(n27), .C1(DATA1[4]), .C2(n141), .A(n143), .ZN(
        n24) );
  INV_X1 U31 ( .A(DATA1[4]), .ZN(n27) );
  OAI22_X1 U32 ( .A1(n28), .A2(n29), .B1(n30), .B2(n31), .ZN(OUT_ALU[3]) );
  AOI21_X1 U33 ( .B1(n5), .B2(n29), .A(n143), .ZN(n30) );
  INV_X1 U34 ( .A(DATA2[3]), .ZN(n29) );
  AOI221_X1 U35 ( .B1(n5), .B2(n31), .C1(DATA1[3]), .C2(n141), .A(n143), .ZN(
        n28) );
  INV_X1 U36 ( .A(DATA1[3]), .ZN(n31) );
  OAI22_X1 U37 ( .A1(n32), .A2(n33), .B1(n34), .B2(n35), .ZN(OUT_ALU[31]) );
  AOI21_X1 U38 ( .B1(n5), .B2(n33), .A(n143), .ZN(n34) );
  INV_X1 U39 ( .A(DATA2[31]), .ZN(n33) );
  AOI221_X1 U40 ( .B1(n5), .B2(n35), .C1(DATA1[31]), .C2(n141), .A(n143), .ZN(
        n32) );
  INV_X1 U41 ( .A(DATA1[31]), .ZN(n35) );
  OAI22_X1 U42 ( .A1(n36), .A2(n37), .B1(n38), .B2(n39), .ZN(OUT_ALU[30]) );
  AOI21_X1 U43 ( .B1(n5), .B2(n37), .A(n143), .ZN(n38) );
  INV_X1 U44 ( .A(DATA2[30]), .ZN(n37) );
  AOI221_X1 U45 ( .B1(n5), .B2(n39), .C1(DATA1[30]), .C2(n141), .A(n143), .ZN(
        n36) );
  INV_X1 U46 ( .A(DATA1[30]), .ZN(n39) );
  OAI22_X1 U47 ( .A1(n40), .A2(n41), .B1(n42), .B2(n43), .ZN(OUT_ALU[2]) );
  AOI21_X1 U48 ( .B1(n5), .B2(n41), .A(n143), .ZN(n42) );
  INV_X1 U49 ( .A(DATA2[2]), .ZN(n41) );
  AOI221_X1 U50 ( .B1(n5), .B2(n43), .C1(DATA1[2]), .C2(n141), .A(n143), .ZN(
        n40) );
  INV_X1 U51 ( .A(DATA1[2]), .ZN(n43) );
  OAI22_X1 U52 ( .A1(n44), .A2(n45), .B1(n46), .B2(n47), .ZN(OUT_ALU[29]) );
  AOI21_X1 U53 ( .B1(n5), .B2(n45), .A(n143), .ZN(n46) );
  INV_X1 U54 ( .A(DATA2[29]), .ZN(n45) );
  AOI221_X1 U55 ( .B1(n5), .B2(n47), .C1(DATA1[29]), .C2(n141), .A(n143), .ZN(
        n44) );
  INV_X1 U56 ( .A(DATA1[29]), .ZN(n47) );
  OAI22_X1 U57 ( .A1(n48), .A2(n49), .B1(n50), .B2(n51), .ZN(OUT_ALU[28]) );
  AOI21_X1 U58 ( .B1(n5), .B2(n49), .A(n143), .ZN(n50) );
  INV_X1 U59 ( .A(DATA2[28]), .ZN(n49) );
  AOI221_X1 U60 ( .B1(n5), .B2(n51), .C1(DATA1[28]), .C2(n141), .A(n143), .ZN(
        n48) );
  INV_X1 U61 ( .A(DATA1[28]), .ZN(n51) );
  OAI22_X1 U62 ( .A1(n52), .A2(n53), .B1(n54), .B2(n55), .ZN(OUT_ALU[27]) );
  AOI21_X1 U63 ( .B1(n5), .B2(n53), .A(n143), .ZN(n54) );
  INV_X1 U64 ( .A(DATA2[27]), .ZN(n53) );
  AOI221_X1 U65 ( .B1(n5), .B2(n55), .C1(DATA1[27]), .C2(n141), .A(n143), .ZN(
        n52) );
  INV_X1 U66 ( .A(DATA1[27]), .ZN(n55) );
  OAI22_X1 U67 ( .A1(n56), .A2(n57), .B1(n58), .B2(n59), .ZN(OUT_ALU[26]) );
  AOI21_X1 U68 ( .B1(n5), .B2(n57), .A(n143), .ZN(n58) );
  INV_X1 U69 ( .A(DATA2[26]), .ZN(n57) );
  AOI221_X1 U70 ( .B1(n5), .B2(n59), .C1(DATA1[26]), .C2(n141), .A(n143), .ZN(
        n56) );
  INV_X1 U71 ( .A(DATA1[26]), .ZN(n59) );
  OAI22_X1 U72 ( .A1(n60), .A2(n61), .B1(n62), .B2(n63), .ZN(OUT_ALU[25]) );
  AOI21_X1 U73 ( .B1(n5), .B2(n61), .A(n143), .ZN(n62) );
  INV_X1 U74 ( .A(DATA2[25]), .ZN(n61) );
  AOI221_X1 U75 ( .B1(n5), .B2(n63), .C1(DATA1[25]), .C2(n141), .A(n143), .ZN(
        n60) );
  INV_X1 U76 ( .A(DATA1[25]), .ZN(n63) );
  OAI22_X1 U77 ( .A1(n64), .A2(n65), .B1(n66), .B2(n67), .ZN(OUT_ALU[24]) );
  AOI21_X1 U78 ( .B1(n5), .B2(n65), .A(n143), .ZN(n66) );
  INV_X1 U79 ( .A(DATA2[24]), .ZN(n65) );
  AOI221_X1 U80 ( .B1(n5), .B2(n67), .C1(DATA1[24]), .C2(n141), .A(n143), .ZN(
        n64) );
  INV_X1 U81 ( .A(DATA1[24]), .ZN(n67) );
  OAI22_X1 U82 ( .A1(n68), .A2(n69), .B1(n70), .B2(n71), .ZN(OUT_ALU[23]) );
  AOI21_X1 U83 ( .B1(n5), .B2(n69), .A(n143), .ZN(n70) );
  INV_X1 U84 ( .A(DATA2[23]), .ZN(n69) );
  AOI221_X1 U85 ( .B1(n5), .B2(n71), .C1(DATA1[23]), .C2(n141), .A(n143), .ZN(
        n68) );
  INV_X1 U86 ( .A(DATA1[23]), .ZN(n71) );
  OAI22_X1 U87 ( .A1(n72), .A2(n73), .B1(n74), .B2(n75), .ZN(OUT_ALU[22]) );
  AOI21_X1 U88 ( .B1(n5), .B2(n73), .A(n143), .ZN(n74) );
  INV_X1 U89 ( .A(DATA2[22]), .ZN(n73) );
  AOI221_X1 U90 ( .B1(n5), .B2(n75), .C1(DATA1[22]), .C2(n141), .A(n143), .ZN(
        n72) );
  INV_X1 U91 ( .A(DATA1[22]), .ZN(n75) );
  OAI22_X1 U92 ( .A1(n76), .A2(n77), .B1(n78), .B2(n79), .ZN(OUT_ALU[21]) );
  AOI21_X1 U93 ( .B1(n5), .B2(n77), .A(n143), .ZN(n78) );
  INV_X1 U94 ( .A(DATA2[21]), .ZN(n77) );
  AOI221_X1 U95 ( .B1(n5), .B2(n79), .C1(DATA1[21]), .C2(n141), .A(n143), .ZN(
        n76) );
  INV_X1 U96 ( .A(DATA1[21]), .ZN(n79) );
  OAI22_X1 U97 ( .A1(n80), .A2(n81), .B1(n82), .B2(n83), .ZN(OUT_ALU[20]) );
  AOI21_X1 U98 ( .B1(n5), .B2(n81), .A(n143), .ZN(n82) );
  INV_X1 U99 ( .A(DATA2[20]), .ZN(n81) );
  AOI221_X1 U100 ( .B1(n5), .B2(n83), .C1(DATA1[20]), .C2(n141), .A(n143), 
        .ZN(n80) );
  INV_X1 U101 ( .A(DATA1[20]), .ZN(n83) );
  OAI22_X1 U102 ( .A1(n84), .A2(n85), .B1(n86), .B2(n87), .ZN(OUT_ALU[1]) );
  AOI21_X1 U103 ( .B1(n5), .B2(n85), .A(n143), .ZN(n86) );
  INV_X1 U104 ( .A(DATA2[1]), .ZN(n85) );
  AOI221_X1 U105 ( .B1(n5), .B2(n87), .C1(DATA1[1]), .C2(n141), .A(n143), .ZN(
        n84) );
  INV_X1 U106 ( .A(DATA1[1]), .ZN(n87) );
  OAI22_X1 U107 ( .A1(n88), .A2(n89), .B1(n90), .B2(n91), .ZN(OUT_ALU[19]) );
  AOI21_X1 U108 ( .B1(n5), .B2(n89), .A(n143), .ZN(n90) );
  INV_X1 U109 ( .A(DATA2[19]), .ZN(n89) );
  AOI221_X1 U110 ( .B1(n5), .B2(n91), .C1(DATA1[19]), .C2(n141), .A(n143), 
        .ZN(n88) );
  INV_X1 U111 ( .A(DATA1[19]), .ZN(n91) );
  OAI22_X1 U112 ( .A1(n92), .A2(n93), .B1(n94), .B2(n95), .ZN(OUT_ALU[18]) );
  AOI21_X1 U113 ( .B1(n5), .B2(n93), .A(n143), .ZN(n94) );
  INV_X1 U114 ( .A(DATA2[18]), .ZN(n93) );
  AOI221_X1 U115 ( .B1(n5), .B2(n95), .C1(DATA1[18]), .C2(n141), .A(n143), 
        .ZN(n92) );
  INV_X1 U116 ( .A(DATA1[18]), .ZN(n95) );
  OAI22_X1 U117 ( .A1(n96), .A2(n97), .B1(n98), .B2(n99), .ZN(OUT_ALU[17]) );
  AOI21_X1 U118 ( .B1(n5), .B2(n97), .A(n143), .ZN(n98) );
  INV_X1 U119 ( .A(DATA2[17]), .ZN(n97) );
  AOI221_X1 U120 ( .B1(n5), .B2(n99), .C1(DATA1[17]), .C2(n141), .A(n143), 
        .ZN(n96) );
  INV_X1 U121 ( .A(DATA1[17]), .ZN(n99) );
  OAI22_X1 U122 ( .A1(n100), .A2(n101), .B1(n102), .B2(n103), .ZN(OUT_ALU[16])
         );
  AOI21_X1 U123 ( .B1(n5), .B2(n101), .A(n143), .ZN(n102) );
  INV_X1 U124 ( .A(DATA2[16]), .ZN(n101) );
  AOI221_X1 U125 ( .B1(n5), .B2(n103), .C1(DATA1[16]), .C2(n141), .A(n143), 
        .ZN(n100) );
  INV_X1 U126 ( .A(DATA1[16]), .ZN(n103) );
  OAI22_X1 U127 ( .A1(n104), .A2(n105), .B1(n106), .B2(n107), .ZN(OUT_ALU[15])
         );
  AOI21_X1 U128 ( .B1(n5), .B2(n105), .A(n143), .ZN(n106) );
  INV_X1 U129 ( .A(DATA2[15]), .ZN(n105) );
  AOI221_X1 U130 ( .B1(n5), .B2(n107), .C1(DATA1[15]), .C2(n141), .A(n143), 
        .ZN(n104) );
  INV_X1 U131 ( .A(DATA1[15]), .ZN(n107) );
  OAI22_X1 U132 ( .A1(n108), .A2(n109), .B1(n110), .B2(n111), .ZN(OUT_ALU[14])
         );
  AOI21_X1 U133 ( .B1(n5), .B2(n109), .A(n143), .ZN(n110) );
  INV_X1 U134 ( .A(DATA2[14]), .ZN(n109) );
  AOI221_X1 U135 ( .B1(n5), .B2(n111), .C1(DATA1[14]), .C2(n141), .A(n143), 
        .ZN(n108) );
  INV_X1 U136 ( .A(DATA1[14]), .ZN(n111) );
  OAI22_X1 U137 ( .A1(n112), .A2(n113), .B1(n114), .B2(n115), .ZN(OUT_ALU[13])
         );
  AOI21_X1 U138 ( .B1(n5), .B2(n113), .A(n143), .ZN(n114) );
  INV_X1 U139 ( .A(DATA2[13]), .ZN(n113) );
  AOI221_X1 U140 ( .B1(n5), .B2(n115), .C1(DATA1[13]), .C2(n141), .A(n143), 
        .ZN(n112) );
  INV_X1 U141 ( .A(DATA1[13]), .ZN(n115) );
  OAI22_X1 U142 ( .A1(n116), .A2(n117), .B1(n118), .B2(n119), .ZN(OUT_ALU[12])
         );
  AOI21_X1 U143 ( .B1(n5), .B2(n117), .A(n143), .ZN(n118) );
  INV_X1 U144 ( .A(DATA2[12]), .ZN(n117) );
  AOI221_X1 U145 ( .B1(n5), .B2(n119), .C1(DATA1[12]), .C2(n141), .A(n143), 
        .ZN(n116) );
  INV_X1 U146 ( .A(DATA1[12]), .ZN(n119) );
  OAI22_X1 U147 ( .A1(n120), .A2(n121), .B1(n122), .B2(n123), .ZN(OUT_ALU[11])
         );
  AOI21_X1 U148 ( .B1(n5), .B2(n121), .A(n143), .ZN(n122) );
  INV_X1 U149 ( .A(DATA2[11]), .ZN(n121) );
  AOI221_X1 U150 ( .B1(n5), .B2(n123), .C1(DATA1[11]), .C2(n141), .A(n143), 
        .ZN(n120) );
  INV_X1 U151 ( .A(DATA1[11]), .ZN(n123) );
  OAI22_X1 U152 ( .A1(n124), .A2(n125), .B1(n126), .B2(n127), .ZN(OUT_ALU[10])
         );
  AOI21_X1 U153 ( .B1(n5), .B2(n125), .A(n143), .ZN(n126) );
  INV_X1 U154 ( .A(DATA2[10]), .ZN(n125) );
  AOI221_X1 U155 ( .B1(n5), .B2(n127), .C1(DATA1[10]), .C2(n141), .A(n143), 
        .ZN(n124) );
  INV_X1 U156 ( .A(DATA1[10]), .ZN(n127) );
  OAI22_X1 U157 ( .A1(n128), .A2(n129), .B1(n130), .B2(n131), .ZN(OUT_ALU[0])
         );
  AOI21_X1 U158 ( .B1(n5), .B2(n129), .A(n143), .ZN(n130) );
  INV_X1 U159 ( .A(DATA2[0]), .ZN(n129) );
  AOI221_X1 U160 ( .B1(n5), .B2(n131), .C1(DATA1[0]), .C2(n141), .A(n143), 
        .ZN(n128) );
  OAI21_X1 U161 ( .B1(FUNC[0]), .B2(n132), .A(n133), .ZN(n6) );
  OR3_X1 U162 ( .A1(n134), .A2(FUNC[3]), .A3(n135), .ZN(n133) );
  AOI21_X1 U163 ( .B1(n135), .B2(FUNC[3]), .A(n134), .ZN(n7) );
  NAND4_X1 U164 ( .A1(FUNC[2]), .A2(FUNC[1]), .A3(n136), .A4(n137), .ZN(n134)
         );
  INV_X1 U165 ( .A(FUNC[5]), .ZN(n137) );
  INV_X1 U166 ( .A(DATA1[0]), .ZN(n131) );
  NAND4_X1 U168 ( .A1(FUNC[3]), .A2(n139), .A3(n135), .A4(n136), .ZN(n138) );
  INV_X1 U169 ( .A(FUNC[4]), .ZN(n136) );
  INV_X1 U170 ( .A(FUNC[0]), .ZN(n135) );
  NAND3_X1 U171 ( .A1(n139), .A2(n140), .A3(FUNC[4]), .ZN(n132) );
  INV_X1 U172 ( .A(FUNC[3]), .ZN(n140) );
  NOR3_X1 U173 ( .A1(FUNC[2]), .A2(FUNC[5]), .A3(FUNC[1]), .ZN(n139) );
  INV_X1 U29 ( .A(n7), .ZN(n25) );
  INV_X2 U167 ( .A(n25), .ZN(n141) );
  NAND2_X4 U174 ( .A1(n132), .A2(n138), .ZN(n5) );
  INV_X1 U175 ( .A(n6), .ZN(n142) );
  INV_X4 U176 ( .A(n142), .ZN(n143) );
  INV_X1 U177 ( .A(DATA2[4]), .ZN(n144) );
endmodule


module comparator ( DATA1, DATA2i, .tipo({\tipo[5] , \tipo[4] , \tipo[3] , 
        \tipo[2] , \tipo[1] , \tipo[0] }), OUTALU );
  input [31:0] DATA1;
  output [31:0] OUTALU;
  input DATA2i, \tipo[5] , \tipo[4] , \tipo[3] , \tipo[2] , \tipo[1] ,
         \tipo[0] ;
  wire   N57, N58, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49;
  wire   [5:0] tipo;
  assign OUTALU[31] = 1'b0;
  assign OUTALU[30] = 1'b0;
  assign OUTALU[29] = 1'b0;
  assign OUTALU[28] = 1'b0;
  assign OUTALU[27] = 1'b0;
  assign OUTALU[26] = 1'b0;
  assign OUTALU[25] = 1'b0;
  assign OUTALU[24] = 1'b0;
  assign OUTALU[23] = 1'b0;
  assign OUTALU[22] = 1'b0;
  assign OUTALU[21] = 1'b0;
  assign OUTALU[20] = 1'b0;
  assign OUTALU[19] = 1'b0;
  assign OUTALU[18] = 1'b0;
  assign OUTALU[17] = 1'b0;
  assign OUTALU[16] = 1'b0;
  assign OUTALU[15] = 1'b0;
  assign OUTALU[14] = 1'b0;
  assign OUTALU[13] = 1'b0;
  assign OUTALU[12] = 1'b0;
  assign OUTALU[11] = 1'b0;
  assign OUTALU[10] = 1'b0;
  assign OUTALU[9] = 1'b0;
  assign OUTALU[8] = 1'b0;
  assign OUTALU[7] = 1'b0;
  assign OUTALU[6] = 1'b0;
  assign OUTALU[5] = 1'b0;
  assign OUTALU[4] = 1'b0;
  assign OUTALU[3] = 1'b0;
  assign OUTALU[2] = 1'b0;
  assign OUTALU[1] = 1'b0;

  DLH_X1 \OUTALU_reg[0]  ( .G(N57), .D(N58), .Q(OUTALU[0]) );
  OAI211_X1 U33 ( .C1(n1), .C2(n2), .A(n3), .B(n4), .ZN(N58) );
  AOI22_X1 U34 ( .A1(n5), .A2(n2), .B1(n6), .B2(n7), .ZN(n4) );
  OAI21_X1 U35 ( .B1(n8), .B2(n9), .A(n10), .ZN(n3) );
  INV_X1 U36 ( .A(DATA2i), .ZN(n2) );
  AOI21_X1 U37 ( .B1(n11), .B2(n7), .A(n12), .ZN(n1) );
  INV_X1 U38 ( .A(n10), .ZN(n7) );
  NOR2_X1 U39 ( .A1(n13), .A2(n14), .ZN(n10) );
  NAND4_X1 U40 ( .A1(n15), .A2(n16), .A3(n17), .A4(n18), .ZN(n14) );
  NOR4_X1 U41 ( .A1(DATA1[23]), .A2(DATA1[22]), .A3(DATA1[21]), .A4(DATA1[20]), 
        .ZN(n18) );
  NOR4_X1 U42 ( .A1(DATA1[1]), .A2(DATA1[19]), .A3(DATA1[18]), .A4(DATA1[17]), 
        .ZN(n17) );
  NOR4_X1 U43 ( .A1(DATA1[16]), .A2(DATA1[15]), .A3(DATA1[14]), .A4(DATA1[13]), 
        .ZN(n16) );
  NOR4_X1 U44 ( .A1(DATA1[12]), .A2(DATA1[11]), .A3(DATA1[10]), .A4(DATA1[0]), 
        .ZN(n15) );
  NAND4_X1 U45 ( .A1(n19), .A2(n20), .A3(n21), .A4(n22), .ZN(n13) );
  NOR4_X1 U46 ( .A1(DATA1[9]), .A2(DATA1[8]), .A3(DATA1[7]), .A4(DATA1[6]), 
        .ZN(n22) );
  NOR4_X1 U47 ( .A1(DATA1[5]), .A2(DATA1[4]), .A3(DATA1[3]), .A4(DATA1[31]), 
        .ZN(n21) );
  NOR4_X1 U48 ( .A1(DATA1[30]), .A2(DATA1[2]), .A3(DATA1[29]), .A4(DATA1[28]), 
        .ZN(n20) );
  NOR4_X1 U49 ( .A1(DATA1[27]), .A2(DATA1[26]), .A3(DATA1[25]), .A4(DATA1[24]), 
        .ZN(n19) );
  OR4_X1 U50 ( .A1(n6), .A2(n5), .A3(n23), .A4(n11), .ZN(N57) );
  OAI21_X1 U51 ( .B1(n24), .B2(n25), .A(n26), .ZN(n11) );
  INV_X1 U52 ( .A(n27), .ZN(n26) );
  AOI21_X1 U53 ( .B1(n28), .B2(n29), .A(n30), .ZN(n27) );
  OR2_X1 U54 ( .A1(n8), .A2(n12), .ZN(n23) );
  OAI221_X1 U55 ( .B1(n31), .B2(n28), .C1(n25), .C2(n32), .A(n33), .ZN(n12) );
  INV_X1 U56 ( .A(n34), .ZN(n33) );
  AOI211_X1 U57 ( .C1(n29), .C2(n35), .A(n36), .B(n37), .ZN(n34) );
  NAND4_X1 U58 ( .A1(tipo[5]), .A2(tipo[4]), .A3(n38), .A4(n39), .ZN(n28) );
  INV_X1 U59 ( .A(tipo[2]), .ZN(n38) );
  OAI21_X1 U60 ( .B1(n40), .B2(n30), .A(n41), .ZN(n8) );
  NAND4_X1 U61 ( .A1(tipo[4]), .A2(tipo[2]), .A3(n42), .A4(n43), .ZN(n41) );
  INV_X1 U62 ( .A(n25), .ZN(n43) );
  NOR2_X1 U63 ( .A1(tipo[5]), .A2(n39), .ZN(n42) );
  OAI221_X1 U64 ( .B1(n44), .B2(n45), .C1(n24), .C2(n31), .A(n46), .ZN(n5) );
  INV_X1 U65 ( .A(n9), .ZN(n46) );
  OAI22_X1 U66 ( .A1(n31), .A2(n32), .B1(n25), .B2(n35), .ZN(n9) );
  NAND2_X1 U67 ( .A1(tipo[1]), .A2(n37), .ZN(n25) );
  AND2_X1 U68 ( .A1(n40), .A2(n29), .ZN(n24) );
  NAND3_X1 U69 ( .A1(n47), .A2(n39), .A3(tipo[5]), .ZN(n29) );
  NAND3_X1 U70 ( .A1(tipo[3]), .A2(n47), .A3(tipo[5]), .ZN(n40) );
  NAND2_X1 U71 ( .A1(tipo[0]), .A2(tipo[2]), .ZN(n45) );
  NAND3_X1 U72 ( .A1(tipo[3]), .A2(n48), .A3(tipo[1]), .ZN(n44) );
  XNOR2_X1 U73 ( .A(n49), .B(tipo[4]), .ZN(n48) );
  OAI22_X1 U74 ( .A1(n35), .A2(n31), .B1(n32), .B2(n30), .ZN(n6) );
  NAND2_X1 U75 ( .A1(n37), .A2(n36), .ZN(n30) );
  INV_X1 U76 ( .A(tipo[0]), .ZN(n37) );
  NAND4_X1 U77 ( .A1(tipo[4]), .A2(tipo[2]), .A3(n39), .A4(n49), .ZN(n32) );
  INV_X1 U78 ( .A(tipo[3]), .ZN(n39) );
  NAND2_X1 U79 ( .A1(tipo[0]), .A2(n36), .ZN(n31) );
  INV_X1 U80 ( .A(tipo[1]), .ZN(n36) );
  NAND3_X1 U81 ( .A1(n47), .A2(n49), .A3(tipo[3]), .ZN(n35) );
  INV_X1 U82 ( .A(tipo[5]), .ZN(n49) );
  NOR2_X1 U83 ( .A1(tipo[4]), .A2(tipo[2]), .ZN(n47) );
endmodule


module SHIFTER_GENERIC_N32_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [3:0] SHMAG;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n1), .Z(B[31]) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n1), .Z(B[30]) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n1), .Z(B[29]) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n1), .Z(B[28]) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n1), .Z(B[27]) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n1), .Z(B[26]) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n1), .Z(B[25])
         );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n1), .Z(B[24])
         );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n1), .Z(B[23])
         );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n1), .Z(B[22])
         );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n1), .Z(B[21])
         );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n1), .Z(B[20])
         );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n2), .Z(B[19])
         );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n2), .Z(B[18])
         );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n2), .Z(B[17])
         );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n2), .Z(B[16])
         );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(SH[3]), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(SH[3]), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(SH[3]), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(SH[3]), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(SH[3]), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(SH[3]), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(SH[3]), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(SH[3]), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(SH[3]), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(SH[3]), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(SH[3]), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(SH[3]), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(SH[3]), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(SH[3]), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(SH[3]), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(SH[3]), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(SH[3]), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(SH[3]), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(SH[2]), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(SH[2]), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(SH[2]), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(SH[2]), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(SH[2]), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(SH[2]), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(SH[2]), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(SH[2]), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(SH[2]), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(SH[2]), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(SH[2]), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(SH[2]), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(SH[1]), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(SH[1]), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(SH[1]), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(SH[1]), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(SH[1]), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(SH[1]), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(SH[1]), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(SH[1]), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(SH[1]), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(SH[1]), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(SH[1]), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(SH[1]), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(SH[0]), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(SH[0]), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(SH[0]), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(SH[0]), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(SH[0]), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  INV_X1 U3 ( .A(n3), .ZN(n1) );
  INV_X1 U4 ( .A(n3), .ZN(n2) );
  INV_X1 U5 ( .A(SH[4]), .ZN(n3) );
  INV_X1 U6 ( .A(SH[4]), .ZN(n4) );
  INV_X1 U7 ( .A(SH[4]), .ZN(n5) );
  AND2_X1 U8 ( .A1(\ML_int[4][9] ), .A2(n5), .ZN(B[9]) );
  AND2_X1 U9 ( .A1(\ML_int[4][8] ), .A2(n5), .ZN(B[8]) );
  NOR2_X1 U10 ( .A1(n2), .A2(n6), .ZN(B[7]) );
  NOR2_X1 U11 ( .A1(n2), .A2(n7), .ZN(B[6]) );
  NOR2_X1 U12 ( .A1(n2), .A2(n8), .ZN(B[5]) );
  NOR2_X1 U13 ( .A1(n2), .A2(n9), .ZN(B[4]) );
  NOR2_X1 U14 ( .A1(n2), .A2(n10), .ZN(B[3]) );
  NOR2_X1 U15 ( .A1(n2), .A2(n11), .ZN(B[2]) );
  NOR2_X1 U16 ( .A1(n2), .A2(n12), .ZN(B[1]) );
  AND2_X1 U17 ( .A1(\ML_int[4][15] ), .A2(n5), .ZN(B[15]) );
  AND2_X1 U18 ( .A1(\ML_int[4][14] ), .A2(n4), .ZN(B[14]) );
  AND2_X1 U19 ( .A1(\ML_int[4][13] ), .A2(n4), .ZN(B[13]) );
  AND2_X1 U20 ( .A1(\ML_int[4][12] ), .A2(n4), .ZN(B[12]) );
  AND2_X1 U21 ( .A1(\ML_int[4][11] ), .A2(n4), .ZN(B[11]) );
  AND2_X1 U22 ( .A1(\ML_int[4][10] ), .A2(n3), .ZN(B[10]) );
  NOR2_X1 U23 ( .A1(n2), .A2(n13), .ZN(B[0]) );
  INV_X1 U24 ( .A(n6), .ZN(\ML_int[4][7] ) );
  NAND2_X1 U25 ( .A1(\ML_int[3][7] ), .A2(SHMAG[3]), .ZN(n6) );
  INV_X1 U26 ( .A(n7), .ZN(\ML_int[4][6] ) );
  NAND2_X1 U27 ( .A1(\ML_int[3][6] ), .A2(SHMAG[3]), .ZN(n7) );
  INV_X1 U28 ( .A(n8), .ZN(\ML_int[4][5] ) );
  NAND2_X1 U29 ( .A1(\ML_int[3][5] ), .A2(SHMAG[3]), .ZN(n8) );
  INV_X1 U30 ( .A(n9), .ZN(\ML_int[4][4] ) );
  NAND2_X1 U31 ( .A1(\ML_int[3][4] ), .A2(SHMAG[3]), .ZN(n9) );
  INV_X1 U32 ( .A(n10), .ZN(\ML_int[4][3] ) );
  NAND2_X1 U33 ( .A1(\ML_int[3][3] ), .A2(SHMAG[3]), .ZN(n10) );
  INV_X1 U34 ( .A(n11), .ZN(\ML_int[4][2] ) );
  NAND2_X1 U35 ( .A1(\ML_int[3][2] ), .A2(SHMAG[3]), .ZN(n11) );
  INV_X1 U36 ( .A(n12), .ZN(\ML_int[4][1] ) );
  NAND2_X1 U37 ( .A1(\ML_int[3][1] ), .A2(SHMAG[3]), .ZN(n12) );
  INV_X1 U38 ( .A(n13), .ZN(\ML_int[4][0] ) );
  NAND2_X1 U39 ( .A1(\ML_int[3][0] ), .A2(SHMAG[3]), .ZN(n13) );
  INV_X1 U40 ( .A(SH[3]), .ZN(SHMAG[3]) );
  AND2_X1 U41 ( .A1(\ML_int[2][3] ), .A2(SHMAG[2]), .ZN(\ML_int[3][3] ) );
  AND2_X1 U42 ( .A1(\ML_int[2][2] ), .A2(SHMAG[2]), .ZN(\ML_int[3][2] ) );
  AND2_X1 U43 ( .A1(\ML_int[2][1] ), .A2(SHMAG[2]), .ZN(\ML_int[3][1] ) );
  AND2_X1 U44 ( .A1(\ML_int[2][0] ), .A2(SHMAG[2]), .ZN(\ML_int[3][0] ) );
  INV_X1 U45 ( .A(SH[2]), .ZN(SHMAG[2]) );
  AND2_X1 U46 ( .A1(\ML_int[1][1] ), .A2(SHMAG[1]), .ZN(\ML_int[2][1] ) );
  AND2_X1 U47 ( .A1(\ML_int[1][0] ), .A2(SHMAG[1]), .ZN(\ML_int[2][0] ) );
  INV_X1 U48 ( .A(SH[1]), .ZN(SHMAG[1]) );
  AND2_X1 U49 ( .A1(A[0]), .A2(SHMAG[0]), .ZN(\ML_int[1][0] ) );
  INV_X1 U50 ( .A(SH[0]), .ZN(SHMAG[0]) );
endmodule


module SHIFTER_GENERIC_N32_DW_sla_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178;
  assign B[0] = \A[0] ;
  assign \A[0]  = A[0];

  NOR2_X2 U2 ( .A1(SH[2]), .A2(SH[3]), .ZN(n76) );
  NAND2_X2 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n27) );
  OAI221_X4 U4 ( .B1(n25), .B2(n169), .C1(n27), .C2(n152), .A(n176), .ZN(n102)
         );
  OAI221_X4 U5 ( .B1(n25), .B2(n164), .C1(n27), .C2(n171), .A(n172), .ZN(n97)
         );
  OAI221_X4 U6 ( .B1(n25), .B2(n162), .C1(n27), .C2(n169), .A(n170), .ZN(n95)
         );
  OAI221_X4 U7 ( .B1(n25), .B2(n153), .C1(n27), .C2(n164), .A(n165), .ZN(n88)
         );
  OAI221_X4 U8 ( .B1(n25), .B2(n150), .C1(n27), .C2(n162), .A(n163), .ZN(n86)
         );
  NAND2_X2 U9 ( .A1(SH[1]), .A2(n178), .ZN(n25) );
  INV_X1 U10 ( .A(n31), .ZN(n1) );
  INV_X2 U11 ( .A(n1), .ZN(n2) );
  INV_X1 U12 ( .A(n30), .ZN(n3) );
  INV_X2 U13 ( .A(n3), .ZN(n4) );
  INV_X1 U14 ( .A(SH[4]), .ZN(n5) );
  INV_X1 U15 ( .A(SH[4]), .ZN(n6) );
  OAI21_X1 U16 ( .B1(SH[4]), .B2(n7), .A(n8), .ZN(B[9]) );
  OAI21_X1 U17 ( .B1(SH[4]), .B2(n9), .A(n8), .ZN(B[8]) );
  OAI21_X1 U18 ( .B1(SH[4]), .B2(n10), .A(n8), .ZN(B[7]) );
  OAI21_X1 U19 ( .B1(SH[4]), .B2(n11), .A(n8), .ZN(B[6]) );
  OAI21_X1 U20 ( .B1(SH[4]), .B2(n12), .A(n8), .ZN(B[5]) );
  OAI21_X1 U21 ( .B1(SH[4]), .B2(n13), .A(n8), .ZN(B[4]) );
  OAI21_X1 U22 ( .B1(SH[4]), .B2(n14), .A(n8), .ZN(B[3]) );
  OAI221_X1 U23 ( .B1(n15), .B2(n16), .C1(n17), .C2(n5), .A(n18), .ZN(B[31])
         );
  AOI222_X1 U24 ( .A1(n19), .A2(n20), .B1(n21), .B2(n22), .C1(n23), .C2(n24), 
        .ZN(n18) );
  OAI221_X1 U25 ( .B1(n25), .B2(n26), .C1(n27), .C2(n28), .A(n29), .ZN(n22) );
  AOI22_X1 U26 ( .A1(A[30]), .A2(n4), .B1(A[31]), .B2(n2), .ZN(n29) );
  INV_X1 U27 ( .A(A[29]), .ZN(n26) );
  OAI221_X1 U28 ( .B1(n32), .B2(n16), .C1(n33), .C2(n5), .A(n34), .ZN(B[30])
         );
  AOI222_X1 U29 ( .A1(n19), .A2(n35), .B1(n21), .B2(n36), .C1(n23), .C2(n37), 
        .ZN(n34) );
  OAI221_X1 U30 ( .B1(n25), .B2(n28), .C1(n27), .C2(n38), .A(n39), .ZN(n36) );
  AOI22_X1 U31 ( .A1(A[29]), .A2(n4), .B1(A[30]), .B2(n2), .ZN(n39) );
  INV_X1 U32 ( .A(A[28]), .ZN(n28) );
  OAI21_X1 U33 ( .B1(SH[4]), .B2(n40), .A(n8), .ZN(B[2]) );
  OAI221_X1 U34 ( .B1(n41), .B2(n16), .C1(n42), .C2(n5), .A(n43), .ZN(B[29])
         );
  AOI222_X1 U35 ( .A1(n19), .A2(n44), .B1(n21), .B2(n45), .C1(n23), .C2(n46), 
        .ZN(n43) );
  OAI221_X1 U36 ( .B1(n25), .B2(n38), .C1(n27), .C2(n47), .A(n48), .ZN(n45) );
  AOI22_X1 U37 ( .A1(A[28]), .A2(n4), .B1(A[29]), .B2(n2), .ZN(n48) );
  INV_X1 U38 ( .A(A[27]), .ZN(n38) );
  OAI221_X1 U39 ( .B1(n49), .B2(n16), .C1(n50), .C2(n5), .A(n51), .ZN(B[28])
         );
  AOI222_X1 U40 ( .A1(n19), .A2(n52), .B1(n21), .B2(n53), .C1(n23), .C2(n54), 
        .ZN(n51) );
  OAI221_X1 U41 ( .B1(n25), .B2(n47), .C1(n27), .C2(n55), .A(n56), .ZN(n53) );
  AOI22_X1 U42 ( .A1(A[27]), .A2(n4), .B1(A[28]), .B2(n2), .ZN(n56) );
  INV_X1 U43 ( .A(A[26]), .ZN(n47) );
  INV_X1 U44 ( .A(n57), .ZN(n21) );
  OAI221_X1 U45 ( .B1(n15), .B2(n57), .C1(n58), .C2(n5), .A(n59), .ZN(B[27])
         );
  AOI222_X1 U46 ( .A1(n60), .A2(n24), .B1(n23), .B2(n20), .C1(n19), .C2(n61), 
        .ZN(n59) );
  INV_X1 U47 ( .A(n62), .ZN(n15) );
  OAI221_X1 U48 ( .B1(n25), .B2(n55), .C1(n27), .C2(n63), .A(n64), .ZN(n62) );
  AOI22_X1 U49 ( .A1(A[26]), .A2(n4), .B1(A[27]), .B2(n2), .ZN(n64) );
  INV_X1 U50 ( .A(A[25]), .ZN(n55) );
  OAI221_X1 U51 ( .B1(n32), .B2(n57), .C1(n65), .C2(n5), .A(n66), .ZN(B[26])
         );
  AOI222_X1 U52 ( .A1(n60), .A2(n37), .B1(n23), .B2(n35), .C1(n19), .C2(n67), 
        .ZN(n66) );
  INV_X1 U53 ( .A(n68), .ZN(n32) );
  OAI221_X1 U54 ( .B1(n25), .B2(n63), .C1(n27), .C2(n69), .A(n70), .ZN(n68) );
  AOI22_X1 U55 ( .A1(A[25]), .A2(n4), .B1(A[26]), .B2(n2), .ZN(n70) );
  INV_X1 U56 ( .A(A[24]), .ZN(n63) );
  OAI221_X1 U57 ( .B1(n41), .B2(n57), .C1(n7), .C2(n5), .A(n71), .ZN(B[25]) );
  AOI222_X1 U58 ( .A1(n60), .A2(n46), .B1(n23), .B2(n44), .C1(n19), .C2(n72), 
        .ZN(n71) );
  AOI221_X1 U59 ( .B1(n73), .B2(n74), .C1(n75), .C2(n76), .A(n77), .ZN(n7) );
  INV_X1 U60 ( .A(n78), .ZN(n77) );
  AOI21_X1 U61 ( .B1(n79), .B2(n80), .A(n81), .ZN(n78) );
  INV_X1 U62 ( .A(n82), .ZN(n41) );
  OAI221_X1 U63 ( .B1(n25), .B2(n69), .C1(n27), .C2(n83), .A(n84), .ZN(n82) );
  AOI22_X1 U64 ( .A1(A[24]), .A2(n4), .B1(A[25]), .B2(n2), .ZN(n84) );
  INV_X1 U65 ( .A(A[23]), .ZN(n69) );
  OAI221_X1 U66 ( .B1(n49), .B2(n57), .C1(n9), .C2(n5), .A(n85), .ZN(B[24]) );
  AOI222_X1 U67 ( .A1(n60), .A2(n54), .B1(n23), .B2(n52), .C1(n19), .C2(n86), 
        .ZN(n85) );
  AOI221_X1 U68 ( .B1(n87), .B2(n74), .C1(n88), .C2(n76), .A(n89), .ZN(n9) );
  INV_X1 U69 ( .A(n90), .ZN(n49) );
  OAI221_X1 U70 ( .B1(n25), .B2(n83), .C1(n27), .C2(n91), .A(n92), .ZN(n90) );
  AOI22_X1 U71 ( .A1(A[23]), .A2(n4), .B1(A[24]), .B2(n2), .ZN(n92) );
  INV_X1 U72 ( .A(A[22]), .ZN(n83) );
  OAI221_X1 U73 ( .B1(n93), .B2(n57), .C1(n10), .C2(n5), .A(n94), .ZN(B[23])
         );
  AOI222_X1 U74 ( .A1(n60), .A2(n20), .B1(n23), .B2(n61), .C1(n19), .C2(n95), 
        .ZN(n94) );
  AOI221_X1 U75 ( .B1(n96), .B2(n74), .C1(n97), .C2(n76), .A(n89), .ZN(n10) );
  INV_X1 U76 ( .A(n24), .ZN(n93) );
  OAI221_X1 U77 ( .B1(n25), .B2(n91), .C1(n27), .C2(n98), .A(n99), .ZN(n24) );
  AOI22_X1 U78 ( .A1(A[22]), .A2(n4), .B1(A[23]), .B2(n2), .ZN(n99) );
  INV_X1 U79 ( .A(A[21]), .ZN(n91) );
  OAI221_X1 U80 ( .B1(n100), .B2(n57), .C1(n11), .C2(n5), .A(n101), .ZN(B[22])
         );
  AOI222_X1 U81 ( .A1(n60), .A2(n35), .B1(n23), .B2(n67), .C1(n19), .C2(n102), 
        .ZN(n101) );
  AOI221_X1 U82 ( .B1(n103), .B2(n74), .C1(n104), .C2(n76), .A(n89), .ZN(n11)
         );
  INV_X1 U83 ( .A(n37), .ZN(n100) );
  OAI221_X1 U84 ( .B1(n25), .B2(n98), .C1(n27), .C2(n105), .A(n106), .ZN(n37)
         );
  AOI22_X1 U85 ( .A1(A[21]), .A2(n4), .B1(A[22]), .B2(n2), .ZN(n106) );
  INV_X1 U86 ( .A(A[20]), .ZN(n98) );
  OAI221_X1 U87 ( .B1(n107), .B2(n57), .C1(n12), .C2(n6), .A(n108), .ZN(B[21])
         );
  AOI222_X1 U88 ( .A1(n60), .A2(n44), .B1(n23), .B2(n72), .C1(n19), .C2(n75), 
        .ZN(n108) );
  AOI221_X1 U89 ( .B1(n80), .B2(n74), .C1(n73), .C2(n76), .A(n89), .ZN(n12) );
  INV_X1 U90 ( .A(n109), .ZN(n89) );
  INV_X1 U91 ( .A(n46), .ZN(n107) );
  OAI221_X1 U92 ( .B1(n25), .B2(n105), .C1(n27), .C2(n110), .A(n111), .ZN(n46)
         );
  AOI22_X1 U93 ( .A1(A[20]), .A2(n4), .B1(A[21]), .B2(n2), .ZN(n111) );
  INV_X1 U94 ( .A(A[19]), .ZN(n105) );
  OAI221_X1 U95 ( .B1(n112), .B2(n57), .C1(n13), .C2(n6), .A(n113), .ZN(B[20])
         );
  AOI222_X1 U96 ( .A1(n60), .A2(n52), .B1(n23), .B2(n86), .C1(n19), .C2(n88), 
        .ZN(n113) );
  AOI21_X1 U97 ( .B1(n87), .B2(n76), .A(n114), .ZN(n13) );
  INV_X1 U98 ( .A(n54), .ZN(n112) );
  OAI221_X1 U99 ( .B1(n25), .B2(n110), .C1(n27), .C2(n115), .A(n116), .ZN(n54)
         );
  AOI22_X1 U100 ( .A1(A[19]), .A2(n4), .B1(A[20]), .B2(n2), .ZN(n116) );
  INV_X1 U101 ( .A(A[18]), .ZN(n110) );
  OAI21_X1 U102 ( .B1(SH[4]), .B2(n117), .A(n8), .ZN(B[1]) );
  OAI221_X1 U103 ( .B1(n118), .B2(n57), .C1(n14), .C2(n6), .A(n119), .ZN(B[19]) );
  AOI222_X1 U104 ( .A1(n60), .A2(n61), .B1(n23), .B2(n95), .C1(n19), .C2(n97), 
        .ZN(n119) );
  AOI21_X1 U105 ( .B1(n96), .B2(n76), .A(n114), .ZN(n14) );
  INV_X1 U106 ( .A(n20), .ZN(n118) );
  OAI221_X1 U107 ( .B1(n25), .B2(n115), .C1(n27), .C2(n120), .A(n121), .ZN(n20) );
  AOI22_X1 U108 ( .A1(A[18]), .A2(n4), .B1(A[19]), .B2(n2), .ZN(n121) );
  INV_X1 U109 ( .A(A[17]), .ZN(n115) );
  OAI221_X1 U110 ( .B1(n122), .B2(n57), .C1(n40), .C2(n6), .A(n123), .ZN(B[18]) );
  AOI222_X1 U111 ( .A1(n60), .A2(n67), .B1(n23), .B2(n102), .C1(n19), .C2(n104), .ZN(n123) );
  AOI21_X1 U112 ( .B1(n103), .B2(n76), .A(n114), .ZN(n40) );
  INV_X1 U113 ( .A(n35), .ZN(n122) );
  OAI221_X1 U114 ( .B1(n25), .B2(n120), .C1(n27), .C2(n124), .A(n125), .ZN(n35) );
  AOI22_X1 U115 ( .A1(A[17]), .A2(n4), .B1(A[18]), .B2(n2), .ZN(n125) );
  INV_X1 U116 ( .A(A[16]), .ZN(n120) );
  OAI221_X1 U117 ( .B1(n126), .B2(n57), .C1(n117), .C2(n6), .A(n127), .ZN(
        B[17]) );
  AOI222_X1 U118 ( .A1(n60), .A2(n72), .B1(n23), .B2(n75), .C1(n19), .C2(n73), 
        .ZN(n127) );
  INV_X1 U119 ( .A(n16), .ZN(n60) );
  AOI21_X1 U120 ( .B1(n80), .B2(n76), .A(n114), .ZN(n117) );
  OAI21_X1 U121 ( .B1(n128), .B2(n129), .A(n109), .ZN(n114) );
  INV_X1 U122 ( .A(n44), .ZN(n126) );
  OAI221_X1 U123 ( .B1(n25), .B2(n124), .C1(n27), .C2(n130), .A(n131), .ZN(n44) );
  AOI22_X1 U124 ( .A1(A[16]), .A2(n4), .B1(A[17]), .B2(n2), .ZN(n131) );
  INV_X1 U125 ( .A(A[15]), .ZN(n124) );
  OAI221_X1 U126 ( .B1(n132), .B2(n16), .C1(n133), .C2(n57), .A(n134), .ZN(
        B[16]) );
  AOI221_X1 U127 ( .B1(n19), .B2(n87), .C1(n23), .C2(n88), .A(n135), .ZN(n134)
         );
  INV_X1 U128 ( .A(n8), .ZN(n135) );
  AND2_X1 U129 ( .A1(n136), .A2(n129), .ZN(n23) );
  AND2_X1 U130 ( .A1(n136), .A2(SH[2]), .ZN(n19) );
  AND2_X1 U131 ( .A1(SH[3]), .A2(n6), .ZN(n136) );
  NAND2_X1 U132 ( .A1(n76), .A2(n5), .ZN(n57) );
  INV_X1 U133 ( .A(n52), .ZN(n133) );
  OAI221_X1 U134 ( .B1(n25), .B2(n130), .C1(n27), .C2(n137), .A(n138), .ZN(n52) );
  AOI22_X1 U135 ( .A1(A[15]), .A2(n4), .B1(A[16]), .B2(n2), .ZN(n138) );
  INV_X1 U136 ( .A(A[14]), .ZN(n130) );
  NAND2_X1 U137 ( .A1(n74), .A2(n5), .ZN(n16) );
  INV_X1 U138 ( .A(n86), .ZN(n132) );
  OAI21_X1 U139 ( .B1(SH[4]), .B2(n17), .A(n8), .ZN(B[15]) );
  AOI221_X1 U140 ( .B1(n95), .B2(n74), .C1(n61), .C2(n76), .A(n139), .ZN(n17)
         );
  INV_X1 U141 ( .A(n140), .ZN(n139) );
  AOI22_X1 U142 ( .A1(n141), .A2(n96), .B1(n79), .B2(n97), .ZN(n140) );
  OAI221_X1 U143 ( .B1(n25), .B2(n137), .C1(n27), .C2(n142), .A(n143), .ZN(n61) );
  AOI22_X1 U144 ( .A1(A[14]), .A2(n4), .B1(A[15]), .B2(n2), .ZN(n143) );
  INV_X1 U145 ( .A(A[13]), .ZN(n137) );
  OAI21_X1 U146 ( .B1(SH[4]), .B2(n33), .A(n8), .ZN(B[14]) );
  AOI221_X1 U147 ( .B1(n102), .B2(n74), .C1(n67), .C2(n76), .A(n144), .ZN(n33)
         );
  INV_X1 U148 ( .A(n145), .ZN(n144) );
  AOI22_X1 U149 ( .A1(n141), .A2(n103), .B1(n79), .B2(n104), .ZN(n145) );
  OAI221_X1 U150 ( .B1(n25), .B2(n142), .C1(n27), .C2(n146), .A(n147), .ZN(n67) );
  AOI22_X1 U151 ( .A1(A[13]), .A2(n4), .B1(A[14]), .B2(n2), .ZN(n147) );
  INV_X1 U152 ( .A(A[12]), .ZN(n142) );
  OAI21_X1 U153 ( .B1(SH[4]), .B2(n42), .A(n8), .ZN(B[13]) );
  AOI221_X1 U154 ( .B1(n80), .B2(n141), .C1(n73), .C2(n79), .A(n148), .ZN(n42)
         );
  INV_X1 U155 ( .A(n149), .ZN(n148) );
  AOI22_X1 U156 ( .A1(n74), .A2(n75), .B1(n76), .B2(n72), .ZN(n149) );
  OAI221_X1 U157 ( .B1(n25), .B2(n146), .C1(n27), .C2(n150), .A(n151), .ZN(n72) );
  AOI22_X1 U158 ( .A1(A[12]), .A2(n4), .B1(A[13]), .B2(n2), .ZN(n151) );
  INV_X1 U159 ( .A(A[11]), .ZN(n146) );
  OAI221_X1 U160 ( .B1(n25), .B2(n152), .C1(n27), .C2(n153), .A(n154), .ZN(n75) );
  AOI22_X1 U161 ( .A1(A[8]), .A2(n4), .B1(A[9]), .B2(n2), .ZN(n154) );
  OAI221_X1 U162 ( .B1(n25), .B2(n155), .C1(n27), .C2(n156), .A(n157), .ZN(n73) );
  AOI22_X1 U163 ( .A1(A[4]), .A2(n4), .B1(A[5]), .B2(n2), .ZN(n157) );
  AND2_X1 U164 ( .A1(SH[2]), .A2(SH[3]), .ZN(n141) );
  MUX2_X1 U165 ( .A(\A[0] ), .B(A[1]), .S(n2), .Z(n80) );
  OAI21_X1 U166 ( .B1(SH[4]), .B2(n50), .A(n8), .ZN(B[12]) );
  AOI221_X1 U167 ( .B1(n88), .B2(n74), .C1(n86), .C2(n76), .A(n158), .ZN(n50)
         );
  INV_X1 U168 ( .A(n159), .ZN(n158) );
  AOI21_X1 U169 ( .B1(n79), .B2(n87), .A(n81), .ZN(n159) );
  OAI221_X1 U170 ( .B1(n25), .B2(n156), .C1(n160), .C2(n27), .A(n161), .ZN(n87) );
  AOI22_X1 U171 ( .A1(n4), .A2(A[3]), .B1(A[4]), .B2(n2), .ZN(n161) );
  INV_X1 U172 ( .A(A[2]), .ZN(n156) );
  AOI22_X1 U173 ( .A1(A[11]), .A2(n4), .B1(A[12]), .B2(n2), .ZN(n163) );
  INV_X1 U174 ( .A(A[10]), .ZN(n150) );
  AOI22_X1 U175 ( .A1(A[7]), .A2(n4), .B1(A[8]), .B2(n2), .ZN(n165) );
  INV_X1 U176 ( .A(A[6]), .ZN(n153) );
  OAI21_X1 U177 ( .B1(SH[4]), .B2(n58), .A(n8), .ZN(B[11]) );
  AOI221_X1 U178 ( .B1(n97), .B2(n74), .C1(n95), .C2(n76), .A(n166), .ZN(n58)
         );
  INV_X1 U179 ( .A(n167), .ZN(n166) );
  AOI21_X1 U180 ( .B1(n79), .B2(n96), .A(n81), .ZN(n167) );
  OAI221_X1 U181 ( .B1(n160), .B2(n25), .C1(n128), .C2(n27), .A(n168), .ZN(n96) );
  AOI22_X1 U182 ( .A1(n4), .A2(A[2]), .B1(A[3]), .B2(n2), .ZN(n168) );
  INV_X1 U183 ( .A(\A[0] ), .ZN(n128) );
  INV_X1 U184 ( .A(A[1]), .ZN(n160) );
  AOI22_X1 U185 ( .A1(A[10]), .A2(n4), .B1(A[11]), .B2(n2), .ZN(n170) );
  INV_X1 U186 ( .A(A[9]), .ZN(n162) );
  AOI22_X1 U187 ( .A1(A[6]), .A2(n4), .B1(A[7]), .B2(n2), .ZN(n172) );
  INV_X1 U188 ( .A(A[5]), .ZN(n164) );
  OAI21_X1 U189 ( .B1(SH[4]), .B2(n65), .A(n8), .ZN(B[10]) );
  NAND2_X1 U190 ( .A1(SH[4]), .A2(\A[0] ), .ZN(n8) );
  AOI221_X1 U191 ( .B1(n104), .B2(n74), .C1(n102), .C2(n76), .A(n173), .ZN(n65) );
  INV_X1 U192 ( .A(n174), .ZN(n173) );
  AOI21_X1 U193 ( .B1(n79), .B2(n103), .A(n81), .ZN(n174) );
  NOR2_X1 U194 ( .A1(n129), .A2(n109), .ZN(n81) );
  NAND2_X1 U195 ( .A1(SH[3]), .A2(\A[0] ), .ZN(n109) );
  INV_X1 U196 ( .A(n175), .ZN(n103) );
  AOI222_X1 U197 ( .A1(n2), .A2(A[2]), .B1(A[1]), .B2(n4), .C1(\A[0] ), .C2(
        SH[1]), .ZN(n175) );
  AND2_X1 U198 ( .A1(SH[3]), .A2(n129), .ZN(n79) );
  AOI22_X1 U199 ( .A1(A[9]), .A2(n4), .B1(A[10]), .B2(n2), .ZN(n176) );
  INV_X1 U200 ( .A(A[7]), .ZN(n152) );
  INV_X1 U201 ( .A(A[8]), .ZN(n169) );
  NOR2_X1 U202 ( .A1(n129), .A2(SH[3]), .ZN(n74) );
  INV_X1 U203 ( .A(SH[2]), .ZN(n129) );
  OAI221_X1 U204 ( .B1(n25), .B2(n171), .C1(n155), .C2(n27), .A(n177), .ZN(
        n104) );
  AOI22_X1 U205 ( .A1(A[5]), .A2(n4), .B1(A[6]), .B2(n2), .ZN(n177) );
  NOR2_X1 U206 ( .A1(SH[0]), .A2(SH[1]), .ZN(n31) );
  NOR2_X1 U207 ( .A1(n178), .A2(SH[1]), .ZN(n30) );
  INV_X1 U208 ( .A(A[3]), .ZN(n155) );
  INV_X1 U209 ( .A(A[4]), .ZN(n171) );
  INV_X1 U210 ( .A(SH[0]), .ZN(n178) );
endmodule


module SHIFTER_GENERIC_N32_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163;

  NOR2_X2 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n51) );
  NOR2_X2 U4 ( .A1(n163), .A2(SH[1]), .ZN(n50) );
  INV_X1 U5 ( .A(SH[4]), .ZN(n1) );
  INV_X1 U6 ( .A(SH[4]), .ZN(n2) );
  OAI221_X1 U7 ( .B1(n3), .B2(n4), .C1(n5), .C2(n1), .A(n6), .ZN(B[9]) );
  AOI222_X1 U8 ( .A1(n7), .A2(n8), .B1(n9), .B2(n10), .C1(n11), .C2(n12), .ZN(
        n6) );
  OAI221_X1 U9 ( .B1(n13), .B2(n4), .C1(n14), .C2(n1), .A(n15), .ZN(B[8]) );
  AOI222_X1 U10 ( .A1(n7), .A2(n16), .B1(n9), .B2(n17), .C1(n11), .C2(n18), 
        .ZN(n15) );
  OAI221_X1 U11 ( .B1(n19), .B2(n4), .C1(n20), .C2(n1), .A(n21), .ZN(B[7]) );
  AOI222_X1 U12 ( .A1(n7), .A2(n22), .B1(n9), .B2(n23), .C1(n11), .C2(n24), 
        .ZN(n21) );
  OAI221_X1 U13 ( .B1(n25), .B2(n4), .C1(n26), .C2(n1), .A(n27), .ZN(B[6]) );
  AOI222_X1 U14 ( .A1(n7), .A2(n28), .B1(n9), .B2(n29), .C1(n11), .C2(n30), 
        .ZN(n27) );
  OAI221_X1 U15 ( .B1(n31), .B2(n4), .C1(n32), .C2(n1), .A(n33), .ZN(B[5]) );
  AOI222_X1 U16 ( .A1(n7), .A2(n34), .B1(n9), .B2(n8), .C1(n11), .C2(n10), 
        .ZN(n33) );
  OAI221_X1 U17 ( .B1(n35), .B2(n4), .C1(n36), .C2(n1), .A(n37), .ZN(B[4]) );
  AOI222_X1 U18 ( .A1(n7), .A2(n38), .B1(n9), .B2(n16), .C1(n11), .C2(n17), 
        .ZN(n37) );
  OAI221_X1 U19 ( .B1(n19), .B2(n39), .C1(n40), .C2(n1), .A(n41), .ZN(B[3]) );
  AOI222_X1 U20 ( .A1(n11), .A2(n23), .B1(n42), .B2(n43), .C1(n9), .C2(n22), 
        .ZN(n41) );
  INV_X1 U21 ( .A(n44), .ZN(n22) );
  OAI221_X1 U22 ( .B1(n45), .B2(n46), .C1(n47), .C2(n48), .A(n49), .ZN(n43) );
  AOI22_X1 U23 ( .A1(A[4]), .A2(n50), .B1(A[3]), .B2(n51), .ZN(n49) );
  AOI221_X1 U24 ( .B1(n52), .B2(A[10]), .C1(n53), .C2(A[9]), .A(n54), .ZN(n19)
         );
  OAI22_X1 U25 ( .A1(n55), .A2(n56), .B1(n57), .B2(n58), .ZN(n54) );
  AND2_X1 U26 ( .A1(n42), .A2(n59), .ZN(B[31]) );
  AND2_X1 U27 ( .A1(n60), .A2(n42), .ZN(B[30]) );
  OAI221_X1 U28 ( .B1(n25), .B2(n39), .C1(n61), .C2(n2), .A(n62), .ZN(B[2]) );
  AOI222_X1 U29 ( .A1(n11), .A2(n29), .B1(n42), .B2(n63), .C1(n9), .C2(n28), 
        .ZN(n62) );
  INV_X1 U30 ( .A(n64), .ZN(n28) );
  OAI221_X1 U31 ( .B1(n45), .B2(n48), .C1(n47), .C2(n65), .A(n66), .ZN(n63) );
  AOI22_X1 U32 ( .A1(A[3]), .A2(n50), .B1(A[2]), .B2(n51), .ZN(n66) );
  AOI221_X1 U33 ( .B1(n52), .B2(A[9]), .C1(n53), .C2(A[8]), .A(n67), .ZN(n25)
         );
  OAI22_X1 U34 ( .A1(n57), .A2(n56), .B1(n46), .B2(n58), .ZN(n67) );
  INV_X1 U35 ( .A(A[7]), .ZN(n57) );
  AND2_X1 U36 ( .A1(n68), .A2(n42), .ZN(B[29]) );
  AND2_X1 U37 ( .A1(n69), .A2(n42), .ZN(B[28]) );
  NOR3_X1 U38 ( .A1(n70), .A2(SH[4]), .A3(SH[3]), .ZN(B[27]) );
  NOR2_X1 U39 ( .A1(SH[4]), .A2(n71), .ZN(B[26]) );
  NOR2_X1 U40 ( .A1(SH[4]), .A2(n5), .ZN(B[25]) );
  AOI22_X1 U41 ( .A1(n72), .A2(n73), .B1(n68), .B2(n74), .ZN(n5) );
  NOR2_X1 U42 ( .A1(SH[4]), .A2(n14), .ZN(B[24]) );
  AOI22_X1 U43 ( .A1(n75), .A2(n73), .B1(n69), .B2(n74), .ZN(n14) );
  NOR2_X1 U44 ( .A1(SH[4]), .A2(n20), .ZN(B[23]) );
  AOI222_X1 U45 ( .A1(n76), .A2(n74), .B1(n59), .B2(n77), .C1(n78), .C2(n73), 
        .ZN(n20) );
  NOR2_X1 U46 ( .A1(SH[4]), .A2(n26), .ZN(B[22]) );
  AOI222_X1 U47 ( .A1(n79), .A2(n74), .B1(n60), .B2(n77), .C1(n80), .C2(n73), 
        .ZN(n26) );
  NOR2_X1 U48 ( .A1(SH[4]), .A2(n32), .ZN(B[21]) );
  AOI222_X1 U49 ( .A1(n72), .A2(n74), .B1(n68), .B2(n77), .C1(n12), .C2(n73), 
        .ZN(n32) );
  NOR2_X1 U50 ( .A1(SH[4]), .A2(n36), .ZN(B[20]) );
  AOI222_X1 U51 ( .A1(n75), .A2(n74), .B1(n69), .B2(n77), .C1(n18), .C2(n73), 
        .ZN(n36) );
  OAI221_X1 U52 ( .B1(n31), .B2(n39), .C1(n81), .C2(n2), .A(n82), .ZN(B[1]) );
  AOI222_X1 U53 ( .A1(n11), .A2(n8), .B1(n42), .B2(n83), .C1(n9), .C2(n34), 
        .ZN(n82) );
  INV_X1 U54 ( .A(n3), .ZN(n34) );
  AOI221_X1 U55 ( .B1(n52), .B2(A[12]), .C1(n53), .C2(A[11]), .A(n84), .ZN(n3)
         );
  OAI22_X1 U56 ( .A1(n85), .A2(n56), .B1(n86), .B2(n58), .ZN(n84) );
  OAI221_X1 U57 ( .B1(n45), .B2(n65), .C1(n47), .C2(n87), .A(n88), .ZN(n83) );
  AOI22_X1 U58 ( .A1(A[2]), .A2(n50), .B1(A[1]), .B2(n51), .ZN(n88) );
  AOI221_X1 U59 ( .B1(n52), .B2(A[8]), .C1(n53), .C2(A[7]), .A(n89), .ZN(n31)
         );
  OAI22_X1 U60 ( .A1(n46), .A2(n56), .B1(n48), .B2(n58), .ZN(n89) );
  INV_X1 U61 ( .A(A[6]), .ZN(n46) );
  NOR2_X1 U62 ( .A1(SH[4]), .A2(n40), .ZN(B[19]) );
  AOI222_X1 U63 ( .A1(n24), .A2(n73), .B1(n78), .B2(n74), .C1(n90), .C2(SH[3]), 
        .ZN(n40) );
  NOR2_X1 U64 ( .A1(SH[4]), .A2(n61), .ZN(B[18]) );
  AOI221_X1 U65 ( .B1(n80), .B2(n74), .C1(n30), .C2(n73), .A(n91), .ZN(n61) );
  INV_X1 U66 ( .A(n92), .ZN(n91) );
  AOI22_X1 U67 ( .A1(n93), .A2(n60), .B1(n77), .B2(n79), .ZN(n92) );
  NOR2_X1 U68 ( .A1(SH[4]), .A2(n81), .ZN(B[17]) );
  AOI221_X1 U69 ( .B1(n12), .B2(n74), .C1(n10), .C2(n73), .A(n94), .ZN(n81) );
  INV_X1 U70 ( .A(n95), .ZN(n94) );
  AOI22_X1 U71 ( .A1(n93), .A2(n68), .B1(n77), .B2(n72), .ZN(n95) );
  NOR2_X1 U72 ( .A1(SH[4]), .A2(n96), .ZN(B[16]) );
  OAI221_X1 U73 ( .B1(n97), .B2(n39), .C1(n98), .C2(n4), .A(n99), .ZN(B[15])
         );
  AOI222_X1 U74 ( .A1(n11), .A2(n76), .B1(n100), .B2(n59), .C1(n9), .C2(n78), 
        .ZN(n99) );
  INV_X1 U75 ( .A(n24), .ZN(n97) );
  OAI221_X1 U76 ( .B1(n101), .B2(n39), .C1(n102), .C2(n4), .A(n103), .ZN(B[14]) );
  AOI222_X1 U77 ( .A1(n11), .A2(n79), .B1(n100), .B2(n60), .C1(n9), .C2(n80), 
        .ZN(n103) );
  INV_X1 U78 ( .A(n29), .ZN(n102) );
  INV_X1 U79 ( .A(n30), .ZN(n101) );
  OAI221_X1 U80 ( .B1(n104), .B2(n39), .C1(n105), .C2(n4), .A(n106), .ZN(B[13]) );
  AOI222_X1 U81 ( .A1(n11), .A2(n72), .B1(n100), .B2(n68), .C1(n9), .C2(n12), 
        .ZN(n106) );
  OAI221_X1 U82 ( .B1(n45), .B2(n107), .C1(n47), .C2(n108), .A(n109), .ZN(n12)
         );
  AOI22_X1 U83 ( .A1(A[22]), .A2(n50), .B1(A[21]), .B2(n51), .ZN(n109) );
  INV_X1 U84 ( .A(A[23]), .ZN(n108) );
  OAI222_X1 U85 ( .A1(n56), .A2(n110), .B1(n47), .B2(n111), .C1(n58), .C2(n112), .ZN(n68) );
  OAI221_X1 U86 ( .B1(n45), .B2(n113), .C1(n47), .C2(n114), .A(n115), .ZN(n72)
         );
  AOI22_X1 U87 ( .A1(A[26]), .A2(n50), .B1(A[25]), .B2(n51), .ZN(n115) );
  INV_X1 U88 ( .A(n8), .ZN(n105) );
  OAI221_X1 U89 ( .B1(n45), .B2(n116), .C1(n47), .C2(n117), .A(n118), .ZN(n8)
         );
  AOI22_X1 U90 ( .A1(A[14]), .A2(n50), .B1(A[13]), .B2(n51), .ZN(n118) );
  INV_X1 U91 ( .A(n10), .ZN(n104) );
  OAI221_X1 U92 ( .B1(n45), .B2(n119), .C1(n47), .C2(n120), .A(n121), .ZN(n10)
         );
  AOI22_X1 U93 ( .A1(A[18]), .A2(n50), .B1(A[17]), .B2(n51), .ZN(n121) );
  INV_X1 U94 ( .A(n122), .ZN(B[12]) );
  AOI221_X1 U95 ( .B1(n17), .B2(n7), .C1(n16), .C2(n42), .A(n123), .ZN(n122)
         );
  INV_X1 U96 ( .A(n124), .ZN(n123) );
  AOI222_X1 U97 ( .A1(n11), .A2(n75), .B1(n100), .B2(n69), .C1(n9), .C2(n18), 
        .ZN(n124) );
  NOR2_X1 U98 ( .A1(n1), .A2(n125), .ZN(n100) );
  OAI221_X1 U99 ( .B1(n98), .B2(n39), .C1(n44), .C2(n4), .A(n126), .ZN(B[11])
         );
  AOI221_X1 U100 ( .B1(n11), .B2(n78), .C1(n9), .C2(n24), .A(n127), .ZN(n126)
         );
  NOR3_X1 U101 ( .A1(n1), .A2(SH[3]), .A3(n70), .ZN(n127) );
  INV_X1 U102 ( .A(n90), .ZN(n70) );
  MUX2_X1 U103 ( .A(n76), .B(n59), .S(SH[2]), .Z(n90) );
  NOR2_X1 U104 ( .A1(n111), .A2(n58), .ZN(n59) );
  OAI221_X1 U105 ( .B1(n45), .B2(n110), .C1(n47), .C2(n112), .A(n128), .ZN(n76) );
  AOI22_X1 U106 ( .A1(A[28]), .A2(n50), .B1(A[27]), .B2(n51), .ZN(n128) );
  OAI221_X1 U107 ( .B1(n119), .B2(n56), .C1(n120), .C2(n58), .A(n129), .ZN(n24) );
  AOI22_X1 U108 ( .A1(A[22]), .A2(n52), .B1(A[21]), .B2(n53), .ZN(n129) );
  OAI221_X1 U109 ( .B1(n45), .B2(n130), .C1(n47), .C2(n131), .A(n132), .ZN(n78) );
  AOI22_X1 U110 ( .A1(A[24]), .A2(n50), .B1(A[23]), .B2(n51), .ZN(n132) );
  AOI221_X1 U111 ( .B1(n52), .B2(A[14]), .C1(n53), .C2(A[13]), .A(n133), .ZN(
        n44) );
  OAI22_X1 U112 ( .A1(n134), .A2(n56), .B1(n135), .B2(n58), .ZN(n133) );
  INV_X1 U113 ( .A(A[12]), .ZN(n134) );
  INV_X1 U114 ( .A(n23), .ZN(n98) );
  OAI221_X1 U115 ( .B1(n45), .B2(n136), .C1(n47), .C2(n137), .A(n138), .ZN(n23) );
  AOI22_X1 U116 ( .A1(A[16]), .A2(n50), .B1(A[15]), .B2(n51), .ZN(n138) );
  OAI221_X1 U117 ( .B1(n64), .B2(n4), .C1(n71), .C2(n2), .A(n139), .ZN(B[10])
         );
  AOI222_X1 U118 ( .A1(n7), .A2(n29), .B1(n9), .B2(n30), .C1(n11), .C2(n80), 
        .ZN(n139) );
  OAI221_X1 U119 ( .B1(n45), .B2(n131), .C1(n47), .C2(n107), .A(n140), .ZN(n80) );
  AOI22_X1 U120 ( .A1(A[23]), .A2(n50), .B1(A[22]), .B2(n51), .ZN(n140) );
  INV_X1 U121 ( .A(A[24]), .ZN(n107) );
  INV_X1 U122 ( .A(A[25]), .ZN(n131) );
  OAI221_X1 U123 ( .B1(n45), .B2(n141), .C1(n119), .C2(n47), .A(n142), .ZN(n30) );
  AOI22_X1 U124 ( .A1(n50), .A2(A[19]), .B1(n51), .B2(A[18]), .ZN(n142) );
  OAI221_X1 U125 ( .B1(n45), .B2(n137), .C1(n47), .C2(n116), .A(n143), .ZN(n29) );
  AOI22_X1 U126 ( .A1(A[15]), .A2(n50), .B1(A[14]), .B2(n51), .ZN(n143) );
  INV_X1 U127 ( .A(A[16]), .ZN(n116) );
  INV_X1 U128 ( .A(A[17]), .ZN(n137) );
  INV_X1 U129 ( .A(n39), .ZN(n7) );
  AOI22_X1 U130 ( .A1(n79), .A2(n73), .B1(n60), .B2(n74), .ZN(n71) );
  OAI22_X1 U131 ( .A1(n58), .A2(n110), .B1(n56), .B2(n111), .ZN(n60) );
  OAI221_X1 U132 ( .B1(n45), .B2(n112), .C1(n47), .C2(n113), .A(n144), .ZN(n79) );
  AOI22_X1 U133 ( .A1(A[27]), .A2(n50), .B1(A[26]), .B2(n51), .ZN(n144) );
  INV_X1 U134 ( .A(A[28]), .ZN(n113) );
  INV_X1 U135 ( .A(A[29]), .ZN(n112) );
  AOI221_X1 U136 ( .B1(n52), .B2(A[13]), .C1(n53), .C2(A[12]), .A(n145), .ZN(
        n64) );
  OAI22_X1 U137 ( .A1(n135), .A2(n56), .B1(n85), .B2(n58), .ZN(n145) );
  INV_X1 U138 ( .A(A[10]), .ZN(n85) );
  INV_X1 U139 ( .A(A[11]), .ZN(n135) );
  OAI221_X1 U140 ( .B1(n35), .B2(n39), .C1(n96), .C2(n1), .A(n146), .ZN(B[0])
         );
  AOI222_X1 U141 ( .A1(n11), .A2(n16), .B1(n42), .B2(n147), .C1(n9), .C2(n38), 
        .ZN(n146) );
  INV_X1 U142 ( .A(n13), .ZN(n38) );
  AOI221_X1 U143 ( .B1(n52), .B2(A[11]), .C1(n53), .C2(A[10]), .A(n148), .ZN(
        n13) );
  OAI22_X1 U144 ( .A1(n86), .A2(n56), .B1(n55), .B2(n58), .ZN(n148) );
  INV_X1 U145 ( .A(A[8]), .ZN(n55) );
  INV_X1 U146 ( .A(A[9]), .ZN(n86) );
  AND2_X1 U147 ( .A1(n149), .A2(n150), .ZN(n9) );
  OAI221_X1 U148 ( .B1(n45), .B2(n87), .C1(n47), .C2(n151), .A(n152), .ZN(n147) );
  AOI22_X1 U149 ( .A1(A[1]), .A2(n50), .B1(A[0]), .B2(n51), .ZN(n152) );
  INV_X1 U150 ( .A(A[2]), .ZN(n151) );
  INV_X1 U151 ( .A(A[3]), .ZN(n87) );
  INV_X1 U152 ( .A(n4), .ZN(n42) );
  NAND2_X1 U153 ( .A1(n73), .A2(n1), .ZN(n4) );
  OAI221_X1 U154 ( .B1(n45), .B2(n117), .C1(n47), .C2(n153), .A(n154), .ZN(n16) );
  AOI22_X1 U155 ( .A1(A[13]), .A2(n50), .B1(A[12]), .B2(n51), .ZN(n154) );
  INV_X1 U156 ( .A(A[14]), .ZN(n153) );
  INV_X1 U157 ( .A(A[15]), .ZN(n117) );
  AND2_X1 U158 ( .A1(SH[2]), .A2(n149), .ZN(n11) );
  NOR2_X1 U159 ( .A1(n155), .A2(SH[4]), .ZN(n149) );
  AOI221_X1 U160 ( .B1(n18), .B2(n74), .C1(n17), .C2(n73), .A(n156), .ZN(n96)
         );
  INV_X1 U161 ( .A(n157), .ZN(n156) );
  AOI22_X1 U162 ( .A1(n93), .A2(n69), .B1(n77), .B2(n75), .ZN(n157) );
  OAI221_X1 U163 ( .B1(n45), .B2(n114), .C1(n47), .C2(n130), .A(n158), .ZN(n75) );
  AOI22_X1 U164 ( .A1(A[25]), .A2(n50), .B1(A[24]), .B2(n51), .ZN(n158) );
  INV_X1 U165 ( .A(A[26]), .ZN(n130) );
  INV_X1 U166 ( .A(A[27]), .ZN(n114) );
  NOR2_X1 U167 ( .A1(n155), .A2(SH[2]), .ZN(n77) );
  OAI221_X1 U168 ( .B1(n45), .B2(n111), .C1(n47), .C2(n110), .A(n159), .ZN(n69) );
  AOI22_X1 U169 ( .A1(A[29]), .A2(n50), .B1(A[28]), .B2(n51), .ZN(n159) );
  INV_X1 U170 ( .A(A[30]), .ZN(n110) );
  INV_X1 U171 ( .A(A[31]), .ZN(n111) );
  NOR2_X1 U172 ( .A1(n150), .A2(n155), .ZN(n93) );
  INV_X1 U173 ( .A(n125), .ZN(n73) );
  NAND2_X1 U174 ( .A1(n150), .A2(n155), .ZN(n125) );
  INV_X1 U175 ( .A(SH[3]), .ZN(n155) );
  OAI221_X1 U176 ( .B1(n45), .B2(n120), .C1(n47), .C2(n136), .A(n160), .ZN(n17) );
  AOI22_X1 U177 ( .A1(A[17]), .A2(n50), .B1(A[16]), .B2(n51), .ZN(n160) );
  INV_X1 U178 ( .A(A[18]), .ZN(n136) );
  INV_X1 U179 ( .A(A[19]), .ZN(n120) );
  OAI221_X1 U180 ( .B1(n56), .B2(n141), .C1(n119), .C2(n58), .A(n161), .ZN(n18) );
  AOI22_X1 U181 ( .A1(A[23]), .A2(n52), .B1(A[22]), .B2(n53), .ZN(n161) );
  INV_X1 U182 ( .A(A[20]), .ZN(n119) );
  INV_X1 U183 ( .A(A[21]), .ZN(n141) );
  NAND2_X1 U184 ( .A1(n74), .A2(n1), .ZN(n39) );
  NOR2_X1 U185 ( .A1(n150), .A2(SH[3]), .ZN(n74) );
  INV_X1 U186 ( .A(SH[2]), .ZN(n150) );
  AOI221_X1 U187 ( .B1(n52), .B2(A[7]), .C1(n53), .C2(A[6]), .A(n162), .ZN(n35) );
  OAI22_X1 U188 ( .A1(n48), .A2(n56), .B1(n65), .B2(n58), .ZN(n162) );
  INV_X1 U189 ( .A(n51), .ZN(n58) );
  INV_X1 U190 ( .A(A[4]), .ZN(n65) );
  INV_X1 U191 ( .A(n50), .ZN(n56) );
  INV_X1 U192 ( .A(A[5]), .ZN(n48) );
  INV_X1 U193 ( .A(n47), .ZN(n53) );
  NAND2_X1 U194 ( .A1(SH[1]), .A2(n163), .ZN(n47) );
  INV_X1 U195 ( .A(SH[0]), .ZN(n163) );
  INV_X1 U196 ( .A(n45), .ZN(n52) );
  NAND2_X1 U197 ( .A1(SH[1]), .A2(SH[0]), .ZN(n45) );
endmodule


module SHIFTER_GENERIC_N32_DW_sra_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  NOR2_X2 U2 ( .A1(n131), .A2(SH[0]), .ZN(n52) );
  AOI221_X4 U3 ( .B1(n52), .B2(A[6]), .C1(n53), .C2(A[7]), .A(n171), .ZN(n35)
         );
  AOI221_X4 U4 ( .B1(n52), .B2(A[14]), .C1(n53), .C2(A[15]), .A(n162), .ZN(
        n135) );
  AOI221_X4 U5 ( .B1(n52), .B2(A[10]), .C1(n53), .C2(A[11]), .A(n158), .ZN(n13) );
  AOI221_X4 U6 ( .B1(n52), .B2(A[12]), .C1(n53), .C2(A[13]), .A(n155), .ZN(n64) );
  AOI221_X4 U7 ( .B1(n52), .B2(A[16]), .C1(n53), .C2(A[17]), .A(n152), .ZN(
        n116) );
  NOR2_X2 U8 ( .A1(n172), .A2(n131), .ZN(n53) );
  NOR2_X2 U9 ( .A1(SH[2]), .A2(SH[3]), .ZN(n75) );
  INV_X1 U10 ( .A(SH[4]), .ZN(n1) );
  INV_X1 U11 ( .A(SH[4]), .ZN(n2) );
  OAI221_X1 U12 ( .B1(n3), .B2(n4), .C1(n5), .C2(n1), .A(n6), .ZN(B[9]) );
  AOI222_X1 U13 ( .A1(n7), .A2(n8), .B1(n9), .B2(n10), .C1(n11), .C2(n12), 
        .ZN(n6) );
  OAI221_X1 U14 ( .B1(n13), .B2(n4), .C1(n14), .C2(n1), .A(n15), .ZN(B[8]) );
  AOI222_X1 U15 ( .A1(n7), .A2(n16), .B1(n9), .B2(n17), .C1(n11), .C2(n18), 
        .ZN(n15) );
  OAI221_X1 U16 ( .B1(n19), .B2(n4), .C1(n20), .C2(n1), .A(n21), .ZN(B[7]) );
  AOI222_X1 U17 ( .A1(n7), .A2(n22), .B1(n9), .B2(n23), .C1(n11), .C2(n24), 
        .ZN(n21) );
  OAI221_X1 U18 ( .B1(n25), .B2(n4), .C1(n26), .C2(n1), .A(n27), .ZN(B[6]) );
  AOI222_X1 U19 ( .A1(n7), .A2(n28), .B1(n9), .B2(n29), .C1(n11), .C2(n30), 
        .ZN(n27) );
  OAI221_X1 U20 ( .B1(n31), .B2(n4), .C1(n32), .C2(n1), .A(n33), .ZN(B[5]) );
  AOI222_X1 U21 ( .A1(n7), .A2(n34), .B1(n9), .B2(n8), .C1(n11), .C2(n10), 
        .ZN(n33) );
  OAI221_X1 U22 ( .B1(n35), .B2(n4), .C1(n36), .C2(n1), .A(n37), .ZN(B[4]) );
  AOI222_X1 U23 ( .A1(n7), .A2(n38), .B1(n9), .B2(n16), .C1(n11), .C2(n17), 
        .ZN(n37) );
  OAI221_X1 U24 ( .B1(n19), .B2(n39), .C1(n40), .C2(n1), .A(n41), .ZN(B[3]) );
  AOI222_X1 U25 ( .A1(n11), .A2(n23), .B1(n42), .B2(n43), .C1(n9), .C2(n22), 
        .ZN(n41) );
  INV_X1 U26 ( .A(n44), .ZN(n22) );
  OAI221_X1 U27 ( .B1(n45), .B2(n46), .C1(n47), .C2(n48), .A(n49), .ZN(n43) );
  AOI22_X1 U28 ( .A1(A[4]), .A2(n50), .B1(A[3]), .B2(n51), .ZN(n49) );
  AOI221_X1 U29 ( .B1(n52), .B2(A[9]), .C1(n53), .C2(A[10]), .A(n54), .ZN(n19)
         );
  OAI22_X1 U30 ( .A1(n55), .A2(n56), .B1(n57), .B2(n58), .ZN(n54) );
  OAI21_X1 U31 ( .B1(SH[4]), .B2(n59), .A(n60), .ZN(B[30]) );
  OAI221_X1 U32 ( .B1(n25), .B2(n39), .C1(n61), .C2(n1), .A(n62), .ZN(B[2]) );
  AOI222_X1 U33 ( .A1(n11), .A2(n29), .B1(n42), .B2(n63), .C1(n9), .C2(n28), 
        .ZN(n62) );
  INV_X1 U34 ( .A(n64), .ZN(n28) );
  OAI221_X1 U35 ( .B1(n45), .B2(n65), .C1(n47), .C2(n46), .A(n66), .ZN(n63) );
  AOI22_X1 U36 ( .A1(A[3]), .A2(n50), .B1(A[2]), .B2(n51), .ZN(n66) );
  AOI221_X1 U37 ( .B1(n52), .B2(A[8]), .C1(n53), .C2(A[9]), .A(n67), .ZN(n25)
         );
  OAI22_X1 U38 ( .A1(n57), .A2(n56), .B1(n48), .B2(n58), .ZN(n67) );
  INV_X1 U39 ( .A(A[7]), .ZN(n57) );
  OAI21_X1 U40 ( .B1(SH[4]), .B2(n68), .A(n60), .ZN(B[29]) );
  OAI21_X1 U41 ( .B1(SH[4]), .B2(n69), .A(n60), .ZN(B[28]) );
  OAI21_X1 U42 ( .B1(SH[4]), .B2(n70), .A(n60), .ZN(B[27]) );
  OAI21_X1 U43 ( .B1(SH[4]), .B2(n71), .A(n60), .ZN(B[26]) );
  OAI21_X1 U44 ( .B1(SH[4]), .B2(n5), .A(n60), .ZN(B[25]) );
  AOI221_X1 U45 ( .B1(n72), .B2(n73), .C1(n74), .C2(n75), .A(n76), .ZN(n5) );
  OAI21_X1 U46 ( .B1(SH[4]), .B2(n14), .A(n60), .ZN(B[24]) );
  AOI221_X1 U47 ( .B1(n77), .B2(n73), .C1(n78), .C2(n75), .A(n76), .ZN(n14) );
  OAI21_X1 U48 ( .B1(SH[4]), .B2(n20), .A(n60), .ZN(B[23]) );
  AOI221_X1 U49 ( .B1(n79), .B2(n73), .C1(n80), .C2(n75), .A(n76), .ZN(n20) );
  OAI21_X1 U50 ( .B1(SH[4]), .B2(n26), .A(n60), .ZN(B[22]) );
  AOI221_X1 U51 ( .B1(n81), .B2(n73), .C1(n82), .C2(n75), .A(n83), .ZN(n26) );
  INV_X1 U52 ( .A(n84), .ZN(n83) );
  AOI21_X1 U53 ( .B1(n85), .B2(n86), .A(n87), .ZN(n84) );
  OAI21_X1 U54 ( .B1(SH[4]), .B2(n32), .A(n60), .ZN(B[21]) );
  AOI221_X1 U55 ( .B1(n74), .B2(n73), .C1(n12), .C2(n75), .A(n88), .ZN(n32) );
  INV_X1 U56 ( .A(n89), .ZN(n88) );
  AOI21_X1 U57 ( .B1(n85), .B2(n72), .A(n87), .ZN(n89) );
  OAI21_X1 U58 ( .B1(SH[4]), .B2(n36), .A(n60), .ZN(B[20]) );
  AOI221_X1 U59 ( .B1(n78), .B2(n73), .C1(n18), .C2(n75), .A(n90), .ZN(n36) );
  INV_X1 U60 ( .A(n91), .ZN(n90) );
  AOI21_X1 U61 ( .B1(n85), .B2(n77), .A(n87), .ZN(n91) );
  OAI221_X1 U62 ( .B1(n31), .B2(n39), .C1(n92), .C2(n1), .A(n93), .ZN(B[1]) );
  AOI222_X1 U63 ( .A1(n11), .A2(n8), .B1(n42), .B2(n94), .C1(n9), .C2(n34), 
        .ZN(n93) );
  INV_X1 U64 ( .A(n3), .ZN(n34) );
  AOI221_X1 U65 ( .B1(n52), .B2(A[11]), .C1(n53), .C2(A[12]), .A(n95), .ZN(n3)
         );
  OAI22_X1 U66 ( .A1(n96), .A2(n56), .B1(n97), .B2(n58), .ZN(n95) );
  OAI221_X1 U67 ( .B1(n45), .B2(n98), .C1(n47), .C2(n65), .A(n99), .ZN(n94) );
  AOI22_X1 U68 ( .A1(A[2]), .A2(n50), .B1(A[1]), .B2(n51), .ZN(n99) );
  INV_X1 U69 ( .A(n100), .ZN(n8) );
  AOI221_X1 U70 ( .B1(n52), .B2(A[7]), .C1(n53), .C2(A[8]), .A(n101), .ZN(n31)
         );
  OAI22_X1 U71 ( .A1(n48), .A2(n56), .B1(n46), .B2(n58), .ZN(n101) );
  INV_X1 U72 ( .A(A[6]), .ZN(n48) );
  OAI21_X1 U73 ( .B1(SH[4]), .B2(n40), .A(n60), .ZN(B[19]) );
  AOI221_X1 U74 ( .B1(n80), .B2(n73), .C1(n24), .C2(n75), .A(n102), .ZN(n40)
         );
  INV_X1 U75 ( .A(n103), .ZN(n102) );
  AOI21_X1 U76 ( .B1(n85), .B2(n79), .A(n87), .ZN(n103) );
  NOR2_X1 U77 ( .A1(n104), .A2(n105), .ZN(n87) );
  OAI21_X1 U78 ( .B1(SH[4]), .B2(n61), .A(n60), .ZN(B[18]) );
  AOI221_X1 U79 ( .B1(n86), .B2(n106), .C1(n81), .C2(n85), .A(n107), .ZN(n61)
         );
  INV_X1 U80 ( .A(n108), .ZN(n107) );
  AOI22_X1 U81 ( .A1(n73), .A2(n82), .B1(n75), .B2(n30), .ZN(n108) );
  OAI21_X1 U82 ( .B1(SH[4]), .B2(n92), .A(n60), .ZN(B[17]) );
  AOI221_X1 U83 ( .B1(n12), .B2(n73), .C1(n10), .C2(n75), .A(n109), .ZN(n92)
         );
  INV_X1 U84 ( .A(n110), .ZN(n109) );
  AOI22_X1 U85 ( .A1(n106), .A2(n72), .B1(n85), .B2(n74), .ZN(n110) );
  OAI21_X1 U86 ( .B1(SH[4]), .B2(n111), .A(n60), .ZN(B[16]) );
  OAI221_X1 U87 ( .B1(n112), .B2(n39), .C1(n113), .C2(n4), .A(n114), .ZN(B[15]) );
  AOI221_X1 U88 ( .B1(n11), .B2(n79), .C1(n9), .C2(n80), .A(n115), .ZN(n114)
         );
  INV_X1 U89 ( .A(n60), .ZN(n115) );
  NAND2_X1 U90 ( .A1(SH[4]), .A2(\A[31] ), .ZN(n60) );
  INV_X1 U91 ( .A(n23), .ZN(n113) );
  INV_X1 U92 ( .A(n24), .ZN(n112) );
  OAI221_X1 U93 ( .B1(n116), .B2(n4), .C1(n59), .C2(n1), .A(n117), .ZN(B[14])
         );
  AOI222_X1 U94 ( .A1(n7), .A2(n30), .B1(n9), .B2(n82), .C1(n11), .C2(n81), 
        .ZN(n117) );
  AOI21_X1 U95 ( .B1(n86), .B2(n75), .A(n118), .ZN(n59) );
  OAI221_X1 U96 ( .B1(n100), .B2(n4), .C1(n68), .C2(n2), .A(n119), .ZN(B[13])
         );
  AOI222_X1 U97 ( .A1(n7), .A2(n10), .B1(n9), .B2(n12), .C1(n11), .C2(n74), 
        .ZN(n119) );
  OAI221_X1 U98 ( .B1(n45), .B2(n120), .C1(n47), .C2(n121), .A(n122), .ZN(n74)
         );
  AOI22_X1 U99 ( .A1(A[26]), .A2(n50), .B1(A[25]), .B2(n51), .ZN(n122) );
  OAI221_X1 U100 ( .B1(n45), .B2(n123), .C1(n47), .C2(n124), .A(n125), .ZN(n12) );
  AOI22_X1 U101 ( .A1(A[22]), .A2(n50), .B1(A[21]), .B2(n51), .ZN(n125) );
  INV_X1 U102 ( .A(A[23]), .ZN(n123) );
  OAI221_X1 U103 ( .B1(n45), .B2(n126), .C1(n47), .C2(n127), .A(n128), .ZN(n10) );
  AOI22_X1 U104 ( .A1(A[18]), .A2(n50), .B1(A[17]), .B2(n51), .ZN(n128) );
  AOI21_X1 U105 ( .B1(n72), .B2(n75), .A(n118), .ZN(n68) );
  OAI222_X1 U106 ( .A1(n58), .A2(n129), .B1(n56), .B2(n130), .C1(n131), .C2(
        n132), .ZN(n72) );
  AOI221_X1 U107 ( .B1(n52), .B2(A[15]), .C1(n53), .C2(A[16]), .A(n133), .ZN(
        n100) );
  INV_X1 U108 ( .A(n134), .ZN(n133) );
  AOI22_X1 U109 ( .A1(A[14]), .A2(n50), .B1(A[13]), .B2(n51), .ZN(n134) );
  OAI221_X1 U110 ( .B1(n135), .B2(n4), .C1(n69), .C2(n2), .A(n136), .ZN(B[12])
         );
  AOI222_X1 U111 ( .A1(n7), .A2(n17), .B1(n9), .B2(n18), .C1(n11), .C2(n78), 
        .ZN(n136) );
  AOI21_X1 U112 ( .B1(n77), .B2(n75), .A(n118), .ZN(n69) );
  OAI221_X1 U113 ( .B1(n44), .B2(n4), .C1(n70), .C2(n2), .A(n137), .ZN(B[11])
         );
  AOI222_X1 U114 ( .A1(n7), .A2(n23), .B1(n9), .B2(n24), .C1(n11), .C2(n80), 
        .ZN(n137) );
  OAI221_X1 U115 ( .B1(n45), .B2(n138), .C1(n47), .C2(n139), .A(n140), .ZN(n80) );
  AOI22_X1 U116 ( .A1(A[24]), .A2(n50), .B1(A[23]), .B2(n51), .ZN(n140) );
  OAI221_X1 U117 ( .B1(n127), .B2(n56), .C1(n126), .C2(n58), .A(n141), .ZN(n24) );
  AOI22_X1 U118 ( .A1(A[21]), .A2(n52), .B1(A[22]), .B2(n53), .ZN(n141) );
  OAI221_X1 U119 ( .B1(n45), .B2(n142), .C1(n47), .C2(n143), .A(n144), .ZN(n23) );
  AOI22_X1 U120 ( .A1(A[16]), .A2(n50), .B1(A[15]), .B2(n51), .ZN(n144) );
  INV_X1 U121 ( .A(A[17]), .ZN(n142) );
  AOI21_X1 U122 ( .B1(n79), .B2(n75), .A(n118), .ZN(n70) );
  OAI21_X1 U123 ( .B1(n105), .B2(n132), .A(n104), .ZN(n118) );
  OAI221_X1 U124 ( .B1(n45), .B2(n129), .C1(n47), .C2(n130), .A(n145), .ZN(n79) );
  AOI22_X1 U125 ( .A1(A[28]), .A2(n50), .B1(A[27]), .B2(n51), .ZN(n145) );
  AOI221_X1 U126 ( .B1(n52), .B2(A[13]), .C1(n53), .C2(A[14]), .A(n146), .ZN(
        n44) );
  OAI22_X1 U127 ( .A1(n147), .A2(n56), .B1(n148), .B2(n58), .ZN(n146) );
  INV_X1 U128 ( .A(A[12]), .ZN(n147) );
  OAI221_X1 U129 ( .B1(n64), .B2(n4), .C1(n71), .C2(n2), .A(n149), .ZN(B[10])
         );
  AOI222_X1 U130 ( .A1(n7), .A2(n29), .B1(n9), .B2(n30), .C1(n11), .C2(n82), 
        .ZN(n149) );
  OAI221_X1 U131 ( .B1(n45), .B2(n124), .C1(n47), .C2(n138), .A(n150), .ZN(n82) );
  AOI22_X1 U132 ( .A1(A[23]), .A2(n50), .B1(A[22]), .B2(n51), .ZN(n150) );
  INV_X1 U133 ( .A(A[25]), .ZN(n138) );
  INV_X1 U134 ( .A(A[24]), .ZN(n124) );
  OAI221_X1 U135 ( .B1(n126), .B2(n56), .C1(n143), .C2(n58), .A(n151), .ZN(n30) );
  AOI22_X1 U136 ( .A1(A[20]), .A2(n52), .B1(A[21]), .B2(n53), .ZN(n151) );
  INV_X1 U137 ( .A(n116), .ZN(n29) );
  INV_X1 U138 ( .A(n153), .ZN(n152) );
  AOI22_X1 U139 ( .A1(A[15]), .A2(n50), .B1(A[14]), .B2(n51), .ZN(n153) );
  INV_X1 U140 ( .A(n39), .ZN(n7) );
  AOI221_X1 U141 ( .B1(n86), .B2(n73), .C1(n81), .C2(n75), .A(n76), .ZN(n71)
         );
  INV_X1 U142 ( .A(n104), .ZN(n76) );
  NAND2_X1 U143 ( .A1(\A[31] ), .A2(SH[3]), .ZN(n104) );
  OAI221_X1 U144 ( .B1(n45), .B2(n121), .C1(n47), .C2(n129), .A(n154), .ZN(n81) );
  AOI22_X1 U145 ( .A1(A[27]), .A2(n50), .B1(A[26]), .B2(n51), .ZN(n154) );
  INV_X1 U146 ( .A(A[29]), .ZN(n129) );
  INV_X1 U147 ( .A(A[28]), .ZN(n121) );
  MUX2_X1 U148 ( .A(A[30]), .B(\A[31] ), .S(n58), .Z(n86) );
  OAI22_X1 U149 ( .A1(n148), .A2(n56), .B1(n96), .B2(n58), .ZN(n155) );
  INV_X1 U150 ( .A(A[10]), .ZN(n96) );
  INV_X1 U151 ( .A(A[11]), .ZN(n148) );
  OAI221_X1 U152 ( .B1(n35), .B2(n39), .C1(n111), .C2(n2), .A(n156), .ZN(B[0])
         );
  AOI222_X1 U153 ( .A1(n11), .A2(n16), .B1(n42), .B2(n157), .C1(n9), .C2(n38), 
        .ZN(n156) );
  INV_X1 U154 ( .A(n13), .ZN(n38) );
  OAI22_X1 U155 ( .A1(n97), .A2(n56), .B1(n55), .B2(n58), .ZN(n158) );
  INV_X1 U156 ( .A(A[8]), .ZN(n55) );
  INV_X1 U157 ( .A(A[9]), .ZN(n97) );
  AND2_X1 U158 ( .A1(n159), .A2(n105), .ZN(n9) );
  OAI221_X1 U159 ( .B1(n45), .B2(n160), .C1(n47), .C2(n98), .A(n161), .ZN(n157) );
  AOI22_X1 U160 ( .A1(A[1]), .A2(n50), .B1(A[0]), .B2(n51), .ZN(n161) );
  INV_X1 U161 ( .A(A[3]), .ZN(n98) );
  INV_X1 U162 ( .A(A[2]), .ZN(n160) );
  INV_X1 U163 ( .A(n4), .ZN(n42) );
  NAND2_X1 U164 ( .A1(n75), .A2(n1), .ZN(n4) );
  INV_X1 U165 ( .A(n135), .ZN(n16) );
  INV_X1 U166 ( .A(n163), .ZN(n162) );
  AOI22_X1 U167 ( .A1(A[13]), .A2(n50), .B1(A[12]), .B2(n51), .ZN(n163) );
  AND2_X1 U168 ( .A1(SH[2]), .A2(n159), .ZN(n11) );
  AND2_X1 U169 ( .A1(SH[3]), .A2(n2), .ZN(n159) );
  AOI221_X1 U170 ( .B1(n18), .B2(n73), .C1(n17), .C2(n75), .A(n164), .ZN(n111)
         );
  INV_X1 U171 ( .A(n165), .ZN(n164) );
  AOI22_X1 U172 ( .A1(n106), .A2(n77), .B1(n85), .B2(n78), .ZN(n165) );
  OAI221_X1 U173 ( .B1(n45), .B2(n139), .C1(n47), .C2(n120), .A(n166), .ZN(n78) );
  AOI22_X1 U174 ( .A1(A[25]), .A2(n50), .B1(A[24]), .B2(n51), .ZN(n166) );
  INV_X1 U175 ( .A(A[27]), .ZN(n120) );
  INV_X1 U176 ( .A(A[26]), .ZN(n139) );
  AND2_X1 U177 ( .A1(SH[3]), .A2(n105), .ZN(n85) );
  OAI221_X1 U178 ( .B1(n45), .B2(n130), .C1(n47), .C2(n132), .A(n167), .ZN(n77) );
  AOI22_X1 U179 ( .A1(A[29]), .A2(n50), .B1(A[28]), .B2(n51), .ZN(n167) );
  INV_X1 U180 ( .A(\A[31] ), .ZN(n132) );
  INV_X1 U181 ( .A(A[30]), .ZN(n130) );
  AND2_X1 U182 ( .A1(SH[2]), .A2(SH[3]), .ZN(n106) );
  OAI221_X1 U183 ( .B1(n45), .B2(n143), .C1(n126), .C2(n47), .A(n168), .ZN(n17) );
  AOI22_X1 U184 ( .A1(A[17]), .A2(n50), .B1(A[16]), .B2(n51), .ZN(n168) );
  INV_X1 U185 ( .A(n58), .ZN(n51) );
  INV_X1 U186 ( .A(n56), .ZN(n50) );
  INV_X1 U187 ( .A(n53), .ZN(n47) );
  INV_X1 U188 ( .A(A[19]), .ZN(n126) );
  INV_X1 U189 ( .A(A[18]), .ZN(n143) );
  INV_X1 U190 ( .A(n52), .ZN(n45) );
  OAI221_X1 U191 ( .B1(n56), .B2(n169), .C1(n127), .C2(n58), .A(n170), .ZN(n18) );
  AOI22_X1 U192 ( .A1(A[22]), .A2(n52), .B1(A[23]), .B2(n53), .ZN(n170) );
  INV_X1 U193 ( .A(A[20]), .ZN(n127) );
  INV_X1 U194 ( .A(A[21]), .ZN(n169) );
  NAND2_X1 U195 ( .A1(n73), .A2(n1), .ZN(n39) );
  NOR2_X1 U196 ( .A1(n105), .A2(SH[3]), .ZN(n73) );
  INV_X1 U197 ( .A(SH[2]), .ZN(n105) );
  OAI22_X1 U198 ( .A1(n46), .A2(n56), .B1(n65), .B2(n58), .ZN(n171) );
  NAND2_X1 U199 ( .A1(n172), .A2(n131), .ZN(n58) );
  INV_X1 U200 ( .A(A[4]), .ZN(n65) );
  NAND2_X1 U201 ( .A1(SH[0]), .A2(n131), .ZN(n56) );
  INV_X1 U202 ( .A(A[5]), .ZN(n46) );
  INV_X1 U203 ( .A(SH[0]), .ZN(n172) );
  INV_X1 U204 ( .A(SH[1]), .ZN(n131) );
endmodule


module SHIFTER_GENERIC_N32_DW_lbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n1,
         n2, n3;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n3), .Z(B[31]) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n3), .Z(B[30]) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n3), .Z(B[29]) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n3), .Z(B[28]) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n3), .Z(B[27]) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n3), .Z(B[26]) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n3), .Z(B[25])
         );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n3), .Z(B[24])
         );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n2), .Z(B[23])
         );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n2), .Z(B[22])
         );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n2), .Z(B[21])
         );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n2), .Z(B[20])
         );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n2), .Z(B[19])
         );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n2), .Z(B[18])
         );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n2), .Z(B[17])
         );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n2), .Z(B[16])
         );
  MUX2_X1 M0_4_15 ( .A(\ML_int[4][15] ), .B(\ML_int[4][31] ), .S(n2), .Z(B[15]) );
  MUX2_X1 M0_4_14 ( .A(\ML_int[4][14] ), .B(\ML_int[4][30] ), .S(n2), .Z(B[14]) );
  MUX2_X1 M0_4_13 ( .A(\ML_int[4][13] ), .B(\ML_int[4][29] ), .S(n2), .Z(B[13]) );
  MUX2_X1 M0_4_12 ( .A(\ML_int[4][12] ), .B(\ML_int[4][28] ), .S(n2), .Z(B[12]) );
  MUX2_X1 M0_4_11 ( .A(\ML_int[4][11] ), .B(\ML_int[4][27] ), .S(n1), .Z(B[11]) );
  MUX2_X1 M0_4_10 ( .A(\ML_int[4][10] ), .B(\ML_int[4][26] ), .S(n1), .Z(B[10]) );
  MUX2_X1 M0_4_9 ( .A(\ML_int[4][9] ), .B(\ML_int[4][25] ), .S(n1), .Z(B[9])
         );
  MUX2_X1 M0_4_8 ( .A(\ML_int[4][8] ), .B(\ML_int[4][24] ), .S(n1), .Z(B[8])
         );
  MUX2_X1 M0_4_7 ( .A(\ML_int[4][7] ), .B(\ML_int[4][23] ), .S(n1), .Z(B[7])
         );
  MUX2_X1 M0_4_6 ( .A(\ML_int[4][6] ), .B(\ML_int[4][22] ), .S(n1), .Z(B[6])
         );
  MUX2_X1 M0_4_5 ( .A(\ML_int[4][5] ), .B(\ML_int[4][21] ), .S(n1), .Z(B[5])
         );
  MUX2_X1 M0_4_4 ( .A(\ML_int[4][4] ), .B(\ML_int[4][20] ), .S(n1), .Z(B[4])
         );
  MUX2_X1 M0_4_3 ( .A(\ML_int[4][3] ), .B(\ML_int[4][19] ), .S(n1), .Z(B[3])
         );
  MUX2_X1 M0_4_2 ( .A(\ML_int[4][2] ), .B(\ML_int[4][18] ), .S(n1), .Z(B[2])
         );
  MUX2_X1 M0_4_1 ( .A(\ML_int[4][1] ), .B(\ML_int[4][17] ), .S(n1), .Z(B[1])
         );
  MUX2_X1 M0_4_0 ( .A(\ML_int[4][0] ), .B(\ML_int[4][16] ), .S(n1), .Z(B[0])
         );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(SH[3]), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(SH[3]), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(SH[3]), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(SH[3]), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(SH[3]), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(SH[3]), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(SH[3]), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(SH[3]), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(SH[3]), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(SH[3]), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(SH[3]), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(SH[3]), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(SH[3]), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(SH[3]), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(SH[3]), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(SH[3]), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(SH[3]), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(SH[3]), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(SH[3]), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(SH[3]), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(SH[3]), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M0_3_7 ( .A(\ML_int[3][7] ), .B(\ML_int[3][31] ), .S(SH[3]), .Z(
        \ML_int[4][7] ) );
  MUX2_X1 M0_3_6 ( .A(\ML_int[3][6] ), .B(\ML_int[3][30] ), .S(SH[3]), .Z(
        \ML_int[4][6] ) );
  MUX2_X1 M0_3_5 ( .A(\ML_int[3][5] ), .B(\ML_int[3][29] ), .S(SH[3]), .Z(
        \ML_int[4][5] ) );
  MUX2_X1 M0_3_4 ( .A(\ML_int[3][4] ), .B(\ML_int[3][28] ), .S(SH[3]), .Z(
        \ML_int[4][4] ) );
  MUX2_X1 M0_3_3 ( .A(\ML_int[3][3] ), .B(\ML_int[3][27] ), .S(SH[3]), .Z(
        \ML_int[4][3] ) );
  MUX2_X1 M0_3_2 ( .A(\ML_int[3][2] ), .B(\ML_int[3][26] ), .S(SH[3]), .Z(
        \ML_int[4][2] ) );
  MUX2_X1 M0_3_1 ( .A(\ML_int[3][1] ), .B(\ML_int[3][25] ), .S(SH[3]), .Z(
        \ML_int[4][1] ) );
  MUX2_X1 M0_3_0 ( .A(\ML_int[3][0] ), .B(\ML_int[3][24] ), .S(SH[3]), .Z(
        \ML_int[4][0] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(SH[2]), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(SH[2]), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(SH[2]), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(SH[2]), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(SH[2]), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(SH[2]), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(SH[2]), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(SH[2]), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(SH[2]), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(SH[2]), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(SH[2]), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(SH[2]), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M0_2_3 ( .A(\ML_int[2][3] ), .B(\ML_int[2][31] ), .S(SH[2]), .Z(
        \ML_int[3][3] ) );
  MUX2_X1 M0_2_2 ( .A(\ML_int[2][2] ), .B(\ML_int[2][30] ), .S(SH[2]), .Z(
        \ML_int[3][2] ) );
  MUX2_X1 M0_2_1 ( .A(\ML_int[2][1] ), .B(\ML_int[2][29] ), .S(SH[2]), .Z(
        \ML_int[3][1] ) );
  MUX2_X1 M0_2_0 ( .A(\ML_int[2][0] ), .B(\ML_int[2][28] ), .S(SH[2]), .Z(
        \ML_int[3][0] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(SH[1]), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(SH[1]), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(SH[1]), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(SH[1]), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(SH[1]), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(SH[1]), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(SH[1]), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(SH[1]), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(SH[1]), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(SH[1]), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(SH[1]), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(SH[1]), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(SH[1]), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(SH[1]), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(SH[1]), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(SH[1]), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(SH[1]), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(SH[1]), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(SH[1]), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(SH[1]), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(SH[1]), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(SH[1]), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(SH[1]), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(SH[1]), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(SH[1]), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(SH[1]), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(SH[1]), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(SH[1]), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(SH[1]), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M0_1_1 ( .A(\ML_int[1][1] ), .B(\ML_int[1][31] ), .S(SH[1]), .Z(
        \ML_int[2][1] ) );
  MUX2_X1 M0_1_0 ( .A(\ML_int[1][0] ), .B(\ML_int[1][30] ), .S(SH[1]), .Z(
        \ML_int[2][0] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(SH[0]), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(SH[0]), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(SH[0]), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(SH[0]), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(SH[0]), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2_X1 M0_0_0 ( .A(A[0]), .B(A[31]), .S(SH[0]), .Z(\ML_int[1][0] ) );
  CLKBUF_X3 U2 ( .A(SH[4]), .Z(n1) );
  CLKBUF_X3 U3 ( .A(SH[4]), .Z(n2) );
  CLKBUF_X3 U4 ( .A(SH[4]), .Z(n3) );
endmodule


module SHIFTER_GENERIC_N32_DW_rbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \MR_int[1][31] , \MR_int[1][30] , \MR_int[1][29] , \MR_int[1][28] ,
         \MR_int[1][27] , \MR_int[1][26] , \MR_int[1][25] , \MR_int[1][24] ,
         \MR_int[1][23] , \MR_int[1][22] , \MR_int[1][21] , \MR_int[1][20] ,
         \MR_int[1][19] , \MR_int[1][18] , \MR_int[1][17] , \MR_int[1][16] ,
         \MR_int[1][15] , \MR_int[1][14] , \MR_int[1][13] , \MR_int[1][12] ,
         \MR_int[1][11] , \MR_int[1][10] , \MR_int[1][9] , \MR_int[1][8] ,
         \MR_int[1][7] , \MR_int[1][6] , \MR_int[1][5] , \MR_int[1][4] ,
         \MR_int[1][3] , \MR_int[1][2] , \MR_int[1][1] , \MR_int[1][0] ,
         \MR_int[2][31] , \MR_int[2][30] , \MR_int[2][29] , \MR_int[2][28] ,
         \MR_int[2][27] , \MR_int[2][26] , \MR_int[2][25] , \MR_int[2][24] ,
         \MR_int[2][23] , \MR_int[2][22] , \MR_int[2][21] , \MR_int[2][20] ,
         \MR_int[2][19] , \MR_int[2][18] , \MR_int[2][17] , \MR_int[2][16] ,
         \MR_int[2][15] , \MR_int[2][14] , \MR_int[2][13] , \MR_int[2][12] ,
         \MR_int[2][11] , \MR_int[2][10] , \MR_int[2][9] , \MR_int[2][8] ,
         \MR_int[2][7] , \MR_int[2][6] , \MR_int[2][5] , \MR_int[2][4] ,
         \MR_int[2][3] , \MR_int[2][2] , \MR_int[2][1] , \MR_int[2][0] ,
         \MR_int[3][31] , \MR_int[3][30] , \MR_int[3][29] , \MR_int[3][28] ,
         \MR_int[3][27] , \MR_int[3][26] , \MR_int[3][25] , \MR_int[3][24] ,
         \MR_int[3][23] , \MR_int[3][22] , \MR_int[3][21] , \MR_int[3][20] ,
         \MR_int[3][19] , \MR_int[3][18] , \MR_int[3][17] , \MR_int[3][16] ,
         \MR_int[3][15] , \MR_int[3][14] , \MR_int[3][13] , \MR_int[3][12] ,
         \MR_int[3][11] , \MR_int[3][10] , \MR_int[3][9] , \MR_int[3][8] ,
         \MR_int[3][7] , \MR_int[3][6] , \MR_int[3][5] , \MR_int[3][4] ,
         \MR_int[3][3] , \MR_int[3][2] , \MR_int[3][1] , \MR_int[3][0] ,
         \MR_int[4][31] , \MR_int[4][30] , \MR_int[4][29] , \MR_int[4][28] ,
         \MR_int[4][27] , \MR_int[4][26] , \MR_int[4][25] , \MR_int[4][24] ,
         \MR_int[4][23] , \MR_int[4][22] , \MR_int[4][21] , \MR_int[4][20] ,
         \MR_int[4][19] , \MR_int[4][18] , \MR_int[4][17] , \MR_int[4][16] ,
         \MR_int[4][15] , \MR_int[4][14] , \MR_int[4][13] , \MR_int[4][12] ,
         \MR_int[4][11] , \MR_int[4][10] , \MR_int[4][9] , \MR_int[4][8] ,
         \MR_int[4][7] , \MR_int[4][6] , \MR_int[4][5] , \MR_int[4][4] ,
         \MR_int[4][3] , \MR_int[4][2] , \MR_int[4][1] , \MR_int[4][0] , n1,
         n2, n3;

  MUX2_X1 M1_4_31 ( .A(\MR_int[4][31] ), .B(\MR_int[4][15] ), .S(n3), .Z(B[31]) );
  MUX2_X1 M1_4_30 ( .A(\MR_int[4][30] ), .B(\MR_int[4][14] ), .S(n3), .Z(B[30]) );
  MUX2_X1 M1_4_29 ( .A(\MR_int[4][29] ), .B(\MR_int[4][13] ), .S(n3), .Z(B[29]) );
  MUX2_X1 M1_4_28 ( .A(\MR_int[4][28] ), .B(\MR_int[4][12] ), .S(n3), .Z(B[28]) );
  MUX2_X1 M1_4_27 ( .A(\MR_int[4][27] ), .B(\MR_int[4][11] ), .S(n3), .Z(B[27]) );
  MUX2_X1 M1_4_26 ( .A(\MR_int[4][26] ), .B(\MR_int[4][10] ), .S(n3), .Z(B[26]) );
  MUX2_X1 M1_4_25 ( .A(\MR_int[4][25] ), .B(\MR_int[4][9] ), .S(n3), .Z(B[25])
         );
  MUX2_X1 M1_4_24 ( .A(\MR_int[4][24] ), .B(\MR_int[4][8] ), .S(n3), .Z(B[24])
         );
  MUX2_X1 M1_4_23 ( .A(\MR_int[4][23] ), .B(\MR_int[4][7] ), .S(n2), .Z(B[23])
         );
  MUX2_X1 M1_4_22 ( .A(\MR_int[4][22] ), .B(\MR_int[4][6] ), .S(n2), .Z(B[22])
         );
  MUX2_X1 M1_4_21 ( .A(\MR_int[4][21] ), .B(\MR_int[4][5] ), .S(n2), .Z(B[21])
         );
  MUX2_X1 M1_4_20 ( .A(\MR_int[4][20] ), .B(\MR_int[4][4] ), .S(n2), .Z(B[20])
         );
  MUX2_X1 M1_4_19 ( .A(\MR_int[4][19] ), .B(\MR_int[4][3] ), .S(n2), .Z(B[19])
         );
  MUX2_X1 M1_4_18 ( .A(\MR_int[4][18] ), .B(\MR_int[4][2] ), .S(n2), .Z(B[18])
         );
  MUX2_X1 M1_4_17 ( .A(\MR_int[4][17] ), .B(\MR_int[4][1] ), .S(n2), .Z(B[17])
         );
  MUX2_X1 M1_4_16 ( .A(\MR_int[4][16] ), .B(\MR_int[4][0] ), .S(n2), .Z(B[16])
         );
  MUX2_X1 M1_4_15 ( .A(\MR_int[4][15] ), .B(\MR_int[4][31] ), .S(n2), .Z(B[15]) );
  MUX2_X1 M1_4_14 ( .A(\MR_int[4][14] ), .B(\MR_int[4][30] ), .S(n2), .Z(B[14]) );
  MUX2_X1 M1_4_13 ( .A(\MR_int[4][13] ), .B(\MR_int[4][29] ), .S(n2), .Z(B[13]) );
  MUX2_X1 M1_4_12 ( .A(\MR_int[4][12] ), .B(\MR_int[4][28] ), .S(n2), .Z(B[12]) );
  MUX2_X1 M1_4_11 ( .A(\MR_int[4][11] ), .B(\MR_int[4][27] ), .S(n1), .Z(B[11]) );
  MUX2_X1 M1_4_10 ( .A(\MR_int[4][10] ), .B(\MR_int[4][26] ), .S(n1), .Z(B[10]) );
  MUX2_X1 M1_4_9 ( .A(\MR_int[4][9] ), .B(\MR_int[4][25] ), .S(n1), .Z(B[9])
         );
  MUX2_X1 M1_4_8 ( .A(\MR_int[4][8] ), .B(\MR_int[4][24] ), .S(n1), .Z(B[8])
         );
  MUX2_X1 M1_4_7 ( .A(\MR_int[4][7] ), .B(\MR_int[4][23] ), .S(n1), .Z(B[7])
         );
  MUX2_X1 M1_4_6 ( .A(\MR_int[4][6] ), .B(\MR_int[4][22] ), .S(n1), .Z(B[6])
         );
  MUX2_X1 M1_4_5 ( .A(\MR_int[4][5] ), .B(\MR_int[4][21] ), .S(n1), .Z(B[5])
         );
  MUX2_X1 M1_4_4 ( .A(\MR_int[4][4] ), .B(\MR_int[4][20] ), .S(n1), .Z(B[4])
         );
  MUX2_X1 M1_4_3 ( .A(\MR_int[4][3] ), .B(\MR_int[4][19] ), .S(n1), .Z(B[3])
         );
  MUX2_X1 M1_4_2 ( .A(\MR_int[4][2] ), .B(\MR_int[4][18] ), .S(n1), .Z(B[2])
         );
  MUX2_X1 M1_4_1 ( .A(\MR_int[4][1] ), .B(\MR_int[4][17] ), .S(n1), .Z(B[1])
         );
  MUX2_X1 M1_4_0 ( .A(\MR_int[4][0] ), .B(\MR_int[4][16] ), .S(n1), .Z(B[0])
         );
  MUX2_X1 M1_3_31_0 ( .A(\MR_int[3][31] ), .B(\MR_int[3][7] ), .S(SH[3]), .Z(
        \MR_int[4][31] ) );
  MUX2_X1 M1_3_30_0 ( .A(\MR_int[3][30] ), .B(\MR_int[3][6] ), .S(SH[3]), .Z(
        \MR_int[4][30] ) );
  MUX2_X1 M1_3_29_0 ( .A(\MR_int[3][29] ), .B(\MR_int[3][5] ), .S(SH[3]), .Z(
        \MR_int[4][29] ) );
  MUX2_X1 M1_3_28_0 ( .A(\MR_int[3][28] ), .B(\MR_int[3][4] ), .S(SH[3]), .Z(
        \MR_int[4][28] ) );
  MUX2_X1 M1_3_27_0 ( .A(\MR_int[3][27] ), .B(\MR_int[3][3] ), .S(SH[3]), .Z(
        \MR_int[4][27] ) );
  MUX2_X1 M1_3_26_0 ( .A(\MR_int[3][26] ), .B(\MR_int[3][2] ), .S(SH[3]), .Z(
        \MR_int[4][26] ) );
  MUX2_X1 M1_3_25_0 ( .A(\MR_int[3][25] ), .B(\MR_int[3][1] ), .S(SH[3]), .Z(
        \MR_int[4][25] ) );
  MUX2_X1 M1_3_24_0 ( .A(\MR_int[3][24] ), .B(\MR_int[3][0] ), .S(SH[3]), .Z(
        \MR_int[4][24] ) );
  MUX2_X1 M1_3_23_0 ( .A(\MR_int[3][23] ), .B(\MR_int[3][31] ), .S(SH[3]), .Z(
        \MR_int[4][23] ) );
  MUX2_X1 M1_3_22_0 ( .A(\MR_int[3][22] ), .B(\MR_int[3][30] ), .S(SH[3]), .Z(
        \MR_int[4][22] ) );
  MUX2_X1 M1_3_21_0 ( .A(\MR_int[3][21] ), .B(\MR_int[3][29] ), .S(SH[3]), .Z(
        \MR_int[4][21] ) );
  MUX2_X1 M1_3_20_0 ( .A(\MR_int[3][20] ), .B(\MR_int[3][28] ), .S(SH[3]), .Z(
        \MR_int[4][20] ) );
  MUX2_X1 M1_3_19_0 ( .A(\MR_int[3][19] ), .B(\MR_int[3][27] ), .S(SH[3]), .Z(
        \MR_int[4][19] ) );
  MUX2_X1 M1_3_18_0 ( .A(\MR_int[3][18] ), .B(\MR_int[3][26] ), .S(SH[3]), .Z(
        \MR_int[4][18] ) );
  MUX2_X1 M1_3_17_0 ( .A(\MR_int[3][17] ), .B(\MR_int[3][25] ), .S(SH[3]), .Z(
        \MR_int[4][17] ) );
  MUX2_X1 M1_3_16_0 ( .A(\MR_int[3][16] ), .B(\MR_int[3][24] ), .S(SH[3]), .Z(
        \MR_int[4][16] ) );
  MUX2_X1 M1_3_15_0 ( .A(\MR_int[3][15] ), .B(\MR_int[3][23] ), .S(SH[3]), .Z(
        \MR_int[4][15] ) );
  MUX2_X1 M1_3_14_0 ( .A(\MR_int[3][14] ), .B(\MR_int[3][22] ), .S(SH[3]), .Z(
        \MR_int[4][14] ) );
  MUX2_X1 M1_3_13_0 ( .A(\MR_int[3][13] ), .B(\MR_int[3][21] ), .S(SH[3]), .Z(
        \MR_int[4][13] ) );
  MUX2_X1 M1_3_12_0 ( .A(\MR_int[3][12] ), .B(\MR_int[3][20] ), .S(SH[3]), .Z(
        \MR_int[4][12] ) );
  MUX2_X1 M1_3_11_0 ( .A(\MR_int[3][11] ), .B(\MR_int[3][19] ), .S(SH[3]), .Z(
        \MR_int[4][11] ) );
  MUX2_X1 M1_3_10_0 ( .A(\MR_int[3][10] ), .B(\MR_int[3][18] ), .S(SH[3]), .Z(
        \MR_int[4][10] ) );
  MUX2_X1 M1_3_9_0 ( .A(\MR_int[3][9] ), .B(\MR_int[3][17] ), .S(SH[3]), .Z(
        \MR_int[4][9] ) );
  MUX2_X1 M1_3_8_0 ( .A(\MR_int[3][8] ), .B(\MR_int[3][16] ), .S(SH[3]), .Z(
        \MR_int[4][8] ) );
  MUX2_X1 M1_3_7 ( .A(\MR_int[3][7] ), .B(\MR_int[3][15] ), .S(SH[3]), .Z(
        \MR_int[4][7] ) );
  MUX2_X1 M1_3_6 ( .A(\MR_int[3][6] ), .B(\MR_int[3][14] ), .S(SH[3]), .Z(
        \MR_int[4][6] ) );
  MUX2_X1 M1_3_5 ( .A(\MR_int[3][5] ), .B(\MR_int[3][13] ), .S(SH[3]), .Z(
        \MR_int[4][5] ) );
  MUX2_X1 M1_3_4 ( .A(\MR_int[3][4] ), .B(\MR_int[3][12] ), .S(SH[3]), .Z(
        \MR_int[4][4] ) );
  MUX2_X1 M1_3_3 ( .A(\MR_int[3][3] ), .B(\MR_int[3][11] ), .S(SH[3]), .Z(
        \MR_int[4][3] ) );
  MUX2_X1 M1_3_2 ( .A(\MR_int[3][2] ), .B(\MR_int[3][10] ), .S(SH[3]), .Z(
        \MR_int[4][2] ) );
  MUX2_X1 M1_3_1 ( .A(\MR_int[3][1] ), .B(\MR_int[3][9] ), .S(SH[3]), .Z(
        \MR_int[4][1] ) );
  MUX2_X1 M1_3_0 ( .A(\MR_int[3][0] ), .B(\MR_int[3][8] ), .S(SH[3]), .Z(
        \MR_int[4][0] ) );
  MUX2_X1 M1_2_31_0 ( .A(\MR_int[2][31] ), .B(\MR_int[2][3] ), .S(SH[2]), .Z(
        \MR_int[3][31] ) );
  MUX2_X1 M1_2_30_0 ( .A(\MR_int[2][30] ), .B(\MR_int[2][2] ), .S(SH[2]), .Z(
        \MR_int[3][30] ) );
  MUX2_X1 M1_2_29_0 ( .A(\MR_int[2][29] ), .B(\MR_int[2][1] ), .S(SH[2]), .Z(
        \MR_int[3][29] ) );
  MUX2_X1 M1_2_28_0 ( .A(\MR_int[2][28] ), .B(\MR_int[2][0] ), .S(SH[2]), .Z(
        \MR_int[3][28] ) );
  MUX2_X1 M1_2_27_0 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(SH[2]), .Z(
        \MR_int[3][27] ) );
  MUX2_X1 M1_2_26_0 ( .A(\MR_int[2][26] ), .B(\MR_int[2][30] ), .S(SH[2]), .Z(
        \MR_int[3][26] ) );
  MUX2_X1 M1_2_25_0 ( .A(\MR_int[2][25] ), .B(\MR_int[2][29] ), .S(SH[2]), .Z(
        \MR_int[3][25] ) );
  MUX2_X1 M1_2_24_0 ( .A(\MR_int[2][24] ), .B(\MR_int[2][28] ), .S(SH[2]), .Z(
        \MR_int[3][24] ) );
  MUX2_X1 M1_2_23_0 ( .A(\MR_int[2][23] ), .B(\MR_int[2][27] ), .S(SH[2]), .Z(
        \MR_int[3][23] ) );
  MUX2_X1 M1_2_22_0 ( .A(\MR_int[2][22] ), .B(\MR_int[2][26] ), .S(SH[2]), .Z(
        \MR_int[3][22] ) );
  MUX2_X1 M1_2_21_0 ( .A(\MR_int[2][21] ), .B(\MR_int[2][25] ), .S(SH[2]), .Z(
        \MR_int[3][21] ) );
  MUX2_X1 M1_2_20_0 ( .A(\MR_int[2][20] ), .B(\MR_int[2][24] ), .S(SH[2]), .Z(
        \MR_int[3][20] ) );
  MUX2_X1 M1_2_19_0 ( .A(\MR_int[2][19] ), .B(\MR_int[2][23] ), .S(SH[2]), .Z(
        \MR_int[3][19] ) );
  MUX2_X1 M1_2_18_0 ( .A(\MR_int[2][18] ), .B(\MR_int[2][22] ), .S(SH[2]), .Z(
        \MR_int[3][18] ) );
  MUX2_X1 M1_2_17_0 ( .A(\MR_int[2][17] ), .B(\MR_int[2][21] ), .S(SH[2]), .Z(
        \MR_int[3][17] ) );
  MUX2_X1 M1_2_16_0 ( .A(\MR_int[2][16] ), .B(\MR_int[2][20] ), .S(SH[2]), .Z(
        \MR_int[3][16] ) );
  MUX2_X1 M1_2_15_0 ( .A(\MR_int[2][15] ), .B(\MR_int[2][19] ), .S(SH[2]), .Z(
        \MR_int[3][15] ) );
  MUX2_X1 M1_2_14_0 ( .A(\MR_int[2][14] ), .B(\MR_int[2][18] ), .S(SH[2]), .Z(
        \MR_int[3][14] ) );
  MUX2_X1 M1_2_13_0 ( .A(\MR_int[2][13] ), .B(\MR_int[2][17] ), .S(SH[2]), .Z(
        \MR_int[3][13] ) );
  MUX2_X1 M1_2_12_0 ( .A(\MR_int[2][12] ), .B(\MR_int[2][16] ), .S(SH[2]), .Z(
        \MR_int[3][12] ) );
  MUX2_X1 M1_2_11_0 ( .A(\MR_int[2][11] ), .B(\MR_int[2][15] ), .S(SH[2]), .Z(
        \MR_int[3][11] ) );
  MUX2_X1 M1_2_10_0 ( .A(\MR_int[2][10] ), .B(\MR_int[2][14] ), .S(SH[2]), .Z(
        \MR_int[3][10] ) );
  MUX2_X1 M1_2_9_0 ( .A(\MR_int[2][9] ), .B(\MR_int[2][13] ), .S(SH[2]), .Z(
        \MR_int[3][9] ) );
  MUX2_X1 M1_2_8_0 ( .A(\MR_int[2][8] ), .B(\MR_int[2][12] ), .S(SH[2]), .Z(
        \MR_int[3][8] ) );
  MUX2_X1 M1_2_7_0 ( .A(\MR_int[2][7] ), .B(\MR_int[2][11] ), .S(SH[2]), .Z(
        \MR_int[3][7] ) );
  MUX2_X1 M1_2_6_0 ( .A(\MR_int[2][6] ), .B(\MR_int[2][10] ), .S(SH[2]), .Z(
        \MR_int[3][6] ) );
  MUX2_X1 M1_2_5_0 ( .A(\MR_int[2][5] ), .B(\MR_int[2][9] ), .S(SH[2]), .Z(
        \MR_int[3][5] ) );
  MUX2_X1 M1_2_4_0 ( .A(\MR_int[2][4] ), .B(\MR_int[2][8] ), .S(SH[2]), .Z(
        \MR_int[3][4] ) );
  MUX2_X1 M1_2_3 ( .A(\MR_int[2][3] ), .B(\MR_int[2][7] ), .S(SH[2]), .Z(
        \MR_int[3][3] ) );
  MUX2_X1 M1_2_2 ( .A(\MR_int[2][2] ), .B(\MR_int[2][6] ), .S(SH[2]), .Z(
        \MR_int[3][2] ) );
  MUX2_X1 M1_2_1 ( .A(\MR_int[2][1] ), .B(\MR_int[2][5] ), .S(SH[2]), .Z(
        \MR_int[3][1] ) );
  MUX2_X1 M1_2_0 ( .A(\MR_int[2][0] ), .B(\MR_int[2][4] ), .S(SH[2]), .Z(
        \MR_int[3][0] ) );
  MUX2_X1 M1_1_31_0 ( .A(\MR_int[1][31] ), .B(\MR_int[1][1] ), .S(SH[1]), .Z(
        \MR_int[2][31] ) );
  MUX2_X1 M1_1_30_0 ( .A(\MR_int[1][30] ), .B(\MR_int[1][0] ), .S(SH[1]), .Z(
        \MR_int[2][30] ) );
  MUX2_X1 M1_1_29_0 ( .A(\MR_int[1][29] ), .B(\MR_int[1][31] ), .S(SH[1]), .Z(
        \MR_int[2][29] ) );
  MUX2_X1 M1_1_28_0 ( .A(\MR_int[1][28] ), .B(\MR_int[1][30] ), .S(SH[1]), .Z(
        \MR_int[2][28] ) );
  MUX2_X1 M1_1_27_0 ( .A(\MR_int[1][27] ), .B(\MR_int[1][29] ), .S(SH[1]), .Z(
        \MR_int[2][27] ) );
  MUX2_X1 M1_1_26_0 ( .A(\MR_int[1][26] ), .B(\MR_int[1][28] ), .S(SH[1]), .Z(
        \MR_int[2][26] ) );
  MUX2_X1 M1_1_25_0 ( .A(\MR_int[1][25] ), .B(\MR_int[1][27] ), .S(SH[1]), .Z(
        \MR_int[2][25] ) );
  MUX2_X1 M1_1_24_0 ( .A(\MR_int[1][24] ), .B(\MR_int[1][26] ), .S(SH[1]), .Z(
        \MR_int[2][24] ) );
  MUX2_X1 M1_1_23_0 ( .A(\MR_int[1][23] ), .B(\MR_int[1][25] ), .S(SH[1]), .Z(
        \MR_int[2][23] ) );
  MUX2_X1 M1_1_22_0 ( .A(\MR_int[1][22] ), .B(\MR_int[1][24] ), .S(SH[1]), .Z(
        \MR_int[2][22] ) );
  MUX2_X1 M1_1_21_0 ( .A(\MR_int[1][21] ), .B(\MR_int[1][23] ), .S(SH[1]), .Z(
        \MR_int[2][21] ) );
  MUX2_X1 M1_1_20_0 ( .A(\MR_int[1][20] ), .B(\MR_int[1][22] ), .S(SH[1]), .Z(
        \MR_int[2][20] ) );
  MUX2_X1 M1_1_19_0 ( .A(\MR_int[1][19] ), .B(\MR_int[1][21] ), .S(SH[1]), .Z(
        \MR_int[2][19] ) );
  MUX2_X1 M1_1_18_0 ( .A(\MR_int[1][18] ), .B(\MR_int[1][20] ), .S(SH[1]), .Z(
        \MR_int[2][18] ) );
  MUX2_X1 M1_1_17_0 ( .A(\MR_int[1][17] ), .B(\MR_int[1][19] ), .S(SH[1]), .Z(
        \MR_int[2][17] ) );
  MUX2_X1 M1_1_16_0 ( .A(\MR_int[1][16] ), .B(\MR_int[1][18] ), .S(SH[1]), .Z(
        \MR_int[2][16] ) );
  MUX2_X1 M1_1_15_0 ( .A(\MR_int[1][15] ), .B(\MR_int[1][17] ), .S(SH[1]), .Z(
        \MR_int[2][15] ) );
  MUX2_X1 M1_1_14_0 ( .A(\MR_int[1][14] ), .B(\MR_int[1][16] ), .S(SH[1]), .Z(
        \MR_int[2][14] ) );
  MUX2_X1 M1_1_13_0 ( .A(\MR_int[1][13] ), .B(\MR_int[1][15] ), .S(SH[1]), .Z(
        \MR_int[2][13] ) );
  MUX2_X1 M1_1_12_0 ( .A(\MR_int[1][12] ), .B(\MR_int[1][14] ), .S(SH[1]), .Z(
        \MR_int[2][12] ) );
  MUX2_X1 M1_1_11_0 ( .A(\MR_int[1][11] ), .B(\MR_int[1][13] ), .S(SH[1]), .Z(
        \MR_int[2][11] ) );
  MUX2_X1 M1_1_10_0 ( .A(\MR_int[1][10] ), .B(\MR_int[1][12] ), .S(SH[1]), .Z(
        \MR_int[2][10] ) );
  MUX2_X1 M1_1_9_0 ( .A(\MR_int[1][9] ), .B(\MR_int[1][11] ), .S(SH[1]), .Z(
        \MR_int[2][9] ) );
  MUX2_X1 M1_1_8_0 ( .A(\MR_int[1][8] ), .B(\MR_int[1][10] ), .S(SH[1]), .Z(
        \MR_int[2][8] ) );
  MUX2_X1 M1_1_7_0 ( .A(\MR_int[1][7] ), .B(\MR_int[1][9] ), .S(SH[1]), .Z(
        \MR_int[2][7] ) );
  MUX2_X1 M1_1_6_0 ( .A(\MR_int[1][6] ), .B(\MR_int[1][8] ), .S(SH[1]), .Z(
        \MR_int[2][6] ) );
  MUX2_X1 M1_1_5_0 ( .A(\MR_int[1][5] ), .B(\MR_int[1][7] ), .S(SH[1]), .Z(
        \MR_int[2][5] ) );
  MUX2_X1 M1_1_4_0 ( .A(\MR_int[1][4] ), .B(\MR_int[1][6] ), .S(SH[1]), .Z(
        \MR_int[2][4] ) );
  MUX2_X1 M1_1_3_0 ( .A(\MR_int[1][3] ), .B(\MR_int[1][5] ), .S(SH[1]), .Z(
        \MR_int[2][3] ) );
  MUX2_X1 M1_1_2_0 ( .A(\MR_int[1][2] ), .B(\MR_int[1][4] ), .S(SH[1]), .Z(
        \MR_int[2][2] ) );
  MUX2_X1 M1_1_1 ( .A(\MR_int[1][1] ), .B(\MR_int[1][3] ), .S(SH[1]), .Z(
        \MR_int[2][1] ) );
  MUX2_X1 M1_1_0 ( .A(\MR_int[1][0] ), .B(\MR_int[1][2] ), .S(SH[1]), .Z(
        \MR_int[2][0] ) );
  MUX2_X1 M1_0_31_0 ( .A(A[31]), .B(A[0]), .S(SH[0]), .Z(\MR_int[1][31] ) );
  MUX2_X1 M1_0_30_0 ( .A(A[30]), .B(A[31]), .S(SH[0]), .Z(\MR_int[1][30] ) );
  MUX2_X1 M1_0_29_0 ( .A(A[29]), .B(A[30]), .S(SH[0]), .Z(\MR_int[1][29] ) );
  MUX2_X1 M1_0_28_0 ( .A(A[28]), .B(A[29]), .S(SH[0]), .Z(\MR_int[1][28] ) );
  MUX2_X1 M1_0_27_0 ( .A(A[27]), .B(A[28]), .S(SH[0]), .Z(\MR_int[1][27] ) );
  MUX2_X1 M1_0_26_0 ( .A(A[26]), .B(A[27]), .S(SH[0]), .Z(\MR_int[1][26] ) );
  MUX2_X1 M1_0_25_0 ( .A(A[25]), .B(A[26]), .S(SH[0]), .Z(\MR_int[1][25] ) );
  MUX2_X1 M1_0_24_0 ( .A(A[24]), .B(A[25]), .S(SH[0]), .Z(\MR_int[1][24] ) );
  MUX2_X1 M1_0_23_0 ( .A(A[23]), .B(A[24]), .S(SH[0]), .Z(\MR_int[1][23] ) );
  MUX2_X1 M1_0_22_0 ( .A(A[22]), .B(A[23]), .S(SH[0]), .Z(\MR_int[1][22] ) );
  MUX2_X1 M1_0_21_0 ( .A(A[21]), .B(A[22]), .S(SH[0]), .Z(\MR_int[1][21] ) );
  MUX2_X1 M1_0_20_0 ( .A(A[20]), .B(A[21]), .S(SH[0]), .Z(\MR_int[1][20] ) );
  MUX2_X1 M1_0_19_0 ( .A(A[19]), .B(A[20]), .S(SH[0]), .Z(\MR_int[1][19] ) );
  MUX2_X1 M1_0_18_0 ( .A(A[18]), .B(A[19]), .S(SH[0]), .Z(\MR_int[1][18] ) );
  MUX2_X1 M1_0_17_0 ( .A(A[17]), .B(A[18]), .S(SH[0]), .Z(\MR_int[1][17] ) );
  MUX2_X1 M1_0_16_0 ( .A(A[16]), .B(A[17]), .S(SH[0]), .Z(\MR_int[1][16] ) );
  MUX2_X1 M1_0_15_0 ( .A(A[15]), .B(A[16]), .S(SH[0]), .Z(\MR_int[1][15] ) );
  MUX2_X1 M1_0_14_0 ( .A(A[14]), .B(A[15]), .S(SH[0]), .Z(\MR_int[1][14] ) );
  MUX2_X1 M1_0_13_0 ( .A(A[13]), .B(A[14]), .S(SH[0]), .Z(\MR_int[1][13] ) );
  MUX2_X1 M1_0_12_0 ( .A(A[12]), .B(A[13]), .S(SH[0]), .Z(\MR_int[1][12] ) );
  MUX2_X1 M1_0_11_0 ( .A(A[11]), .B(A[12]), .S(SH[0]), .Z(\MR_int[1][11] ) );
  MUX2_X1 M1_0_10_0 ( .A(A[10]), .B(A[11]), .S(SH[0]), .Z(\MR_int[1][10] ) );
  MUX2_X1 M1_0_9_0 ( .A(A[9]), .B(A[10]), .S(SH[0]), .Z(\MR_int[1][9] ) );
  MUX2_X1 M1_0_8_0 ( .A(A[8]), .B(A[9]), .S(SH[0]), .Z(\MR_int[1][8] ) );
  MUX2_X1 M1_0_7_0 ( .A(A[7]), .B(A[8]), .S(SH[0]), .Z(\MR_int[1][7] ) );
  MUX2_X1 M1_0_6_0 ( .A(A[6]), .B(A[7]), .S(SH[0]), .Z(\MR_int[1][6] ) );
  MUX2_X1 M1_0_5_0 ( .A(A[5]), .B(A[6]), .S(SH[0]), .Z(\MR_int[1][5] ) );
  MUX2_X1 M1_0_4_0 ( .A(A[4]), .B(A[5]), .S(SH[0]), .Z(\MR_int[1][4] ) );
  MUX2_X1 M1_0_3_0 ( .A(A[3]), .B(A[4]), .S(SH[0]), .Z(\MR_int[1][3] ) );
  MUX2_X1 M1_0_2_0 ( .A(A[2]), .B(A[3]), .S(SH[0]), .Z(\MR_int[1][2] ) );
  MUX2_X1 M1_0_1_0 ( .A(A[1]), .B(A[2]), .S(SH[0]), .Z(\MR_int[1][1] ) );
  MUX2_X1 M1_0_0 ( .A(A[0]), .B(A[1]), .S(SH[0]), .Z(\MR_int[1][0] ) );
  CLKBUF_X3 U2 ( .A(SH[4]), .Z(n1) );
  CLKBUF_X3 U3 ( .A(SH[4]), .Z(n2) );
  CLKBUF_X3 U4 ( .A(SH[4]), .Z(n3) );
endmodule


module SHIFTER_GENERIC_N32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE, 
        OUTPUT );
  input [31:0] A;
  input [4:0] B;
  output [31:0] OUTPUT;
  input LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n1;

  NAND2_X1 U13 ( .A1(n19), .A2(n20), .ZN(OUTPUT[9]) );
  AOI222_X1 U14 ( .A1(N211), .A2(n21), .B1(N114), .B2(n22), .C1(N146), .C2(n23), .ZN(n20) );
  AOI222_X1 U15 ( .A1(N48), .A2(n24), .B1(N243), .B2(n25), .C1(N16), .C2(n26), 
        .ZN(n19) );
  NAND2_X1 U16 ( .A1(n27), .A2(n28), .ZN(OUTPUT[8]) );
  AOI222_X1 U17 ( .A1(N210), .A2(n21), .B1(N113), .B2(n22), .C1(N145), .C2(n23), .ZN(n28) );
  AOI222_X1 U18 ( .A1(N47), .A2(n24), .B1(N242), .B2(n25), .C1(N15), .C2(n26), 
        .ZN(n27) );
  NAND2_X1 U19 ( .A1(n29), .A2(n30), .ZN(OUTPUT[7]) );
  AOI222_X1 U20 ( .A1(N209), .A2(n21), .B1(N112), .B2(n22), .C1(N144), .C2(n23), .ZN(n30) );
  AOI222_X1 U21 ( .A1(N46), .A2(n24), .B1(N241), .B2(n25), .C1(N14), .C2(n26), 
        .ZN(n29) );
  NAND2_X1 U22 ( .A1(n31), .A2(n32), .ZN(OUTPUT[6]) );
  AOI222_X1 U23 ( .A1(N208), .A2(n21), .B1(N111), .B2(n22), .C1(N143), .C2(n23), .ZN(n32) );
  AOI222_X1 U24 ( .A1(N45), .A2(n24), .B1(N240), .B2(n25), .C1(N13), .C2(n26), 
        .ZN(n31) );
  NAND2_X1 U25 ( .A1(n33), .A2(n34), .ZN(OUTPUT[5]) );
  AOI222_X1 U26 ( .A1(N207), .A2(n21), .B1(N110), .B2(n22), .C1(N142), .C2(n23), .ZN(n34) );
  AOI222_X1 U27 ( .A1(N44), .A2(n24), .B1(N239), .B2(n25), .C1(N12), .C2(n26), 
        .ZN(n33) );
  NAND2_X1 U28 ( .A1(n35), .A2(n36), .ZN(OUTPUT[4]) );
  AOI222_X1 U29 ( .A1(N206), .A2(n21), .B1(N109), .B2(n22), .C1(N141), .C2(n23), .ZN(n36) );
  AOI222_X1 U30 ( .A1(N43), .A2(n24), .B1(N238), .B2(n25), .C1(N11), .C2(n26), 
        .ZN(n35) );
  NAND2_X1 U31 ( .A1(n37), .A2(n38), .ZN(OUTPUT[3]) );
  AOI222_X1 U32 ( .A1(N205), .A2(n21), .B1(N108), .B2(n22), .C1(N140), .C2(n23), .ZN(n38) );
  AOI222_X1 U33 ( .A1(N42), .A2(n24), .B1(N237), .B2(n25), .C1(N10), .C2(n26), 
        .ZN(n37) );
  NAND2_X1 U34 ( .A1(n39), .A2(n40), .ZN(OUTPUT[31]) );
  AOI222_X1 U35 ( .A1(N233), .A2(n21), .B1(N136), .B2(n22), .C1(N168), .C2(n23), .ZN(n40) );
  AOI222_X1 U36 ( .A1(N70), .A2(n24), .B1(N265), .B2(n25), .C1(N38), .C2(n26), 
        .ZN(n39) );
  NAND2_X1 U37 ( .A1(n41), .A2(n42), .ZN(OUTPUT[30]) );
  AOI222_X1 U38 ( .A1(N232), .A2(n21), .B1(N135), .B2(n22), .C1(N167), .C2(n23), .ZN(n42) );
  AOI222_X1 U39 ( .A1(N69), .A2(n24), .B1(N264), .B2(n25), .C1(N37), .C2(n26), 
        .ZN(n41) );
  NAND2_X1 U40 ( .A1(n43), .A2(n44), .ZN(OUTPUT[2]) );
  AOI222_X1 U41 ( .A1(N204), .A2(n21), .B1(N107), .B2(n22), .C1(N139), .C2(n23), .ZN(n44) );
  AOI222_X1 U42 ( .A1(N41), .A2(n24), .B1(N236), .B2(n25), .C1(N9), .C2(n26), 
        .ZN(n43) );
  NAND2_X1 U43 ( .A1(n45), .A2(n46), .ZN(OUTPUT[29]) );
  AOI222_X1 U44 ( .A1(N231), .A2(n21), .B1(N134), .B2(n22), .C1(N166), .C2(n23), .ZN(n46) );
  AOI222_X1 U45 ( .A1(N68), .A2(n24), .B1(N263), .B2(n25), .C1(N36), .C2(n26), 
        .ZN(n45) );
  NAND2_X1 U46 ( .A1(n47), .A2(n48), .ZN(OUTPUT[28]) );
  AOI222_X1 U47 ( .A1(N230), .A2(n21), .B1(N133), .B2(n22), .C1(N165), .C2(n23), .ZN(n48) );
  AOI222_X1 U48 ( .A1(N67), .A2(n24), .B1(N262), .B2(n25), .C1(N35), .C2(n26), 
        .ZN(n47) );
  NAND2_X1 U49 ( .A1(n49), .A2(n50), .ZN(OUTPUT[27]) );
  AOI222_X1 U50 ( .A1(N229), .A2(n21), .B1(N132), .B2(n22), .C1(N164), .C2(n23), .ZN(n50) );
  AOI222_X1 U51 ( .A1(N66), .A2(n24), .B1(N261), .B2(n25), .C1(N34), .C2(n26), 
        .ZN(n49) );
  NAND2_X1 U52 ( .A1(n51), .A2(n52), .ZN(OUTPUT[26]) );
  AOI222_X1 U53 ( .A1(N228), .A2(n21), .B1(N131), .B2(n22), .C1(N163), .C2(n23), .ZN(n52) );
  AOI222_X1 U54 ( .A1(N65), .A2(n24), .B1(N260), .B2(n25), .C1(N33), .C2(n26), 
        .ZN(n51) );
  NAND2_X1 U55 ( .A1(n53), .A2(n54), .ZN(OUTPUT[25]) );
  AOI222_X1 U56 ( .A1(N227), .A2(n21), .B1(N130), .B2(n22), .C1(N162), .C2(n23), .ZN(n54) );
  AOI222_X1 U57 ( .A1(N64), .A2(n24), .B1(N259), .B2(n25), .C1(N32), .C2(n26), 
        .ZN(n53) );
  NAND2_X1 U58 ( .A1(n55), .A2(n56), .ZN(OUTPUT[24]) );
  AOI222_X1 U59 ( .A1(N226), .A2(n21), .B1(N129), .B2(n22), .C1(N161), .C2(n23), .ZN(n56) );
  AOI222_X1 U60 ( .A1(N63), .A2(n24), .B1(N258), .B2(n25), .C1(N31), .C2(n26), 
        .ZN(n55) );
  NAND2_X1 U61 ( .A1(n57), .A2(n58), .ZN(OUTPUT[23]) );
  AOI222_X1 U62 ( .A1(N225), .A2(n21), .B1(N128), .B2(n22), .C1(N160), .C2(n23), .ZN(n58) );
  AOI222_X1 U63 ( .A1(N62), .A2(n24), .B1(N257), .B2(n25), .C1(N30), .C2(n26), 
        .ZN(n57) );
  NAND2_X1 U64 ( .A1(n59), .A2(n60), .ZN(OUTPUT[22]) );
  AOI222_X1 U65 ( .A1(N224), .A2(n21), .B1(N127), .B2(n22), .C1(N159), .C2(n23), .ZN(n60) );
  AOI222_X1 U66 ( .A1(N61), .A2(n24), .B1(N256), .B2(n25), .C1(N29), .C2(n26), 
        .ZN(n59) );
  NAND2_X1 U67 ( .A1(n61), .A2(n62), .ZN(OUTPUT[21]) );
  AOI222_X1 U68 ( .A1(N223), .A2(n21), .B1(N126), .B2(n22), .C1(N158), .C2(n23), .ZN(n62) );
  AOI222_X1 U69 ( .A1(N60), .A2(n24), .B1(N255), .B2(n25), .C1(N28), .C2(n26), 
        .ZN(n61) );
  NAND2_X1 U70 ( .A1(n63), .A2(n64), .ZN(OUTPUT[20]) );
  AOI222_X1 U71 ( .A1(N222), .A2(n21), .B1(N125), .B2(n22), .C1(N157), .C2(n23), .ZN(n64) );
  AOI222_X1 U72 ( .A1(N59), .A2(n24), .B1(N254), .B2(n25), .C1(N27), .C2(n26), 
        .ZN(n63) );
  NAND2_X1 U73 ( .A1(n65), .A2(n66), .ZN(OUTPUT[1]) );
  AOI222_X1 U74 ( .A1(N203), .A2(n21), .B1(N106), .B2(n22), .C1(N138), .C2(n23), .ZN(n66) );
  AOI222_X1 U75 ( .A1(N40), .A2(n24), .B1(N235), .B2(n25), .C1(N8), .C2(n26), 
        .ZN(n65) );
  NAND2_X1 U76 ( .A1(n67), .A2(n68), .ZN(OUTPUT[19]) );
  AOI222_X1 U77 ( .A1(N221), .A2(n21), .B1(N124), .B2(n22), .C1(N156), .C2(n23), .ZN(n68) );
  AOI222_X1 U78 ( .A1(N58), .A2(n24), .B1(N253), .B2(n25), .C1(N26), .C2(n26), 
        .ZN(n67) );
  NAND2_X1 U79 ( .A1(n69), .A2(n70), .ZN(OUTPUT[18]) );
  AOI222_X1 U80 ( .A1(N220), .A2(n21), .B1(N123), .B2(n22), .C1(N155), .C2(n23), .ZN(n70) );
  AOI222_X1 U81 ( .A1(N57), .A2(n24), .B1(N252), .B2(n25), .C1(N25), .C2(n26), 
        .ZN(n69) );
  NAND2_X1 U82 ( .A1(n71), .A2(n72), .ZN(OUTPUT[17]) );
  AOI222_X1 U83 ( .A1(N219), .A2(n21), .B1(N122), .B2(n22), .C1(N154), .C2(n23), .ZN(n72) );
  AOI222_X1 U84 ( .A1(N56), .A2(n24), .B1(N251), .B2(n25), .C1(N24), .C2(n26), 
        .ZN(n71) );
  NAND2_X1 U85 ( .A1(n73), .A2(n74), .ZN(OUTPUT[16]) );
  AOI222_X1 U86 ( .A1(N218), .A2(n21), .B1(N121), .B2(n22), .C1(N153), .C2(n23), .ZN(n74) );
  AOI222_X1 U87 ( .A1(N55), .A2(n24), .B1(N250), .B2(n25), .C1(N23), .C2(n26), 
        .ZN(n73) );
  NAND2_X1 U88 ( .A1(n75), .A2(n76), .ZN(OUTPUT[15]) );
  AOI222_X1 U89 ( .A1(N217), .A2(n21), .B1(N120), .B2(n22), .C1(N152), .C2(n23), .ZN(n76) );
  AOI222_X1 U90 ( .A1(N54), .A2(n24), .B1(N249), .B2(n25), .C1(N22), .C2(n26), 
        .ZN(n75) );
  NAND2_X1 U91 ( .A1(n77), .A2(n78), .ZN(OUTPUT[14]) );
  AOI222_X1 U92 ( .A1(N216), .A2(n21), .B1(N119), .B2(n22), .C1(N151), .C2(n23), .ZN(n78) );
  AOI222_X1 U93 ( .A1(N53), .A2(n24), .B1(N248), .B2(n25), .C1(N21), .C2(n26), 
        .ZN(n77) );
  NAND2_X1 U94 ( .A1(n79), .A2(n80), .ZN(OUTPUT[13]) );
  AOI222_X1 U95 ( .A1(N215), .A2(n21), .B1(N118), .B2(n22), .C1(N150), .C2(n23), .ZN(n80) );
  AOI222_X1 U96 ( .A1(N52), .A2(n24), .B1(N247), .B2(n25), .C1(N20), .C2(n26), 
        .ZN(n79) );
  NAND2_X1 U97 ( .A1(n81), .A2(n82), .ZN(OUTPUT[12]) );
  AOI222_X1 U98 ( .A1(N214), .A2(n21), .B1(N117), .B2(n22), .C1(N149), .C2(n23), .ZN(n82) );
  AOI222_X1 U99 ( .A1(N51), .A2(n24), .B1(N246), .B2(n25), .C1(N19), .C2(n26), 
        .ZN(n81) );
  NAND2_X1 U100 ( .A1(n83), .A2(n84), .ZN(OUTPUT[11]) );
  AOI222_X1 U101 ( .A1(N213), .A2(n21), .B1(N116), .B2(n22), .C1(N148), .C2(
        n23), .ZN(n84) );
  AOI222_X1 U102 ( .A1(N50), .A2(n24), .B1(N245), .B2(n25), .C1(N18), .C2(n26), 
        .ZN(n83) );
  NAND2_X1 U103 ( .A1(n85), .A2(n86), .ZN(OUTPUT[10]) );
  AOI222_X1 U104 ( .A1(N212), .A2(n21), .B1(N115), .B2(n22), .C1(N147), .C2(
        n23), .ZN(n86) );
  AOI222_X1 U105 ( .A1(N49), .A2(n24), .B1(N244), .B2(n25), .C1(N17), .C2(n26), 
        .ZN(n85) );
  NAND2_X1 U106 ( .A1(n87), .A2(n88), .ZN(OUTPUT[0]) );
  AOI222_X1 U107 ( .A1(N202), .A2(n21), .B1(N105), .B2(n22), .C1(N137), .C2(
        n23), .ZN(n88) );
  NOR2_X1 U111 ( .A1(n92), .A2(LOGIC_ARITH), .ZN(n91) );
  INV_X1 U112 ( .A(SHIFT_ROTATE), .ZN(n92) );
  AOI222_X1 U113 ( .A1(N39), .A2(n24), .B1(N234), .B2(n25), .C1(N7), .C2(n26), 
        .ZN(n87) );
  AND2_X1 U116 ( .A1(LOGIC_ARITH), .A2(SHIFT_ROTATE), .ZN(n89) );
  INV_X1 U118 ( .A(LEFT_RIGHT), .ZN(n90) );
  SHIFTER_GENERIC_N32_DW01_ash_0 sll_49 ( .A(A), .DATA_TC(1'b0), .SH({n1, 
        B[3:0]}), .SH_TC(1'b0), .B({N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234}) );
  SHIFTER_GENERIC_N32_DW_sla_0 sla_47 ( .A(A), .SH({n1, B[3:0]}), .SH_TC(1'b0), 
        .B({N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, 
        N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, 
        N210, N209, N208, N207, N206, N205, N204, N203, N202}) );
  SHIFTER_GENERIC_N32_DW_rash_0 srl_42 ( .A(A), .DATA_TC(1'b0), .SH({n1, 
        B[3:0]}), .SH_TC(1'b0), .B({N168, N167, N166, N165, N164, N163, N162, 
        N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, 
        N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, 
        N137}) );
  SHIFTER_GENERIC_N32_DW_sra_0 sra_40 ( .A(A), .SH({n1, B[3:0]}), .SH_TC(1'b0), 
        .B({N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, 
        N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, 
        N113, N112, N111, N110, N109, N108, N107, N106, N105}) );
  SHIFTER_GENERIC_N32_DW_lbsh_0 rol_33 ( .A(A), .SH({n1, B[3:0]}), .SH_TC(1'b0), .B({N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39}) );
  SHIFTER_GENERIC_N32_DW_rbsh_0 ror_31 ( .A(A), .SH({n1, B[3:0]}), .SH_TC(1'b0), .B({N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7}) );
  AND2_X2 U5 ( .A1(n89), .A2(n90), .ZN(n23) );
  AND2_X2 U6 ( .A1(n91), .A2(n90), .ZN(n22) );
  AND2_X2 U7 ( .A1(LEFT_RIGHT), .A2(n89), .ZN(n25) );
  AND2_X2 U8 ( .A1(LEFT_RIGHT), .A2(n91), .ZN(n21) );
  NOR2_X4 U9 ( .A1(n90), .A2(SHIFT_ROTATE), .ZN(n24) );
  NOR2_X4 U10 ( .A1(LEFT_RIGHT), .A2(SHIFT_ROTATE), .ZN(n26) );
  BUF_X4 U108 ( .A(B[4]), .Z(n1) );
endmodule


module G_0 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n1) );
endmodule


module G_43 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_0 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_0 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_43 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_0 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_52 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_42 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_42 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_42 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_42 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_42 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_41 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_41 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_41 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_41 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_41 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_40 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_40 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_40 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_40 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_40 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_39 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_39 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_39 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_39 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_39 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_38 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_38 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_38 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_38 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_38 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_37 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_37 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_37 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_37 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_37 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_36 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_36 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_36 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_36 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_36 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_35 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_35 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_35 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_35 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_35 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_34 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_34 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_34 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_34 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_34 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_33 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_33 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_33 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_33 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_33 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_32 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_32 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_32 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_32 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_32 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_31 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_31 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_31 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_31 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_31 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_30 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_30 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_30 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_30 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_30 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_29 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_29 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_29 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_29 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_29 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_28 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_28 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_28 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_28 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_28 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_27 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_27 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_27 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_27 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_27 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_26 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_26 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_26 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_26 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_26 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_25 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_25 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_25 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_25 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_25 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_24 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_24 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_24 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_24 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_24 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_23 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_23 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_23 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_23 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_23 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_22 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_22 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_22 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_22 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_22 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_21 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_21 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_21 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_21 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_21 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_20 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_20 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_20 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_20 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_20 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_19 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_19 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_19 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_19 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_19 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_18 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_18 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_18 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_18 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_18 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_17 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_17 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_17 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_17 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_17 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_16 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_16 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_16 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_16 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_16 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_15 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_15 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_15 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_15 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_15 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_14 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_14 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_14 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_14 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_14 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_13 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_13 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_13 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_13 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_13 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_51 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_12 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_12 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_12 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_12 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_12 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_11 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_11 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_11 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_11 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_11 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_10 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_10 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_10 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_10 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_10 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_9 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_9 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_9 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_9 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_9 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_8 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_8 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_8 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_8 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_8 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_7 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_7 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_7 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_7 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_7 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_6 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_6 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_6 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_6 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_6 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_50 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_5 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_5 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_5 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_5 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_5 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_4 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_4 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_4 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_4 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_4 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_3 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_3 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_3 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_3 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_3 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_49 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_48 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_2 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_2 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_2 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_2 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_2 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_1 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module P_1 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_1 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_1 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_1 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_47 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_46 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_45 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_44 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   \gi[32][4] , \gi[32][3] , \gi[32][2] , \gi[32][1] , \gi[32][0] ,
         \gi[31][0] , \gi[30][0] , \gi[29][0] , \gi[28][4] , \gi[28][2] ,
         \gi[28][1] , \gi[28][0] , \gi[27][0] , \gi[26][0] , \gi[25][0] ,
         \gi[24][3] , \gi[24][2] , \gi[24][1] , \gi[24][0] , \gi[23][0] ,
         \gi[22][0] , \gi[21][0] , \gi[20][2] , \gi[20][1] , \gi[20][0] ,
         \gi[19][0] , \gi[18][0] , \gi[17][0] , \gi[16][3] , \gi[16][2] ,
         \gi[16][1] , \gi[16][0] , \gi[15][0] , \gi[14][0] , \gi[13][0] ,
         \gi[12][2] , \gi[12][1] , \gi[12][0] , \gi[11][0] , \gi[10][0] ,
         \gi[9][0] , \gi[8][2] , \gi[8][1] , \gi[8][0] , \gi[7][0] ,
         \gi[6][0] , \gi[5][0] , \gi[4][1] , \gi[4][0] , \gi[3][0] ,
         \gi[2][1] , \gi[2][0] , \gi[1][0] , \gi[0][0] , \pi[32][4] ,
         \pi[32][3] , \pi[32][2] , \pi[32][1] , \pi[32][0] , \pi[31][0] ,
         \pi[30][0] , \pi[29][0] , \pi[28][4] , \pi[28][2] , \pi[28][1] ,
         \pi[28][0] , \pi[27][0] , \pi[26][0] , \pi[25][0] , \pi[24][3] ,
         \pi[24][2] , \pi[24][1] , \pi[24][0] , \pi[23][0] , \pi[22][0] ,
         \pi[21][0] , \pi[20][2] , \pi[20][1] , \pi[20][0] , \pi[19][0] ,
         \pi[18][0] , \pi[17][0] , \pi[16][3] , \pi[16][2] , \pi[16][1] ,
         \pi[16][0] , \pi[15][0] , \pi[14][0] , \pi[13][0] , \pi[12][2] ,
         \pi[12][1] , \pi[12][0] , \pi[11][0] , \pi[10][0] , \pi[9][0] ,
         \pi[8][2] , \pi[8][1] , \pi[8][0] , \pi[7][0] , \pi[6][0] ,
         \pi[5][0] , \pi[4][1] , \pi[4][0] , \pi[3][0] , \pi[2][0] ,
         \pi[0][0] ;

  XOR2_X1 U2 ( .A(B[8]), .B(A[8]), .Z(\pi[9][0] ) );
  XOR2_X1 U3 ( .A(B[7]), .B(A[7]), .Z(\pi[8][0] ) );
  XOR2_X1 U4 ( .A(B[6]), .B(A[6]), .Z(\pi[7][0] ) );
  XOR2_X1 U5 ( .A(B[5]), .B(A[5]), .Z(\pi[6][0] ) );
  XOR2_X1 U6 ( .A(B[4]), .B(A[4]), .Z(\pi[5][0] ) );
  XOR2_X1 U7 ( .A(B[3]), .B(A[3]), .Z(\pi[4][0] ) );
  XOR2_X1 U8 ( .A(B[2]), .B(A[2]), .Z(\pi[3][0] ) );
  XOR2_X1 U9 ( .A(B[31]), .B(A[31]), .Z(\pi[32][0] ) );
  XOR2_X1 U10 ( .A(B[30]), .B(A[30]), .Z(\pi[31][0] ) );
  XOR2_X1 U11 ( .A(B[29]), .B(A[29]), .Z(\pi[30][0] ) );
  XOR2_X1 U12 ( .A(B[1]), .B(A[1]), .Z(\pi[2][0] ) );
  XOR2_X1 U13 ( .A(B[28]), .B(A[28]), .Z(\pi[29][0] ) );
  XOR2_X1 U14 ( .A(B[27]), .B(A[27]), .Z(\pi[28][0] ) );
  XOR2_X1 U15 ( .A(B[26]), .B(A[26]), .Z(\pi[27][0] ) );
  XOR2_X1 U16 ( .A(B[25]), .B(A[25]), .Z(\pi[26][0] ) );
  XOR2_X1 U17 ( .A(B[24]), .B(A[24]), .Z(\pi[25][0] ) );
  XOR2_X1 U18 ( .A(B[23]), .B(A[23]), .Z(\pi[24][0] ) );
  XOR2_X1 U19 ( .A(B[22]), .B(A[22]), .Z(\pi[23][0] ) );
  XOR2_X1 U20 ( .A(B[21]), .B(A[21]), .Z(\pi[22][0] ) );
  XOR2_X1 U21 ( .A(B[20]), .B(A[20]), .Z(\pi[21][0] ) );
  XOR2_X1 U22 ( .A(B[19]), .B(A[19]), .Z(\pi[20][0] ) );
  XOR2_X1 U23 ( .A(B[18]), .B(A[18]), .Z(\pi[19][0] ) );
  XOR2_X1 U24 ( .A(B[17]), .B(A[17]), .Z(\pi[18][0] ) );
  XOR2_X1 U25 ( .A(B[16]), .B(A[16]), .Z(\pi[17][0] ) );
  XOR2_X1 U26 ( .A(B[15]), .B(A[15]), .Z(\pi[16][0] ) );
  XOR2_X1 U27 ( .A(B[14]), .B(A[14]), .Z(\pi[15][0] ) );
  XOR2_X1 U28 ( .A(B[13]), .B(A[13]), .Z(\pi[14][0] ) );
  XOR2_X1 U29 ( .A(B[12]), .B(A[12]), .Z(\pi[13][0] ) );
  XOR2_X1 U30 ( .A(B[11]), .B(A[11]), .Z(\pi[12][0] ) );
  XOR2_X1 U31 ( .A(B[10]), .B(A[10]), .Z(\pi[11][0] ) );
  XOR2_X1 U32 ( .A(B[9]), .B(A[9]), .Z(\pi[10][0] ) );
  XOR2_X1 U33 ( .A(B[0]), .B(A[0]), .Z(\pi[0][0] ) );
  AND2_X1 U34 ( .A1(B[8]), .A2(A[8]), .ZN(\gi[9][0] ) );
  AND2_X1 U35 ( .A1(B[7]), .A2(A[7]), .ZN(\gi[8][0] ) );
  AND2_X1 U36 ( .A1(B[6]), .A2(A[6]), .ZN(\gi[7][0] ) );
  AND2_X1 U37 ( .A1(B[5]), .A2(A[5]), .ZN(\gi[6][0] ) );
  AND2_X1 U38 ( .A1(B[4]), .A2(A[4]), .ZN(\gi[5][0] ) );
  AND2_X1 U39 ( .A1(B[3]), .A2(A[3]), .ZN(\gi[4][0] ) );
  AND2_X1 U40 ( .A1(B[2]), .A2(A[2]), .ZN(\gi[3][0] ) );
  AND2_X1 U41 ( .A1(B[31]), .A2(A[31]), .ZN(\gi[32][0] ) );
  AND2_X1 U42 ( .A1(B[30]), .A2(A[30]), .ZN(\gi[31][0] ) );
  AND2_X1 U43 ( .A1(B[29]), .A2(A[29]), .ZN(\gi[30][0] ) );
  AND2_X1 U44 ( .A1(B[1]), .A2(A[1]), .ZN(\gi[2][0] ) );
  AND2_X1 U45 ( .A1(B[28]), .A2(A[28]), .ZN(\gi[29][0] ) );
  AND2_X1 U46 ( .A1(B[27]), .A2(A[27]), .ZN(\gi[28][0] ) );
  AND2_X1 U47 ( .A1(B[26]), .A2(A[26]), .ZN(\gi[27][0] ) );
  AND2_X1 U48 ( .A1(B[25]), .A2(A[25]), .ZN(\gi[26][0] ) );
  AND2_X1 U49 ( .A1(B[24]), .A2(A[24]), .ZN(\gi[25][0] ) );
  AND2_X1 U50 ( .A1(B[23]), .A2(A[23]), .ZN(\gi[24][0] ) );
  AND2_X1 U51 ( .A1(B[22]), .A2(A[22]), .ZN(\gi[23][0] ) );
  AND2_X1 U52 ( .A1(B[21]), .A2(A[21]), .ZN(\gi[22][0] ) );
  AND2_X1 U53 ( .A1(B[20]), .A2(A[20]), .ZN(\gi[21][0] ) );
  AND2_X1 U54 ( .A1(B[19]), .A2(A[19]), .ZN(\gi[20][0] ) );
  AND2_X1 U55 ( .A1(B[18]), .A2(A[18]), .ZN(\gi[19][0] ) );
  AND2_X1 U56 ( .A1(B[17]), .A2(A[17]), .ZN(\gi[18][0] ) );
  AND2_X1 U57 ( .A1(B[16]), .A2(A[16]), .ZN(\gi[17][0] ) );
  AND2_X1 U58 ( .A1(B[15]), .A2(A[15]), .ZN(\gi[16][0] ) );
  AND2_X1 U59 ( .A1(B[14]), .A2(A[14]), .ZN(\gi[15][0] ) );
  AND2_X1 U60 ( .A1(B[13]), .A2(A[13]), .ZN(\gi[14][0] ) );
  AND2_X1 U61 ( .A1(B[12]), .A2(A[12]), .ZN(\gi[13][0] ) );
  AND2_X1 U62 ( .A1(B[11]), .A2(A[11]), .ZN(\gi[12][0] ) );
  AND2_X1 U63 ( .A1(B[10]), .A2(A[10]), .ZN(\gi[11][0] ) );
  AND2_X1 U64 ( .A1(B[9]), .A2(A[9]), .ZN(\gi[10][0] ) );
  AND2_X1 U65 ( .A1(B[0]), .A2(A[0]), .ZN(\gi[0][0] ) );
  G_0 g_port0_0_1 ( .G1(\gi[0][0] ), .P(\pi[0][0] ), .G2(Cin), .Co(\gi[1][0] )
         );
  PG_0 pg_port2_1_1 ( .G1(\gi[1][0] ), .P1(1'b0), .G2(\gi[0][0] ), .P2(
        \pi[0][0] ) );
  G_52 g_port1_1_2 ( .G1(\gi[2][0] ), .P(\pi[2][0] ), .G2(\gi[1][0] ), .Co(
        \gi[2][1] ) );
  PG_42 pg_port2_1_3 ( .G1(\gi[3][0] ), .P1(\pi[3][0] ), .G2(\gi[2][0] ), .P2(
        \pi[2][0] ) );
  PG_41 pg_port2_1_4 ( .G1(\gi[4][0] ), .P1(\pi[4][0] ), .G2(\gi[3][0] ), .P2(
        \pi[3][0] ), .gout(\gi[4][1] ), .pout(\pi[4][1] ) );
  PG_40 pg_port2_1_5 ( .G1(\gi[5][0] ), .P1(\pi[5][0] ), .G2(\gi[4][0] ), .P2(
        \pi[4][0] ) );
  PG_39 pg_port2_1_6 ( .G1(\gi[6][0] ), .P1(\pi[6][0] ), .G2(\gi[5][0] ), .P2(
        \pi[5][0] ) );
  PG_38 pg_port2_1_7 ( .G1(\gi[7][0] ), .P1(\pi[7][0] ), .G2(\gi[6][0] ), .P2(
        \pi[6][0] ) );
  PG_37 pg_port2_1_8 ( .G1(\gi[8][0] ), .P1(\pi[8][0] ), .G2(\gi[7][0] ), .P2(
        \pi[7][0] ), .gout(\gi[8][1] ), .pout(\pi[8][1] ) );
  PG_36 pg_port2_1_9 ( .G1(\gi[9][0] ), .P1(\pi[9][0] ), .G2(\gi[8][0] ), .P2(
        \pi[8][0] ) );
  PG_35 pg_port2_1_10 ( .G1(\gi[10][0] ), .P1(\pi[10][0] ), .G2(\gi[9][0] ), 
        .P2(\pi[9][0] ) );
  PG_34 pg_port2_1_11 ( .G1(\gi[11][0] ), .P1(\pi[11][0] ), .G2(\gi[10][0] ), 
        .P2(\pi[10][0] ) );
  PG_33 pg_port2_1_12 ( .G1(\gi[12][0] ), .P1(\pi[12][0] ), .G2(\gi[11][0] ), 
        .P2(\pi[11][0] ), .gout(\gi[12][1] ), .pout(\pi[12][1] ) );
  PG_32 pg_port2_1_13 ( .G1(\gi[13][0] ), .P1(\pi[13][0] ), .G2(\gi[12][0] ), 
        .P2(\pi[12][0] ) );
  PG_31 pg_port2_1_14 ( .G1(\gi[14][0] ), .P1(\pi[14][0] ), .G2(\gi[13][0] ), 
        .P2(\pi[13][0] ) );
  PG_30 pg_port2_1_15 ( .G1(\gi[15][0] ), .P1(\pi[15][0] ), .G2(\gi[14][0] ), 
        .P2(\pi[14][0] ) );
  PG_29 pg_port2_1_16 ( .G1(\gi[16][0] ), .P1(\pi[16][0] ), .G2(\gi[15][0] ), 
        .P2(\pi[15][0] ), .gout(\gi[16][1] ), .pout(\pi[16][1] ) );
  PG_28 pg_port2_1_17 ( .G1(\gi[17][0] ), .P1(\pi[17][0] ), .G2(\gi[16][0] ), 
        .P2(\pi[16][0] ) );
  PG_27 pg_port2_1_18 ( .G1(\gi[18][0] ), .P1(\pi[18][0] ), .G2(\gi[17][0] ), 
        .P2(\pi[17][0] ) );
  PG_26 pg_port2_1_19 ( .G1(\gi[19][0] ), .P1(\pi[19][0] ), .G2(\gi[18][0] ), 
        .P2(\pi[18][0] ) );
  PG_25 pg_port2_1_20 ( .G1(\gi[20][0] ), .P1(\pi[20][0] ), .G2(\gi[19][0] ), 
        .P2(\pi[19][0] ), .gout(\gi[20][1] ), .pout(\pi[20][1] ) );
  PG_24 pg_port2_1_21 ( .G1(\gi[21][0] ), .P1(\pi[21][0] ), .G2(\gi[20][0] ), 
        .P2(\pi[20][0] ) );
  PG_23 pg_port2_1_22 ( .G1(\gi[22][0] ), .P1(\pi[22][0] ), .G2(\gi[21][0] ), 
        .P2(\pi[21][0] ) );
  PG_22 pg_port2_1_23 ( .G1(\gi[23][0] ), .P1(\pi[23][0] ), .G2(\gi[22][0] ), 
        .P2(\pi[22][0] ) );
  PG_21 pg_port2_1_24 ( .G1(\gi[24][0] ), .P1(\pi[24][0] ), .G2(\gi[23][0] ), 
        .P2(\pi[23][0] ), .gout(\gi[24][1] ), .pout(\pi[24][1] ) );
  PG_20 pg_port2_1_25 ( .G1(\gi[25][0] ), .P1(\pi[25][0] ), .G2(\gi[24][0] ), 
        .P2(\pi[24][0] ) );
  PG_19 pg_port2_1_26 ( .G1(\gi[26][0] ), .P1(\pi[26][0] ), .G2(\gi[25][0] ), 
        .P2(\pi[25][0] ) );
  PG_18 pg_port2_1_27 ( .G1(\gi[27][0] ), .P1(\pi[27][0] ), .G2(\gi[26][0] ), 
        .P2(\pi[26][0] ) );
  PG_17 pg_port2_1_28 ( .G1(\gi[28][0] ), .P1(\pi[28][0] ), .G2(\gi[27][0] ), 
        .P2(\pi[27][0] ), .gout(\gi[28][1] ), .pout(\pi[28][1] ) );
  PG_16 pg_port2_1_29 ( .G1(\gi[29][0] ), .P1(\pi[29][0] ), .G2(\gi[28][0] ), 
        .P2(\pi[28][0] ) );
  PG_15 pg_port2_1_30 ( .G1(\gi[30][0] ), .P1(\pi[30][0] ), .G2(\gi[29][0] ), 
        .P2(\pi[29][0] ) );
  PG_14 pg_port2_1_31 ( .G1(\gi[31][0] ), .P1(\pi[31][0] ), .G2(\gi[30][0] ), 
        .P2(\pi[30][0] ) );
  PG_13 pg_port2_1_32 ( .G1(\gi[32][0] ), .P1(\pi[32][0] ), .G2(\gi[31][0] ), 
        .P2(\pi[31][0] ), .gout(\gi[32][1] ), .pout(\pi[32][1] ) );
  G_51 g_port_0 ( .G1(\gi[4][1] ), .P(\pi[4][1] ), .G2(\gi[2][1] ), .Co(Co[0])
         );
  PG_12 pg_port2_0_1_2 ( .G1(\gi[8][1] ), .P1(\pi[8][1] ), .G2(\gi[4][1] ), 
        .P2(\pi[4][1] ), .gout(\gi[8][2] ), .pout(\pi[8][2] ) );
  PG_11 pg_port2_0_2_3 ( .G1(\gi[12][1] ), .P1(\pi[12][1] ), .G2(\gi[8][1] ), 
        .P2(\pi[8][1] ), .gout(\gi[12][2] ), .pout(\pi[12][2] ) );
  PG_10 pg_port2_0_3_4 ( .G1(\gi[16][1] ), .P1(\pi[16][1] ), .G2(\gi[12][1] ), 
        .P2(\pi[12][1] ), .gout(\gi[16][2] ), .pout(\pi[16][2] ) );
  PG_9 pg_port2_0_4_5 ( .G1(\gi[20][1] ), .P1(\pi[20][1] ), .G2(\gi[16][1] ), 
        .P2(\pi[16][1] ), .gout(\gi[20][2] ), .pout(\pi[20][2] ) );
  PG_8 pg_port2_0_5_6 ( .G1(\gi[24][1] ), .P1(\pi[24][1] ), .G2(\gi[20][1] ), 
        .P2(\pi[20][1] ), .gout(\gi[24][2] ), .pout(\pi[24][2] ) );
  PG_7 pg_port2_0_6_7 ( .G1(\gi[28][1] ), .P1(\pi[28][1] ), .G2(\gi[24][1] ), 
        .P2(\pi[24][1] ), .gout(\gi[28][2] ), .pout(\pi[28][2] ) );
  PG_6 pg_port2_0_7_8 ( .G1(\gi[32][1] ), .P1(\pi[32][1] ), .G2(\gi[28][1] ), 
        .P2(\pi[28][1] ), .gout(\gi[32][2] ), .pout(\pi[32][2] ) );
  G_50 g_port_1_2 ( .G1(\gi[8][2] ), .P(\pi[8][2] ), .G2(Co[0]), .Co(Co[1]) );
  PG_5 pg_port2_1_1_4 ( .G1(\gi[16][2] ), .P1(\pi[16][2] ), .G2(\gi[12][2] ), 
        .P2(\pi[12][2] ), .gout(\gi[16][3] ), .pout(\pi[16][3] ) );
  PG_4 pg_port2_1_2_6 ( .G1(\gi[24][2] ), .P1(\pi[24][2] ), .G2(\gi[20][2] ), 
        .P2(\pi[20][2] ), .gout(\gi[24][3] ), .pout(\pi[24][3] ) );
  PG_3 pg_port2_1_3_8 ( .G1(\gi[32][2] ), .P1(\pi[32][2] ), .G2(\gi[28][2] ), 
        .P2(\pi[28][2] ), .gout(\gi[32][3] ), .pout(\pi[32][3] ) );
  G_49 g_port_2_3 ( .G1(\gi[12][2] ), .P(\pi[12][2] ), .G2(Co[1]), .Co(Co[2])
         );
  G_48 g_port_2_4 ( .G1(\gi[16][3] ), .P(\pi[16][3] ), .G2(Co[1]), .Co(Co[3])
         );
  PG_2 pg_port2_2_1_7 ( .G1(\gi[28][2] ), .P1(\pi[28][2] ), .G2(\gi[24][3] ), 
        .P2(\pi[24][3] ), .gout(\gi[28][4] ), .pout(\pi[28][4] ) );
  PG_1 pg_port2_2_1_8 ( .G1(\gi[32][3] ), .P1(\pi[32][3] ), .G2(\gi[24][3] ), 
        .P2(\pi[24][3] ), .gout(\gi[32][4] ), .pout(\pi[32][4] ) );
  G_47 g_port_3_5 ( .G1(\gi[20][2] ), .P(\pi[20][2] ), .G2(Co[3]), .Co(Co[4])
         );
  G_46 g_port_3_6 ( .G1(\gi[24][3] ), .P(\pi[24][3] ), .G2(Co[3]), .Co(Co[5])
         );
  G_45 g_port_3_7 ( .G1(\gi[28][4] ), .P(\pi[28][4] ), .G2(Co[3]), .Co(Co[6])
         );
  G_44 g_port_3_8 ( .G1(\gi[32][4] ), .P(\pi[32][4] ), .G2(Co[3]), .Co(Co[7])
         );
endmodule


module RCA_NBIT4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_32 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_32 UIV ( .A(S), .Y(SB) );
  ND2_96 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_95 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_94 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31 UIV ( .A(S), .Y(SB) );
  ND2_93 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_92 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_91 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30 UIV ( .A(S), .Y(SB) );
  ND2_90 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_89 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_88 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_29 UIV ( .A(S), .Y(SB) );
  ND2_87 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_86 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_85 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_32 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_29 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_0 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_28 UIV ( .A(S), .Y(SB) );
  ND2_84 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_83 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_82 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_27 UIV ( .A(S), .Y(SB) );
  ND2_81 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_80 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_79 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_26 UIV ( .A(S), .Y(SB) );
  ND2_78 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_77 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_76 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_25 UIV ( .A(S), .Y(SB) );
  ND2_75 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_74 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_73 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_28 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_27 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_26 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_25 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_7 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_24 UIV ( .A(S), .Y(SB) );
  ND2_72 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_71 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_70 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_23 UIV ( .A(S), .Y(SB) );
  ND2_69 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_68 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_67 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_22 UIV ( .A(S), .Y(SB) );
  ND2_66 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_65 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_64 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_21 UIV ( .A(S), .Y(SB) );
  ND2_63 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_62 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_61 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_24 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_23 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_22 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_21 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_6 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_20 UIV ( .A(S), .Y(SB) );
  ND2_60 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_59 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_58 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_19 UIV ( .A(S), .Y(SB) );
  ND2_57 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_56 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_55 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_18 UIV ( .A(S), .Y(SB) );
  ND2_54 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_53 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_52 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_17 UIV ( .A(S), .Y(SB) );
  ND2_51 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_50 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_49 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_20 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_19 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_18 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_17 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_5 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_16 UIV ( .A(S), .Y(SB) );
  ND2_48 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_47 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_46 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_15 UIV ( .A(S), .Y(SB) );
  ND2_45 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_44 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_43 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_14 UIV ( .A(S), .Y(SB) );
  ND2_42 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_41 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_40 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_13 UIV ( .A(S), .Y(SB) );
  ND2_39 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_38 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_37 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_16 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_15 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_14 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_13 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_4 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_12 UIV ( .A(S), .Y(SB) );
  ND2_36 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_35 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_34 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_11 UIV ( .A(S), .Y(SB) );
  ND2_33 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_32 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_31 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_10 UIV ( .A(S), .Y(SB) );
  ND2_30 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_29 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_28 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_9 UIV ( .A(S), .Y(SB) );
  ND2_27 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_26 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_25 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_12 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_11 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_10 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_9 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_3 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_8 UIV ( .A(S), .Y(SB) );
  ND2_24 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_23 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_22 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_7 UIV ( .A(S), .Y(SB) );
  ND2_21 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_20 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_19 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_6 UIV ( .A(S), .Y(SB) );
  ND2_18 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_17 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_16 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_5 UIV ( .A(S), .Y(SB) );
  ND2_15 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_14 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_13 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_8 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_7 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_6 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_5 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_2 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_4 UIV ( .A(S), .Y(SB) );
  ND2_12 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_11 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_10 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_3 UIV ( .A(S), .Y(SB) );
  ND2_9 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_8 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_7 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_2 UIV ( .A(S), .Y(SB) );
  ND2_6 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_5 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_4 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_1 UIV ( .A(S), .Y(SB) );
  ND2_3 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_2 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_1 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_4 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_3 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_2 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_1 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_1 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSB_NBIT4_0 CSBI_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSB_NBIT4_7 CSBI_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSB_NBIT4_6 CSBI_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  CSB_NBIT4_5 CSBI_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(S[15:12]) );
  CSB_NBIT4_4 CSBI_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(S[19:16]) );
  CSB_NBIT4_3 CSBI_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(S[23:20]) );
  CSB_NBIT4_2 CSBI_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(S[27:24]) );
  CSB_NBIT4_1 CSBI_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28]) );
endmodule


module P4_ADDER_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [6:0] Cout_gen;

  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 carry_logic ( .A(A), .B(B), .Cin(Cin), 
        .Co({Cout, Cout_gen}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 sum_logic ( .A(A), .B(B), .Ci({
        Cout_gen, Cin}), .S(S) );
endmodule


module ALU_N32 ( CLK, .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , 
        \FUNC[1] , \FUNC[0] }), DATA1, DATA2, OUT_ALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUT_ALU;
  input CLK, \FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   Cout_i, \OUTPUT3[0] , LOGIC_ARITH_i, LEFT_RIGHT_i, Cin_i, N139, N140,
         N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151,
         N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162,
         N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173,
         N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184,
         N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159;
  wire   [5:0] FUNC;
  wire   [31:0] OUTPUT_alu_i;
  wire   [31:0] OUTPUT4;
  wire   [31:0] OUTPUT2;
  wire   [31:0] OUTPUT1;
  wire   [31:0] data1i;
  wire   [31:0] data2i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  DLH_X1 Cin_i_reg ( .G(n155), .D(N140), .Q(Cin_i) );
  DLH_X1 \data2i_reg[31]  ( .G(n155), .D(N205), .Q(data2i[31]) );
  DLH_X1 \data2i_reg[30]  ( .G(n155), .D(N204), .Q(data2i[30]) );
  DLH_X1 \data2i_reg[29]  ( .G(n155), .D(N203), .Q(data2i[29]) );
  DLH_X1 \data2i_reg[28]  ( .G(n155), .D(N202), .Q(data2i[28]) );
  DLH_X1 \data2i_reg[27]  ( .G(n155), .D(N201), .Q(data2i[27]) );
  DLH_X1 \data2i_reg[26]  ( .G(n155), .D(N200), .Q(data2i[26]) );
  DLH_X1 \data2i_reg[25]  ( .G(n155), .D(N199), .Q(data2i[25]) );
  DLH_X1 \data2i_reg[24]  ( .G(n155), .D(N198), .Q(data2i[24]) );
  DLH_X1 \data2i_reg[23]  ( .G(n155), .D(N197), .Q(data2i[23]) );
  DLH_X1 \data2i_reg[22]  ( .G(n155), .D(N196), .Q(data2i[22]) );
  DLH_X1 \data2i_reg[21]  ( .G(n155), .D(N195), .Q(data2i[21]) );
  DLH_X1 \data2i_reg[20]  ( .G(n155), .D(N194), .Q(data2i[20]) );
  DLH_X1 \data2i_reg[19]  ( .G(n155), .D(N193), .Q(data2i[19]) );
  DLH_X1 \data2i_reg[18]  ( .G(n155), .D(N192), .Q(data2i[18]) );
  DLH_X1 \data2i_reg[17]  ( .G(n155), .D(N191), .Q(data2i[17]) );
  DLH_X1 \data2i_reg[16]  ( .G(n155), .D(N190), .Q(data2i[16]) );
  DLH_X1 \data2i_reg[15]  ( .G(n155), .D(N189), .Q(data2i[15]) );
  DLH_X1 \data2i_reg[14]  ( .G(n155), .D(N188), .Q(data2i[14]) );
  DLH_X1 \data2i_reg[13]  ( .G(n155), .D(N187), .Q(data2i[13]) );
  DLH_X1 \data2i_reg[12]  ( .G(n155), .D(N186), .Q(data2i[12]) );
  DLH_X1 \data2i_reg[11]  ( .G(n155), .D(N185), .Q(data2i[11]) );
  DLH_X1 \data2i_reg[10]  ( .G(n155), .D(N184), .Q(data2i[10]) );
  DLH_X1 \data2i_reg[9]  ( .G(n155), .D(N183), .Q(data2i[9]) );
  DLH_X1 \data2i_reg[8]  ( .G(n155), .D(N182), .Q(data2i[8]) );
  DLH_X1 \data2i_reg[7]  ( .G(n155), .D(N181), .Q(data2i[7]) );
  DLH_X1 \data2i_reg[6]  ( .G(n155), .D(N180), .Q(data2i[6]) );
  DLH_X1 \data2i_reg[5]  ( .G(n155), .D(N179), .Q(data2i[5]) );
  DLH_X1 \data2i_reg[4]  ( .G(n155), .D(N178), .Q(data2i[4]) );
  DLH_X1 \data2i_reg[3]  ( .G(n155), .D(N177), .Q(data2i[3]) );
  DLH_X1 \data2i_reg[2]  ( .G(n155), .D(N176), .Q(data2i[2]) );
  DLH_X1 \data2i_reg[1]  ( .G(n155), .D(N175), .Q(data2i[1]) );
  DLH_X1 \data2i_reg[0]  ( .G(n155), .D(N174), .Q(data2i[0]) );
  DLH_X1 \data1i_reg[31]  ( .G(n155), .D(DATA1[31]), .Q(data1i[31]) );
  DLH_X1 \data1i_reg[30]  ( .G(n155), .D(DATA1[30]), .Q(data1i[30]) );
  DLH_X1 \data1i_reg[29]  ( .G(n155), .D(DATA1[29]), .Q(data1i[29]) );
  DLH_X1 \data1i_reg[28]  ( .G(n155), .D(DATA1[28]), .Q(data1i[28]) );
  DLH_X1 \data1i_reg[27]  ( .G(n155), .D(DATA1[27]), .Q(data1i[27]) );
  DLH_X1 \data1i_reg[26]  ( .G(n155), .D(DATA1[26]), .Q(data1i[26]) );
  DLH_X1 \data1i_reg[25]  ( .G(n155), .D(DATA1[25]), .Q(data1i[25]) );
  DLH_X1 \data1i_reg[24]  ( .G(n155), .D(DATA1[24]), .Q(data1i[24]) );
  DLH_X1 \data1i_reg[23]  ( .G(n155), .D(DATA1[23]), .Q(data1i[23]) );
  DLH_X1 \data1i_reg[22]  ( .G(n155), .D(DATA1[22]), .Q(data1i[22]) );
  DLH_X1 \data1i_reg[21]  ( .G(n155), .D(DATA1[21]), .Q(data1i[21]) );
  DLH_X1 \data1i_reg[20]  ( .G(n155), .D(DATA1[20]), .Q(data1i[20]) );
  DLH_X1 \data1i_reg[19]  ( .G(n155), .D(DATA1[19]), .Q(data1i[19]) );
  DLH_X1 \data1i_reg[18]  ( .G(n155), .D(DATA1[18]), .Q(data1i[18]) );
  DLH_X1 \data1i_reg[17]  ( .G(n155), .D(DATA1[17]), .Q(data1i[17]) );
  DLH_X1 \data1i_reg[16]  ( .G(n155), .D(DATA1[16]), .Q(data1i[16]) );
  DLH_X1 \data1i_reg[15]  ( .G(n155), .D(DATA1[15]), .Q(data1i[15]) );
  DLH_X1 \data1i_reg[14]  ( .G(n155), .D(DATA1[14]), .Q(data1i[14]) );
  DLH_X1 \data1i_reg[13]  ( .G(n155), .D(DATA1[13]), .Q(data1i[13]) );
  DLH_X1 \data1i_reg[12]  ( .G(n155), .D(DATA1[12]), .Q(data1i[12]) );
  DLH_X1 \data1i_reg[11]  ( .G(n155), .D(DATA1[11]), .Q(data1i[11]) );
  DLH_X1 \data1i_reg[10]  ( .G(n155), .D(DATA1[10]), .Q(data1i[10]) );
  DLH_X1 \data1i_reg[9]  ( .G(n155), .D(DATA1[9]), .Q(data1i[9]) );
  DLH_X1 \data1i_reg[8]  ( .G(n155), .D(DATA1[8]), .Q(data1i[8]) );
  DLH_X1 \data1i_reg[7]  ( .G(n155), .D(DATA1[7]), .Q(data1i[7]) );
  DLH_X1 \data1i_reg[6]  ( .G(n155), .D(DATA1[6]), .Q(data1i[6]) );
  DLH_X1 \data1i_reg[5]  ( .G(n155), .D(DATA1[5]), .Q(data1i[5]) );
  DLH_X1 \data1i_reg[4]  ( .G(n155), .D(DATA1[4]), .Q(data1i[4]) );
  DLH_X1 \data1i_reg[3]  ( .G(n155), .D(DATA1[3]), .Q(data1i[3]) );
  DLH_X1 \data1i_reg[2]  ( .G(n155), .D(DATA1[2]), .Q(data1i[2]) );
  DLH_X1 \data1i_reg[1]  ( .G(n155), .D(DATA1[1]), .Q(data1i[1]) );
  DLH_X1 \data1i_reg[0]  ( .G(n155), .D(DATA1[0]), .Q(data1i[0]) );
  DLH_X1 LOGIC_ARITH_i_reg ( .G(n159), .D(N207), .Q(LOGIC_ARITH_i) );
  DLH_X1 LEFT_RIGHT_i_reg ( .G(n159), .D(N207), .Q(LEFT_RIGHT_i) );
  DLH_X1 \OUTPUT_alu_i_reg[0]  ( .G(N141), .D(N142), .Q(OUTPUT_alu_i[0]) );
  DFF_X1 \OUT_ALU_reg[0]  ( .D(OUTPUT_alu_i[0]), .CK(CLK), .Q(OUT_ALU[0]) );
  DLH_X1 \OUTPUT_alu_i_reg[1]  ( .G(N141), .D(N143), .Q(OUTPUT_alu_i[1]) );
  DFF_X1 \OUT_ALU_reg[1]  ( .D(OUTPUT_alu_i[1]), .CK(CLK), .Q(OUT_ALU[1]) );
  DLH_X1 \OUTPUT_alu_i_reg[2]  ( .G(N141), .D(N144), .Q(OUTPUT_alu_i[2]) );
  DFF_X1 \OUT_ALU_reg[2]  ( .D(OUTPUT_alu_i[2]), .CK(CLK), .Q(OUT_ALU[2]) );
  DLH_X1 \OUTPUT_alu_i_reg[3]  ( .G(N141), .D(N145), .Q(OUTPUT_alu_i[3]) );
  DFF_X1 \OUT_ALU_reg[3]  ( .D(OUTPUT_alu_i[3]), .CK(CLK), .Q(OUT_ALU[3]) );
  DLH_X1 \OUTPUT_alu_i_reg[4]  ( .G(N141), .D(N146), .Q(OUTPUT_alu_i[4]) );
  DFF_X1 \OUT_ALU_reg[4]  ( .D(OUTPUT_alu_i[4]), .CK(CLK), .Q(OUT_ALU[4]) );
  DLH_X1 \OUTPUT_alu_i_reg[5]  ( .G(N141), .D(N147), .Q(OUTPUT_alu_i[5]) );
  DFF_X1 \OUT_ALU_reg[5]  ( .D(OUTPUT_alu_i[5]), .CK(CLK), .Q(OUT_ALU[5]) );
  DLH_X1 \OUTPUT_alu_i_reg[6]  ( .G(N141), .D(N148), .Q(OUTPUT_alu_i[6]) );
  DFF_X1 \OUT_ALU_reg[6]  ( .D(OUTPUT_alu_i[6]), .CK(CLK), .Q(OUT_ALU[6]) );
  DLH_X1 \OUTPUT_alu_i_reg[7]  ( .G(N141), .D(N149), .Q(OUTPUT_alu_i[7]) );
  DFF_X1 \OUT_ALU_reg[7]  ( .D(OUTPUT_alu_i[7]), .CK(CLK), .Q(OUT_ALU[7]) );
  DLH_X1 \OUTPUT_alu_i_reg[8]  ( .G(N141), .D(N150), .Q(OUTPUT_alu_i[8]) );
  DFF_X1 \OUT_ALU_reg[8]  ( .D(OUTPUT_alu_i[8]), .CK(CLK), .Q(OUT_ALU[8]) );
  DLH_X1 \OUTPUT_alu_i_reg[9]  ( .G(N141), .D(N151), .Q(OUTPUT_alu_i[9]) );
  DFF_X1 \OUT_ALU_reg[9]  ( .D(OUTPUT_alu_i[9]), .CK(CLK), .Q(OUT_ALU[9]) );
  DLH_X1 \OUTPUT_alu_i_reg[10]  ( .G(N141), .D(N152), .Q(OUTPUT_alu_i[10]) );
  DFF_X1 \OUT_ALU_reg[10]  ( .D(OUTPUT_alu_i[10]), .CK(CLK), .Q(OUT_ALU[10])
         );
  DLH_X1 \OUTPUT_alu_i_reg[11]  ( .G(N141), .D(N153), .Q(OUTPUT_alu_i[11]) );
  DFF_X1 \OUT_ALU_reg[11]  ( .D(OUTPUT_alu_i[11]), .CK(CLK), .Q(OUT_ALU[11])
         );
  DLH_X1 \OUTPUT_alu_i_reg[12]  ( .G(N141), .D(N154), .Q(OUTPUT_alu_i[12]) );
  DFF_X1 \OUT_ALU_reg[12]  ( .D(OUTPUT_alu_i[12]), .CK(CLK), .Q(OUT_ALU[12])
         );
  DLH_X1 \OUTPUT_alu_i_reg[13]  ( .G(N141), .D(N155), .Q(OUTPUT_alu_i[13]) );
  DFF_X1 \OUT_ALU_reg[13]  ( .D(OUTPUT_alu_i[13]), .CK(CLK), .Q(OUT_ALU[13])
         );
  DLH_X1 \OUTPUT_alu_i_reg[14]  ( .G(N141), .D(N156), .Q(OUTPUT_alu_i[14]) );
  DFF_X1 \OUT_ALU_reg[14]  ( .D(OUTPUT_alu_i[14]), .CK(CLK), .Q(OUT_ALU[14])
         );
  DLH_X1 \OUTPUT_alu_i_reg[15]  ( .G(N141), .D(N157), .Q(OUTPUT_alu_i[15]) );
  DFF_X1 \OUT_ALU_reg[15]  ( .D(OUTPUT_alu_i[15]), .CK(CLK), .Q(OUT_ALU[15])
         );
  DLH_X1 \OUTPUT_alu_i_reg[16]  ( .G(N141), .D(N158), .Q(OUTPUT_alu_i[16]) );
  DFF_X1 \OUT_ALU_reg[16]  ( .D(OUTPUT_alu_i[16]), .CK(CLK), .Q(OUT_ALU[16])
         );
  DLH_X1 \OUTPUT_alu_i_reg[17]  ( .G(N141), .D(N159), .Q(OUTPUT_alu_i[17]) );
  DFF_X1 \OUT_ALU_reg[17]  ( .D(OUTPUT_alu_i[17]), .CK(CLK), .Q(OUT_ALU[17])
         );
  DLH_X1 \OUTPUT_alu_i_reg[18]  ( .G(N141), .D(N160), .Q(OUTPUT_alu_i[18]) );
  DFF_X1 \OUT_ALU_reg[18]  ( .D(OUTPUT_alu_i[18]), .CK(CLK), .Q(OUT_ALU[18])
         );
  DLH_X1 \OUTPUT_alu_i_reg[19]  ( .G(N141), .D(N161), .Q(OUTPUT_alu_i[19]) );
  DFF_X1 \OUT_ALU_reg[19]  ( .D(OUTPUT_alu_i[19]), .CK(CLK), .Q(OUT_ALU[19])
         );
  DLH_X1 \OUTPUT_alu_i_reg[20]  ( .G(N141), .D(N162), .Q(OUTPUT_alu_i[20]) );
  DFF_X1 \OUT_ALU_reg[20]  ( .D(OUTPUT_alu_i[20]), .CK(CLK), .Q(OUT_ALU[20])
         );
  DLH_X1 \OUTPUT_alu_i_reg[21]  ( .G(N141), .D(N163), .Q(OUTPUT_alu_i[21]) );
  DFF_X1 \OUT_ALU_reg[21]  ( .D(OUTPUT_alu_i[21]), .CK(CLK), .Q(OUT_ALU[21])
         );
  DLH_X1 \OUTPUT_alu_i_reg[22]  ( .G(N141), .D(N164), .Q(OUTPUT_alu_i[22]) );
  DFF_X1 \OUT_ALU_reg[22]  ( .D(OUTPUT_alu_i[22]), .CK(CLK), .Q(OUT_ALU[22])
         );
  DLH_X1 \OUTPUT_alu_i_reg[23]  ( .G(N141), .D(N165), .Q(OUTPUT_alu_i[23]) );
  DFF_X1 \OUT_ALU_reg[23]  ( .D(OUTPUT_alu_i[23]), .CK(CLK), .Q(OUT_ALU[23])
         );
  DLH_X1 \OUTPUT_alu_i_reg[24]  ( .G(N141), .D(N166), .Q(OUTPUT_alu_i[24]) );
  DFF_X1 \OUT_ALU_reg[24]  ( .D(OUTPUT_alu_i[24]), .CK(CLK), .Q(OUT_ALU[24])
         );
  DLH_X1 \OUTPUT_alu_i_reg[25]  ( .G(N141), .D(N167), .Q(OUTPUT_alu_i[25]) );
  DFF_X1 \OUT_ALU_reg[25]  ( .D(OUTPUT_alu_i[25]), .CK(CLK), .Q(OUT_ALU[25])
         );
  DLH_X1 \OUTPUT_alu_i_reg[26]  ( .G(N141), .D(N168), .Q(OUTPUT_alu_i[26]) );
  DFF_X1 \OUT_ALU_reg[26]  ( .D(OUTPUT_alu_i[26]), .CK(CLK), .Q(OUT_ALU[26])
         );
  DLH_X1 \OUTPUT_alu_i_reg[27]  ( .G(N141), .D(N169), .Q(OUTPUT_alu_i[27]) );
  DFF_X1 \OUT_ALU_reg[27]  ( .D(OUTPUT_alu_i[27]), .CK(CLK), .Q(OUT_ALU[27])
         );
  DLH_X1 \OUTPUT_alu_i_reg[28]  ( .G(N141), .D(N170), .Q(OUTPUT_alu_i[28]) );
  DFF_X1 \OUT_ALU_reg[28]  ( .D(OUTPUT_alu_i[28]), .CK(CLK), .Q(OUT_ALU[28])
         );
  DLH_X1 \OUTPUT_alu_i_reg[29]  ( .G(N141), .D(N171), .Q(OUTPUT_alu_i[29]) );
  DFF_X1 \OUT_ALU_reg[29]  ( .D(OUTPUT_alu_i[29]), .CK(CLK), .Q(OUT_ALU[29])
         );
  DLH_X1 \OUTPUT_alu_i_reg[30]  ( .G(N141), .D(N172), .Q(OUTPUT_alu_i[30]) );
  DFF_X1 \OUT_ALU_reg[30]  ( .D(OUTPUT_alu_i[30]), .CK(CLK), .Q(OUT_ALU[30])
         );
  DLH_X1 \OUTPUT_alu_i_reg[31]  ( .G(N141), .D(N173), .Q(OUTPUT_alu_i[31]) );
  DFF_X1 \OUT_ALU_reg[31]  ( .D(OUTPUT_alu_i[31]), .CK(CLK), .Q(OUT_ALU[31])
         );
  INV_X1 U4 ( .A(n1), .ZN(N207) );
  OAI22_X1 U5 ( .A1(DATA2[31]), .A2(n157), .B1(n3), .B2(n4), .ZN(N205) );
  INV_X1 U6 ( .A(DATA2[31]), .ZN(n4) );
  OAI22_X1 U7 ( .A1(DATA2[30]), .A2(n157), .B1(n3), .B2(n5), .ZN(N204) );
  INV_X1 U8 ( .A(DATA2[30]), .ZN(n5) );
  OAI22_X1 U9 ( .A1(DATA2[29]), .A2(n157), .B1(n3), .B2(n6), .ZN(N203) );
  INV_X1 U10 ( .A(DATA2[29]), .ZN(n6) );
  OAI22_X1 U11 ( .A1(DATA2[28]), .A2(n157), .B1(n3), .B2(n7), .ZN(N202) );
  INV_X1 U12 ( .A(DATA2[28]), .ZN(n7) );
  OAI22_X1 U13 ( .A1(DATA2[27]), .A2(n157), .B1(n3), .B2(n8), .ZN(N201) );
  INV_X1 U14 ( .A(DATA2[27]), .ZN(n8) );
  OAI22_X1 U15 ( .A1(DATA2[26]), .A2(n157), .B1(n3), .B2(n9), .ZN(N200) );
  INV_X1 U16 ( .A(DATA2[26]), .ZN(n9) );
  OAI22_X1 U17 ( .A1(DATA2[25]), .A2(n157), .B1(n3), .B2(n10), .ZN(N199) );
  INV_X1 U18 ( .A(DATA2[25]), .ZN(n10) );
  OAI22_X1 U19 ( .A1(DATA2[24]), .A2(n157), .B1(n3), .B2(n11), .ZN(N198) );
  INV_X1 U20 ( .A(DATA2[24]), .ZN(n11) );
  OAI22_X1 U21 ( .A1(DATA2[23]), .A2(n157), .B1(n3), .B2(n12), .ZN(N197) );
  INV_X1 U22 ( .A(DATA2[23]), .ZN(n12) );
  OAI22_X1 U23 ( .A1(DATA2[22]), .A2(n157), .B1(n3), .B2(n13), .ZN(N196) );
  INV_X1 U24 ( .A(DATA2[22]), .ZN(n13) );
  OAI22_X1 U25 ( .A1(DATA2[21]), .A2(n157), .B1(n3), .B2(n14), .ZN(N195) );
  INV_X1 U26 ( .A(DATA2[21]), .ZN(n14) );
  OAI22_X1 U27 ( .A1(DATA2[20]), .A2(n157), .B1(n3), .B2(n15), .ZN(N194) );
  INV_X1 U28 ( .A(DATA2[20]), .ZN(n15) );
  OAI22_X1 U29 ( .A1(DATA2[19]), .A2(n157), .B1(n3), .B2(n16), .ZN(N193) );
  INV_X1 U30 ( .A(DATA2[19]), .ZN(n16) );
  OAI22_X1 U31 ( .A1(DATA2[18]), .A2(n157), .B1(n3), .B2(n17), .ZN(N192) );
  INV_X1 U32 ( .A(DATA2[18]), .ZN(n17) );
  OAI22_X1 U33 ( .A1(DATA2[17]), .A2(n157), .B1(n3), .B2(n18), .ZN(N191) );
  INV_X1 U34 ( .A(DATA2[17]), .ZN(n18) );
  OAI22_X1 U35 ( .A1(DATA2[16]), .A2(n157), .B1(n3), .B2(n19), .ZN(N190) );
  INV_X1 U36 ( .A(DATA2[16]), .ZN(n19) );
  OAI22_X1 U37 ( .A1(DATA2[15]), .A2(n157), .B1(n3), .B2(n20), .ZN(N189) );
  INV_X1 U38 ( .A(DATA2[15]), .ZN(n20) );
  OAI22_X1 U39 ( .A1(DATA2[14]), .A2(n157), .B1(n3), .B2(n21), .ZN(N188) );
  INV_X1 U40 ( .A(DATA2[14]), .ZN(n21) );
  OAI22_X1 U41 ( .A1(DATA2[13]), .A2(n157), .B1(n3), .B2(n22), .ZN(N187) );
  INV_X1 U42 ( .A(DATA2[13]), .ZN(n22) );
  OAI22_X1 U43 ( .A1(DATA2[12]), .A2(n157), .B1(n3), .B2(n23), .ZN(N186) );
  INV_X1 U44 ( .A(DATA2[12]), .ZN(n23) );
  OAI22_X1 U45 ( .A1(DATA2[11]), .A2(n157), .B1(n3), .B2(n24), .ZN(N185) );
  INV_X1 U46 ( .A(DATA2[11]), .ZN(n24) );
  OAI22_X1 U47 ( .A1(DATA2[10]), .A2(n157), .B1(n3), .B2(n25), .ZN(N184) );
  INV_X1 U48 ( .A(DATA2[10]), .ZN(n25) );
  OAI22_X1 U49 ( .A1(DATA2[9]), .A2(n157), .B1(n3), .B2(n26), .ZN(N183) );
  INV_X1 U50 ( .A(DATA2[9]), .ZN(n26) );
  OAI22_X1 U51 ( .A1(DATA2[8]), .A2(n157), .B1(n3), .B2(n27), .ZN(N182) );
  INV_X1 U52 ( .A(DATA2[8]), .ZN(n27) );
  OAI22_X1 U53 ( .A1(DATA2[7]), .A2(n157), .B1(n3), .B2(n28), .ZN(N181) );
  INV_X1 U54 ( .A(DATA2[7]), .ZN(n28) );
  OAI22_X1 U55 ( .A1(DATA2[6]), .A2(n157), .B1(n3), .B2(n29), .ZN(N180) );
  INV_X1 U56 ( .A(DATA2[6]), .ZN(n29) );
  OAI22_X1 U57 ( .A1(DATA2[5]), .A2(n157), .B1(n3), .B2(n30), .ZN(N179) );
  INV_X1 U58 ( .A(DATA2[5]), .ZN(n30) );
  OAI22_X1 U59 ( .A1(DATA2[4]), .A2(n157), .B1(n3), .B2(n31), .ZN(N178) );
  INV_X1 U60 ( .A(DATA2[4]), .ZN(n31) );
  OAI22_X1 U61 ( .A1(DATA2[3]), .A2(n157), .B1(n3), .B2(n32), .ZN(N177) );
  INV_X1 U62 ( .A(DATA2[3]), .ZN(n32) );
  OAI22_X1 U63 ( .A1(DATA2[2]), .A2(n157), .B1(n3), .B2(n33), .ZN(N176) );
  INV_X1 U64 ( .A(DATA2[2]), .ZN(n33) );
  OAI22_X1 U65 ( .A1(DATA2[1]), .A2(n157), .B1(n3), .B2(n34), .ZN(N175) );
  INV_X1 U66 ( .A(DATA2[1]), .ZN(n34) );
  OAI22_X1 U67 ( .A1(DATA2[0]), .A2(n157), .B1(n3), .B2(n35), .ZN(N174) );
  INV_X1 U68 ( .A(DATA2[0]), .ZN(n35) );
  NAND2_X1 U70 ( .A1(n37), .A2(n38), .ZN(N173) );
  AOI22_X1 U71 ( .A1(OUTPUT2[31]), .A2(n39), .B1(OUTPUT4[31]), .B2(n153), .ZN(
        n38) );
  NAND2_X1 U73 ( .A1(n42), .A2(n43), .ZN(N172) );
  AOI22_X1 U74 ( .A1(OUTPUT2[30]), .A2(n39), .B1(OUTPUT4[30]), .B2(n153), .ZN(
        n43) );
  NAND2_X1 U76 ( .A1(n44), .A2(n45), .ZN(N171) );
  AOI22_X1 U77 ( .A1(OUTPUT2[29]), .A2(n39), .B1(OUTPUT4[29]), .B2(n153), .ZN(
        n45) );
  NAND2_X1 U79 ( .A1(n46), .A2(n47), .ZN(N170) );
  AOI22_X1 U80 ( .A1(OUTPUT2[28]), .A2(n39), .B1(OUTPUT4[28]), .B2(n153), .ZN(
        n47) );
  NAND2_X1 U82 ( .A1(n48), .A2(n49), .ZN(N169) );
  AOI22_X1 U83 ( .A1(OUTPUT2[27]), .A2(n39), .B1(OUTPUT4[27]), .B2(n153), .ZN(
        n49) );
  NAND2_X1 U85 ( .A1(n50), .A2(n51), .ZN(N168) );
  AOI22_X1 U86 ( .A1(OUTPUT2[26]), .A2(n39), .B1(OUTPUT4[26]), .B2(n153), .ZN(
        n51) );
  NAND2_X1 U88 ( .A1(n52), .A2(n53), .ZN(N167) );
  AOI22_X1 U89 ( .A1(OUTPUT2[25]), .A2(n39), .B1(OUTPUT4[25]), .B2(n153), .ZN(
        n53) );
  NAND2_X1 U91 ( .A1(n54), .A2(n55), .ZN(N166) );
  AOI22_X1 U92 ( .A1(OUTPUT2[24]), .A2(n39), .B1(OUTPUT4[24]), .B2(n153), .ZN(
        n55) );
  NAND2_X1 U94 ( .A1(n56), .A2(n57), .ZN(N165) );
  AOI22_X1 U95 ( .A1(OUTPUT2[23]), .A2(n39), .B1(OUTPUT4[23]), .B2(n153), .ZN(
        n57) );
  NAND2_X1 U97 ( .A1(n58), .A2(n59), .ZN(N164) );
  AOI22_X1 U98 ( .A1(OUTPUT2[22]), .A2(n39), .B1(OUTPUT4[22]), .B2(n153), .ZN(
        n59) );
  NAND2_X1 U100 ( .A1(n60), .A2(n61), .ZN(N163) );
  AOI22_X1 U101 ( .A1(OUTPUT2[21]), .A2(n39), .B1(OUTPUT4[21]), .B2(n153), 
        .ZN(n61) );
  NAND2_X1 U103 ( .A1(n62), .A2(n63), .ZN(N162) );
  AOI22_X1 U104 ( .A1(OUTPUT2[20]), .A2(n39), .B1(OUTPUT4[20]), .B2(n153), 
        .ZN(n63) );
  NAND2_X1 U106 ( .A1(n64), .A2(n65), .ZN(N161) );
  AOI22_X1 U107 ( .A1(OUTPUT2[19]), .A2(n39), .B1(OUTPUT4[19]), .B2(n153), 
        .ZN(n65) );
  NAND2_X1 U109 ( .A1(n66), .A2(n67), .ZN(N160) );
  AOI22_X1 U110 ( .A1(OUTPUT2[18]), .A2(n39), .B1(OUTPUT4[18]), .B2(n153), 
        .ZN(n67) );
  NAND2_X1 U112 ( .A1(n68), .A2(n69), .ZN(N159) );
  AOI22_X1 U113 ( .A1(OUTPUT2[17]), .A2(n39), .B1(OUTPUT4[17]), .B2(n153), 
        .ZN(n69) );
  NAND2_X1 U115 ( .A1(n70), .A2(n71), .ZN(N158) );
  AOI22_X1 U116 ( .A1(OUTPUT2[16]), .A2(n39), .B1(OUTPUT4[16]), .B2(n153), 
        .ZN(n71) );
  NAND2_X1 U118 ( .A1(n72), .A2(n73), .ZN(N157) );
  AOI22_X1 U119 ( .A1(OUTPUT2[15]), .A2(n39), .B1(OUTPUT4[15]), .B2(n153), 
        .ZN(n73) );
  NAND2_X1 U121 ( .A1(n74), .A2(n75), .ZN(N156) );
  AOI22_X1 U122 ( .A1(OUTPUT2[14]), .A2(n39), .B1(OUTPUT4[14]), .B2(n153), 
        .ZN(n75) );
  NAND2_X1 U124 ( .A1(n76), .A2(n77), .ZN(N155) );
  AOI22_X1 U125 ( .A1(OUTPUT2[13]), .A2(n39), .B1(OUTPUT4[13]), .B2(n153), 
        .ZN(n77) );
  NAND2_X1 U127 ( .A1(n78), .A2(n79), .ZN(N154) );
  AOI22_X1 U128 ( .A1(OUTPUT2[12]), .A2(n39), .B1(OUTPUT4[12]), .B2(n153), 
        .ZN(n79) );
  NAND2_X1 U130 ( .A1(n80), .A2(n81), .ZN(N153) );
  AOI22_X1 U131 ( .A1(OUTPUT2[11]), .A2(n39), .B1(OUTPUT4[11]), .B2(n153), 
        .ZN(n81) );
  NAND2_X1 U133 ( .A1(n82), .A2(n83), .ZN(N152) );
  AOI22_X1 U134 ( .A1(OUTPUT2[10]), .A2(n39), .B1(OUTPUT4[10]), .B2(n153), 
        .ZN(n83) );
  NAND2_X1 U136 ( .A1(n84), .A2(n85), .ZN(N151) );
  AOI22_X1 U137 ( .A1(OUTPUT2[9]), .A2(n39), .B1(OUTPUT4[9]), .B2(n153), .ZN(
        n85) );
  NAND2_X1 U139 ( .A1(n86), .A2(n87), .ZN(N150) );
  AOI22_X1 U140 ( .A1(OUTPUT2[8]), .A2(n39), .B1(OUTPUT4[8]), .B2(n153), .ZN(
        n87) );
  NAND2_X1 U142 ( .A1(n88), .A2(n89), .ZN(N149) );
  AOI22_X1 U143 ( .A1(OUTPUT2[7]), .A2(n39), .B1(OUTPUT4[7]), .B2(n153), .ZN(
        n89) );
  NAND2_X1 U145 ( .A1(n90), .A2(n91), .ZN(N148) );
  AOI22_X1 U146 ( .A1(OUTPUT2[6]), .A2(n39), .B1(OUTPUT4[6]), .B2(n153), .ZN(
        n91) );
  NAND2_X1 U148 ( .A1(n92), .A2(n93), .ZN(N147) );
  AOI22_X1 U149 ( .A1(OUTPUT2[5]), .A2(n39), .B1(OUTPUT4[5]), .B2(n153), .ZN(
        n93) );
  NAND2_X1 U151 ( .A1(n94), .A2(n95), .ZN(N146) );
  AOI22_X1 U152 ( .A1(OUTPUT2[4]), .A2(n39), .B1(OUTPUT4[4]), .B2(n153), .ZN(
        n95) );
  NAND2_X1 U154 ( .A1(n96), .A2(n97), .ZN(N145) );
  AOI22_X1 U155 ( .A1(OUTPUT2[3]), .A2(n39), .B1(OUTPUT4[3]), .B2(n153), .ZN(
        n97) );
  NAND2_X1 U157 ( .A1(n98), .A2(n99), .ZN(N144) );
  AOI22_X1 U158 ( .A1(OUTPUT2[2]), .A2(n39), .B1(OUTPUT4[2]), .B2(n153), .ZN(
        n99) );
  NAND2_X1 U160 ( .A1(n100), .A2(n101), .ZN(N143) );
  AOI22_X1 U161 ( .A1(OUTPUT2[1]), .A2(n39), .B1(OUTPUT4[1]), .B2(n153), .ZN(
        n101) );
  NAND2_X1 U163 ( .A1(n102), .A2(n103), .ZN(N142) );
  AOI22_X1 U164 ( .A1(OUTPUT2[0]), .A2(n39), .B1(OUTPUT4[0]), .B2(n153), .ZN(
        n103) );
  AOI22_X1 U165 ( .A1(\OUTPUT3[0] ), .A2(n41), .B1(OUTPUT1[0]), .B2(n159), 
        .ZN(n102) );
  OR3_X1 U166 ( .A1(n155), .A2(n159), .A3(n153), .ZN(N141) );
  OAI221_X1 U167 ( .B1(n104), .B2(n105), .C1(n106), .C2(n107), .A(n108), .ZN(
        n40) );
  INV_X1 U168 ( .A(n109), .ZN(n108) );
  OAI22_X1 U169 ( .A1(n110), .A2(n111), .B1(n112), .B2(n113), .ZN(n109) );
  INV_X1 U170 ( .A(n114), .ZN(n111) );
  OAI211_X1 U171 ( .C1(n115), .C2(n116), .A(n117), .B(n1), .ZN(N206) );
  NAND2_X1 U172 ( .A1(n118), .A2(n119), .ZN(n1) );
  OAI21_X1 U173 ( .B1(n120), .B2(n119), .A(n121), .ZN(n117) );
  NAND2_X1 U174 ( .A1(n122), .A2(n112), .ZN(n119) );
  NAND2_X1 U175 ( .A1(n123), .A2(n124), .ZN(n112) );
  NOR3_X1 U176 ( .A1(n125), .A2(FUNC[3]), .A3(n126), .ZN(n120) );
  INV_X1 U177 ( .A(n157), .ZN(N140) );
  NOR3_X1 U178 ( .A1(n127), .A2(n128), .A3(n41), .ZN(n2) );
  OR2_X1 U179 ( .A1(n39), .A2(n41), .ZN(N139) );
  OAI221_X1 U180 ( .B1(n116), .B2(n105), .C1(n106), .C2(n129), .A(n130), .ZN(
        n41) );
  AOI221_X1 U181 ( .B1(n131), .B2(n114), .C1(n132), .C2(n133), .A(n134), .ZN(
        n130) );
  NOR3_X1 U182 ( .A1(n135), .A2(n113), .A3(n136), .ZN(n134) );
  NAND2_X1 U183 ( .A1(n137), .A2(n138), .ZN(n132) );
  NAND2_X1 U184 ( .A1(n106), .A2(n139), .ZN(n114) );
  OAI211_X1 U185 ( .C1(n136), .C2(n126), .A(n105), .B(n115), .ZN(n131) );
  INV_X1 U186 ( .A(n140), .ZN(n126) );
  NAND2_X1 U187 ( .A1(n141), .A2(n142), .ZN(n105) );
  OAI221_X1 U189 ( .B1(n113), .B2(n107), .C1(n116), .C2(n122), .A(n143), .ZN(
        n36) );
  AOI222_X1 U190 ( .A1(n144), .A2(n133), .B1(n121), .B2(n145), .C1(n146), .C2(
        n147), .ZN(n143) );
  NAND4_X1 U191 ( .A1(n110), .A2(n148), .A3(n115), .A4(n122), .ZN(n147) );
  NAND2_X1 U192 ( .A1(n149), .A2(n124), .ZN(n115) );
  NAND3_X1 U193 ( .A1(n138), .A2(n137), .A3(n148), .ZN(n145) );
  NAND3_X1 U194 ( .A1(n124), .A2(n150), .A3(FUNC[2]), .ZN(n137) );
  NAND2_X1 U195 ( .A1(n141), .A2(n140), .ZN(n138) );
  INV_X1 U196 ( .A(n106), .ZN(n121) );
  NAND2_X1 U197 ( .A1(FUNC[0]), .A2(FUNC[1]), .ZN(n106) );
  NAND2_X1 U198 ( .A1(n113), .A2(n139), .ZN(n133) );
  INV_X1 U199 ( .A(n129), .ZN(n144) );
  NAND2_X1 U200 ( .A1(n149), .A2(n140), .ZN(n129) );
  NOR2_X1 U201 ( .A1(n135), .A2(FUNC[4]), .ZN(n140) );
  NAND2_X1 U202 ( .A1(n142), .A2(n123), .ZN(n122) );
  INV_X1 U203 ( .A(n136), .ZN(n123) );
  NAND2_X1 U204 ( .A1(n150), .A2(n125), .ZN(n136) );
  AND2_X1 U205 ( .A1(n116), .A2(n104), .ZN(n113) );
  INV_X1 U206 ( .A(n146), .ZN(n104) );
  NOR2_X1 U207 ( .A1(FUNC[1]), .A2(FUNC[0]), .ZN(n146) );
  AOI21_X1 U208 ( .B1(n110), .B2(n148), .A(n116), .ZN(n128) );
  NAND2_X1 U209 ( .A1(FUNC[0]), .A2(n151), .ZN(n116) );
  NAND3_X1 U210 ( .A1(n142), .A2(n150), .A3(FUNC[2]), .ZN(n110) );
  AOI21_X1 U211 ( .B1(n148), .B2(n107), .A(n139), .ZN(n127) );
  INV_X1 U212 ( .A(n118), .ZN(n139) );
  NOR2_X1 U213 ( .A1(n151), .A2(FUNC[0]), .ZN(n118) );
  INV_X1 U214 ( .A(FUNC[1]), .ZN(n151) );
  NAND2_X1 U215 ( .A1(n149), .A2(n142), .ZN(n107) );
  NOR2_X1 U216 ( .A1(FUNC[5]), .A2(FUNC[4]), .ZN(n142) );
  NOR2_X1 U217 ( .A1(n150), .A2(n125), .ZN(n149) );
  INV_X1 U218 ( .A(FUNC[2]), .ZN(n125) );
  NAND2_X1 U219 ( .A1(n141), .A2(n124), .ZN(n148) );
  AND2_X1 U220 ( .A1(FUNC[4]), .A2(n135), .ZN(n124) );
  INV_X1 U221 ( .A(FUNC[5]), .ZN(n135) );
  NOR2_X1 U222 ( .A1(n150), .A2(FUNC[2]), .ZN(n141) );
  INV_X1 U223 ( .A(FUNC[3]), .ZN(n150) );
  logic_N32 log ( .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , 
        \FUNC[0] }), .DATA1(DATA1), .DATA2(DATA2), .OUT_ALU(OUTPUT4) );
  comparator comp ( .DATA1(OUTPUT2), .DATA2i(Cout_i), .tipo({\FUNC[5] , 
        \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }), .OUTALU({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, \OUTPUT3[0] }) );
  SHIFTER_GENERIC_N32 shifter ( .A(DATA1), .B(DATA2[4:0]), .LOGIC_ARITH(
        LOGIC_ARITH_i), .LEFT_RIGHT(LEFT_RIGHT_i), .SHIFT_ROTATE(1'b1), 
        .OUTPUT(OUTPUT1) );
  P4_ADDER_NBIT32 adder ( .A(data1i), .B(data2i), .Cin(Cin_i), .S(OUTPUT2), 
        .Cout(Cout_i) );
  INV_X2 U69 ( .A(n36), .ZN(n3) );
  OR3_X2 U72 ( .A1(n127), .A2(n128), .A3(n36), .ZN(n39) );
  INV_X1 U75 ( .A(n40), .ZN(n152) );
  INV_X2 U78 ( .A(n152), .ZN(n153) );
  INV_X1 U81 ( .A(N139), .ZN(n154) );
  INV_X2 U84 ( .A(n154), .ZN(n155) );
  INV_X1 U87 ( .A(n2), .ZN(n156) );
  INV_X2 U90 ( .A(n156), .ZN(n157) );
  INV_X1 U93 ( .A(N206), .ZN(n158) );
  INV_X4 U96 ( .A(n158), .ZN(n159) );
  NAND2_X2 U99 ( .A1(OUTPUT1[31]), .A2(n159), .ZN(n37) );
  NAND2_X2 U102 ( .A1(OUTPUT1[30]), .A2(n159), .ZN(n42) );
  NAND2_X2 U105 ( .A1(OUTPUT1[29]), .A2(n159), .ZN(n44) );
  NAND2_X2 U108 ( .A1(OUTPUT1[28]), .A2(n159), .ZN(n46) );
  NAND2_X2 U111 ( .A1(OUTPUT1[27]), .A2(n159), .ZN(n48) );
  NAND2_X2 U114 ( .A1(OUTPUT1[26]), .A2(n159), .ZN(n50) );
  NAND2_X2 U117 ( .A1(OUTPUT1[25]), .A2(n159), .ZN(n52) );
  NAND2_X2 U120 ( .A1(OUTPUT1[24]), .A2(n159), .ZN(n54) );
  NAND2_X2 U123 ( .A1(OUTPUT1[23]), .A2(n159), .ZN(n56) );
  NAND2_X2 U126 ( .A1(OUTPUT1[22]), .A2(n159), .ZN(n58) );
  NAND2_X2 U129 ( .A1(OUTPUT1[21]), .A2(n159), .ZN(n60) );
  NAND2_X2 U132 ( .A1(OUTPUT1[20]), .A2(n159), .ZN(n62) );
  NAND2_X2 U135 ( .A1(OUTPUT1[19]), .A2(n159), .ZN(n64) );
  NAND2_X2 U138 ( .A1(OUTPUT1[18]), .A2(n159), .ZN(n66) );
  NAND2_X2 U141 ( .A1(OUTPUT1[17]), .A2(n159), .ZN(n68) );
  NAND2_X2 U144 ( .A1(OUTPUT1[16]), .A2(n159), .ZN(n70) );
  NAND2_X2 U147 ( .A1(OUTPUT1[15]), .A2(n159), .ZN(n72) );
  NAND2_X2 U150 ( .A1(OUTPUT1[14]), .A2(n159), .ZN(n74) );
  NAND2_X2 U153 ( .A1(OUTPUT1[13]), .A2(n159), .ZN(n76) );
  NAND2_X2 U156 ( .A1(OUTPUT1[12]), .A2(n159), .ZN(n78) );
  NAND2_X2 U159 ( .A1(OUTPUT1[11]), .A2(n159), .ZN(n80) );
  NAND2_X2 U162 ( .A1(OUTPUT1[10]), .A2(n159), .ZN(n82) );
  NAND2_X2 U188 ( .A1(OUTPUT1[9]), .A2(n159), .ZN(n84) );
  NAND2_X2 U224 ( .A1(OUTPUT1[8]), .A2(n159), .ZN(n86) );
  NAND2_X2 U225 ( .A1(OUTPUT1[7]), .A2(n159), .ZN(n88) );
  NAND2_X2 U226 ( .A1(OUTPUT1[6]), .A2(n159), .ZN(n90) );
  NAND2_X2 U227 ( .A1(OUTPUT1[5]), .A2(n159), .ZN(n92) );
  NAND2_X2 U228 ( .A1(OUTPUT1[4]), .A2(n159), .ZN(n94) );
  NAND2_X2 U229 ( .A1(OUTPUT1[3]), .A2(n159), .ZN(n96) );
  NAND2_X2 U230 ( .A1(OUTPUT1[2]), .A2(n159), .ZN(n98) );
  NAND2_X2 U231 ( .A1(OUTPUT1[1]), .A2(n159), .ZN(n100) );
endmodule


module zero_eval_NBIT32 ( \input , res );
  input [31:0] \input ;
  output res;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(res) );
  NAND4_X1 U2 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NOR4_X1 U3 ( .A1(\input [23]), .A2(\input [22]), .A3(\input [21]), .A4(
        \input [20]), .ZN(n6) );
  NOR4_X1 U4 ( .A1(\input [1]), .A2(\input [19]), .A3(\input [18]), .A4(
        \input [17]), .ZN(n5) );
  NOR4_X1 U5 ( .A1(\input [16]), .A2(\input [15]), .A3(\input [14]), .A4(
        \input [13]), .ZN(n4) );
  NOR4_X1 U6 ( .A1(\input [12]), .A2(\input [11]), .A3(\input [10]), .A4(
        \input [0]), .ZN(n3) );
  NAND4_X1 U7 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NOR4_X1 U8 ( .A1(\input [9]), .A2(\input [8]), .A3(\input [7]), .A4(
        \input [6]), .ZN(n10) );
  NOR4_X1 U9 ( .A1(\input [5]), .A2(\input [4]), .A3(\input [3]), .A4(
        \input [31]), .ZN(n9) );
  NOR4_X1 U10 ( .A1(\input [30]), .A2(\input [2]), .A3(\input [29]), .A4(
        \input [28]), .ZN(n8) );
  NOR4_X1 U11 ( .A1(\input [27]), .A2(\input [26]), .A3(\input [25]), .A4(
        \input [24]), .ZN(n7) );
endmodule


module COND_BT_NBIT32 ( ZERO_BIT, OPCODE_0, branch_op, con_sign );
  input ZERO_BIT, OPCODE_0, branch_op;
  output con_sign;
  wire   n1;

  AND2_X1 U2 ( .A1(branch_op), .A2(n1), .ZN(con_sign) );
  XOR2_X1 U3 ( .A(ZERO_BIT), .B(OPCODE_0), .Z(n1) );
endmodule


module IV_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_480 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_479 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_478 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_160 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_160 UIV ( .A(S), .Y(SB) );
  ND2_480 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_479 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_478 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_477 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_476 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_475 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_159 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_159 UIV ( .A(S), .Y(SB) );
  ND2_477 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_476 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_475 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_474 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_473 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_472 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_158 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_158 UIV ( .A(S), .Y(SB) );
  ND2_474 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_473 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_472 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_471 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_470 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_469 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_157 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_157 UIV ( .A(S), .Y(SB) );
  ND2_471 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_470 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_469 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_468 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_467 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_466 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_156 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_156 UIV ( .A(S), .Y(SB) );
  ND2_468 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_467 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_466 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_465 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_464 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_463 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_155 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_155 UIV ( .A(S), .Y(SB) );
  ND2_465 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_464 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_463 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_462 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_461 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_460 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_154 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_154 UIV ( .A(S), .Y(SB) );
  ND2_462 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_461 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_460 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_459 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_458 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_457 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_153 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_153 UIV ( .A(S), .Y(SB) );
  ND2_459 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_458 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_457 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_456 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_455 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_454 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_152 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_152 UIV ( .A(S), .Y(SB) );
  ND2_456 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_455 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_454 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_453 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_452 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_451 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_151 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_151 UIV ( .A(S), .Y(SB) );
  ND2_453 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_452 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_451 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_450 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_449 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_448 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_150 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_150 UIV ( .A(S), .Y(SB) );
  ND2_450 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_449 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_448 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_447 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_446 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_445 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_149 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_149 UIV ( .A(S), .Y(SB) );
  ND2_447 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_446 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_445 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_444 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_443 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_442 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_148 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_148 UIV ( .A(S), .Y(SB) );
  ND2_444 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_443 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_442 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_441 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_440 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_439 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_147 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_147 UIV ( .A(S), .Y(SB) );
  ND2_441 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_440 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_439 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_438 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_437 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_436 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_146 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_146 UIV ( .A(S), .Y(SB) );
  ND2_438 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_437 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_436 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_435 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_434 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_433 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_145 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_145 UIV ( .A(S), .Y(SB) );
  ND2_435 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_434 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_433 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_432 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_431 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_430 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_144 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_144 UIV ( .A(S), .Y(SB) );
  ND2_432 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_431 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_430 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_429 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_428 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_427 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_143 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_143 UIV ( .A(S), .Y(SB) );
  ND2_429 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_428 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_427 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_426 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_425 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_424 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_142 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_142 UIV ( .A(S), .Y(SB) );
  ND2_426 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_425 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_424 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_423 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_422 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_421 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_141 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_141 UIV ( .A(S), .Y(SB) );
  ND2_423 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_422 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_421 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_420 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_419 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_418 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_140 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_140 UIV ( .A(S), .Y(SB) );
  ND2_420 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_419 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_418 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_417 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_416 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_415 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_139 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_139 UIV ( .A(S), .Y(SB) );
  ND2_417 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_416 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_415 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_414 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_413 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_412 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_138 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_138 UIV ( .A(S), .Y(SB) );
  ND2_414 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_413 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_412 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_411 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_410 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_409 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_137 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_137 UIV ( .A(S), .Y(SB) );
  ND2_411 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_410 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_409 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_408 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_407 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_406 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_136 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_136 UIV ( .A(S), .Y(SB) );
  ND2_408 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_407 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_406 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_405 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_404 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_403 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_135 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_135 UIV ( .A(S), .Y(SB) );
  ND2_405 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_404 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_403 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_402 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_401 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_400 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_134 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_134 UIV ( .A(S), .Y(SB) );
  ND2_402 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_401 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_400 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_399 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_398 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_397 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_133 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_133 UIV ( .A(S), .Y(SB) );
  ND2_399 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_398 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_397 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_396 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_395 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_394 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_132 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_132 UIV ( .A(S), .Y(SB) );
  ND2_396 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_395 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_394 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_393 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_392 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_391 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_131 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_131 UIV ( .A(S), .Y(SB) );
  ND2_393 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_392 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_391 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_390 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_389 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_388 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_130 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_130 UIV ( .A(S), .Y(SB) );
  ND2_390 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_389 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_388 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_387 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_386 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_385 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_129 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_129 UIV ( .A(S), .Y(SB) );
  ND2_387 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_386 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_385 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_160 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_159 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_158 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_157 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_156 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_155 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_154 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_153 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_152 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_151 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_150 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_149 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_148 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_147 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_146 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_145 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_144 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_143 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_142 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_141 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_140 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_139 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_138 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_137 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_136 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_135 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_134 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_133 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_132 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_131 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_130 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_129 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module FF_6 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n5, n6, n7, n8;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n8), .A2(n7), .ZN(n5) );
  INV_X1 U4 ( .A(RESET), .ZN(n7) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n6), .ZN(n8) );
  INV_X1 U6 ( .A(EN), .ZN(n6) );
endmodule


module regFFD_NBIT32_5 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module FF_5 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n5, n6, n7, n8;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n8), .A2(n7), .ZN(n5) );
  INV_X1 U4 ( .A(RESET), .ZN(n7) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n6), .ZN(n8) );
  INV_X1 U6 ( .A(EN), .ZN(n6) );
endmodule


module regFFD_NBIT32_4 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT5_2 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \Q_reg[4]  ( .D(n16), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n21) );
  DFFR_X1 \Q_reg[3]  ( .D(n17), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n22) );
  DFFR_X1 \Q_reg[2]  ( .D(n18), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n23) );
  DFFR_X1 \Q_reg[1]  ( .D(n19), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n24) );
  DFFR_X1 \Q_reg[0]  ( .D(n20), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n25) );
  OAI21_X1 U2 ( .B1(n25), .B2(ENABLE), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(ENABLE), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(ENABLE), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(ENABLE), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(ENABLE), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n26) );
endmodule


module FF_4 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n4, n5;

  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n4), .ZN(n5) );
  INV_X1 U6 ( .A(EN), .ZN(n4) );
  SDFF_X1 Q_reg ( .D(RESET), .SI(1'b0), .SE(n5), .CK(CLK), .Q(Q) );
endmodule


module regFFD_NBIT6_1 ( CK, RESET, ENABLE, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET, ENABLE;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36;

  DFFR_X1 \Q_reg[5]  ( .D(n19), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n25) );
  DFFR_X1 \Q_reg[4]  ( .D(n20), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n26) );
  DFFR_X1 \Q_reg[3]  ( .D(n21), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n27) );
  DFFR_X1 \Q_reg[2]  ( .D(n22), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n28) );
  DFFR_X1 \Q_reg[1]  ( .D(n23), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n29) );
  DFFR_X1 \Q_reg[0]  ( .D(n24), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n30) );
  OAI21_X1 U2 ( .B1(n30), .B2(ENABLE), .A(n36), .ZN(n24) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n36) );
  OAI21_X1 U4 ( .B1(n29), .B2(ENABLE), .A(n35), .ZN(n23) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n35) );
  OAI21_X1 U6 ( .B1(n28), .B2(ENABLE), .A(n34), .ZN(n22) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n34) );
  OAI21_X1 U8 ( .B1(n27), .B2(ENABLE), .A(n33), .ZN(n21) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n33) );
  OAI21_X1 U10 ( .B1(n26), .B2(ENABLE), .A(n32), .ZN(n20) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n32) );
  OAI21_X1 U12 ( .B1(n25), .B2(ENABLE), .A(n31), .ZN(n19) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n31) );
endmodule


module IV_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_384 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_383 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_382 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_128 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_128 UIV ( .A(S), .Y(SB) );
  ND2_384 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_383 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_382 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_381 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_380 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_379 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_127 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_127 UIV ( .A(S), .Y(SB) );
  ND2_381 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_380 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_379 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_378 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_377 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_376 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_126 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_126 UIV ( .A(S), .Y(SB) );
  ND2_378 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_377 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_376 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_375 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_374 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_373 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_125 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_125 UIV ( .A(S), .Y(SB) );
  ND2_375 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_374 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_373 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_372 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_371 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_370 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_124 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_124 UIV ( .A(S), .Y(SB) );
  ND2_372 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_371 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_370 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_369 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_368 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_367 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_123 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_123 UIV ( .A(S), .Y(SB) );
  ND2_369 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_368 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_367 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_366 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_365 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_364 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_122 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_122 UIV ( .A(S), .Y(SB) );
  ND2_366 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_365 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_364 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_363 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_362 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_361 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_121 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_121 UIV ( .A(S), .Y(SB) );
  ND2_363 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_362 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_361 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_360 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_359 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_358 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_120 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_120 UIV ( .A(S), .Y(SB) );
  ND2_360 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_359 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_358 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_357 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_356 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_355 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_119 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_119 UIV ( .A(S), .Y(SB) );
  ND2_357 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_356 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_355 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_354 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_353 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_352 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_118 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_118 UIV ( .A(S), .Y(SB) );
  ND2_354 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_353 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_352 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_351 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_350 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_349 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_117 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_117 UIV ( .A(S), .Y(SB) );
  ND2_351 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_350 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_349 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_348 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_347 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_346 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_116 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_116 UIV ( .A(S), .Y(SB) );
  ND2_348 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_347 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_346 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_345 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_344 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_343 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_115 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_115 UIV ( .A(S), .Y(SB) );
  ND2_345 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_344 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_343 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_342 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_341 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_340 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_114 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_114 UIV ( .A(S), .Y(SB) );
  ND2_342 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_341 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_340 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_339 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_338 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_337 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_113 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_113 UIV ( .A(S), .Y(SB) );
  ND2_339 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_338 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_337 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_336 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_335 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_334 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_112 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_112 UIV ( .A(S), .Y(SB) );
  ND2_336 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_335 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_334 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_333 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_332 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_331 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_111 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_111 UIV ( .A(S), .Y(SB) );
  ND2_333 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_332 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_331 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_330 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_329 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_328 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_110 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_110 UIV ( .A(S), .Y(SB) );
  ND2_330 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_329 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_328 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_327 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_326 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_325 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_109 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_109 UIV ( .A(S), .Y(SB) );
  ND2_327 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_326 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_325 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_324 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_323 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_322 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_108 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_108 UIV ( .A(S), .Y(SB) );
  ND2_324 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_323 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_322 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_321 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_320 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_319 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_107 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_107 UIV ( .A(S), .Y(SB) );
  ND2_321 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_320 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_319 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_318 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_317 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_316 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_106 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_106 UIV ( .A(S), .Y(SB) );
  ND2_318 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_317 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_316 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_315 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_314 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_313 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_105 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_105 UIV ( .A(S), .Y(SB) );
  ND2_315 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_314 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_313 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_312 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_311 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_310 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_104 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_104 UIV ( .A(S), .Y(SB) );
  ND2_312 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_311 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_310 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_309 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_308 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_307 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_103 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_103 UIV ( .A(S), .Y(SB) );
  ND2_309 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_308 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_307 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_306 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_305 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_304 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_102 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_102 UIV ( .A(S), .Y(SB) );
  ND2_306 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_305 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_304 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_303 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_302 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_301 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_101 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_101 UIV ( .A(S), .Y(SB) );
  ND2_303 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_302 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_301 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_300 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_299 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_298 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_100 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_100 UIV ( .A(S), .Y(SB) );
  ND2_300 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_299 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_298 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_297 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_296 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_295 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_99 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_99 UIV ( .A(S), .Y(SB) );
  ND2_297 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_296 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_295 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_294 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_293 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_292 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_98 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_98 UIV ( .A(S), .Y(SB) );
  ND2_294 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_293 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_292 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_291 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_290 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_289 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_97 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_97 UIV ( .A(S), .Y(SB) );
  ND2_291 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_290 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_289 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_128 gen1_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_127 gen1_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_126 gen1_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_125 gen1_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_124 gen1_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_123 gen1_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_122 gen1_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_121 gen1_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_120 gen1_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_119 gen1_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_118 gen1_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_117 gen1_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_116 gen1_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_115 gen1_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_114 gen1_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_113 gen1_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_112 gen1_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_111 gen1_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_110 gen1_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_109 gen1_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_108 gen1_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_107 gen1_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_106 gen1_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_105 gen1_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_104 gen1_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_103 gen1_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_102 gen1_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_101 gen1_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_100 gen1_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_99 gen1_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_98 gen1_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_97 gen1_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  CLKBUF_X3 U1 ( .A(SEL), .Z(n1) );
  CLKBUF_X3 U2 ( .A(SEL), .Z(n2) );
  CLKBUF_X3 U3 ( .A(SEL), .Z(n3) );
endmodule


module load_data ( data_in, signed_val, load_op, load_type, data_out );
  input [31:0] data_in;
  input [1:0] load_type;
  output [31:0] data_out;
  input signed_val, load_op;
  wire   N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30;

  DLH_X1 \data_out_reg[31]  ( .G(load_op), .D(N67), .Q(data_out[31]) );
  DLH_X1 \data_out_reg[30]  ( .G(load_op), .D(N66), .Q(data_out[30]) );
  DLH_X1 \data_out_reg[29]  ( .G(load_op), .D(N65), .Q(data_out[29]) );
  DLH_X1 \data_out_reg[28]  ( .G(load_op), .D(N64), .Q(data_out[28]) );
  DLH_X1 \data_out_reg[27]  ( .G(load_op), .D(N63), .Q(data_out[27]) );
  DLH_X1 \data_out_reg[26]  ( .G(load_op), .D(N62), .Q(data_out[26]) );
  DLH_X1 \data_out_reg[25]  ( .G(load_op), .D(N61), .Q(data_out[25]) );
  DLH_X1 \data_out_reg[24]  ( .G(load_op), .D(N60), .Q(data_out[24]) );
  DLH_X1 \data_out_reg[23]  ( .G(load_op), .D(N59), .Q(data_out[23]) );
  DLH_X1 \data_out_reg[22]  ( .G(load_op), .D(N58), .Q(data_out[22]) );
  DLH_X1 \data_out_reg[21]  ( .G(load_op), .D(N57), .Q(data_out[21]) );
  DLH_X1 \data_out_reg[20]  ( .G(load_op), .D(N56), .Q(data_out[20]) );
  DLH_X1 \data_out_reg[19]  ( .G(load_op), .D(N55), .Q(data_out[19]) );
  DLH_X1 \data_out_reg[18]  ( .G(load_op), .D(N54), .Q(data_out[18]) );
  DLH_X1 \data_out_reg[17]  ( .G(load_op), .D(N53), .Q(data_out[17]) );
  DLH_X1 \data_out_reg[16]  ( .G(load_op), .D(N52), .Q(data_out[16]) );
  DLH_X1 \data_out_reg[15]  ( .G(load_op), .D(N51), .Q(data_out[15]) );
  DLH_X1 \data_out_reg[14]  ( .G(load_op), .D(N50), .Q(data_out[14]) );
  DLH_X1 \data_out_reg[13]  ( .G(load_op), .D(N49), .Q(data_out[13]) );
  DLH_X1 \data_out_reg[12]  ( .G(load_op), .D(N48), .Q(data_out[12]) );
  DLH_X1 \data_out_reg[11]  ( .G(load_op), .D(N47), .Q(data_out[11]) );
  DLH_X1 \data_out_reg[10]  ( .G(load_op), .D(N46), .Q(data_out[10]) );
  DLH_X1 \data_out_reg[9]  ( .G(load_op), .D(N45), .Q(data_out[9]) );
  DLH_X1 \data_out_reg[8]  ( .G(load_op), .D(N44), .Q(data_out[8]) );
  DLH_X1 \data_out_reg[7]  ( .G(load_op), .D(N43), .Q(data_out[7]) );
  DLH_X1 \data_out_reg[6]  ( .G(load_op), .D(N42), .Q(data_out[6]) );
  DLH_X1 \data_out_reg[5]  ( .G(load_op), .D(N41), .Q(data_out[5]) );
  DLH_X1 \data_out_reg[4]  ( .G(load_op), .D(N40), .Q(data_out[4]) );
  DLH_X1 \data_out_reg[3]  ( .G(load_op), .D(N39), .Q(data_out[3]) );
  DLH_X1 \data_out_reg[2]  ( .G(load_op), .D(N38), .Q(data_out[2]) );
  DLH_X1 \data_out_reg[1]  ( .G(load_op), .D(N37), .Q(data_out[1]) );
  DLH_X1 \data_out_reg[0]  ( .G(load_op), .D(N36), .Q(data_out[0]) );
  OAI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(N67) );
  NAND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(N66) );
  NAND2_X1 U4 ( .A1(data_in[30]), .A2(n5), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n3), .A2(n6), .ZN(N65) );
  NAND2_X1 U6 ( .A1(data_in[29]), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n3), .A2(n7), .ZN(N64) );
  NAND2_X1 U8 ( .A1(data_in[28]), .A2(n5), .ZN(n7) );
  NAND2_X1 U9 ( .A1(n3), .A2(n8), .ZN(N63) );
  NAND2_X1 U10 ( .A1(data_in[27]), .A2(n5), .ZN(n8) );
  NAND2_X1 U11 ( .A1(n3), .A2(n9), .ZN(N62) );
  NAND2_X1 U12 ( .A1(data_in[26]), .A2(n5), .ZN(n9) );
  NAND2_X1 U13 ( .A1(n3), .A2(n10), .ZN(N61) );
  NAND2_X1 U14 ( .A1(data_in[25]), .A2(n5), .ZN(n10) );
  NAND2_X1 U15 ( .A1(n3), .A2(n11), .ZN(N60) );
  NAND2_X1 U16 ( .A1(data_in[24]), .A2(n5), .ZN(n11) );
  NAND2_X1 U17 ( .A1(n3), .A2(n12), .ZN(N59) );
  NAND2_X1 U18 ( .A1(data_in[23]), .A2(n5), .ZN(n12) );
  NAND2_X1 U19 ( .A1(n3), .A2(n13), .ZN(N58) );
  NAND2_X1 U20 ( .A1(data_in[22]), .A2(n5), .ZN(n13) );
  NAND2_X1 U21 ( .A1(n3), .A2(n14), .ZN(N57) );
  NAND2_X1 U22 ( .A1(data_in[21]), .A2(n5), .ZN(n14) );
  NAND2_X1 U23 ( .A1(n3), .A2(n15), .ZN(N56) );
  NAND2_X1 U24 ( .A1(data_in[20]), .A2(n5), .ZN(n15) );
  NAND2_X1 U25 ( .A1(n3), .A2(n16), .ZN(N55) );
  NAND2_X1 U26 ( .A1(data_in[19]), .A2(n5), .ZN(n16) );
  NAND2_X1 U27 ( .A1(n3), .A2(n17), .ZN(N54) );
  NAND2_X1 U28 ( .A1(data_in[18]), .A2(n5), .ZN(n17) );
  NAND2_X1 U29 ( .A1(n3), .A2(n18), .ZN(N53) );
  NAND2_X1 U30 ( .A1(data_in[17]), .A2(n5), .ZN(n18) );
  NAND2_X1 U31 ( .A1(n3), .A2(n19), .ZN(N52) );
  NAND2_X1 U32 ( .A1(data_in[16]), .A2(n5), .ZN(n19) );
  INV_X1 U33 ( .A(n1), .ZN(n5) );
  NAND2_X1 U34 ( .A1(load_type[1]), .A2(load_type[0]), .ZN(n1) );
  NAND2_X1 U35 ( .A1(n3), .A2(n20), .ZN(N51) );
  NAND2_X1 U36 ( .A1(data_in[15]), .A2(load_type[0]), .ZN(n20) );
  NAND2_X1 U37 ( .A1(n3), .A2(n21), .ZN(N50) );
  NAND2_X1 U38 ( .A1(data_in[14]), .A2(load_type[0]), .ZN(n21) );
  NAND2_X1 U39 ( .A1(n3), .A2(n22), .ZN(N49) );
  NAND2_X1 U40 ( .A1(data_in[13]), .A2(load_type[0]), .ZN(n22) );
  NAND2_X1 U41 ( .A1(n3), .A2(n23), .ZN(N48) );
  NAND2_X1 U42 ( .A1(data_in[12]), .A2(load_type[0]), .ZN(n23) );
  NAND2_X1 U43 ( .A1(n3), .A2(n24), .ZN(N47) );
  NAND2_X1 U44 ( .A1(data_in[11]), .A2(load_type[0]), .ZN(n24) );
  NAND2_X1 U45 ( .A1(n3), .A2(n25), .ZN(N46) );
  NAND2_X1 U46 ( .A1(data_in[10]), .A2(load_type[0]), .ZN(n25) );
  NAND2_X1 U47 ( .A1(n3), .A2(n26), .ZN(N45) );
  NAND2_X1 U48 ( .A1(data_in[9]), .A2(load_type[0]), .ZN(n26) );
  NAND2_X1 U49 ( .A1(n3), .A2(n27), .ZN(N44) );
  NAND2_X1 U50 ( .A1(data_in[8]), .A2(load_type[0]), .ZN(n27) );
  OR3_X1 U51 ( .A1(signed_val), .A2(n2), .A3(n28), .ZN(n3) );
  INV_X1 U52 ( .A(data_in[31]), .ZN(n2) );
  AND2_X1 U53 ( .A1(data_in[7]), .A2(n29), .ZN(N43) );
  AND2_X1 U54 ( .A1(data_in[6]), .A2(n29), .ZN(N42) );
  AND2_X1 U55 ( .A1(data_in[5]), .A2(n29), .ZN(N41) );
  AND2_X1 U56 ( .A1(data_in[4]), .A2(n29), .ZN(N40) );
  AND2_X1 U57 ( .A1(data_in[3]), .A2(n29), .ZN(N39) );
  AND2_X1 U58 ( .A1(data_in[2]), .A2(n29), .ZN(N38) );
  AND2_X1 U59 ( .A1(data_in[1]), .A2(n29), .ZN(N37) );
  AND2_X1 U60 ( .A1(data_in[0]), .A2(n29), .ZN(N36) );
  NAND2_X1 U61 ( .A1(n30), .A2(n28), .ZN(n29) );
  OR2_X1 U62 ( .A1(load_type[1]), .A2(load_type[0]), .ZN(n28) );
  INV_X1 U63 ( .A(load_type[0]), .ZN(n30) );
endmodule


module regFFD_NBIT32_3 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT32_2 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module regFFD_NBIT5_1 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \Q_reg[4]  ( .D(n16), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n21) );
  DFFR_X1 \Q_reg[3]  ( .D(n17), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n22) );
  DFFR_X1 \Q_reg[2]  ( .D(n18), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n23) );
  DFFR_X1 \Q_reg[1]  ( .D(n19), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n24) );
  DFFR_X1 \Q_reg[0]  ( .D(n20), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n25) );
  OAI21_X1 U2 ( .B1(n25), .B2(ENABLE), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(ENABLE), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(ENABLE), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(ENABLE), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(ENABLE), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n26) );
endmodule


module FF_3 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n5, n6, n7, n8;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n8), .A2(n7), .ZN(n5) );
  INV_X1 U4 ( .A(RESET), .ZN(n7) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n6), .ZN(n8) );
  INV_X1 U6 ( .A(EN), .ZN(n6) );
endmodule


module FF_2 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n5, n6, n7, n8;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n8), .A2(n7), .ZN(n5) );
  INV_X1 U4 ( .A(RESET), .ZN(n7) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n6), .ZN(n8) );
  INV_X1 U6 ( .A(EN), .ZN(n6) );
endmodule


module FF_1 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n11, n5, n7, n8, n9, n10;

  DFF_X1 Q_reg ( .D(n7), .CK(CLK), .Q(n11) );
  NOR2_X1 U3 ( .A1(n10), .A2(n9), .ZN(n7) );
  INV_X1 U4 ( .A(RESET), .ZN(n9) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(Q), .B2(n8), .ZN(n10) );
  INV_X1 U6 ( .A(EN), .ZN(n8) );
  INV_X1 U7 ( .A(n11), .ZN(n5) );
  INV_X4 U8 ( .A(n5), .ZN(Q) );
endmodule


module regFFD_NBIT32_1 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192;

  DFFR_X1 \Q_reg[31]  ( .D(n97), .CK(CK), .RN(RESET), .Q(Q[31]), .QN(n129) );
  DFFR_X1 \Q_reg[30]  ( .D(n98), .CK(CK), .RN(RESET), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n99), .CK(CK), .RN(RESET), .Q(Q[29]), .QN(n131) );
  DFFR_X1 \Q_reg[28]  ( .D(n100), .CK(CK), .RN(RESET), .Q(Q[28]), .QN(n132) );
  DFFR_X1 \Q_reg[27]  ( .D(n101), .CK(CK), .RN(RESET), .Q(Q[27]), .QN(n133) );
  DFFR_X1 \Q_reg[26]  ( .D(n102), .CK(CK), .RN(RESET), .Q(Q[26]), .QN(n134) );
  DFFR_X1 \Q_reg[25]  ( .D(n103), .CK(CK), .RN(RESET), .Q(Q[25]), .QN(n135) );
  DFFR_X1 \Q_reg[24]  ( .D(n104), .CK(CK), .RN(RESET), .Q(Q[24]), .QN(n136) );
  DFFR_X1 \Q_reg[23]  ( .D(n105), .CK(CK), .RN(RESET), .Q(Q[23]), .QN(n137) );
  DFFR_X1 \Q_reg[22]  ( .D(n106), .CK(CK), .RN(RESET), .Q(Q[22]), .QN(n138) );
  DFFR_X1 \Q_reg[21]  ( .D(n107), .CK(CK), .RN(RESET), .Q(Q[21]), .QN(n139) );
  DFFR_X1 \Q_reg[20]  ( .D(n108), .CK(CK), .RN(RESET), .Q(Q[20]), .QN(n140) );
  DFFR_X1 \Q_reg[19]  ( .D(n109), .CK(CK), .RN(RESET), .Q(Q[19]), .QN(n141) );
  DFFR_X1 \Q_reg[18]  ( .D(n110), .CK(CK), .RN(RESET), .Q(Q[18]), .QN(n142) );
  DFFR_X1 \Q_reg[17]  ( .D(n111), .CK(CK), .RN(RESET), .Q(Q[17]), .QN(n143) );
  DFFR_X1 \Q_reg[16]  ( .D(n112), .CK(CK), .RN(RESET), .Q(Q[16]), .QN(n144) );
  DFFR_X1 \Q_reg[15]  ( .D(n113), .CK(CK), .RN(RESET), .Q(Q[15]), .QN(n145) );
  DFFR_X1 \Q_reg[14]  ( .D(n114), .CK(CK), .RN(RESET), .Q(Q[14]), .QN(n146) );
  DFFR_X1 \Q_reg[13]  ( .D(n115), .CK(CK), .RN(RESET), .Q(Q[13]), .QN(n147) );
  DFFR_X1 \Q_reg[12]  ( .D(n116), .CK(CK), .RN(RESET), .Q(Q[12]), .QN(n148) );
  DFFR_X1 \Q_reg[11]  ( .D(n117), .CK(CK), .RN(RESET), .Q(Q[11]), .QN(n149) );
  DFFR_X1 \Q_reg[10]  ( .D(n118), .CK(CK), .RN(RESET), .Q(Q[10]), .QN(n150) );
  DFFR_X1 \Q_reg[9]  ( .D(n119), .CK(CK), .RN(RESET), .Q(Q[9]), .QN(n151) );
  DFFR_X1 \Q_reg[8]  ( .D(n120), .CK(CK), .RN(RESET), .Q(Q[8]), .QN(n152) );
  DFFR_X1 \Q_reg[7]  ( .D(n121), .CK(CK), .RN(RESET), .Q(Q[7]), .QN(n153) );
  DFFR_X1 \Q_reg[6]  ( .D(n122), .CK(CK), .RN(RESET), .Q(Q[6]), .QN(n154) );
  DFFR_X1 \Q_reg[5]  ( .D(n123), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n155) );
  DFFR_X1 \Q_reg[4]  ( .D(n124), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n156) );
  DFFR_X1 \Q_reg[3]  ( .D(n125), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n157) );
  DFFR_X1 \Q_reg[2]  ( .D(n126), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n158) );
  DFFR_X1 \Q_reg[1]  ( .D(n127), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n159) );
  DFFR_X1 \Q_reg[0]  ( .D(n128), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n160) );
  OAI21_X1 U2 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n192) );
  OAI21_X1 U4 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U6 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U8 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U10 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U12 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U14 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U15 ( .A1(D[6]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U16 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U17 ( .A1(D[7]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U18 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U19 ( .A1(D[8]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U20 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U21 ( .A1(D[9]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U22 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U23 ( .A1(D[10]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U24 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U25 ( .A1(D[11]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U26 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U27 ( .A1(D[12]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U28 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U29 ( .A1(D[13]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U30 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U31 ( .A1(D[14]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U32 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U33 ( .A1(D[15]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U34 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U35 ( .A1(D[16]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U36 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U37 ( .A1(D[17]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U38 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U39 ( .A1(D[18]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U40 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U41 ( .A1(D[19]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U42 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U43 ( .A1(D[20]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U44 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U45 ( .A1(D[21]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U46 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U47 ( .A1(D[22]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U48 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U49 ( .A1(D[23]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U50 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U51 ( .A1(D[24]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U52 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U53 ( .A1(D[25]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U54 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U55 ( .A1(D[26]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U56 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U57 ( .A1(D[27]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U58 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U59 ( .A1(D[28]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U60 ( .B1(n131), .B2(ENABLE), .A(n163), .ZN(n99) );
  NAND2_X1 U61 ( .A1(D[29]), .A2(ENABLE), .ZN(n163) );
  OAI21_X1 U62 ( .B1(n130), .B2(ENABLE), .A(n162), .ZN(n98) );
  NAND2_X1 U63 ( .A1(D[30]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U64 ( .B1(n129), .B2(ENABLE), .A(n161), .ZN(n97) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(ENABLE), .ZN(n161) );
endmodule


module IV_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_288 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_287 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_286 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_96 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_96 UIV ( .A(S), .Y(SB) );
  ND2_288 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_287 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_286 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_285 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_284 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_283 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_95 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_95 UIV ( .A(S), .Y(SB) );
  ND2_285 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_284 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_283 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_282 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_281 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_280 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_94 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_94 UIV ( .A(S), .Y(SB) );
  ND2_282 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_281 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_280 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_279 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_278 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_277 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_93 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_93 UIV ( .A(S), .Y(SB) );
  ND2_279 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_278 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_277 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_276 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_275 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_274 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_92 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_92 UIV ( .A(S), .Y(SB) );
  ND2_276 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_275 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_274 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_273 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_272 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_271 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_91 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_91 UIV ( .A(S), .Y(SB) );
  ND2_273 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_272 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_271 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_270 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_269 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_268 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_90 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_90 UIV ( .A(S), .Y(SB) );
  ND2_270 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_269 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_268 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_267 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_266 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_265 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_89 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_89 UIV ( .A(S), .Y(SB) );
  ND2_267 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_266 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_265 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_264 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_263 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_262 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_88 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_88 UIV ( .A(S), .Y(SB) );
  ND2_264 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_263 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_262 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_261 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_260 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_259 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_87 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_87 UIV ( .A(S), .Y(SB) );
  ND2_261 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_260 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_259 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_258 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_257 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_256 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_86 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_86 UIV ( .A(S), .Y(SB) );
  ND2_258 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_257 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_256 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_255 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_254 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_253 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_85 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_85 UIV ( .A(S), .Y(SB) );
  ND2_255 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_254 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_253 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_252 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_251 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_250 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_84 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_84 UIV ( .A(S), .Y(SB) );
  ND2_252 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_251 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_250 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_249 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_248 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_247 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_83 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_83 UIV ( .A(S), .Y(SB) );
  ND2_249 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_248 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_247 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_246 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_245 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_244 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_82 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_82 UIV ( .A(S), .Y(SB) );
  ND2_246 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_245 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_244 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_243 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_242 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_241 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_81 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_81 UIV ( .A(S), .Y(SB) );
  ND2_243 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_242 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_241 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_240 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_239 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_238 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_80 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_80 UIV ( .A(S), .Y(SB) );
  ND2_240 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_239 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_238 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_237 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_236 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_235 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_79 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_79 UIV ( .A(S), .Y(SB) );
  ND2_237 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_236 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_235 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_234 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_233 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_232 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_78 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_78 UIV ( .A(S), .Y(SB) );
  ND2_234 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_233 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_232 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_231 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_230 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_229 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_77 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_77 UIV ( .A(S), .Y(SB) );
  ND2_231 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_230 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_229 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_228 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_227 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_226 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_76 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_76 UIV ( .A(S), .Y(SB) );
  ND2_228 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_227 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_226 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_225 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_224 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_223 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_75 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_75 UIV ( .A(S), .Y(SB) );
  ND2_225 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_224 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_223 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_222 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_221 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_220 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_74 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_74 UIV ( .A(S), .Y(SB) );
  ND2_222 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_221 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_220 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_219 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_218 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_217 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_73 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_73 UIV ( .A(S), .Y(SB) );
  ND2_219 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_218 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_217 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_216 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_215 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_214 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_72 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_72 UIV ( .A(S), .Y(SB) );
  ND2_216 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_215 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_214 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_213 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_212 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_211 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_71 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_71 UIV ( .A(S), .Y(SB) );
  ND2_213 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_212 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_211 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_210 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_209 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_208 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_70 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_70 UIV ( .A(S), .Y(SB) );
  ND2_210 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_209 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_208 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_207 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_206 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_205 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_69 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_69 UIV ( .A(S), .Y(SB) );
  ND2_207 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_206 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_205 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_204 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_203 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_202 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_68 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_68 UIV ( .A(S), .Y(SB) );
  ND2_204 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_203 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_202 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_201 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_200 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_199 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_67 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_67 UIV ( .A(S), .Y(SB) );
  ND2_201 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_200 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_199 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_198 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_197 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_196 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_66 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_66 UIV ( .A(S), .Y(SB) );
  ND2_198 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_197 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_196 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_195 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_194 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_193 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_65 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_65 UIV ( .A(S), .Y(SB) );
  ND2_195 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_194 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_193 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_96 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_95 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_94 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_93 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_92 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_91 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_90 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_89 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_88 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_87 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_86 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_85 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_84 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_83 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_82 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_81 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_80 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_79 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_78 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_77 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_76 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_75 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_74 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_73 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_72 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_71 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_70 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_69 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_68 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_67 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_66 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_65 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_192 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_64 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_64 UIV ( .A(S), .Y(SB) );
  ND2_192 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_191 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_190 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_63 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_63 UIV ( .A(S), .Y(SB) );
  ND2_189 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_188 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_187 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_62 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_62 UIV ( .A(S), .Y(SB) );
  ND2_186 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_185 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_184 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_61 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_61 UIV ( .A(S), .Y(SB) );
  ND2_183 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_182 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_181 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_60 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_60 UIV ( .A(S), .Y(SB) );
  ND2_180 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_179 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_178 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_59 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_59 UIV ( .A(S), .Y(SB) );
  ND2_177 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_176 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_175 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_58 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_58 UIV ( .A(S), .Y(SB) );
  ND2_174 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_173 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_172 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_57 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_57 UIV ( .A(S), .Y(SB) );
  ND2_171 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_170 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_169 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_56 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_56 UIV ( .A(S), .Y(SB) );
  ND2_168 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_167 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_166 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_55 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_55 UIV ( .A(S), .Y(SB) );
  ND2_165 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_164 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_163 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_54 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_54 UIV ( .A(S), .Y(SB) );
  ND2_162 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_161 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_160 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_53 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_53 UIV ( .A(S), .Y(SB) );
  ND2_159 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_158 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_157 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_52 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_52 UIV ( .A(S), .Y(SB) );
  ND2_156 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_155 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_154 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_51 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_51 UIV ( .A(S), .Y(SB) );
  ND2_153 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_152 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_151 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_50 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_50 UIV ( .A(S), .Y(SB) );
  ND2_150 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_149 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_148 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_49 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_49 UIV ( .A(S), .Y(SB) );
  ND2_147 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_146 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_145 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_48 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_48 UIV ( .A(S), .Y(SB) );
  ND2_144 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_143 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_142 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_47 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_47 UIV ( .A(S), .Y(SB) );
  ND2_141 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_140 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_139 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_46 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_46 UIV ( .A(S), .Y(SB) );
  ND2_138 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_137 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_136 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_45 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_45 UIV ( .A(S), .Y(SB) );
  ND2_135 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_134 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_133 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_44 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_44 UIV ( .A(S), .Y(SB) );
  ND2_132 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_131 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_130 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_43 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_43 UIV ( .A(S), .Y(SB) );
  ND2_129 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_128 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_127 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_42 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_42 UIV ( .A(S), .Y(SB) );
  ND2_126 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_125 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_124 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_41 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_41 UIV ( .A(S), .Y(SB) );
  ND2_123 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_122 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_121 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_40 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_40 UIV ( .A(S), .Y(SB) );
  ND2_120 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_119 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_118 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_39 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_39 UIV ( .A(S), .Y(SB) );
  ND2_117 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_116 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_115 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_38 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_38 UIV ( .A(S), .Y(SB) );
  ND2_114 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_113 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_112 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_37 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_37 UIV ( .A(S), .Y(SB) );
  ND2_111 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_110 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_109 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_36 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_36 UIV ( .A(S), .Y(SB) );
  ND2_108 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_107 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_106 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_35 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_35 UIV ( .A(S), .Y(SB) );
  ND2_105 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_104 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_103 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_34 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_34 UIV ( .A(S), .Y(SB) );
  ND2_102 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_101 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_100 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;
  wire   N1;
  assign Y = N1;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(N1) );
endmodule


module MUX21_33 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_33 UIV ( .A(S), .Y(SB) );
  ND2_99 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_98 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_97 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_64 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_63 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_62 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_61 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_60 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_59 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_58 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_57 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_56 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_55 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_54 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_53 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_52 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_51 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_50 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_49 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_48 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_47 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_46 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_45 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_44 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_43 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_42 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_41 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_40 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_39 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_38 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_37 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_36 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_35 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_34 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_33 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[31]), .B(A[31]), .Z(SUM[31]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module DATAPTH_NBIT32_REG_BIT5 ( CLK, RST, PC, IR, PC_OUT, NPC_LATCH_EN, 
        ir_LATCH_EN, signed_op, RF1, RF2, WF1, regImm_LATCH_EN, S1, S2, EN2, 
        lhi_sel, jump_en, branch_cond, sb_op, RM, WM, EN3, S3, 
    .instruction_alu({\instruction_alu[5] , \instruction_alu[4] , 
        \instruction_alu[3] , \instruction_alu[2] , \instruction_alu[1] , 
        \instruction_alu[0] }), DATA_MEM_ADDR, DATA_MEM_IN, DATA_MEM_OUT, 
        DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM );
  input [31:0] PC;
  input [31:0] IR;
  output [31:0] PC_OUT;
  output [31:0] DATA_MEM_ADDR;
  output [31:0] DATA_MEM_IN;
  input [31:0] DATA_MEM_OUT;
  input CLK, RST, NPC_LATCH_EN, ir_LATCH_EN, signed_op, RF1, RF2, WF1,
         regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond, sb_op,
         RM, WM, EN3, S3, \instruction_alu[5] , \instruction_alu[4] ,
         \instruction_alu[3] , \instruction_alu[2] , \instruction_alu[1] ,
         \instruction_alu[0] ;
  output DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM;
  wire   RM, WM, sel_npc, wr_signal, wr_signal_wb, signed_op_ex, wr_signal_exe,
         is_zero, cond, signed_op_mem, cond_mem, wr_signal_mem, sel_saved_reg,
         N14, wr_signal_mem1, sel_saved_reg_wb, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45;
  wire   [5:0] instruction_alu;
  wire   [31:0] PC_fetch0;
  wire   [31:0] NPC;
  wire   [31:0] NPC_fetch1;
  wire   [31:0] PC_fetch1;
  wire   [31:0] PC_OUT_i;
  wire   [31:0] NPC_fetch;
  wire   [31:0] PC_fetch;
  wire   [31:0] ir_fetch;
  wire   [31:0] NPC_Dec;
  wire   [31:0] IR_Dec;
  wire   [4:0] RS1;
  wire   [4:0] RS2;
  wire   [4:0] RD;
  wire   [31:0] Imm;
  wire   [4:0] RD_wb;
  wire   [31:0] OUT_data;
  wire   [31:0] regA;
  wire   [31:0] regB;
  wire   [31:0] NPC_ex;
  wire   [31:0] regA_ex;
  wire   [31:0] regB_ex;
  wire   [31:0] Imm_ex;
  wire   [4:0] RD_ex;
  wire   [5:0] IR_26_ex;
  wire   [31:0] LHI_ex;
  wire   [31:0] input1_ALU;
  wire   [31:0] input2_ALU;
  wire   [31:0] ALU_out;
  wire   [31:0] ALU_ex;
  wire   [31:0] NPC_mem;
  wire   [31:0] regB_mem;
  wire   [4:0] RD_mem;
  wire   [5:0] IR_26_mem;
  wire   [31:0] LMD_out;
  wire   [31:0] ALU_wb;
  wire   [31:0] LMD_wb;
  wire   [31:0] NPC_wb;
  assign DATA_MEM_RM = RM;
  assign DATA_MEM_WM = WM;

  DLH_X1 \DATA_MEM_ADDR_reg[31]  ( .G(N14), .D(ALU_ex[31]), .Q(
        DATA_MEM_ADDR[31]) );
  DLH_X1 \DATA_MEM_ADDR_reg[30]  ( .G(N14), .D(ALU_ex[30]), .Q(
        DATA_MEM_ADDR[30]) );
  DLH_X1 \DATA_MEM_ADDR_reg[29]  ( .G(N14), .D(ALU_ex[29]), .Q(
        DATA_MEM_ADDR[29]) );
  DLH_X1 \DATA_MEM_ADDR_reg[28]  ( .G(N14), .D(ALU_ex[28]), .Q(
        DATA_MEM_ADDR[28]) );
  DLH_X1 \DATA_MEM_ADDR_reg[27]  ( .G(N14), .D(ALU_ex[27]), .Q(
        DATA_MEM_ADDR[27]) );
  DLH_X1 \DATA_MEM_ADDR_reg[26]  ( .G(N14), .D(ALU_ex[26]), .Q(
        DATA_MEM_ADDR[26]) );
  DLH_X1 \DATA_MEM_ADDR_reg[25]  ( .G(N14), .D(ALU_ex[25]), .Q(
        DATA_MEM_ADDR[25]) );
  DLH_X1 \DATA_MEM_ADDR_reg[24]  ( .G(N14), .D(ALU_ex[24]), .Q(
        DATA_MEM_ADDR[24]) );
  DLH_X1 \DATA_MEM_ADDR_reg[23]  ( .G(N14), .D(ALU_ex[23]), .Q(
        DATA_MEM_ADDR[23]) );
  DLH_X1 \DATA_MEM_ADDR_reg[22]  ( .G(N14), .D(ALU_ex[22]), .Q(
        DATA_MEM_ADDR[22]) );
  DLH_X1 \DATA_MEM_ADDR_reg[21]  ( .G(N14), .D(ALU_ex[21]), .Q(
        DATA_MEM_ADDR[21]) );
  DLH_X1 \DATA_MEM_ADDR_reg[20]  ( .G(N14), .D(ALU_ex[20]), .Q(
        DATA_MEM_ADDR[20]) );
  DLH_X1 \DATA_MEM_ADDR_reg[19]  ( .G(N14), .D(ALU_ex[19]), .Q(
        DATA_MEM_ADDR[19]) );
  DLH_X1 \DATA_MEM_ADDR_reg[18]  ( .G(N14), .D(ALU_ex[18]), .Q(
        DATA_MEM_ADDR[18]) );
  DLH_X1 \DATA_MEM_ADDR_reg[17]  ( .G(N14), .D(ALU_ex[17]), .Q(
        DATA_MEM_ADDR[17]) );
  DLH_X1 \DATA_MEM_ADDR_reg[16]  ( .G(N14), .D(ALU_ex[16]), .Q(
        DATA_MEM_ADDR[16]) );
  DLH_X1 \DATA_MEM_ADDR_reg[15]  ( .G(N14), .D(ALU_ex[15]), .Q(
        DATA_MEM_ADDR[15]) );
  DLH_X1 \DATA_MEM_ADDR_reg[14]  ( .G(N14), .D(ALU_ex[14]), .Q(
        DATA_MEM_ADDR[14]) );
  DLH_X1 \DATA_MEM_ADDR_reg[13]  ( .G(N14), .D(ALU_ex[13]), .Q(
        DATA_MEM_ADDR[13]) );
  DLH_X1 \DATA_MEM_ADDR_reg[12]  ( .G(N14), .D(ALU_ex[12]), .Q(
        DATA_MEM_ADDR[12]) );
  DLH_X1 \DATA_MEM_ADDR_reg[11]  ( .G(N14), .D(ALU_ex[11]), .Q(
        DATA_MEM_ADDR[11]) );
  DLH_X1 \DATA_MEM_ADDR_reg[10]  ( .G(N14), .D(ALU_ex[10]), .Q(
        DATA_MEM_ADDR[10]) );
  DLH_X1 \DATA_MEM_ADDR_reg[9]  ( .G(N14), .D(ALU_ex[9]), .Q(DATA_MEM_ADDR[9])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[8]  ( .G(N14), .D(ALU_ex[8]), .Q(DATA_MEM_ADDR[8])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[7]  ( .G(N14), .D(ALU_ex[7]), .Q(DATA_MEM_ADDR[7])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[6]  ( .G(N14), .D(ALU_ex[6]), .Q(DATA_MEM_ADDR[6])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[5]  ( .G(N14), .D(ALU_ex[5]), .Q(DATA_MEM_ADDR[5])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[4]  ( .G(N14), .D(ALU_ex[4]), .Q(DATA_MEM_ADDR[4])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[3]  ( .G(N14), .D(ALU_ex[3]), .Q(DATA_MEM_ADDR[3])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[2]  ( .G(N14), .D(ALU_ex[2]), .Q(DATA_MEM_ADDR[2])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[1]  ( .G(N14), .D(ALU_ex[1]), .Q(DATA_MEM_ADDR[1])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[0]  ( .G(N14), .D(ALU_ex[0]), .Q(DATA_MEM_ADDR[0])
         );
  NOR2_X1 U3 ( .A1(n1), .A2(jump_en), .ZN(wr_signal_mem1) );
  INV_X1 U4 ( .A(wr_signal_mem), .ZN(n1) );
  INV_X1 U5 ( .A(n2), .ZN(wr_signal) );
  OAI33_X1 U6 ( .A1(n3), .A2(n42), .A3(n45), .B1(n4), .B2(n5), .B3(n6), .ZN(n2) );
  XOR2_X1 U7 ( .A(IR_Dec[27]), .B(n40), .Z(n6) );
  INV_X1 U8 ( .A(n42), .ZN(n5) );
  NAND3_X1 U9 ( .A1(n7), .A2(n8), .A3(n45), .ZN(n4) );
  NAND2_X1 U10 ( .A1(n9), .A2(n10), .ZN(n3) );
  INV_X1 U11 ( .A(IR_Dec[27]), .ZN(n10) );
  OAI33_X1 U12 ( .A1(n8), .A2(n11), .A3(n7), .B1(n12), .B2(n13), .B3(n14), 
        .ZN(n9) );
  OR4_X1 U13 ( .A1(IR_Dec[11]), .A2(IR_Dec[10]), .A3(IR_Dec[0]), .A4(n15), 
        .ZN(n14) );
  OR4_X1 U14 ( .A1(IR_Dec[13]), .A2(IR_Dec[12]), .A3(IR_Dec[15]), .A4(
        IR_Dec[14]), .ZN(n15) );
  OR4_X1 U15 ( .A1(IR_Dec[18]), .A2(IR_Dec[17]), .A3(IR_Dec[16]), .A4(n16), 
        .ZN(n13) );
  OR4_X1 U16 ( .A1(IR_Dec[1]), .A2(IR_Dec[19]), .A3(IR_Dec[21]), .A4(
        IR_Dec[20]), .ZN(n16) );
  NAND4_X1 U17 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .ZN(n12) );
  NOR4_X1 U18 ( .A1(IR_Dec[9]), .A2(IR_Dec[8]), .A3(IR_Dec[7]), .A4(IR_Dec[6]), 
        .ZN(n20) );
  NOR4_X1 U19 ( .A1(IR_Dec[5]), .A2(IR_Dec[4]), .A3(IR_Dec[3]), .A4(n43), .ZN(
        n19) );
  NOR4_X1 U20 ( .A1(IR_Dec[2]), .A2(IR_Dec[28]), .A3(IR_Dec[26]), .A4(
        IR_Dec[25]), .ZN(n18) );
  NOR3_X1 U21 ( .A1(IR_Dec[22]), .A2(IR_Dec[24]), .A3(IR_Dec[23]), .ZN(n17) );
  INV_X1 U22 ( .A(IR_Dec[28]), .ZN(n7) );
  INV_X1 U23 ( .A(n40), .ZN(n11) );
  INV_X1 U24 ( .A(n41), .ZN(n8) );
  AND2_X1 U25 ( .A1(IR_26_mem[0]), .A2(jump_en), .ZN(sel_saved_reg) );
  OR2_X1 U26 ( .A1(cond_mem), .A2(jump_en), .ZN(sel_npc) );
  NAND4_X1 U27 ( .A1(IR_26_mem[2]), .A2(IR_26_mem[0]), .A3(IR_26_mem[4]), .A4(
        n21), .ZN(N14) );
  NOR3_X1 U28 ( .A1(IR_26_mem[1]), .A2(IR_26_mem[5]), .A3(IR_26_mem[3]), .ZN(
        n21) );
  AND2_X1 U29 ( .A1(regB_mem[9]), .A2(n22), .ZN(DATA_MEM_IN[9]) );
  AND2_X1 U30 ( .A1(regB_mem[8]), .A2(n22), .ZN(DATA_MEM_IN[8]) );
  INV_X1 U31 ( .A(n23), .ZN(DATA_MEM_IN[7]) );
  AOI22_X1 U32 ( .A1(n22), .A2(regB_mem[7]), .B1(regB_mem[31]), .B2(sb_op), 
        .ZN(n23) );
  INV_X1 U33 ( .A(n24), .ZN(DATA_MEM_IN[6]) );
  AOI22_X1 U34 ( .A1(n22), .A2(regB_mem[6]), .B1(sb_op), .B2(regB_mem[30]), 
        .ZN(n24) );
  INV_X1 U35 ( .A(n25), .ZN(DATA_MEM_IN[5]) );
  AOI22_X1 U36 ( .A1(n22), .A2(regB_mem[5]), .B1(sb_op), .B2(regB_mem[29]), 
        .ZN(n25) );
  INV_X1 U37 ( .A(n26), .ZN(DATA_MEM_IN[4]) );
  AOI22_X1 U38 ( .A1(n22), .A2(regB_mem[4]), .B1(sb_op), .B2(regB_mem[28]), 
        .ZN(n26) );
  INV_X1 U39 ( .A(n27), .ZN(DATA_MEM_IN[3]) );
  AOI22_X1 U40 ( .A1(n22), .A2(regB_mem[3]), .B1(sb_op), .B2(regB_mem[27]), 
        .ZN(n27) );
  AND2_X1 U41 ( .A1(n22), .A2(regB_mem[31]), .ZN(DATA_MEM_IN[31]) );
  AND2_X1 U42 ( .A1(n22), .A2(regB_mem[30]), .ZN(DATA_MEM_IN[30]) );
  INV_X1 U43 ( .A(n28), .ZN(DATA_MEM_IN[2]) );
  AOI22_X1 U44 ( .A1(n22), .A2(regB_mem[2]), .B1(sb_op), .B2(regB_mem[26]), 
        .ZN(n28) );
  AND2_X1 U45 ( .A1(n22), .A2(regB_mem[29]), .ZN(DATA_MEM_IN[29]) );
  AND2_X1 U46 ( .A1(n22), .A2(regB_mem[28]), .ZN(DATA_MEM_IN[28]) );
  AND2_X1 U47 ( .A1(n22), .A2(regB_mem[27]), .ZN(DATA_MEM_IN[27]) );
  AND2_X1 U48 ( .A1(n22), .A2(regB_mem[26]), .ZN(DATA_MEM_IN[26]) );
  AND2_X1 U49 ( .A1(n22), .A2(regB_mem[25]), .ZN(DATA_MEM_IN[25]) );
  AND2_X1 U50 ( .A1(n22), .A2(regB_mem[24]), .ZN(DATA_MEM_IN[24]) );
  AND2_X1 U51 ( .A1(regB_mem[23]), .A2(n22), .ZN(DATA_MEM_IN[23]) );
  AND2_X1 U52 ( .A1(regB_mem[22]), .A2(n22), .ZN(DATA_MEM_IN[22]) );
  AND2_X1 U53 ( .A1(regB_mem[21]), .A2(n22), .ZN(DATA_MEM_IN[21]) );
  AND2_X1 U54 ( .A1(regB_mem[20]), .A2(n22), .ZN(DATA_MEM_IN[20]) );
  INV_X1 U55 ( .A(n29), .ZN(DATA_MEM_IN[1]) );
  AOI22_X1 U56 ( .A1(sb_op), .A2(regB_mem[25]), .B1(n22), .B2(regB_mem[1]), 
        .ZN(n29) );
  AND2_X1 U57 ( .A1(regB_mem[19]), .A2(n22), .ZN(DATA_MEM_IN[19]) );
  AND2_X1 U58 ( .A1(regB_mem[18]), .A2(n22), .ZN(DATA_MEM_IN[18]) );
  AND2_X1 U59 ( .A1(regB_mem[17]), .A2(n22), .ZN(DATA_MEM_IN[17]) );
  AND2_X1 U60 ( .A1(regB_mem[16]), .A2(n22), .ZN(DATA_MEM_IN[16]) );
  AND2_X1 U61 ( .A1(regB_mem[15]), .A2(n22), .ZN(DATA_MEM_IN[15]) );
  AND2_X1 U62 ( .A1(regB_mem[14]), .A2(n22), .ZN(DATA_MEM_IN[14]) );
  AND2_X1 U63 ( .A1(regB_mem[13]), .A2(n22), .ZN(DATA_MEM_IN[13]) );
  AND2_X1 U64 ( .A1(regB_mem[12]), .A2(n22), .ZN(DATA_MEM_IN[12]) );
  AND2_X1 U65 ( .A1(regB_mem[11]), .A2(n22), .ZN(DATA_MEM_IN[11]) );
  AND2_X1 U66 ( .A1(regB_mem[10]), .A2(n22), .ZN(DATA_MEM_IN[10]) );
  INV_X1 U67 ( .A(n30), .ZN(DATA_MEM_IN[0]) );
  AOI22_X1 U68 ( .A1(sb_op), .A2(regB_mem[24]), .B1(n22), .B2(regB_mem[0]), 
        .ZN(n30) );
  INV_X1 U69 ( .A(sb_op), .ZN(n22) );
  OR4_X1 U70 ( .A1(n31), .A2(n32), .A3(WM), .A4(RM), .ZN(DATA_MEM_ENABLE) );
  NOR4_X1 U71 ( .A1(instruction_alu[4]), .A2(n33), .A3(n34), .A4(n35), .ZN(n32) );
  INV_X1 U72 ( .A(instruction_alu[5]), .ZN(n35) );
  INV_X1 U73 ( .A(instruction_alu[3]), .ZN(n34) );
  AOI22_X1 U74 ( .A1(n36), .A2(instruction_alu[1]), .B1(instruction_alu[2]), 
        .B2(n37), .ZN(n33) );
  INV_X1 U75 ( .A(instruction_alu[1]), .ZN(n37) );
  NOR2_X1 U76 ( .A1(instruction_alu[2]), .A2(n38), .ZN(n36) );
  NOR4_X1 U77 ( .A1(n39), .A2(n38), .A3(instruction_alu[5]), .A4(
        instruction_alu[3]), .ZN(n31) );
  INV_X1 U78 ( .A(instruction_alu[0]), .ZN(n38) );
  NAND3_X1 U79 ( .A1(instruction_alu[2]), .A2(instruction_alu[1]), .A3(
        instruction_alu[4]), .ZN(n39) );
  regFFD_NBIT32_0 pipeline_PCING ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(PC), .Q(PC_fetch0) );
  regFFD_NBIT32_18 pipeline_fetch1_NPC ( .CK(CLK), .RESET(RST), .ENABLE(
        NPC_LATCH_EN), .D(NPC), .Q(NPC_fetch1) );
  regFFD_NBIT32_17 pipeline_fetch1_PC ( .CK(CLK), .RESET(RST), .ENABLE(
        ir_LATCH_EN), .D(PC_fetch0), .Q(PC_fetch1) );
  MUX21_GENERIC_NBIT32_0 MUX_PC1 ( .A(PC_OUT_i), .B(NPC_fetch1), .SEL(sel_npc), 
        .Y(PC_OUT) );
  regFFD_NBIT32_16 pipeline_fetch_NPC ( .CK(CLK), .RESET(RST), .ENABLE(
        NPC_LATCH_EN), .D(NPC_fetch1), .Q(NPC_fetch) );
  regFFD_NBIT32_15 pipeline_fetch_PC ( .CK(CLK), .RESET(RST), .ENABLE(
        ir_LATCH_EN), .D(PC_fetch1), .Q(PC_fetch) );
  regFFD_NBIT32_14 pipeline_fetch_ir ( .CK(CLK), .RESET(RST), .ENABLE(
        ir_LATCH_EN), .D(IR), .Q(ir_fetch) );
  regFFD_NBIT32_13 pipeline_newpc1 ( .CK(CLK), .RESET(RST), .ENABLE(
        NPC_LATCH_EN), .D(NPC_fetch), .Q(NPC_Dec) );
  regFFD_NBIT32_12 pipeline_pc1 ( .CK(CLK), .RESET(RST), .ENABLE(ir_LATCH_EN), 
        .D(PC_fetch) );
  regFFD_NBIT32_11 pipeline_IR1 ( .CK(CLK), .RESET(RST), .ENABLE(ir_LATCH_EN), 
        .D(ir_fetch), .Q(IR_Dec) );
  IR_DECODE_NBIT32_opBIT6_regBIT5 IR_OP ( .CLK(CLK), .IR_26(IR_Dec[25:0]), 
        .OPCODE(IR_Dec[31:26]), .is_signed(signed_op), .RS1(RS1), .RS2(RS2), 
        .RD(RD), .IMMEDIATE(Imm) );
  register_file RF ( .CLK(CLK), .RESET(RST), .ENABLE(1'b1), .RD1(RF1), .RD2(
        RF2), .WR(WF1), .ADD_WR(RD_wb), .ADD_RD1(RS1), .ADD_RD2(RS2), .DATAIN(
        OUT_data), .OUT1(regA), .OUT2(regB), .wr_signal(wr_signal_wb) );
  FF_0 pipeline_sign2 ( .CLK(CLK), .RESET(RST), .EN(1'b1), .D(signed_op), .Q(
        signed_op_ex) );
  regFFD_NBIT32_10 pipeline_newpc2 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(
        NPC_Dec), .Q(NPC_ex) );
  regFFD_NBIT32_9 pipeline_A2 ( .CK(CLK), .RESET(RST), .ENABLE(RF1), .D(regA), 
        .Q(regA_ex) );
  regFFD_NBIT32_8 pipeline_B2 ( .CK(CLK), .RESET(RST), .ENABLE(RF2), .D(regB), 
        .Q(regB_ex) );
  regFFD_NBIT32_7 pipeline_IMM2 ( .CK(CLK), .RESET(RST), .ENABLE(
        regImm_LATCH_EN), .D(Imm), .Q(Imm_ex) );
  regFFD_NBIT5_0 pipeline_RD2 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(RD), 
        .Q(RD_ex) );
  FF_7 pipeline_wr_signal ( .CLK(CLK), .RESET(RST), .EN(1'b1), .D(wr_signal), 
        .Q(wr_signal_exe) );
  regFFD_NBIT6_0 pipeline_IR2 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D({n42, 
        n44, n45, IR_Dec[28:27], n40}), .Q(IR_26_ex) );
  regFFD_NBIT32_6 pipeline_LHI2 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D({
        Imm[15:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Q(LHI_ex) );
  MUX21_GENERIC_NBIT32_6 MUX_ALU_A ( .A(NPC_ex), .B(regA_ex), .SEL(S1), .Y(
        input1_ALU) );
  MUX21_GENERIC_NBIT32_5 MUX_ALU_B ( .A(Imm_ex), .B(regB_ex), .SEL(S2), .Y(
        input2_ALU) );
  ALU_N32 ALU_OP ( .CLK(CLK), .FUNC({\instruction_alu[5] , 
        \instruction_alu[4] , \instruction_alu[3] , \instruction_alu[2] , 
        \instruction_alu[1] , \instruction_alu[0] }), .DATA1(input1_ALU), 
        .DATA2(input2_ALU), .OUT_ALU(ALU_out) );
  zero_eval_NBIT32 ZERO_OP ( .\input (regA_ex), .res(is_zero) );
  COND_BT_NBIT32 COND_OP ( .ZERO_BIT(is_zero), .OPCODE_0(IR_26_ex[0]), 
        .branch_op(branch_cond), .con_sign(cond) );
  MUX21_GENERIC_NBIT32_4 MUX_alu_out ( .A(LHI_ex), .B(ALU_out), .SEL(lhi_sel), 
        .Y(ALU_ex) );
  FF_6 pipeline_sign3 ( .CLK(CLK), .RESET(RST), .EN(1'b1), .D(signed_op_ex), 
        .Q(signed_op_mem) );
  regFFD_NBIT32_5 pipeline_newpc3 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(
        NPC_ex), .Q(NPC_mem) );
  FF_5 pipeline_cond3 ( .CLK(CLK), .RESET(RST), .EN(1'b1), .D(cond), .Q(
        cond_mem) );
  regFFD_NBIT32_4 pipeline_B3 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(
        regB_ex), .Q(regB_mem) );
  regFFD_NBIT5_2 pipeline_RD3 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(RD_ex), .Q(RD_mem) );
  FF_4 pipeline_wr_signal2 ( .CLK(CLK), .RESET(RST), .EN(1'b1), .D(
        wr_signal_exe), .Q(wr_signal_mem) );
  regFFD_NBIT6_1 pipeline_IR3 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(
        IR_26_ex), .Q(IR_26_mem) );
  MUX21_GENERIC_NBIT32_3 MUX_PC ( .A(ALU_ex), .B(NPC_mem), .SEL(sel_npc), .Y(
        PC_OUT_i) );
  load_data LOAD_DATA_OUT ( .data_in(DATA_MEM_OUT), .signed_val(signed_op_mem), 
        .load_op(RM), .load_type(IR_26_mem[1:0]), .data_out(LMD_out) );
  regFFD_NBIT32_3 pipeline_alu4 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(
        ALU_ex), .Q(ALU_wb) );
  regFFD_NBIT32_2 pipeline_LMD4 ( .CK(CLK), .RESET(RST), .ENABLE(RM), .D(
        LMD_out), .Q(LMD_wb) );
  regFFD_NBIT5_1 pipeline_RD4 ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(
        RD_mem), .Q(RD_wb) );
  FF_3 pipeline_wr_signal3 ( .CLK(CLK), .RESET(RST), .EN(1'b1), .D(
        wr_signal_mem1), .Q(wr_signal_wb) );
  FF_2 pipeline_WM ( .CLK(CLK), .RESET(RST), .EN(1'b1), .D(WM) );
  FF_1 pipeline_JAL ( .CLK(CLK), .RESET(RST), .EN(1'b1), .D(sel_saved_reg), 
        .Q(sel_saved_reg_wb) );
  regFFD_NBIT32_1 pipeline_NPC_wb ( .CK(CLK), .RESET(RST), .ENABLE(1'b1), .D(
        NPC_mem), .Q(NPC_wb) );
  MUX21_GENERIC_NBIT32_2 MUX_WB ( .A(ALU_wb), .B(LMD_wb), .SEL(S3), .Y(
        OUT_data) );
  MUX21_GENERIC_NBIT32_1 MUX_jal ( .A(NPC_wb), .B(OUT_data), .SEL(
        sel_saved_reg_wb) );
  DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 add_254 ( .A(PC_fetch0), .SUM(NPC) );
  CLKBUF_X1 U80 ( .A(IR_Dec[26]), .Z(n40) );
  CLKBUF_X1 U81 ( .A(IR_Dec[30]), .Z(n41) );
  CLKBUF_X1 U82 ( .A(IR_Dec[31]), .Z(n42) );
  INV_X1 U83 ( .A(n8), .ZN(n43) );
  INV_X1 U84 ( .A(n8), .ZN(n44) );
  CLKBUF_X1 U85 ( .A(IR_Dec[29]), .Z(n45) );
endmodule


module DLX_IR_SIZE32_PC_SIZE32 ( CLK, RST, IRAM_ADDRESS, IRAM_ISSUE, 
        IRAM_READY, IRAM_DATA, DRAM_ADDRESS, DRAM_ISSUE, DRAM_READNOTWRITE, 
        DRAM_READY, DRAM_DATA );
  output [31:0] IRAM_ADDRESS;
  input [63:0] IRAM_DATA;
  output [31:0] DRAM_ADDRESS;
  inout [63:0] DRAM_DATA;
  input CLK, RST, IRAM_READY, DRAM_READY;
  output IRAM_ISSUE, DRAM_ISSUE, DRAM_READNOTWRITE;
  wire   N9, signed_unsigned_i, lhi_sel_i, sb_op_i, DATA_MEM_WM_i;
  wire   [31:0] IR;
  wire   [31:0] PC;
  wire   [5:0] ALU_OPCODE_i;
  wire   [31:0] DATA_MEM_IN_i;
  wire   [31:0] dram_data_i;
  tri   [63:0] DRAM_DATA;
  assign IRAM_ADDRESS[31] = 1'b0;
  assign IRAM_ADDRESS[30] = 1'b0;
  assign IRAM_ADDRESS[29] = 1'b0;
  assign IRAM_ADDRESS[28] = 1'b0;
  assign IRAM_ADDRESS[27] = 1'b0;
  assign IRAM_ADDRESS[26] = 1'b0;
  assign IRAM_ADDRESS[25] = 1'b0;
  assign IRAM_ADDRESS[24] = 1'b0;
  assign IRAM_ADDRESS[23] = 1'b0;
  assign IRAM_ADDRESS[22] = 1'b0;
  assign IRAM_ADDRESS[21] = 1'b0;
  assign IRAM_ADDRESS[20] = 1'b0;
  assign IRAM_ADDRESS[19] = 1'b0;
  assign IRAM_ADDRESS[18] = 1'b0;
  assign IRAM_ADDRESS[17] = 1'b0;
  assign IRAM_ADDRESS[16] = 1'b0;
  assign IRAM_ADDRESS[15] = 1'b0;
  assign IRAM_ADDRESS[14] = 1'b0;
  assign IRAM_ADDRESS[13] = 1'b0;
  assign IRAM_ADDRESS[12] = 1'b0;
  assign IRAM_ADDRESS[11] = 1'b0;
  assign IRAM_ADDRESS[10] = 1'b0;
  assign IRAM_ADDRESS[9] = 1'b0;
  assign IRAM_ADDRESS[8] = 1'b0;
  assign IRAM_ADDRESS[7] = 1'b0;
  assign IRAM_ADDRESS[6] = 1'b0;
  assign IRAM_ADDRESS[5] = 1'b0;
  assign IRAM_ADDRESS[4] = 1'b0;
  assign IRAM_ADDRESS[3] = 1'b0;
  assign IRAM_ADDRESS[2] = 1'b0;
  assign IRAM_ADDRESS[1] = 1'b0;
  assign IRAM_ADDRESS[0] = 1'b0;

  DFF_X1 DRAM_READNOTWRITE_reg ( .D(N9), .CK(CLK), .Q(DRAM_READNOTWRITE) );
  TBUF_X2 \DRAM_DATA_tri[0]  ( .A(DATA_MEM_IN_i[0]), .EN(N9), .Z(DRAM_DATA[0])
         );
  TBUF_X2 \DRAM_DATA_tri[1]  ( .A(DATA_MEM_IN_i[1]), .EN(N9), .Z(DRAM_DATA[1])
         );
  TBUF_X2 \DRAM_DATA_tri[2]  ( .A(DATA_MEM_IN_i[2]), .EN(N9), .Z(DRAM_DATA[2])
         );
  TBUF_X2 \DRAM_DATA_tri[3]  ( .A(DATA_MEM_IN_i[3]), .EN(N9), .Z(DRAM_DATA[3])
         );
  TBUF_X2 \DRAM_DATA_tri[4]  ( .A(DATA_MEM_IN_i[4]), .EN(N9), .Z(DRAM_DATA[4])
         );
  TBUF_X2 \DRAM_DATA_tri[5]  ( .A(DATA_MEM_IN_i[5]), .EN(N9), .Z(DRAM_DATA[5])
         );
  TBUF_X2 \DRAM_DATA_tri[6]  ( .A(DATA_MEM_IN_i[6]), .EN(N9), .Z(DRAM_DATA[6])
         );
  TBUF_X2 \DRAM_DATA_tri[7]  ( .A(DATA_MEM_IN_i[7]), .EN(N9), .Z(DRAM_DATA[7])
         );
  TBUF_X2 \DRAM_DATA_tri[8]  ( .A(DATA_MEM_IN_i[8]), .EN(N9), .Z(DRAM_DATA[8])
         );
  TBUF_X2 \DRAM_DATA_tri[9]  ( .A(DATA_MEM_IN_i[9]), .EN(N9), .Z(DRAM_DATA[9])
         );
  TBUF_X2 \DRAM_DATA_tri[10]  ( .A(DATA_MEM_IN_i[10]), .EN(N9), .Z(
        DRAM_DATA[10]) );
  TBUF_X2 \DRAM_DATA_tri[11]  ( .A(DATA_MEM_IN_i[11]), .EN(N9), .Z(
        DRAM_DATA[11]) );
  TBUF_X2 \DRAM_DATA_tri[12]  ( .A(DATA_MEM_IN_i[12]), .EN(N9), .Z(
        DRAM_DATA[12]) );
  TBUF_X2 \DRAM_DATA_tri[13]  ( .A(DATA_MEM_IN_i[13]), .EN(N9), .Z(
        DRAM_DATA[13]) );
  TBUF_X2 \DRAM_DATA_tri[14]  ( .A(DATA_MEM_IN_i[14]), .EN(N9), .Z(
        DRAM_DATA[14]) );
  TBUF_X2 \DRAM_DATA_tri[15]  ( .A(DATA_MEM_IN_i[15]), .EN(N9), .Z(
        DRAM_DATA[15]) );
  TBUF_X2 \DRAM_DATA_tri[16]  ( .A(DATA_MEM_IN_i[16]), .EN(N9), .Z(
        DRAM_DATA[16]) );
  TBUF_X2 \DRAM_DATA_tri[17]  ( .A(DATA_MEM_IN_i[17]), .EN(N9), .Z(
        DRAM_DATA[17]) );
  TBUF_X2 \DRAM_DATA_tri[18]  ( .A(DATA_MEM_IN_i[18]), .EN(N9), .Z(
        DRAM_DATA[18]) );
  TBUF_X2 \DRAM_DATA_tri[19]  ( .A(DATA_MEM_IN_i[19]), .EN(N9), .Z(
        DRAM_DATA[19]) );
  TBUF_X2 \DRAM_DATA_tri[20]  ( .A(DATA_MEM_IN_i[20]), .EN(N9), .Z(
        DRAM_DATA[20]) );
  TBUF_X2 \DRAM_DATA_tri[21]  ( .A(DATA_MEM_IN_i[21]), .EN(N9), .Z(
        DRAM_DATA[21]) );
  TBUF_X2 \DRAM_DATA_tri[22]  ( .A(DATA_MEM_IN_i[22]), .EN(N9), .Z(
        DRAM_DATA[22]) );
  TBUF_X2 \DRAM_DATA_tri[23]  ( .A(DATA_MEM_IN_i[23]), .EN(N9), .Z(
        DRAM_DATA[23]) );
  TBUF_X2 \DRAM_DATA_tri[24]  ( .A(DATA_MEM_IN_i[24]), .EN(N9), .Z(
        DRAM_DATA[24]) );
  TBUF_X2 \DRAM_DATA_tri[25]  ( .A(DATA_MEM_IN_i[25]), .EN(N9), .Z(
        DRAM_DATA[25]) );
  TBUF_X2 \DRAM_DATA_tri[26]  ( .A(DATA_MEM_IN_i[26]), .EN(N9), .Z(
        DRAM_DATA[26]) );
  TBUF_X2 \DRAM_DATA_tri[27]  ( .A(DATA_MEM_IN_i[27]), .EN(N9), .Z(
        DRAM_DATA[27]) );
  TBUF_X2 \DRAM_DATA_tri[28]  ( .A(DATA_MEM_IN_i[28]), .EN(N9), .Z(
        DRAM_DATA[28]) );
  TBUF_X2 \DRAM_DATA_tri[29]  ( .A(DATA_MEM_IN_i[29]), .EN(N9), .Z(
        DRAM_DATA[29]) );
  TBUF_X2 \DRAM_DATA_tri[30]  ( .A(DATA_MEM_IN_i[30]), .EN(N9), .Z(
        DRAM_DATA[30]) );
  TBUF_X2 \DRAM_DATA_tri[31]  ( .A(DATA_MEM_IN_i[31]), .EN(N9), .Z(
        DRAM_DATA[31]) );
  TBUF_X2 \DRAM_DATA_tri[32]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[32]) );
  TBUF_X2 \DRAM_DATA_tri[33]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[33]) );
  TBUF_X2 \DRAM_DATA_tri[34]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[34]) );
  TBUF_X2 \DRAM_DATA_tri[35]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[35]) );
  TBUF_X2 \DRAM_DATA_tri[36]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[36]) );
  TBUF_X2 \DRAM_DATA_tri[37]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[37]) );
  TBUF_X2 \DRAM_DATA_tri[38]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[38]) );
  TBUF_X2 \DRAM_DATA_tri[39]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[39]) );
  TBUF_X2 \DRAM_DATA_tri[40]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[40]) );
  TBUF_X2 \DRAM_DATA_tri[41]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[41]) );
  TBUF_X2 \DRAM_DATA_tri[42]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[42]) );
  TBUF_X2 \DRAM_DATA_tri[43]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[43]) );
  TBUF_X2 \DRAM_DATA_tri[44]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[44]) );
  TBUF_X2 \DRAM_DATA_tri[45]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[45]) );
  TBUF_X2 \DRAM_DATA_tri[46]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[46]) );
  TBUF_X2 \DRAM_DATA_tri[47]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[47]) );
  TBUF_X2 \DRAM_DATA_tri[48]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[48]) );
  TBUF_X2 \DRAM_DATA_tri[49]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[49]) );
  TBUF_X2 \DRAM_DATA_tri[50]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[50]) );
  TBUF_X2 \DRAM_DATA_tri[51]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[51]) );
  TBUF_X2 \DRAM_DATA_tri[52]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[52]) );
  TBUF_X2 \DRAM_DATA_tri[53]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[53]) );
  TBUF_X2 \DRAM_DATA_tri[54]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[54]) );
  TBUF_X2 \DRAM_DATA_tri[55]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[55]) );
  TBUF_X2 \DRAM_DATA_tri[56]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[56]) );
  TBUF_X2 \DRAM_DATA_tri[57]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[57]) );
  TBUF_X2 \DRAM_DATA_tri[58]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[58]) );
  TBUF_X2 \DRAM_DATA_tri[59]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[59]) );
  TBUF_X2 \DRAM_DATA_tri[60]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[60]) );
  TBUF_X2 \DRAM_DATA_tri[61]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[61]) );
  TBUF_X2 \DRAM_DATA_tri[62]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[62]) );
  TBUF_X2 \DRAM_DATA_tri[63]  ( .A(1'b0), .EN(N9), .Z(DRAM_DATA[63]) );
  AND2_X1 U166 ( .A1(N9), .A2(DRAM_DATA[41]), .ZN(dram_data_i[9]) );
  AND2_X1 U167 ( .A1(DRAM_DATA[40]), .A2(N9), .ZN(dram_data_i[8]) );
  AND2_X1 U168 ( .A1(DRAM_DATA[39]), .A2(N9), .ZN(dram_data_i[7]) );
  AND2_X1 U169 ( .A1(DRAM_DATA[38]), .A2(N9), .ZN(dram_data_i[6]) );
  AND2_X1 U170 ( .A1(DRAM_DATA[37]), .A2(N9), .ZN(dram_data_i[5]) );
  AND2_X1 U171 ( .A1(DRAM_DATA[36]), .A2(N9), .ZN(dram_data_i[4]) );
  AND2_X1 U172 ( .A1(DRAM_DATA[35]), .A2(N9), .ZN(dram_data_i[3]) );
  AND2_X1 U173 ( .A1(DRAM_DATA[63]), .A2(N9), .ZN(dram_data_i[31]) );
  AND2_X1 U174 ( .A1(DRAM_DATA[62]), .A2(N9), .ZN(dram_data_i[30]) );
  AND2_X1 U175 ( .A1(DRAM_DATA[34]), .A2(N9), .ZN(dram_data_i[2]) );
  AND2_X1 U176 ( .A1(DRAM_DATA[61]), .A2(N9), .ZN(dram_data_i[29]) );
  AND2_X1 U177 ( .A1(DRAM_DATA[60]), .A2(N9), .ZN(dram_data_i[28]) );
  AND2_X1 U178 ( .A1(DRAM_DATA[59]), .A2(N9), .ZN(dram_data_i[27]) );
  AND2_X1 U179 ( .A1(DRAM_DATA[58]), .A2(N9), .ZN(dram_data_i[26]) );
  AND2_X1 U180 ( .A1(DRAM_DATA[57]), .A2(N9), .ZN(dram_data_i[25]) );
  AND2_X1 U181 ( .A1(DRAM_DATA[56]), .A2(N9), .ZN(dram_data_i[24]) );
  AND2_X1 U182 ( .A1(DRAM_DATA[55]), .A2(N9), .ZN(dram_data_i[23]) );
  AND2_X1 U183 ( .A1(DRAM_DATA[54]), .A2(N9), .ZN(dram_data_i[22]) );
  AND2_X1 U184 ( .A1(DRAM_DATA[53]), .A2(N9), .ZN(dram_data_i[21]) );
  AND2_X1 U185 ( .A1(DRAM_DATA[52]), .A2(N9), .ZN(dram_data_i[20]) );
  AND2_X1 U186 ( .A1(DRAM_DATA[33]), .A2(N9), .ZN(dram_data_i[1]) );
  AND2_X1 U187 ( .A1(DRAM_DATA[51]), .A2(N9), .ZN(dram_data_i[19]) );
  AND2_X1 U188 ( .A1(DRAM_DATA[50]), .A2(N9), .ZN(dram_data_i[18]) );
  AND2_X1 U189 ( .A1(DRAM_DATA[49]), .A2(N9), .ZN(dram_data_i[17]) );
  AND2_X1 U190 ( .A1(DRAM_DATA[48]), .A2(N9), .ZN(dram_data_i[16]) );
  AND2_X1 U191 ( .A1(DRAM_DATA[47]), .A2(N9), .ZN(dram_data_i[15]) );
  AND2_X1 U192 ( .A1(DRAM_DATA[46]), .A2(N9), .ZN(dram_data_i[14]) );
  AND2_X1 U193 ( .A1(DRAM_DATA[45]), .A2(N9), .ZN(dram_data_i[13]) );
  AND2_X1 U194 ( .A1(DRAM_DATA[44]), .A2(N9), .ZN(dram_data_i[12]) );
  AND2_X1 U195 ( .A1(DRAM_DATA[43]), .A2(N9), .ZN(dram_data_i[11]) );
  AND2_X1 U196 ( .A1(DRAM_DATA[42]), .A2(N9), .ZN(dram_data_i[10]) );
  AND2_X1 U197 ( .A1(DRAM_DATA[32]), .A2(N9), .ZN(dram_data_i[0]) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 CU_I ( 
        .Clk(CLK), .Rst(RST), .IR_IN({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .ALU_OPCODE(ALU_OPCODE_i), .signed_unsigned(signed_unsigned_i), 
        .lhi_sel(lhi_sel_i), .sb_op(sb_op_i) );
  DATAPTH_NBIT32_REG_BIT5 DTPTH_I ( .CLK(CLK), .RST(RST), .PC({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IR({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .NPC_LATCH_EN(1'b0), .ir_LATCH_EN(1'b0), 
        .signed_op(signed_unsigned_i), .RF1(1'b0), .RF2(1'b0), .WF1(1'b0), 
        .regImm_LATCH_EN(1'b0), .S1(1'b0), .S2(1'b0), .EN2(1'b0), .lhi_sel(
        lhi_sel_i), .jump_en(1'b0), .branch_cond(1'b0), .sb_op(sb_op_i), .RM(
        1'b0), .WM(1'b0), .EN3(1'b0), .S3(1'b0), .instruction_alu(ALU_OPCODE_i), .DATA_MEM_ADDR(DRAM_ADDRESS), .DATA_MEM_IN(DATA_MEM_IN_i), .DATA_MEM_OUT(
        dram_data_i), .DATA_MEM_ENABLE(DRAM_ISSUE), .DATA_MEM_WM(DATA_MEM_WM_i) );
  INV_X8 U198 ( .A(DATA_MEM_WM_i), .ZN(N9) );
endmodule




    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_3 ( 
        A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106;

  CLKBUF_X1 U2 ( .A(A[7]), .Z(n1) );
  NAND2_X1 U3 ( .A1(A[7]), .A2(A[6]), .ZN(n2) );
  AND2_X1 U4 ( .A1(n69), .A2(n37), .ZN(n28) );
  AND2_X1 U5 ( .A1(n69), .A2(n6), .ZN(n57) );
  BUF_X1 U6 ( .A(A[1]), .Z(n8) );
  AND2_X1 U7 ( .A1(A[12]), .A2(n21), .ZN(n3) );
  AND2_X1 U8 ( .A1(A[20]), .A2(A[21]), .ZN(n4) );
  AND2_X1 U9 ( .A1(A[24]), .A2(A[25]), .ZN(n5) );
  NOR2_X1 U10 ( .A1(n85), .A2(n86), .ZN(n6) );
  XOR2_X1 U11 ( .A(A[22]), .B(n7), .Z(SUM[22]) );
  AND2_X1 U12 ( .A1(n88), .A2(n4), .ZN(n7) );
  NOR2_X1 U13 ( .A1(n65), .A2(n2), .ZN(n9) );
  CLKBUF_X1 U14 ( .A(A[0]), .Z(n10) );
  INV_X1 U15 ( .A(n87), .ZN(n11) );
  CLKBUF_X1 U16 ( .A(A[11]), .Z(n12) );
  INV_X1 U17 ( .A(n74), .ZN(n13) );
  CLKBUF_X1 U18 ( .A(n92), .Z(n14) );
  CLKBUF_X1 U19 ( .A(A[9]), .Z(n15) );
  CLKBUF_X1 U20 ( .A(A[10]), .Z(n16) );
  XNOR2_X1 U21 ( .A(n81), .B(n17), .ZN(SUM[28]) );
  NOR2_X1 U22 ( .A1(n27), .A2(n59), .ZN(n17) );
  INV_X1 U23 ( .A(A[28]), .ZN(n81) );
  XOR2_X1 U24 ( .A(A[21]), .B(n18), .Z(SUM[21]) );
  AND2_X1 U25 ( .A1(n88), .A2(A[20]), .ZN(n18) );
  XOR2_X1 U26 ( .A(A[25]), .B(n19), .Z(SUM[25]) );
  AND2_X1 U27 ( .A1(A[24]), .A2(n44), .ZN(n19) );
  CLKBUF_X1 U28 ( .A(A[15]), .Z(n20) );
  CLKBUF_X1 U29 ( .A(A[13]), .Z(n21) );
  AND2_X1 U30 ( .A1(n53), .A2(n3), .ZN(n22) );
  XOR2_X1 U31 ( .A(n1), .B(n23), .Z(SUM[7]) );
  AND2_X1 U32 ( .A1(n70), .A2(n45), .ZN(n23) );
  BUF_X1 U33 ( .A(A[3]), .Z(n34) );
  XOR2_X1 U34 ( .A(A[26]), .B(n24), .Z(SUM[26]) );
  AND2_X1 U35 ( .A1(n44), .A2(n5), .ZN(n24) );
  CLKBUF_X1 U36 ( .A(A[8]), .Z(n25) );
  BUF_X1 U37 ( .A(A[2]), .Z(n40) );
  NAND4_X1 U38 ( .A1(A[15]), .A2(A[13]), .A3(A[12]), .A4(A[14]), .ZN(n26) );
  INV_X1 U39 ( .A(n28), .ZN(n93) );
  NAND2_X1 U40 ( .A1(n57), .A2(n56), .ZN(n27) );
  AND2_X1 U41 ( .A1(n5), .A2(A[26]), .ZN(n29) );
  XOR2_X1 U42 ( .A(A[27]), .B(n30), .Z(SUM[27]) );
  AND2_X1 U43 ( .A1(n44), .A2(n29), .ZN(n30) );
  NAND4_X1 U44 ( .A1(A[9]), .A2(A[10]), .A3(A[11]), .A4(A[8]), .ZN(n31) );
  NOR2_X1 U45 ( .A1(n27), .A2(n32), .ZN(n78) );
  OR2_X1 U46 ( .A1(n59), .A2(n79), .ZN(n32) );
  CLKBUF_X1 U47 ( .A(n10), .Z(n33) );
  AND2_X1 U48 ( .A1(n35), .A2(n36), .ZN(n80) );
  NOR2_X1 U49 ( .A1(n84), .A2(n59), .ZN(n35) );
  AND2_X1 U50 ( .A1(A[28]), .A2(A[29]), .ZN(n36) );
  AND2_X1 U51 ( .A1(n102), .A2(n103), .ZN(n69) );
  NOR2_X1 U52 ( .A1(n31), .A2(n26), .ZN(n37) );
  OR2_X1 U53 ( .A1(n81), .A2(n59), .ZN(n38) );
  XOR2_X1 U54 ( .A(A[19]), .B(n39), .Z(SUM[19]) );
  AND2_X1 U55 ( .A1(n91), .A2(A[18]), .ZN(n39) );
  CLKBUF_X1 U56 ( .A(A[5]), .Z(n41) );
  NAND2_X1 U57 ( .A1(A[3]), .A2(A[2]), .ZN(n42) );
  NAND2_X1 U58 ( .A1(n53), .A2(n3), .ZN(n97) );
  XOR2_X1 U59 ( .A(A[17]), .B(n43), .Z(SUM[17]) );
  AND2_X1 U60 ( .A1(n28), .A2(A[16]), .ZN(n43) );
  AND2_X1 U61 ( .A1(n57), .A2(n56), .ZN(n44) );
  CLKBUF_X1 U62 ( .A(A[6]), .Z(n45) );
  AND2_X1 U63 ( .A1(n11), .A2(n4), .ZN(n46) );
  CLKBUF_X1 U64 ( .A(A[14]), .Z(n47) );
  CLKBUF_X1 U65 ( .A(A[4]), .Z(n48) );
  CLKBUF_X1 U66 ( .A(A[12]), .Z(n49) );
  CLKBUF_X1 U67 ( .A(n67), .Z(n50) );
  INV_X1 U68 ( .A(n53), .ZN(n99) );
  AND2_X1 U69 ( .A1(n9), .A2(n68), .ZN(n67) );
  CLKBUF_X1 U70 ( .A(n104), .Z(n51) );
  CLKBUF_X1 U71 ( .A(n25), .Z(n52) );
  AND2_X2 U72 ( .A1(n67), .A2(n55), .ZN(n53) );
  NOR2_X1 U73 ( .A1(n89), .A2(n90), .ZN(n54) );
  AND4_X1 U74 ( .A1(n12), .A2(A[10]), .A3(A[9]), .A4(n25), .ZN(n55) );
  AND2_X1 U75 ( .A1(n54), .A2(n37), .ZN(n56) );
  NAND2_X1 U76 ( .A1(n57), .A2(n56), .ZN(n84) );
  NAND2_X1 U77 ( .A1(n69), .A2(n58), .ZN(n87) );
  AND2_X1 U78 ( .A1(n94), .A2(n54), .ZN(n58) );
  OR2_X1 U79 ( .A1(n82), .A2(n83), .ZN(n59) );
  XOR2_X1 U80 ( .A(n20), .B(n60), .Z(SUM[15]) );
  AND2_X1 U81 ( .A1(n47), .A2(n22), .ZN(n60) );
  XOR2_X1 U82 ( .A(n78), .B(A[31]), .Z(SUM[31]) );
  XOR2_X1 U83 ( .A(n61), .B(A[23]), .Z(SUM[23]) );
  AND2_X1 U84 ( .A1(n46), .A2(A[22]), .ZN(n61) );
  XNOR2_X1 U85 ( .A(n47), .B(n97), .ZN(SUM[14]) );
  XNOR2_X1 U86 ( .A(n14), .B(A[18]), .ZN(SUM[18]) );
  XNOR2_X1 U87 ( .A(n16), .B(n101), .ZN(SUM[10]) );
  XNOR2_X1 U88 ( .A(n62), .B(A[29]), .ZN(SUM[29]) );
  OR2_X1 U89 ( .A1(n38), .A2(n27), .ZN(n62) );
  XOR2_X1 U90 ( .A(n80), .B(A[30]), .Z(SUM[30]) );
  XNOR2_X1 U91 ( .A(n49), .B(n99), .ZN(SUM[12]) );
  XOR2_X1 U92 ( .A(n15), .B(n63), .Z(SUM[9]) );
  AND2_X1 U93 ( .A1(n52), .A2(n50), .ZN(n63) );
  XOR2_X1 U94 ( .A(n12), .B(n64), .Z(SUM[11]) );
  AND2_X1 U95 ( .A1(n100), .A2(n16), .ZN(n64) );
  OR2_X1 U96 ( .A1(n65), .A2(n72), .ZN(n71) );
  NAND2_X1 U97 ( .A1(A[5]), .A2(A[4]), .ZN(n65) );
  XNOR2_X1 U98 ( .A(n41), .B(n73), .ZN(SUM[5]) );
  INV_X1 U99 ( .A(n72), .ZN(n74) );
  XOR2_X1 U100 ( .A(n52), .B(n50), .Z(SUM[8]) );
  INV_X1 U101 ( .A(n51), .ZN(n76) );
  XNOR2_X1 U102 ( .A(A[24]), .B(n84), .ZN(SUM[24]) );
  XNOR2_X1 U103 ( .A(A[16]), .B(n93), .ZN(SUM[16]) );
  XNOR2_X1 U104 ( .A(n34), .B(n75), .ZN(SUM[3]) );
  CLKBUF_X1 U105 ( .A(n40), .Z(n66) );
  NOR2_X1 U106 ( .A1(n95), .A2(n96), .ZN(n94) );
  NAND4_X1 U107 ( .A1(A[9]), .A2(A[10]), .A3(A[11]), .A4(A[8]), .ZN(n95) );
  NOR2_X1 U108 ( .A1(n104), .A2(n42), .ZN(n68) );
  XNOR2_X1 U109 ( .A(n45), .B(n71), .ZN(SUM[6]) );
  NOR2_X1 U110 ( .A1(n65), .A2(n106), .ZN(n102) );
  NAND2_X1 U111 ( .A1(n48), .A2(n74), .ZN(n73) );
  NOR2_X1 U112 ( .A1(n77), .A2(n105), .ZN(n103) );
  XNOR2_X1 U113 ( .A(n87), .B(A[20]), .ZN(SUM[20]) );
  INV_X1 U114 ( .A(n87), .ZN(n88) );
  XNOR2_X1 U115 ( .A(n66), .B(n51), .ZN(SUM[2]) );
  NAND2_X1 U116 ( .A1(n66), .A2(n76), .ZN(n75) );
  INV_X1 U117 ( .A(n33), .ZN(SUM[0]) );
  NAND2_X1 U118 ( .A1(A[1]), .A2(A[0]), .ZN(n77) );
  NAND4_X1 U119 ( .A1(n10), .A2(n40), .A3(n8), .A4(n34), .ZN(n72) );
  INV_X1 U120 ( .A(n71), .ZN(n70) );
  XNOR2_X1 U121 ( .A(n13), .B(n48), .ZN(SUM[4]) );
  NAND3_X1 U122 ( .A1(A[30]), .A2(A[29]), .A3(A[28]), .ZN(n79) );
  NAND2_X1 U123 ( .A1(A[24]), .A2(A[25]), .ZN(n83) );
  NAND2_X1 U124 ( .A1(A[27]), .A2(A[26]), .ZN(n82) );
  NAND2_X1 U125 ( .A1(A[20]), .A2(A[21]), .ZN(n86) );
  NAND2_X1 U126 ( .A1(A[23]), .A2(A[22]), .ZN(n85) );
  NAND2_X1 U127 ( .A1(A[16]), .A2(A[17]), .ZN(n90) );
  NAND2_X1 U128 ( .A1(A[19]), .A2(A[18]), .ZN(n89) );
  XOR2_X1 U129 ( .A(n8), .B(n33), .Z(SUM[1]) );
  INV_X1 U130 ( .A(n92), .ZN(n91) );
  NAND3_X1 U131 ( .A1(n28), .A2(A[17]), .A3(A[16]), .ZN(n92) );
  NAND4_X1 U132 ( .A1(A[12]), .A2(A[14]), .A3(A[13]), .A4(A[15]), .ZN(n96) );
  XNOR2_X1 U133 ( .A(n21), .B(n98), .ZN(SUM[13]) );
  NAND2_X1 U134 ( .A1(n53), .A2(n49), .ZN(n98) );
  INV_X1 U135 ( .A(n101), .ZN(n100) );
  NAND3_X1 U136 ( .A1(n67), .A2(n15), .A3(n25), .ZN(n101) );
  NAND2_X1 U137 ( .A1(A[3]), .A2(A[2]), .ZN(n105) );
  NAND2_X1 U138 ( .A1(A[1]), .A2(A[0]), .ZN(n104) );
  NAND2_X1 U139 ( .A1(A[7]), .A2(A[6]), .ZN(n106) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 ( 
        A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75;

  AND2_X1 U2 ( .A1(A[20]), .A2(A[21]), .ZN(n1) );
  BUF_X1 U3 ( .A(n14), .Z(n2) );
  NAND2_X1 U4 ( .A1(n3), .A2(n4), .ZN(n41) );
  AND2_X1 U5 ( .A1(n25), .A2(n26), .ZN(n3) );
  NOR2_X1 U6 ( .A1(n46), .A2(n47), .ZN(n4) );
  XOR2_X1 U7 ( .A(A[25]), .B(n5), .Z(SUM[25]) );
  AND2_X1 U8 ( .A1(A[24]), .A2(n3), .ZN(n5) );
  CLKBUF_X1 U9 ( .A(A[2]), .Z(n6) );
  INV_X1 U10 ( .A(n2), .ZN(n68) );
  INV_X1 U11 ( .A(n63), .ZN(n7) );
  AND2_X1 U12 ( .A1(n30), .A2(n8), .ZN(n25) );
  NOR2_X1 U13 ( .A1(n19), .A2(n7), .ZN(n8) );
  INV_X1 U14 ( .A(n30), .ZN(n9) );
  CLKBUF_X1 U15 ( .A(A[5]), .Z(n10) );
  NOR2_X1 U16 ( .A1(n31), .A2(n19), .ZN(n14) );
  AND2_X1 U17 ( .A1(n25), .A2(n26), .ZN(n11) );
  XOR2_X1 U18 ( .A(A[15]), .B(n12), .Z(SUM[15]) );
  AND2_X1 U19 ( .A1(n66), .A2(A[14]), .ZN(n12) );
  INV_X1 U20 ( .A(SUM[0]), .ZN(n13) );
  NOR2_X1 U21 ( .A1(n31), .A2(n19), .ZN(n15) );
  CLKBUF_X1 U22 ( .A(A[4]), .Z(n16) );
  AND2_X1 U23 ( .A1(n55), .A2(n1), .ZN(n51) );
  AND4_X1 U24 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(n17) );
  AND4_X1 U25 ( .A1(A[1]), .A2(A[2]), .A3(A[3]), .A4(A[0]), .ZN(n28) );
  NAND2_X1 U26 ( .A1(n25), .A2(n26), .ZN(n18) );
  NOR2_X1 U27 ( .A1(n49), .A2(n50), .ZN(n48) );
  XOR2_X1 U28 ( .A(n23), .B(A[18]), .Z(SUM[18]) );
  XOR2_X1 U29 ( .A(n22), .B(A[10]), .Z(SUM[10]) );
  OR2_X1 U30 ( .A1(n70), .A2(n71), .ZN(n19) );
  NOR2_X1 U31 ( .A1(n74), .A2(n75), .ZN(n73) );
  XNOR2_X1 U32 ( .A(A[14]), .B(n67), .ZN(SUM[14]) );
  XNOR2_X1 U33 ( .A(n18), .B(A[24]), .ZN(SUM[24]) );
  XNOR2_X1 U34 ( .A(n6), .B(n38), .ZN(SUM[2]) );
  XNOR2_X1 U35 ( .A(A[17]), .B(n61), .ZN(SUM[17]) );
  XNOR2_X1 U36 ( .A(A[21]), .B(n54), .ZN(SUM[21]) );
  NAND2_X1 U37 ( .A1(A[20]), .A2(n55), .ZN(n54) );
  XNOR2_X1 U38 ( .A(A[13]), .B(n69), .ZN(SUM[13]) );
  NAND2_X1 U39 ( .A1(A[12]), .A2(n2), .ZN(n69) );
  XNOR2_X1 U40 ( .A(n10), .B(n35), .ZN(SUM[5]) );
  XNOR2_X1 U41 ( .A(n20), .B(A[26]), .ZN(SUM[26]) );
  NAND3_X1 U42 ( .A1(A[24]), .A2(A[25]), .A3(n11), .ZN(n20) );
  XOR2_X1 U43 ( .A(n44), .B(A[29]), .Z(SUM[29]) );
  NOR2_X1 U44 ( .A1(n64), .A2(n65), .ZN(n63) );
  XOR2_X1 U45 ( .A(A[27]), .B(n21), .Z(SUM[27]) );
  AND2_X1 U46 ( .A1(n27), .A2(A[26]), .ZN(n21) );
  XNOR2_X1 U47 ( .A(A[6]), .B(n34), .ZN(SUM[6]) );
  XOR2_X1 U48 ( .A(n16), .B(n17), .Z(SUM[4]) );
  XOR2_X1 U49 ( .A(n42), .B(A[30]), .Z(SUM[30]) );
  XOR2_X1 U50 ( .A(n39), .B(A[31]), .Z(SUM[31]) );
  XNOR2_X1 U51 ( .A(A[9]), .B(n29), .ZN(SUM[9]) );
  NAND2_X1 U52 ( .A1(A[8]), .A2(n30), .ZN(n29) );
  XNOR2_X1 U53 ( .A(A[3]), .B(n36), .ZN(SUM[3]) );
  NAND2_X1 U54 ( .A1(n6), .A2(n37), .ZN(n36) );
  INV_X1 U55 ( .A(n38), .ZN(n37) );
  AND3_X1 U56 ( .A1(A[8]), .A2(A[9]), .A3(n30), .ZN(n22) );
  AND3_X1 U57 ( .A1(A[16]), .A2(A[17]), .A3(n62), .ZN(n23) );
  INV_X1 U58 ( .A(A[28]), .ZN(n45) );
  NAND2_X1 U59 ( .A1(A[16]), .A2(n62), .ZN(n61) );
  NAND2_X1 U60 ( .A1(n62), .A2(n56), .ZN(n53) );
  XNOR2_X1 U61 ( .A(A[22]), .B(n52), .ZN(SUM[22]) );
  XOR2_X1 U62 ( .A(A[23]), .B(n24), .Z(SUM[23]) );
  AND2_X1 U63 ( .A1(n51), .A2(A[22]), .ZN(n24) );
  AND2_X1 U64 ( .A1(n48), .A2(n56), .ZN(n26) );
  XNOR2_X1 U65 ( .A(A[28]), .B(n41), .ZN(SUM[28]) );
  NOR2_X1 U66 ( .A1(n41), .A2(n45), .ZN(n44) );
  NOR2_X1 U67 ( .A1(n41), .A2(n43), .ZN(n42) );
  NOR2_X1 U68 ( .A1(n40), .A2(n41), .ZN(n39) );
  NAND2_X1 U69 ( .A1(n15), .A2(n63), .ZN(n60) );
  AND3_X1 U70 ( .A1(A[24]), .A2(A[25]), .A3(n11), .ZN(n27) );
  NOR2_X1 U71 ( .A1(n57), .A2(n58), .ZN(n56) );
  XNOR2_X1 U72 ( .A(n60), .B(A[16]), .ZN(SUM[16]) );
  XNOR2_X1 U73 ( .A(A[12]), .B(n68), .ZN(SUM[12]) );
  INV_X1 U74 ( .A(n60), .ZN(n62) );
  XNOR2_X1 U75 ( .A(A[20]), .B(n53), .ZN(SUM[20]) );
  XNOR2_X1 U76 ( .A(A[8]), .B(n9), .ZN(SUM[8]) );
  INV_X1 U77 ( .A(n53), .ZN(n55) );
  INV_X1 U78 ( .A(n31), .ZN(n30) );
  NAND2_X1 U79 ( .A1(n16), .A2(n17), .ZN(n35) );
  NAND2_X1 U80 ( .A1(n73), .A2(n28), .ZN(n31) );
  INV_X1 U81 ( .A(A[0]), .ZN(SUM[0]) );
  NAND2_X1 U82 ( .A1(A[1]), .A2(n13), .ZN(n38) );
  XNOR2_X1 U83 ( .A(A[7]), .B(n32), .ZN(SUM[7]) );
  NAND2_X1 U84 ( .A1(n33), .A2(A[6]), .ZN(n32) );
  INV_X1 U85 ( .A(n34), .ZN(n33) );
  NAND3_X1 U86 ( .A1(A[4]), .A2(n10), .A3(n17), .ZN(n34) );
  NAND3_X1 U87 ( .A1(A[30]), .A2(A[29]), .A3(A[28]), .ZN(n40) );
  NAND2_X1 U88 ( .A1(A[28]), .A2(A[29]), .ZN(n43) );
  NAND2_X1 U89 ( .A1(A[24]), .A2(A[25]), .ZN(n47) );
  NAND2_X1 U90 ( .A1(A[27]), .A2(A[26]), .ZN(n46) );
  NAND2_X1 U91 ( .A1(A[20]), .A2(A[21]), .ZN(n50) );
  NAND2_X1 U92 ( .A1(A[23]), .A2(A[22]), .ZN(n49) );
  NAND3_X1 U93 ( .A1(A[20]), .A2(A[21]), .A3(n55), .ZN(n52) );
  NAND2_X1 U94 ( .A1(A[16]), .A2(A[17]), .ZN(n58) );
  NAND2_X1 U95 ( .A1(A[19]), .A2(A[18]), .ZN(n57) );
  XOR2_X1 U96 ( .A(A[1]), .B(n13), .Z(SUM[1]) );
  XNOR2_X1 U97 ( .A(A[19]), .B(n59), .ZN(SUM[19]) );
  NAND2_X1 U98 ( .A1(n23), .A2(A[18]), .ZN(n59) );
  NAND2_X1 U99 ( .A1(A[12]), .A2(A[13]), .ZN(n65) );
  NAND2_X1 U100 ( .A1(A[15]), .A2(A[14]), .ZN(n64) );
  INV_X1 U101 ( .A(n67), .ZN(n66) );
  NAND3_X1 U102 ( .A1(A[12]), .A2(A[13]), .A3(n14), .ZN(n67) );
  NAND2_X1 U103 ( .A1(A[8]), .A2(A[9]), .ZN(n71) );
  NAND2_X1 U104 ( .A1(A[11]), .A2(A[10]), .ZN(n70) );
  XNOR2_X1 U105 ( .A(A[11]), .B(n72), .ZN(SUM[11]) );
  NAND2_X1 U106 ( .A1(n22), .A2(A[10]), .ZN(n72) );
  NAND2_X1 U107 ( .A1(A[4]), .A2(A[5]), .ZN(n75) );
  NAND2_X1 U108 ( .A1(A[7]), .A2(A[6]), .ZN(n74) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 ( 
        A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;

  AND3_X1 U2 ( .A1(A[24]), .A2(A[25]), .A3(n9), .ZN(n1) );
  OR2_X1 U3 ( .A1(n43), .A2(n44), .ZN(n2) );
  NOR2_X1 U4 ( .A1(n52), .A2(n8), .ZN(n7) );
  NAND2_X1 U5 ( .A1(n3), .A2(n4), .ZN(n40) );
  AND2_X1 U6 ( .A1(n54), .A2(n55), .ZN(n3) );
  NOR2_X1 U7 ( .A1(n2), .A2(n8), .ZN(n4) );
  NOR2_X1 U8 ( .A1(n40), .A2(n10), .ZN(n9) );
  NOR2_X1 U9 ( .A1(n31), .A2(n32), .ZN(n30) );
  NOR2_X1 U10 ( .A1(n56), .A2(n57), .ZN(n55) );
  NAND2_X1 U11 ( .A1(n17), .A2(n59), .ZN(n13) );
  NOR2_X1 U12 ( .A1(n60), .A2(n61), .ZN(n59) );
  XNOR2_X1 U13 ( .A(A[6]), .B(n16), .ZN(SUM[6]) );
  XNOR2_X1 U14 ( .A(A[14]), .B(n51), .ZN(SUM[14]) );
  XNOR2_X1 U15 ( .A(A[22]), .B(n39), .ZN(SUM[22]) );
  XOR2_X1 U16 ( .A(n6), .B(A[10]), .Z(SUM[10]) );
  XOR2_X1 U17 ( .A(n26), .B(A[30]), .Z(SUM[30]) );
  XOR2_X1 U18 ( .A(n5), .B(A[18]), .Z(SUM[18]) );
  XOR2_X1 U19 ( .A(n1), .B(A[26]), .Z(SUM[26]) );
  XOR2_X1 U20 ( .A(A[16]), .B(n7), .Z(SUM[16]) );
  INV_X1 U21 ( .A(n22), .ZN(n21) );
  XOR2_X1 U22 ( .A(n23), .B(A[31]), .Z(SUM[31]) );
  XOR2_X1 U23 ( .A(n28), .B(A[29]), .Z(SUM[29]) );
  XNOR2_X1 U24 ( .A(A[5]), .B(n18), .ZN(SUM[5]) );
  NAND2_X1 U25 ( .A1(A[4]), .A2(n17), .ZN(n18) );
  XNOR2_X1 U26 ( .A(A[9]), .B(n12), .ZN(SUM[9]) );
  NAND2_X1 U27 ( .A1(A[8]), .A2(n54), .ZN(n12) );
  XNOR2_X1 U28 ( .A(A[13]), .B(n53), .ZN(SUM[13]) );
  NAND2_X1 U29 ( .A1(A[12]), .A2(n3), .ZN(n53) );
  XNOR2_X1 U30 ( .A(A[17]), .B(n46), .ZN(SUM[17]) );
  NAND2_X1 U31 ( .A1(A[16]), .A2(n7), .ZN(n46) );
  XNOR2_X1 U32 ( .A(A[21]), .B(n41), .ZN(SUM[21]) );
  NAND2_X1 U33 ( .A1(A[20]), .A2(n42), .ZN(n41) );
  XNOR2_X1 U34 ( .A(A[25]), .B(n34), .ZN(SUM[25]) );
  AND3_X1 U35 ( .A1(A[16]), .A2(A[17]), .A3(n7), .ZN(n5) );
  AND3_X1 U36 ( .A1(A[8]), .A2(A[9]), .A3(n54), .ZN(n6) );
  INV_X1 U37 ( .A(A[28]), .ZN(n29) );
  OR2_X1 U38 ( .A1(n47), .A2(n48), .ZN(n8) );
  NAND2_X1 U39 ( .A1(n54), .A2(n55), .ZN(n52) );
  XNOR2_X1 U40 ( .A(A[3]), .B(n20), .ZN(SUM[3]) );
  NAND2_X1 U41 ( .A1(A[24]), .A2(n9), .ZN(n34) );
  INV_X1 U42 ( .A(n9), .ZN(n33) );
  OR2_X1 U43 ( .A1(n35), .A2(n36), .ZN(n10) );
  XNOR2_X1 U44 ( .A(A[20]), .B(n40), .ZN(SUM[20]) );
  INV_X1 U45 ( .A(n40), .ZN(n42) );
  XNOR2_X1 U46 ( .A(A[12]), .B(n52), .ZN(SUM[12]) );
  XOR2_X1 U47 ( .A(A[27]), .B(n11), .Z(SUM[27]) );
  AND2_X1 U48 ( .A1(n1), .A2(A[26]), .ZN(n11) );
  XNOR2_X1 U49 ( .A(A[8]), .B(n13), .ZN(SUM[8]) );
  XNOR2_X1 U50 ( .A(A[24]), .B(n33), .ZN(SUM[24]) );
  NAND2_X1 U51 ( .A1(n9), .A2(n30), .ZN(n25) );
  XNOR2_X1 U52 ( .A(A[2]), .B(n22), .ZN(SUM[2]) );
  XNOR2_X1 U53 ( .A(A[28]), .B(n25), .ZN(SUM[28]) );
  NAND2_X1 U54 ( .A1(A[2]), .A2(n21), .ZN(n20) );
  NOR2_X1 U55 ( .A1(n25), .A2(n29), .ZN(n28) );
  NOR2_X1 U56 ( .A1(n25), .A2(n27), .ZN(n26) );
  NOR2_X1 U57 ( .A1(n24), .A2(n25), .ZN(n23) );
  INV_X1 U58 ( .A(A[0]), .ZN(SUM[0]) );
  NAND2_X1 U59 ( .A1(A[1]), .A2(A[0]), .ZN(n22) );
  NAND4_X1 U60 ( .A1(A[0]), .A2(A[2]), .A3(A[1]), .A4(A[3]), .ZN(n19) );
  XNOR2_X1 U61 ( .A(A[7]), .B(n14), .ZN(SUM[7]) );
  NAND2_X1 U62 ( .A1(n15), .A2(A[6]), .ZN(n14) );
  INV_X1 U63 ( .A(n16), .ZN(n15) );
  NAND3_X1 U64 ( .A1(A[4]), .A2(A[5]), .A3(n17), .ZN(n16) );
  XNOR2_X1 U65 ( .A(A[4]), .B(n19), .ZN(SUM[4]) );
  NAND3_X1 U66 ( .A1(A[30]), .A2(A[29]), .A3(A[28]), .ZN(n24) );
  NAND2_X1 U67 ( .A1(A[28]), .A2(A[29]), .ZN(n27) );
  NAND2_X1 U68 ( .A1(A[24]), .A2(A[25]), .ZN(n32) );
  NAND2_X1 U69 ( .A1(A[27]), .A2(A[26]), .ZN(n31) );
  NAND2_X1 U70 ( .A1(A[20]), .A2(A[21]), .ZN(n36) );
  NAND2_X1 U71 ( .A1(A[23]), .A2(A[22]), .ZN(n35) );
  XNOR2_X1 U72 ( .A(A[23]), .B(n37), .ZN(SUM[23]) );
  NAND2_X1 U73 ( .A1(n38), .A2(A[22]), .ZN(n37) );
  INV_X1 U74 ( .A(n39), .ZN(n38) );
  NAND3_X1 U75 ( .A1(A[20]), .A2(A[21]), .A3(n42), .ZN(n39) );
  NAND2_X1 U76 ( .A1(A[16]), .A2(A[17]), .ZN(n44) );
  NAND2_X1 U77 ( .A1(A[19]), .A2(A[18]), .ZN(n43) );
  XOR2_X1 U78 ( .A(A[1]), .B(A[0]), .Z(SUM[1]) );
  XNOR2_X1 U79 ( .A(A[19]), .B(n45), .ZN(SUM[19]) );
  NAND2_X1 U80 ( .A1(n5), .A2(A[18]), .ZN(n45) );
  NAND2_X1 U81 ( .A1(A[12]), .A2(A[13]), .ZN(n48) );
  NAND2_X1 U82 ( .A1(A[15]), .A2(A[14]), .ZN(n47) );
  XNOR2_X1 U83 ( .A(A[15]), .B(n49), .ZN(SUM[15]) );
  NAND2_X1 U84 ( .A1(n50), .A2(A[14]), .ZN(n49) );
  INV_X1 U85 ( .A(n51), .ZN(n50) );
  NAND3_X1 U86 ( .A1(A[12]), .A2(A[13]), .A3(n3), .ZN(n51) );
  NAND2_X1 U87 ( .A1(A[8]), .A2(A[9]), .ZN(n57) );
  NAND2_X1 U88 ( .A1(A[11]), .A2(A[10]), .ZN(n56) );
  XNOR2_X1 U89 ( .A(A[11]), .B(n58), .ZN(SUM[11]) );
  NAND2_X1 U90 ( .A1(n6), .A2(A[10]), .ZN(n58) );
  INV_X1 U91 ( .A(n13), .ZN(n54) );
  NAND2_X1 U92 ( .A1(A[4]), .A2(A[5]), .ZN(n61) );
  NAND2_X1 U93 ( .A1(A[7]), .A2(A[6]), .ZN(n60) );
  INV_X1 U94 ( .A(n19), .ZN(n17) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 ( 
        Clk, Rst, IR_IN, IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, 
        RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
        EQ_COND, .ALU_OPCODE({\ALU_OPCODE[5] , \ALU_OPCODE[4] , 
        \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), 
        signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
        WB_MUX_SEL, RF_WE, lhi_sel, sb_op, s_trap, s_ret );
  input [31:0] IR_IN;
  input Clk, Rst;
  output IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN,
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND,
         \ALU_OPCODE[5] , \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] ,
         \ALU_OPCODE[1] , \ALU_OPCODE[0] , signed_unsigned, DRAM_WE,
         LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE, lhi_sel, sb_op,
         s_trap, s_ret;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274,
         N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         signed_unsigned_i, N550, N551, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n336, n339, n340, n343, n344, n345, n377, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n335, n337, n338, n341, n342,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n378, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549;
  wire   [5:0] ALU_OPCODE;
  wire   [5:0] aluOpcode1;
  wire   [5:0] aluOpcode2;
  wire   [31:0] iterator_trap;
  wire   [31:0] iterator_ret;
  wire   [31:0] iterator1;
  wire   [5:0] aluOpcode_i;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];
  assign IR_LATCH_EN = 1'b0;
  assign NPC_LATCH_EN = 1'b0;
  assign RegA_LATCH_EN = 1'b0;
  assign RegB_LATCH_EN = 1'b0;
  assign RegIMM_LATCH_EN = 1'b0;
  assign MUXA_SEL = 1'b0;
  assign MUXB_SEL = 1'b0;
  assign ALU_OUTREG_EN = 1'b0;
  assign EQ_COND = 1'b0;
  assign DRAM_WE = 1'b0;
  assign LMD_LATCH_EN = 1'b0;
  assign JUMP_EN = 1'b0;
  assign PC_LATCH_EN = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign RF_WE = 1'b0;

  DFFR_X1 \aluOpcode1_reg[5]  ( .D(aluOpcode_i[5]), .CK(Clk), .RN(n64), .Q(
        aluOpcode1[5]) );
  DFFR_X1 \aluOpcode1_reg[4]  ( .D(aluOpcode_i[4]), .CK(Clk), .RN(n63), .Q(
        aluOpcode1[4]) );
  DFFR_X1 \aluOpcode1_reg[3]  ( .D(aluOpcode_i[3]), .CK(Clk), .RN(n63), .Q(
        aluOpcode1[3]) );
  DFFR_X1 \aluOpcode1_reg[2]  ( .D(aluOpcode_i[2]), .CK(Clk), .RN(n63), .Q(
        aluOpcode1[2]) );
  DFFR_X1 \aluOpcode1_reg[1]  ( .D(aluOpcode_i[1]), .CK(Clk), .RN(n63), .Q(
        aluOpcode1[1]) );
  DFFR_X1 \aluOpcode1_reg[0]  ( .D(aluOpcode_i[0]), .CK(Clk), .RN(n63), .Q(
        aluOpcode1[0]) );
  DFFR_X1 \aluOpcode2_reg[5]  ( .D(aluOpcode1[5]), .CK(Clk), .RN(n63), .Q(
        aluOpcode2[5]) );
  DFFR_X1 \aluOpcode2_reg[4]  ( .D(aluOpcode1[4]), .CK(Clk), .RN(n63), .Q(
        aluOpcode2[4]) );
  DFFR_X1 \aluOpcode2_reg[3]  ( .D(aluOpcode1[3]), .CK(Clk), .RN(n63), .Q(
        aluOpcode2[3]) );
  DFFR_X1 \aluOpcode2_reg[2]  ( .D(aluOpcode1[2]), .CK(Clk), .RN(n63), .Q(
        aluOpcode2[2]) );
  DFFR_X1 \aluOpcode2_reg[1]  ( .D(aluOpcode1[1]), .CK(Clk), .RN(n64), .Q(
        aluOpcode2[1]) );
  DFFR_X1 \aluOpcode2_reg[0]  ( .D(aluOpcode1[0]), .CK(Clk), .RN(n64), .Q(
        aluOpcode2[0]) );
  DFFR_X1 \aluOpcode3_reg[5]  ( .D(aluOpcode2[5]), .CK(Clk), .RN(n64), .Q(
        ALU_OPCODE[5]) );
  DFFR_X1 \aluOpcode3_reg[4]  ( .D(aluOpcode2[4]), .CK(Clk), .RN(n64), .Q(
        ALU_OPCODE[4]) );
  DFFR_X1 \aluOpcode3_reg[3]  ( .D(aluOpcode2[3]), .CK(Clk), .RN(n64), .Q(
        ALU_OPCODE[3]) );
  DFFR_X1 \aluOpcode3_reg[2]  ( .D(aluOpcode2[2]), .CK(Clk), .RN(n64), .Q(
        ALU_OPCODE[2]) );
  DFFR_X1 \aluOpcode3_reg[1]  ( .D(aluOpcode2[1]), .CK(Clk), .RN(n64), .Q(
        ALU_OPCODE[1]) );
  DFFR_X1 \aluOpcode3_reg[0]  ( .D(aluOpcode2[0]), .CK(Clk), .RN(n64), .Q(
        ALU_OPCODE[0]) );
  DFF_X1 \iterator_ret_reg[26]  ( .D(n439), .CK(Clk), .Q(iterator_ret[26]), 
        .QN(n329) );
  DFF_X1 \iterator_ret_reg[20]  ( .D(n433), .CK(Clk), .Q(iterator_ret[20]), 
        .QN(n323) );
  DFF_X1 \iterator_ret_reg[19]  ( .D(n432), .CK(Clk), .Q(iterator_ret[19]), 
        .QN(n322) );
  DFF_X1 \iterator_ret_reg[16]  ( .D(n429), .CK(Clk), .Q(iterator_ret[16]), 
        .QN(n319) );
  DFF_X1 \iterator_ret_reg[14]  ( .D(n427), .CK(Clk), .Q(iterator_ret[14]), 
        .QN(n317) );
  DFF_X1 \iterator_ret_reg[8]  ( .D(n421), .CK(Clk), .Q(iterator_ret[8]), .QN(
        n311) );
  DFF_X1 \iterator_ret_reg[7]  ( .D(n420), .CK(Clk), .Q(iterator_ret[7]), .QN(
        n310) );
  DFF_X1 \iterator1_reg[30]  ( .D(n519), .CK(Clk), .Q(iterator1[30]), .QN(n133) );
  DFF_X1 \iterator1_reg[29]  ( .D(n520), .CK(Clk), .Q(iterator1[29]), .QN(n131) );
  DFF_X1 \iterator1_reg[28]  ( .D(n521), .CK(Clk), .Q(iterator1[28]), .QN(n129) );
  DFF_X1 \iterator1_reg[27]  ( .D(n522), .CK(Clk), .Q(iterator1[27]), .QN(n127) );
  DFF_X1 \iterator1_reg[26]  ( .D(n523), .CK(Clk), .Q(iterator1[26]), .QN(n125) );
  DFF_X1 \iterator1_reg[25]  ( .D(n524), .CK(Clk), .Q(iterator1[25]), .QN(n123) );
  DFF_X1 \iterator1_reg[24]  ( .D(n525), .CK(Clk), .Q(iterator1[24]), .QN(n121) );
  DFF_X1 \iterator1_reg[23]  ( .D(n526), .CK(Clk), .Q(iterator1[23]), .QN(n119) );
  DFF_X1 \iterator1_reg[22]  ( .D(n527), .CK(Clk), .Q(iterator1[22]), .QN(n117) );
  DFF_X1 \iterator1_reg[21]  ( .D(n528), .CK(Clk), .Q(iterator1[21]), .QN(n115) );
  DFF_X1 \iterator1_reg[20]  ( .D(n529), .CK(Clk), .Q(iterator1[20]), .QN(n113) );
  DFF_X1 \iterator1_reg[19]  ( .D(n530), .CK(Clk), .Q(iterator1[19]), .QN(n111) );
  DFF_X1 \iterator1_reg[18]  ( .D(n531), .CK(Clk), .Q(iterator1[18]), .QN(n109) );
  DFF_X1 \iterator1_reg[17]  ( .D(n532), .CK(Clk), .Q(iterator1[17]), .QN(n107) );
  DFF_X1 \iterator1_reg[16]  ( .D(n533), .CK(Clk), .Q(iterator1[16]), .QN(n105) );
  DFF_X1 \iterator1_reg[15]  ( .D(n534), .CK(Clk), .Q(iterator1[15]), .QN(n103) );
  DFF_X1 \iterator1_reg[14]  ( .D(n535), .CK(Clk), .Q(iterator1[14]), .QN(n101) );
  DFF_X1 \iterator1_reg[13]  ( .D(n536), .CK(Clk), .Q(iterator1[13]), .QN(n99)
         );
  DFF_X1 \iterator1_reg[12]  ( .D(n537), .CK(Clk), .Q(iterator1[12]), .QN(n97)
         );
  DFF_X1 \iterator1_reg[11]  ( .D(n538), .CK(Clk), .Q(iterator1[11]), .QN(n95)
         );
  DFF_X1 \iterator1_reg[10]  ( .D(n539), .CK(Clk), .Q(iterator1[10]), .QN(n93)
         );
  DFF_X1 \iterator1_reg[9]  ( .D(n540), .CK(Clk), .Q(iterator1[9]), .QN(n91)
         );
  DFF_X1 \iterator1_reg[8]  ( .D(n541), .CK(Clk), .Q(iterator1[8]), .QN(n89)
         );
  DFF_X1 \iterator1_reg[7]  ( .D(n542), .CK(Clk), .Q(iterator1[7]), .QN(n87)
         );
  DFF_X1 \iterator1_reg[6]  ( .D(n543), .CK(Clk), .Q(iterator1[6]), .QN(n85)
         );
  DFF_X1 \iterator1_reg[5]  ( .D(n544), .CK(Clk), .Q(iterator1[5]), .QN(n83)
         );
  DFF_X1 \iterator1_reg[4]  ( .D(n545), .CK(Clk), .Q(iterator1[4]), .QN(n81)
         );
  DFF_X1 \iterator1_reg[31]  ( .D(n549), .CK(Clk), .Q(iterator1[31]), .QN(n76)
         );
  DFF_X1 sb_op_reg ( .D(n345), .CK(Clk), .Q(sb_op) );
  DLH_X1 signed_unsigned_i_reg ( .G(N550), .D(N551), .Q(signed_unsigned_i) );
  DFF_X1 signed_unsigned_1_reg ( .D(n344), .CK(Clk), .Q(n249) );
  DFF_X1 signed_unsigned_2_reg ( .D(n343), .CK(Clk), .Q(signed_unsigned) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_3 add_239 ( 
        .A(iterator_ret), .SUM({N176, N175, N174, N173, N172, N171, N170, N169, 
        N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, 
        N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145}) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 add_217 ( 
        .A(iterator_trap), .SUM({N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34}) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 add_258 ( 
        .A(iterator1), .SUM({N284, N283, N282, N281, N280, N279, N278, N277, 
        N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253}) );
  DFF_X1 \iterator_ret_reg[21]  ( .D(n434), .CK(Clk), .Q(iterator_ret[21]), 
        .QN(n324) );
  DFF_X1 \iterator_ret_reg[24]  ( .D(n437), .CK(Clk), .Q(iterator_ret[24]), 
        .QN(n327) );
  DFF_X1 lhi_sel_reg ( .D(n377), .CK(Clk), .Q(lhi_sel), .QN(n336) );
  DFF_X1 \iterator1_reg[3]  ( .D(n546), .CK(Clk), .Q(iterator1[3]), .QN(n40)
         );
  DFF_X1 \iterator1_reg[2]  ( .D(n547), .CK(Clk), .Q(iterator1[2]), .QN(n41)
         );
  DFF_X1 \iterator1_reg[1]  ( .D(n548), .CK(Clk), .Q(iterator1[1]), .QN(n42)
         );
  DFF_X1 \iterator1_reg[0]  ( .D(n518), .CK(Clk), .Q(iterator1[0]), .QN(n43)
         );
  DFF_X1 s_ret_reg ( .D(n379), .CK(Clk), .Q(s_ret), .QN(n340) );
  DFF_X1 \iterator_trap_reg[0]  ( .D(n381), .CK(Clk), .Q(iterator_trap[0]), 
        .QN(n271) );
  DFF_X1 \iterator_trap_reg[29]  ( .D(n410), .CK(Clk), .Q(iterator_trap[29]), 
        .QN(n300) );
  DFF_X1 \iterator_trap_reg[6]  ( .D(n387), .CK(Clk), .Q(iterator_trap[6]), 
        .QN(n277) );
  DFF_X1 \iterator_trap_reg[17]  ( .D(n398), .CK(Clk), .Q(iterator_trap[17]), 
        .QN(n288) );
  DFF_X1 \iterator_trap_reg[13]  ( .D(n394), .CK(Clk), .Q(iterator_trap[13]), 
        .QN(n284) );
  DFF_X1 \iterator_trap_reg[9]  ( .D(n390), .CK(Clk), .Q(iterator_trap[9]), 
        .QN(n280) );
  DFF_X1 \iterator_trap_reg[30]  ( .D(n411), .CK(Clk), .Q(iterator_trap[30]), 
        .QN(n301) );
  DFF_X1 \iterator_trap_reg[26]  ( .D(n407), .CK(Clk), .Q(iterator_trap[26]), 
        .QN(n297) );
  DFF_X1 sig1_reg ( .D(n446), .CK(Clk), .Q(n188), .QN(n517) );
  DFF_X1 s_trap_reg ( .D(n380), .CK(Clk), .Q(s_trap), .QN(n339) );
  DFF_X1 sig2_reg ( .D(n445), .CK(Clk), .Q(n140) );
  DFF_X1 \iterator_ret_reg[0]  ( .D(n413), .CK(Clk), .Q(iterator_ret[0]), .QN(
        n303) );
  DFF_X1 \iterator_ret_reg[29]  ( .D(n442), .CK(Clk), .Q(iterator_ret[29]), 
        .QN(n332) );
  DFF_X1 \iterator_ret_reg[27]  ( .D(n440), .CK(Clk), .Q(iterator_ret[27]), 
        .QN(n330) );
  DFF_X1 \iterator_ret_reg[30]  ( .D(n443), .CK(Clk), .Q(iterator_ret[30]), 
        .QN(n333) );
  DFF_X1 \iterator_ret_reg[22]  ( .D(n435), .CK(Clk), .Q(iterator_ret[22]), 
        .QN(n325) );
  DFF_X1 \iterator_trap_reg[18]  ( .D(n399), .CK(Clk), .Q(iterator_trap[18]), 
        .QN(n289) );
  DFF_X1 \iterator_trap_reg[14]  ( .D(n395), .CK(Clk), .Q(iterator_trap[14]), 
        .QN(n285) );
  DFF_X1 \iterator_trap_reg[22]  ( .D(n403), .CK(Clk), .Q(iterator_trap[22]), 
        .QN(n293) );
  DFF_X1 \iterator_trap_reg[21]  ( .D(n402), .CK(Clk), .Q(iterator_trap[21]), 
        .QN(n292) );
  DFF_X1 \iterator_ret_reg[23]  ( .D(n436), .CK(Clk), .Q(iterator_ret[23]), 
        .QN(n326) );
  DFF_X1 \iterator_ret_reg[18]  ( .D(n431), .CK(Clk), .Q(iterator_ret[18]), 
        .QN(n321) );
  DFF_X1 \iterator_ret_reg[17]  ( .D(n430), .CK(Clk), .Q(iterator_ret[17]), 
        .QN(n320) );
  DFF_X1 \iterator_ret_reg[15]  ( .D(n428), .CK(Clk), .Q(iterator_ret[15]), 
        .QN(n318) );
  DFF_X1 \iterator_ret_reg[13]  ( .D(n426), .CK(Clk), .Q(iterator_ret[13]), 
        .QN(n316) );
  DFF_X1 \iterator_ret_reg[12]  ( .D(n425), .CK(Clk), .Q(iterator_ret[12]), 
        .QN(n315) );
  DFF_X1 \iterator_ret_reg[10]  ( .D(n423), .CK(Clk), .Q(iterator_ret[10]), 
        .QN(n313) );
  DFF_X1 \iterator_ret_reg[9]  ( .D(n422), .CK(Clk), .Q(iterator_ret[9]), .QN(
        n312) );
  DFF_X1 \iterator_ret_reg[11]  ( .D(n424), .CK(Clk), .Q(iterator_ret[11]), 
        .QN(n314) );
  DFF_X1 \iterator_trap_reg[4]  ( .D(n385), .CK(Clk), .Q(iterator_trap[4]), 
        .QN(n275) );
  DFF_X1 \iterator_trap_reg[10]  ( .D(n391), .CK(Clk), .Q(iterator_trap[10]), 
        .QN(n281) );
  DFF_X1 \iterator_trap_reg[27]  ( .D(n408), .CK(Clk), .Q(iterator_trap[27]), 
        .QN(n298) );
  DFF_X1 \iterator_trap_reg[23]  ( .D(n404), .CK(Clk), .Q(iterator_trap[23]), 
        .QN(n294) );
  DFF_X1 \iterator_trap_reg[20]  ( .D(n401), .CK(Clk), .Q(iterator_trap[20]), 
        .QN(n291) );
  DFF_X1 \iterator_trap_reg[19]  ( .D(n400), .CK(Clk), .Q(iterator_trap[19]), 
        .QN(n290) );
  DFF_X1 \iterator_ret_reg[2]  ( .D(n415), .CK(Clk), .Q(iterator_ret[2]), .QN(
        n305) );
  DFF_X1 \iterator_ret_reg[31]  ( .D(n444), .CK(Clk), .Q(iterator_ret[31]), 
        .QN(n334) );
  DFF_X1 \iterator_ret_reg[6]  ( .D(n419), .CK(Clk), .Q(iterator_ret[6]), .QN(
        n309) );
  DFF_X1 \iterator_ret_reg[5]  ( .D(n418), .CK(Clk), .Q(iterator_ret[5]), .QN(
        n308) );
  DFF_X1 \iterator_ret_reg[4]  ( .D(n417), .CK(Clk), .Q(iterator_ret[4]), .QN(
        n307) );
  DFF_X1 \iterator_ret_reg[3]  ( .D(n416), .CK(Clk), .Q(iterator_ret[3]), .QN(
        n306) );
  DFF_X1 \iterator_ret_reg[1]  ( .D(n414), .CK(Clk), .Q(iterator_ret[1]), .QN(
        n304) );
  DFF_X1 \iterator_trap_reg[2]  ( .D(n383), .CK(Clk), .Q(iterator_trap[2]), 
        .QN(n273) );
  DFF_X1 \iterator_trap_reg[1]  ( .D(n382), .CK(Clk), .Q(iterator_trap[1]), 
        .QN(n272) );
  DFF_X1 \iterator_trap_reg[31]  ( .D(n412), .CK(Clk), .Q(iterator_trap[31]), 
        .QN(n302) );
  DFF_X1 \iterator_trap_reg[7]  ( .D(n388), .CK(Clk), .Q(iterator_trap[7]), 
        .QN(n278) );
  DFF_X1 \iterator_trap_reg[5]  ( .D(n386), .CK(Clk), .Q(iterator_trap[5]), 
        .QN(n276) );
  DFF_X1 \iterator_trap_reg[3]  ( .D(n384), .CK(Clk), .Q(iterator_trap[3]), 
        .QN(n274) );
  DFF_X1 \iterator_trap_reg[24]  ( .D(n405), .CK(Clk), .Q(iterator_trap[24]), 
        .QN(n295) );
  DFF_X1 \iterator_trap_reg[16]  ( .D(n397), .CK(Clk), .Q(iterator_trap[16]), 
        .QN(n287) );
  DFF_X1 \iterator_trap_reg[15]  ( .D(n396), .CK(Clk), .Q(iterator_trap[15]), 
        .QN(n286) );
  DFF_X1 \iterator_trap_reg[12]  ( .D(n393), .CK(Clk), .Q(iterator_trap[12]), 
        .QN(n283) );
  DFF_X1 \iterator_trap_reg[11]  ( .D(n392), .CK(Clk), .Q(iterator_trap[11]), 
        .QN(n282) );
  DFF_X1 \iterator_trap_reg[8]  ( .D(n389), .CK(Clk), .Q(iterator_trap[8]), 
        .QN(n279) );
  DFF_X1 \iterator_trap_reg[28]  ( .D(n409), .CK(Clk), .Q(iterator_trap[28]), 
        .QN(n299) );
  DFF_X1 \iterator_trap_reg[25]  ( .D(n406), .CK(Clk), .Q(iterator_trap[25]), 
        .QN(n296) );
  DFF_X1 \iterator_ret_reg[28]  ( .D(n441), .CK(Clk), .Q(iterator_ret[28]), 
        .QN(n331) );
  DFF_X1 \iterator_ret_reg[25]  ( .D(n438), .CK(Clk), .Q(iterator_ret[25]), 
        .QN(n328) );
  AND3_X2 U3 ( .A1(n27), .A2(n146), .A3(n147), .ZN(n45) );
  AND2_X2 U4 ( .A1(n152), .A2(n55), .ZN(n1) );
  INV_X1 U5 ( .A(n1), .ZN(n186) );
  CLKBUF_X1 U6 ( .A(N163), .Z(n2) );
  AND2_X1 U7 ( .A1(n196), .A2(n60), .ZN(n31) );
  AND2_X1 U8 ( .A1(n32), .A2(n194), .ZN(n3) );
  OR2_X1 U9 ( .A1(N54), .A2(N52), .ZN(n4) );
  BUF_X1 U10 ( .A(n185), .Z(n55) );
  OR2_X1 U11 ( .A1(n199), .A2(n198), .ZN(n5) );
  INV_X1 U12 ( .A(n31), .ZN(n6) );
  OR2_X1 U13 ( .A1(N162), .A2(N165), .ZN(n7) );
  CLKBUF_X1 U14 ( .A(N175), .Z(n8) );
  INV_X1 U15 ( .A(n26), .ZN(n61) );
  CLKBUF_X1 U16 ( .A(N166), .Z(n9) );
  CLKBUF_X1 U17 ( .A(N168), .Z(n10) );
  AND2_X1 U18 ( .A1(n33), .A2(n148), .ZN(n11) );
  CLKBUF_X1 U19 ( .A(n38), .Z(n12) );
  CLKBUF_X1 U20 ( .A(N57), .Z(n13) );
  OR2_X1 U21 ( .A1(N59), .A2(N58), .ZN(n14) );
  CLKBUF_X1 U22 ( .A(N164), .Z(n15) );
  NAND2_X1 U23 ( .A1(n45), .A2(n11), .ZN(n16) );
  AND2_X1 U24 ( .A1(n17), .A2(n180), .ZN(n146) );
  NOR3_X1 U25 ( .A1(N173), .A2(N170), .A3(N171), .ZN(n17) );
  INV_X1 U26 ( .A(N61), .ZN(n18) );
  BUF_X1 U27 ( .A(n45), .Z(n37) );
  NOR3_X1 U28 ( .A1(N55), .A2(N53), .A3(n4), .ZN(n190) );
  NOR3_X1 U29 ( .A1(N164), .A2(N163), .A3(n7), .ZN(n144) );
  INV_X1 U30 ( .A(n31), .ZN(n19) );
  INV_X1 U31 ( .A(n31), .ZN(n20) );
  NOR3_X1 U32 ( .A1(n233), .A2(n230), .A3(n5), .ZN(n195) );
  AND2_X1 U33 ( .A1(n184), .A2(n46), .ZN(n21) );
  INV_X1 U34 ( .A(n25), .ZN(n22) );
  INV_X1 U35 ( .A(n25), .ZN(n62) );
  INV_X1 U36 ( .A(n26), .ZN(n23) );
  NAND2_X1 U37 ( .A1(n140), .A2(n187), .ZN(n24) );
  NAND2_X1 U38 ( .A1(n24), .A2(n34), .ZN(n445) );
  AND2_X1 U39 ( .A1(n196), .A2(n60), .ZN(n25) );
  AND2_X1 U40 ( .A1(n196), .A2(n60), .ZN(n26) );
  AND2_X1 U41 ( .A1(n144), .A2(n145), .ZN(n27) );
  NOR3_X1 U42 ( .A1(N57), .A2(N56), .A3(n14), .ZN(n191) );
  NAND2_X1 U43 ( .A1(n45), .A2(n11), .ZN(n184) );
  INV_X1 U44 ( .A(n26), .ZN(n28) );
  AND2_X1 U45 ( .A1(n16), .A2(n46), .ZN(n151) );
  NAND3_X1 U46 ( .A1(n21), .A2(n33), .A3(n37), .ZN(n29) );
  INV_X1 U47 ( .A(n36), .ZN(n30) );
  BUF_X1 U48 ( .A(n137), .Z(n48) );
  BUF_X1 U49 ( .A(n137), .Z(n47) );
  BUF_X1 U50 ( .A(n137), .Z(n49) );
  INV_X1 U51 ( .A(n36), .ZN(n56) );
  BUF_X1 U52 ( .A(n138), .Z(n50) );
  BUF_X1 U53 ( .A(n138), .Z(n51) );
  BUF_X1 U54 ( .A(n138), .Z(n52) );
  BUF_X1 U55 ( .A(n238), .Z(n58) );
  BUF_X1 U56 ( .A(n185), .Z(n54) );
  BUF_X1 U57 ( .A(n185), .Z(n53) );
  BUF_X1 U58 ( .A(n238), .Z(n59) );
  BUF_X1 U59 ( .A(n238), .Z(n60) );
  AND2_X1 U60 ( .A1(n193), .A2(n192), .ZN(n32) );
  AND2_X1 U61 ( .A1(n143), .A2(n142), .ZN(n33) );
  BUF_X1 U62 ( .A(Rst), .Z(n64) );
  BUF_X1 U63 ( .A(Rst), .Z(n63) );
  BUF_X1 U64 ( .A(Rst), .Z(n65) );
  INV_X1 U65 ( .A(n39), .ZN(n34) );
  INV_X1 U66 ( .A(n1), .ZN(n35) );
  AND2_X1 U67 ( .A1(n29), .A2(n55), .ZN(n36) );
  AND2_X1 U68 ( .A1(n29), .A2(n55), .ZN(n39) );
  INV_X1 U69 ( .A(n12), .ZN(n234) );
  AND2_X1 U70 ( .A1(n191), .A2(n190), .ZN(n38) );
  NAND3_X1 U71 ( .A1(n195), .A2(n3), .A3(n38), .ZN(n196) );
  NAND4_X1 U72 ( .A1(n224), .A2(n225), .A3(n226), .A4(n223), .ZN(n44) );
  NOR3_X1 U73 ( .A1(n150), .A2(n149), .A3(N146), .ZN(n46) );
  INV_X1 U74 ( .A(n39), .ZN(n57) );
  NAND2_X1 U75 ( .A1(IR_IN_26), .A2(IR_IN_27), .ZN(n495) );
  INV_X1 U76 ( .A(n495), .ZN(n241) );
  INV_X1 U77 ( .A(IR_IN_28), .ZN(n244) );
  INV_X1 U78 ( .A(n491), .ZN(n245) );
  NAND3_X1 U79 ( .A1(n374), .A2(n244), .A3(n245), .ZN(n246) );
  NAND3_X1 U80 ( .A1(n457), .A2(n374), .A3(n244), .ZN(n247) );
  INV_X1 U81 ( .A(IR_IN_31), .ZN(n242) );
  INV_X1 U82 ( .A(IR_IN_30), .ZN(n243) );
  NAND4_X1 U83 ( .A1(IR_IN_29), .A2(IR_IN_28), .A3(n242), .A4(n243), .ZN(n460)
         );
  INV_X1 U84 ( .A(n460), .ZN(n240) );
  NAND3_X1 U85 ( .A1(n65), .A2(n241), .A3(n240), .ZN(n136) );
  INV_X1 U86 ( .A(n136), .ZN(n137) );
  INV_X1 U87 ( .A(N274), .ZN(n116) );
  INV_X1 U88 ( .A(N273), .ZN(n114) );
  INV_X1 U89 ( .A(N272), .ZN(n112) );
  INV_X1 U90 ( .A(N271), .ZN(n110) );
  NAND4_X1 U91 ( .A1(n116), .A2(n114), .A3(n112), .A4(n110), .ZN(n69) );
  INV_X1 U92 ( .A(N278), .ZN(n124) );
  INV_X1 U93 ( .A(N277), .ZN(n122) );
  INV_X1 U94 ( .A(N276), .ZN(n120) );
  INV_X1 U95 ( .A(N275), .ZN(n118) );
  NAND4_X1 U96 ( .A1(n124), .A2(n122), .A3(n120), .A4(n118), .ZN(n68) );
  INV_X1 U97 ( .A(N282), .ZN(n132) );
  INV_X1 U98 ( .A(N281), .ZN(n130) );
  INV_X1 U99 ( .A(N280), .ZN(n128) );
  INV_X1 U100 ( .A(N279), .ZN(n126) );
  NAND4_X1 U101 ( .A1(n132), .A2(n130), .A3(n128), .A4(n126), .ZN(n67) );
  INV_X1 U102 ( .A(N284), .ZN(n77) );
  INV_X1 U103 ( .A(N283), .ZN(n134) );
  NAND4_X1 U104 ( .A1(N254), .A2(N253), .A3(n77), .A4(n134), .ZN(n66) );
  NOR4_X1 U105 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .ZN(n75) );
  INV_X1 U106 ( .A(N258), .ZN(n84) );
  INV_X1 U107 ( .A(N257), .ZN(n82) );
  INV_X1 U108 ( .A(N256), .ZN(n80) );
  INV_X1 U109 ( .A(N255), .ZN(n79) );
  NAND4_X1 U110 ( .A1(n84), .A2(n82), .A3(n80), .A4(n79), .ZN(n73) );
  INV_X1 U111 ( .A(N262), .ZN(n92) );
  INV_X1 U112 ( .A(N261), .ZN(n90) );
  INV_X1 U113 ( .A(N260), .ZN(n88) );
  INV_X1 U114 ( .A(N259), .ZN(n86) );
  NAND4_X1 U115 ( .A1(n92), .A2(n90), .A3(n88), .A4(n86), .ZN(n72) );
  INV_X1 U116 ( .A(N266), .ZN(n100) );
  INV_X1 U117 ( .A(N265), .ZN(n98) );
  INV_X1 U118 ( .A(N264), .ZN(n96) );
  INV_X1 U119 ( .A(N263), .ZN(n94) );
  NAND4_X1 U120 ( .A1(n100), .A2(n98), .A3(n96), .A4(n94), .ZN(n71) );
  INV_X1 U121 ( .A(N270), .ZN(n108) );
  INV_X1 U122 ( .A(N269), .ZN(n106) );
  INV_X1 U123 ( .A(N268), .ZN(n104) );
  INV_X1 U124 ( .A(N267), .ZN(n102) );
  NAND4_X1 U125 ( .A1(n108), .A2(n106), .A3(n104), .A4(n102), .ZN(n70) );
  NOR4_X1 U126 ( .A1(n73), .A2(n72), .A3(n71), .A4(n70), .ZN(n74) );
  NAND2_X1 U127 ( .A1(n75), .A2(n74), .ZN(n135) );
  NAND2_X1 U128 ( .A1(n49), .A2(n135), .ZN(n138) );
  OAI22_X1 U129 ( .A1(n50), .A2(n77), .B1(n49), .B2(n76), .ZN(n549) );
  INV_X1 U130 ( .A(N254), .ZN(n78) );
  OAI22_X1 U131 ( .A1(n78), .A2(n52), .B1(n49), .B2(n42), .ZN(n548) );
  OAI22_X1 U132 ( .A1(n50), .A2(n79), .B1(n49), .B2(n41), .ZN(n547) );
  OAI22_X1 U133 ( .A1(n51), .A2(n80), .B1(n49), .B2(n40), .ZN(n546) );
  OAI22_X1 U134 ( .A1(n51), .A2(n82), .B1(n49), .B2(n81), .ZN(n545) );
  OAI22_X1 U135 ( .A1(n50), .A2(n84), .B1(n49), .B2(n83), .ZN(n544) );
  OAI22_X1 U136 ( .A1(n51), .A2(n86), .B1(n49), .B2(n85), .ZN(n543) );
  OAI22_X1 U137 ( .A1(n50), .A2(n88), .B1(n49), .B2(n87), .ZN(n542) );
  OAI22_X1 U138 ( .A1(n50), .A2(n90), .B1(n48), .B2(n89), .ZN(n541) );
  OAI22_X1 U139 ( .A1(n50), .A2(n92), .B1(n48), .B2(n91), .ZN(n540) );
  OAI22_X1 U140 ( .A1(n50), .A2(n94), .B1(n48), .B2(n93), .ZN(n539) );
  OAI22_X1 U141 ( .A1(n51), .A2(n96), .B1(n48), .B2(n95), .ZN(n538) );
  OAI22_X1 U142 ( .A1(n50), .A2(n98), .B1(n48), .B2(n97), .ZN(n537) );
  OAI22_X1 U143 ( .A1(n51), .A2(n100), .B1(n48), .B2(n99), .ZN(n536) );
  OAI22_X1 U144 ( .A1(n50), .A2(n102), .B1(n48), .B2(n101), .ZN(n535) );
  OAI22_X1 U145 ( .A1(n51), .A2(n104), .B1(n48), .B2(n103), .ZN(n534) );
  OAI22_X1 U146 ( .A1(n51), .A2(n106), .B1(n48), .B2(n105), .ZN(n533) );
  OAI22_X1 U147 ( .A1(n50), .A2(n108), .B1(n48), .B2(n107), .ZN(n532) );
  OAI22_X1 U148 ( .A1(n51), .A2(n110), .B1(n48), .B2(n109), .ZN(n531) );
  OAI22_X1 U149 ( .A1(n52), .A2(n112), .B1(n48), .B2(n111), .ZN(n530) );
  OAI22_X1 U150 ( .A1(n52), .A2(n114), .B1(n47), .B2(n113), .ZN(n529) );
  OAI22_X1 U151 ( .A1(n52), .A2(n116), .B1(n47), .B2(n115), .ZN(n528) );
  OAI22_X1 U152 ( .A1(n52), .A2(n118), .B1(n47), .B2(n117), .ZN(n527) );
  OAI22_X1 U153 ( .A1(n50), .A2(n120), .B1(n47), .B2(n119), .ZN(n526) );
  OAI22_X1 U154 ( .A1(n52), .A2(n122), .B1(n47), .B2(n121), .ZN(n525) );
  OAI22_X1 U155 ( .A1(n52), .A2(n124), .B1(n47), .B2(n123), .ZN(n524) );
  OAI22_X1 U156 ( .A1(n52), .A2(n126), .B1(n47), .B2(n125), .ZN(n523) );
  OAI22_X1 U157 ( .A1(n52), .A2(n128), .B1(n47), .B2(n127), .ZN(n522) );
  OAI22_X1 U158 ( .A1(n51), .A2(n130), .B1(n47), .B2(n129), .ZN(n521) );
  OAI22_X1 U159 ( .A1(n51), .A2(n132), .B1(n47), .B2(n131), .ZN(n520) );
  OAI22_X1 U160 ( .A1(n51), .A2(n134), .B1(n47), .B2(n133), .ZN(n519) );
  OAI22_X1 U161 ( .A1(n136), .A2(n135), .B1(n336), .B2(n64), .ZN(n377) );
  INV_X1 U162 ( .A(N253), .ZN(n139) );
  OAI22_X1 U163 ( .A1(n139), .A2(n52), .B1(n47), .B2(n43), .ZN(n518) );
  INV_X1 U164 ( .A(n247), .ZN(n141) );
  OAI21_X1 U165 ( .B1(n141), .B2(n140), .A(n64), .ZN(n187) );
  INV_X1 U166 ( .A(n187), .ZN(n185) );
  INV_X1 U167 ( .A(N153), .ZN(n161) );
  INV_X1 U168 ( .A(N152), .ZN(n160) );
  INV_X1 U169 ( .A(N151), .ZN(n159) );
  INV_X1 U170 ( .A(N150), .ZN(n158) );
  NAND4_X1 U171 ( .A1(n161), .A2(n160), .A3(n159), .A4(n158), .ZN(n150) );
  INV_X1 U172 ( .A(N149), .ZN(n157) );
  INV_X1 U173 ( .A(N148), .ZN(n156) );
  NAND2_X1 U174 ( .A1(n157), .A2(n156), .ZN(n149) );
  NOR4_X1 U175 ( .A1(N160), .A2(N159), .A3(N158), .A4(N161), .ZN(n143) );
  NOR4_X1 U176 ( .A1(N154), .A2(N155), .A3(N156), .A4(N157), .ZN(n142) );
  NOR4_X1 U177 ( .A1(n150), .A2(n149), .A3(N145), .A4(N146), .ZN(n148) );
  INV_X1 U178 ( .A(N147), .ZN(n155) );
  NOR4_X1 U179 ( .A1(N174), .A2(N175), .A3(N176), .A4(n155), .ZN(n147) );
  NOR4_X1 U180 ( .A1(N168), .A2(N167), .A3(N166), .A4(N169), .ZN(n145) );
  NAND3_X1 U181 ( .A1(n151), .A2(n33), .A3(n37), .ZN(n152) );
  INV_X1 U182 ( .A(N176), .ZN(n153) );
  OAI22_X1 U183 ( .A1(n56), .A2(n153), .B1(n334), .B2(n55), .ZN(n444) );
  INV_X1 U184 ( .A(N146), .ZN(n154) );
  OAI22_X1 U185 ( .A1(n30), .A2(n154), .B1(n304), .B2(n55), .ZN(n414) );
  OAI22_X1 U186 ( .A1(n155), .A2(n57), .B1(n305), .B2(n55), .ZN(n415) );
  OAI22_X1 U187 ( .A1(n56), .A2(n156), .B1(n306), .B2(n55), .ZN(n416) );
  OAI22_X1 U188 ( .A1(n56), .A2(n157), .B1(n307), .B2(n55), .ZN(n417) );
  OAI22_X1 U189 ( .A1(n30), .A2(n158), .B1(n308), .B2(n55), .ZN(n418) );
  OAI22_X1 U190 ( .A1(n30), .A2(n159), .B1(n309), .B2(n55), .ZN(n419) );
  OAI22_X1 U191 ( .A1(n30), .A2(n160), .B1(n310), .B2(n54), .ZN(n420) );
  OAI22_X1 U192 ( .A1(n30), .A2(n161), .B1(n311), .B2(n54), .ZN(n421) );
  INV_X1 U193 ( .A(N154), .ZN(n162) );
  OAI22_X1 U194 ( .A1(n35), .A2(n162), .B1(n312), .B2(n54), .ZN(n422) );
  INV_X1 U195 ( .A(N155), .ZN(n163) );
  OAI22_X1 U196 ( .A1(n186), .A2(n163), .B1(n313), .B2(n54), .ZN(n423) );
  INV_X1 U197 ( .A(N156), .ZN(n164) );
  OAI22_X1 U198 ( .A1(n35), .A2(n164), .B1(n314), .B2(n54), .ZN(n424) );
  INV_X1 U199 ( .A(N157), .ZN(n165) );
  OAI22_X1 U200 ( .A1(n35), .A2(n165), .B1(n315), .B2(n54), .ZN(n425) );
  INV_X1 U201 ( .A(N158), .ZN(n166) );
  OAI22_X1 U202 ( .A1(n186), .A2(n166), .B1(n316), .B2(n54), .ZN(n426) );
  INV_X1 U203 ( .A(N159), .ZN(n167) );
  OAI22_X1 U204 ( .A1(n56), .A2(n167), .B1(n317), .B2(n54), .ZN(n427) );
  INV_X1 U205 ( .A(N160), .ZN(n168) );
  OAI22_X1 U206 ( .A1(n35), .A2(n168), .B1(n318), .B2(n54), .ZN(n428) );
  INV_X1 U207 ( .A(N161), .ZN(n169) );
  OAI22_X1 U208 ( .A1(n34), .A2(n169), .B1(n319), .B2(n54), .ZN(n429) );
  INV_X1 U209 ( .A(N162), .ZN(n170) );
  OAI22_X1 U210 ( .A1(n35), .A2(n170), .B1(n320), .B2(n54), .ZN(n430) );
  INV_X1 U211 ( .A(n2), .ZN(n171) );
  OAI22_X1 U212 ( .A1(n186), .A2(n171), .B1(n321), .B2(n53), .ZN(n431) );
  INV_X1 U213 ( .A(n15), .ZN(n172) );
  OAI22_X1 U214 ( .A1(n34), .A2(n172), .B1(n322), .B2(n53), .ZN(n432) );
  INV_X1 U215 ( .A(N165), .ZN(n173) );
  OAI22_X1 U216 ( .A1(n56), .A2(n173), .B1(n323), .B2(n53), .ZN(n433) );
  INV_X1 U217 ( .A(n9), .ZN(n174) );
  OAI22_X1 U218 ( .A1(n34), .A2(n174), .B1(n324), .B2(n53), .ZN(n434) );
  INV_X1 U219 ( .A(N167), .ZN(n175) );
  OAI22_X1 U220 ( .A1(n57), .A2(n175), .B1(n325), .B2(n53), .ZN(n435) );
  INV_X1 U221 ( .A(n10), .ZN(n176) );
  OAI22_X1 U222 ( .A1(n186), .A2(n176), .B1(n326), .B2(n54), .ZN(n436) );
  INV_X1 U223 ( .A(N169), .ZN(n177) );
  OAI22_X1 U224 ( .A1(n56), .A2(n177), .B1(n327), .B2(n53), .ZN(n437) );
  INV_X1 U225 ( .A(N170), .ZN(n178) );
  OAI22_X1 U226 ( .A1(n34), .A2(n178), .B1(n328), .B2(n53), .ZN(n438) );
  INV_X1 U227 ( .A(N171), .ZN(n179) );
  OAI22_X1 U228 ( .A1(n30), .A2(n179), .B1(n329), .B2(n53), .ZN(n439) );
  INV_X1 U229 ( .A(N172), .ZN(n180) );
  OAI22_X1 U230 ( .A1(n57), .A2(n180), .B1(n330), .B2(n53), .ZN(n440) );
  INV_X1 U231 ( .A(N173), .ZN(n181) );
  OAI22_X1 U232 ( .A1(n34), .A2(n181), .B1(n331), .B2(n53), .ZN(n441) );
  INV_X1 U233 ( .A(N174), .ZN(n182) );
  OAI22_X1 U234 ( .A1(n57), .A2(n182), .B1(n332), .B2(n53), .ZN(n442) );
  INV_X1 U235 ( .A(n8), .ZN(n183) );
  OAI22_X1 U236 ( .A1(n57), .A2(n183), .B1(n333), .B2(n53), .ZN(n443) );
  OAI22_X1 U237 ( .A1(n187), .A2(n16), .B1(n340), .B2(n64), .ZN(n379) );
  MUX2_X1 U238 ( .A(n187), .B(n1), .S(n303), .Z(n413) );
  INV_X1 U239 ( .A(n246), .ZN(n189) );
  OAI21_X1 U240 ( .B1(n189), .B2(n188), .A(n64), .ZN(n239) );
  INV_X1 U241 ( .A(n239), .ZN(n238) );
  INV_X1 U242 ( .A(N63), .ZN(n226) );
  INV_X1 U243 ( .A(N62), .ZN(n225) );
  INV_X1 U244 ( .A(N61), .ZN(n224) );
  INV_X1 U245 ( .A(N60), .ZN(n223) );
  NAND4_X1 U246 ( .A1(n226), .A2(n225), .A3(n18), .A4(n223), .ZN(n233) );
  INV_X1 U247 ( .A(N65), .ZN(n197) );
  INV_X1 U248 ( .A(N64), .ZN(n227) );
  NAND2_X1 U249 ( .A1(n197), .A2(n227), .ZN(n230) );
  INV_X1 U250 ( .A(N35), .ZN(n198) );
  INV_X1 U251 ( .A(N36), .ZN(n199) );
  NOR4_X1 U252 ( .A1(N51), .A2(N49), .A3(N50), .A4(N48), .ZN(n193) );
  NOR4_X1 U253 ( .A1(N44), .A2(N45), .A3(N46), .A4(N47), .ZN(n192) );
  INV_X1 U254 ( .A(N43), .ZN(n206) );
  INV_X1 U255 ( .A(N42), .ZN(n205) );
  INV_X1 U256 ( .A(N41), .ZN(n204) );
  INV_X1 U257 ( .A(N40), .ZN(n203) );
  NAND4_X1 U258 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(n229) );
  INV_X1 U259 ( .A(N39), .ZN(n202) );
  INV_X1 U260 ( .A(N38), .ZN(n201) );
  NAND2_X1 U261 ( .A1(n202), .A2(n201), .ZN(n228) );
  NOR4_X1 U262 ( .A1(n229), .A2(n228), .A3(N34), .A4(N37), .ZN(n194) );
  OAI22_X1 U263 ( .A1(n61), .A2(n197), .B1(n302), .B2(n60), .ZN(n412) );
  OAI22_X1 U264 ( .A1(n198), .A2(n20), .B1(n272), .B2(n60), .ZN(n382) );
  OAI22_X1 U265 ( .A1(n199), .A2(n6), .B1(n273), .B2(n60), .ZN(n383) );
  INV_X1 U266 ( .A(N37), .ZN(n200) );
  OAI22_X1 U267 ( .A1(n23), .A2(n200), .B1(n274), .B2(n60), .ZN(n384) );
  OAI22_X1 U268 ( .A1(n20), .A2(n201), .B1(n275), .B2(n60), .ZN(n385) );
  OAI22_X1 U269 ( .A1(n61), .A2(n202), .B1(n276), .B2(n60), .ZN(n386) );
  OAI22_X1 U270 ( .A1(n22), .A2(n203), .B1(n277), .B2(n60), .ZN(n387) );
  OAI22_X1 U271 ( .A1(n23), .A2(n204), .B1(n278), .B2(n60), .ZN(n388) );
  OAI22_X1 U272 ( .A1(n61), .A2(n205), .B1(n279), .B2(n59), .ZN(n389) );
  OAI22_X1 U273 ( .A1(n62), .A2(n206), .B1(n280), .B2(n59), .ZN(n390) );
  INV_X1 U274 ( .A(N44), .ZN(n207) );
  OAI22_X1 U275 ( .A1(n19), .A2(n207), .B1(n281), .B2(n59), .ZN(n391) );
  INV_X1 U276 ( .A(N45), .ZN(n208) );
  OAI22_X1 U277 ( .A1(n28), .A2(n208), .B1(n282), .B2(n59), .ZN(n392) );
  INV_X1 U278 ( .A(N46), .ZN(n209) );
  OAI22_X1 U279 ( .A1(n23), .A2(n209), .B1(n283), .B2(n59), .ZN(n393) );
  INV_X1 U280 ( .A(N47), .ZN(n210) );
  OAI22_X1 U281 ( .A1(n22), .A2(n210), .B1(n284), .B2(n59), .ZN(n394) );
  INV_X1 U282 ( .A(N48), .ZN(n211) );
  OAI22_X1 U283 ( .A1(n62), .A2(n211), .B1(n285), .B2(n59), .ZN(n395) );
  INV_X1 U284 ( .A(N49), .ZN(n212) );
  OAI22_X1 U285 ( .A1(n28), .A2(n212), .B1(n286), .B2(n59), .ZN(n396) );
  INV_X1 U286 ( .A(N50), .ZN(n213) );
  OAI22_X1 U287 ( .A1(n61), .A2(n213), .B1(n287), .B2(n59), .ZN(n397) );
  INV_X1 U288 ( .A(N51), .ZN(n214) );
  OAI22_X1 U289 ( .A1(n22), .A2(n214), .B1(n288), .B2(n59), .ZN(n398) );
  INV_X1 U290 ( .A(N52), .ZN(n215) );
  OAI22_X1 U291 ( .A1(n6), .A2(n215), .B1(n289), .B2(n59), .ZN(n399) );
  INV_X1 U292 ( .A(N53), .ZN(n216) );
  OAI22_X1 U293 ( .A1(n20), .A2(n216), .B1(n290), .B2(n58), .ZN(n400) );
  INV_X1 U294 ( .A(N54), .ZN(n217) );
  OAI22_X1 U295 ( .A1(n19), .A2(n217), .B1(n291), .B2(n58), .ZN(n401) );
  INV_X1 U296 ( .A(N55), .ZN(n218) );
  OAI22_X1 U297 ( .A1(n22), .A2(n218), .B1(n292), .B2(n58), .ZN(n402) );
  INV_X1 U298 ( .A(N56), .ZN(n219) );
  OAI22_X1 U299 ( .A1(n19), .A2(n219), .B1(n293), .B2(n58), .ZN(n403) );
  INV_X1 U300 ( .A(n13), .ZN(n220) );
  OAI22_X1 U301 ( .A1(n19), .A2(n220), .B1(n294), .B2(n58), .ZN(n404) );
  INV_X1 U302 ( .A(N58), .ZN(n221) );
  OAI22_X1 U303 ( .A1(n28), .A2(n221), .B1(n295), .B2(n59), .ZN(n405) );
  INV_X1 U304 ( .A(N59), .ZN(n222) );
  OAI22_X1 U305 ( .A1(n23), .A2(n222), .B1(n296), .B2(n58), .ZN(n406) );
  OAI22_X1 U306 ( .A1(n62), .A2(n223), .B1(n297), .B2(n58), .ZN(n407) );
  OAI22_X1 U307 ( .A1(n20), .A2(n224), .B1(n298), .B2(n58), .ZN(n408) );
  OAI22_X1 U308 ( .A1(n28), .A2(n225), .B1(n299), .B2(n58), .ZN(n409) );
  OAI22_X1 U309 ( .A1(n6), .A2(n226), .B1(n300), .B2(n58), .ZN(n410) );
  OAI22_X1 U310 ( .A1(n62), .A2(n227), .B1(n301), .B2(n58), .ZN(n411) );
  NOR4_X1 U311 ( .A1(n229), .A2(n228), .A3(N37), .A4(N35), .ZN(n236) );
  INV_X1 U312 ( .A(n230), .ZN(n231) );
  NAND4_X1 U313 ( .A1(N34), .A2(N36), .A3(n58), .A4(n231), .ZN(n232) );
  NOR3_X1 U314 ( .A1(n234), .A2(n44), .A3(n232), .ZN(n235) );
  NAND3_X1 U315 ( .A1(n236), .A2(n32), .A3(n235), .ZN(n237) );
  OAI21_X1 U316 ( .B1(n339), .B2(n65), .A(n237), .ZN(n380) );
  OAI21_X1 U317 ( .B1(n517), .B2(n60), .A(n6), .ZN(n446) );
  MUX2_X1 U318 ( .A(n239), .B(n25), .S(n271), .Z(n381) );
  MUX2_X1 U319 ( .A(sb_op), .B(n248), .S(n63), .Z(n345) );
  MUX2_X1 U320 ( .A(n249), .B(signed_unsigned_i), .S(n63), .Z(n344) );
  MUX2_X1 U321 ( .A(signed_unsigned), .B(n249), .S(n63), .Z(n343) );
  INV_X1 U322 ( .A(n250), .ZN(aluOpcode_i[5]) );
  AOI211_X1 U323 ( .C1(n241), .C2(n251), .A(n252), .B(n253), .ZN(n250) );
  OAI211_X1 U324 ( .C1(n254), .C2(n255), .A(n246), .B(n247), .ZN(n253) );
  AND4_X1 U325 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(n255) );
  OR2_X1 U326 ( .A1(n260), .A2(n261), .ZN(n257) );
  NAND4_X1 U327 ( .A1(n246), .A2(n262), .A3(n247), .A4(n263), .ZN(
        aluOpcode_i[4]) );
  AOI211_X1 U328 ( .C1(n264), .C2(n265), .A(n266), .B(n267), .ZN(n263) );
  INV_X1 U329 ( .A(n268), .ZN(n267) );
  OAI21_X1 U330 ( .B1(n269), .B2(n270), .A(n335), .ZN(n265) );
  NAND4_X1 U331 ( .A1(n337), .A2(n338), .A3(n341), .A4(n342), .ZN(
        aluOpcode_i[3]) );
  AOI211_X1 U332 ( .C1(n264), .C2(n346), .A(n347), .B(n348), .ZN(n342) );
  OAI221_X1 U333 ( .B1(n349), .B2(n269), .C1(n350), .C2(n351), .A(n335), .ZN(
        n346) );
  NAND4_X1 U334 ( .A1(n352), .A2(n353), .A3(n354), .A4(n355), .ZN(
        aluOpcode_i[2]) );
  AOI211_X1 U335 ( .C1(n356), .C2(n245), .A(n357), .B(n358), .ZN(n355) );
  INV_X1 U336 ( .A(n359), .ZN(n358) );
  AOI21_X1 U337 ( .B1(n264), .B2(n360), .A(n361), .ZN(n354) );
  OAI221_X1 U338 ( .B1(n261), .B2(n362), .C1(n363), .C2(n349), .A(n364), .ZN(
        n360) );
  NAND4_X1 U339 ( .A1(n365), .A2(n337), .A3(n366), .A4(n367), .ZN(
        aluOpcode_i[1]) );
  AOI221_X1 U340 ( .B1(n264), .B2(n368), .C1(n251), .C2(n369), .A(n370), .ZN(
        n367) );
  NAND3_X1 U341 ( .A1(n246), .A2(n352), .A3(n371), .ZN(n370) );
  INV_X1 U342 ( .A(n248), .ZN(n371) );
  NAND3_X1 U343 ( .A1(n372), .A2(n264), .A3(n373), .ZN(n352) );
  INV_X1 U344 ( .A(n375), .ZN(n369) );
  OAI21_X1 U345 ( .B1(n363), .B2(n260), .A(n376), .ZN(n368) );
  AOI22_X1 U346 ( .A1(n378), .A2(n245), .B1(n447), .B2(n241), .ZN(n366) );
  AOI22_X1 U347 ( .A1(n448), .A2(n264), .B1(n449), .B2(n356), .ZN(n337) );
  INV_X1 U348 ( .A(n450), .ZN(n365) );
  NAND4_X1 U349 ( .A1(n451), .A2(n452), .A3(n453), .A4(n454), .ZN(
        aluOpcode_i[0]) );
  AOI221_X1 U350 ( .B1(n251), .B2(n449), .C1(n455), .C2(n245), .A(n450), .ZN(
        n454) );
  NAND4_X1 U351 ( .A1(n341), .A2(n247), .A3(n456), .A4(n353), .ZN(n450) );
  AOI21_X1 U352 ( .B1(n264), .B2(n458), .A(n459), .ZN(n453) );
  AOI21_X1 U353 ( .B1(n460), .B2(n461), .A(n462), .ZN(n459) );
  NAND4_X1 U354 ( .A1(n256), .A2(n463), .A3(n464), .A4(n465), .ZN(n458) );
  AOI21_X1 U355 ( .B1(n466), .B2(n467), .A(n468), .ZN(n465) );
  INV_X1 U356 ( .A(n469), .ZN(n464) );
  AOI21_X1 U357 ( .B1(n470), .B2(n349), .A(n269), .ZN(n469) );
  INV_X1 U358 ( .A(n467), .ZN(n349) );
  NAND2_X1 U359 ( .A1(n270), .A2(n260), .ZN(n467) );
  NAND3_X1 U360 ( .A1(IR_IN_31), .A2(IR_IN_30), .A3(n471), .ZN(n452) );
  OAI21_X1 U361 ( .B1(n378), .B2(n356), .A(n457), .ZN(n451) );
  NAND4_X1 U362 ( .A1(n341), .A2(n472), .A3(n473), .A4(n262), .ZN(N551) );
  OAI211_X1 U363 ( .C1(n474), .C2(n475), .A(n244), .B(n476), .ZN(n473) );
  NOR2_X1 U364 ( .A1(n477), .A2(n462), .ZN(n475) );
  NOR4_X1 U365 ( .A1(IR_IN_31), .A2(IR_IN_30), .A3(n478), .A4(n479), .ZN(n474)
         );
  AOI21_X1 U366 ( .B1(n480), .B2(n481), .A(n482), .ZN(n478) );
  INV_X1 U367 ( .A(n266), .ZN(n472) );
  AOI21_X1 U368 ( .B1(n240), .B2(n457), .A(n361), .ZN(n341) );
  NAND4_X1 U369 ( .A1(n483), .A2(n484), .A3(n485), .A4(n486), .ZN(N550) );
  NOR3_X1 U370 ( .A1(n487), .A2(n266), .A3(n357), .ZN(n486) );
  OAI211_X1 U371 ( .C1(n460), .C2(n479), .A(n268), .B(n488), .ZN(n357) );
  AOI221_X1 U372 ( .B1(n251), .B2(n241), .C1(n356), .C2(n489), .A(n348), .ZN(
        n488) );
  AOI22_X1 U373 ( .A1(n245), .A2(n447), .B1(n490), .B2(n378), .ZN(n268) );
  NOR3_X1 U374 ( .A1(n476), .A2(n244), .A3(n477), .ZN(n378) );
  OAI211_X1 U375 ( .C1(n460), .C2(n491), .A(n338), .B(n492), .ZN(n266) );
  AOI221_X1 U376 ( .B1(n251), .B2(n457), .C1(n489), .C2(n487), .A(n493), .ZN(
        n492) );
  INV_X1 U377 ( .A(n353), .ZN(n493) );
  NAND3_X1 U378 ( .A1(IR_IN_31), .A2(n241), .A3(n494), .ZN(n353) );
  INV_X1 U379 ( .A(n496), .ZN(n251) );
  AOI21_X1 U395 ( .B1(n245), .B2(n356), .A(n497), .ZN(n338) );
  NOR3_X1 U396 ( .A1(n495), .A2(IR_IN_30), .A3(n498), .ZN(n497) );
  NAND2_X1 U397 ( .A1(n460), .A2(n496), .ZN(n487) );
  NAND2_X1 U398 ( .A1(n374), .A2(IR_IN_28), .ZN(n496) );
  NOR2_X1 U399 ( .A1(n477), .A2(IR_IN_29), .ZN(n374) );
  AOI21_X1 U400 ( .B1(n264), .B2(n499), .A(n252), .ZN(n485) );
  OR3_X1 U401 ( .A1(n361), .A2(n500), .A3(n347), .ZN(n252) );
  OAI211_X1 U402 ( .C1(n375), .C2(n461), .A(n456), .B(n359), .ZN(n347) );
  AOI21_X1 U403 ( .B1(IR_IN_31), .B2(n348), .A(n248), .ZN(n359) );
  NOR4_X1 U404 ( .A1(n242), .A2(n498), .A3(n479), .A4(IR_IN_30), .ZN(n248) );
  AND2_X1 U405 ( .A1(n455), .A2(n490), .ZN(n348) );
  NAND2_X1 U406 ( .A1(n479), .A2(n491), .ZN(n490) );
  INV_X1 U407 ( .A(n457), .ZN(n479) );
  NOR3_X1 U408 ( .A1(IR_IN_29), .A2(IR_IN_30), .A3(n244), .ZN(n455) );
  NAND3_X1 U409 ( .A1(IR_IN_31), .A2(n457), .A3(n494), .ZN(n456) );
  INV_X1 U410 ( .A(n447), .ZN(n461) );
  NOR2_X1 U411 ( .A1(n498), .A2(n477), .ZN(n447) );
  NAND2_X1 U412 ( .A1(IR_IN_30), .A2(n242), .ZN(n477) );
  NOR2_X1 U413 ( .A1(n449), .A2(n457), .ZN(n375) );
  INV_X1 U414 ( .A(n262), .ZN(n500) );
  OAI211_X1 U415 ( .C1(n501), .C2(n471), .A(IR_IN_30), .B(IR_IN_31), .ZN(n262)
         );
  NOR3_X1 U416 ( .A1(n476), .A2(n244), .A3(n491), .ZN(n471) );
  NAND2_X1 U417 ( .A1(IR_IN_26), .A2(n502), .ZN(n491) );
  INV_X1 U418 ( .A(IR_IN_29), .ZN(n476) );
  NOR2_X1 U419 ( .A1(n495), .A2(n498), .ZN(n501) );
  NOR4_X1 U420 ( .A1(n462), .A2(n242), .A3(n498), .A4(n243), .ZN(n361) );
  NAND4_X1 U421 ( .A1(n260), .A2(n270), .A3(n335), .A4(n503), .ZN(n499) );
  NOR2_X1 U422 ( .A1(n482), .A2(n448), .ZN(n503) );
  OAI22_X1 U423 ( .A1(n269), .A2(n470), .B1(n470), .B2(n504), .ZN(n448) );
  NAND3_X1 U424 ( .A1(n505), .A2(n506), .A3(IR_IN[2]), .ZN(n470) );
  INV_X1 U425 ( .A(n507), .ZN(n269) );
  OAI211_X1 U426 ( .C1(n363), .C2(n351), .A(n256), .B(n376), .ZN(n482) );
  AOI211_X1 U427 ( .C1(n507), .C2(n480), .A(n468), .B(n508), .ZN(n376) );
  OAI21_X1 U428 ( .B1(n362), .B2(n504), .A(n258), .ZN(n508) );
  NAND4_X1 U429 ( .A1(n481), .A2(IR_IN[4]), .A3(n505), .A4(n509), .ZN(n258) );
  INV_X1 U430 ( .A(n372), .ZN(n504) );
  OAI211_X1 U431 ( .C1(n350), .C2(n362), .A(n364), .B(n259), .ZN(n468) );
  NAND4_X1 U432 ( .A1(IR_IN[4]), .A2(IR_IN[2]), .A3(n507), .A4(n505), .ZN(n259) );
  NAND2_X1 U433 ( .A1(n373), .A2(n507), .ZN(n364) );
  INV_X1 U434 ( .A(n351), .ZN(n373) );
  INV_X1 U435 ( .A(n510), .ZN(n362) );
  NOR2_X1 U436 ( .A1(n511), .A2(IR_IN[1]), .ZN(n507) );
  NAND4_X1 U437 ( .A1(n466), .A2(IR_IN[4]), .A3(n505), .A4(n509), .ZN(n256) );
  NAND2_X1 U438 ( .A1(n512), .A2(IR_IN[2]), .ZN(n351) );
  INV_X1 U439 ( .A(n513), .ZN(n335) );
  OAI21_X1 U440 ( .B1(n363), .B2(n260), .A(n463), .ZN(n513) );
  OAI21_X1 U441 ( .B1(n480), .B2(n510), .A(n481), .ZN(n463) );
  INV_X1 U442 ( .A(n261), .ZN(n481) );
  NAND2_X1 U443 ( .A1(IR_IN[1]), .A2(IR_IN[0]), .ZN(n261) );
  NOR4_X1 U444 ( .A1(n509), .A2(IR_IN[3]), .A3(IR_IN[4]), .A4(IR_IN[5]), .ZN(
        n510) );
  INV_X1 U445 ( .A(n270), .ZN(n480) );
  NOR2_X1 U446 ( .A1(n466), .A2(n372), .ZN(n363) );
  NOR2_X1 U447 ( .A1(IR_IN[0]), .A2(IR_IN[1]), .ZN(n372) );
  INV_X1 U448 ( .A(n350), .ZN(n466) );
  NAND2_X1 U449 ( .A1(IR_IN[1]), .A2(n511), .ZN(n350) );
  INV_X1 U450 ( .A(IR_IN[0]), .ZN(n511) );
  NAND2_X1 U451 ( .A1(n512), .A2(n509), .ZN(n270) );
  NOR3_X1 U452 ( .A1(IR_IN[3]), .A2(IR_IN[4]), .A3(n514), .ZN(n512) );
  INV_X1 U453 ( .A(IR_IN[5]), .ZN(n514) );
  NAND3_X1 U454 ( .A1(n509), .A2(n506), .A3(n505), .ZN(n260) );
  AND2_X1 U455 ( .A1(IR_IN[5]), .A2(IR_IN[3]), .ZN(n505) );
  INV_X1 U456 ( .A(IR_IN[4]), .ZN(n506) );
  INV_X1 U457 ( .A(IR_IN[2]), .ZN(n509) );
  INV_X1 U458 ( .A(n254), .ZN(n264) );
  NAND4_X1 U459 ( .A1(n494), .A2(n457), .A3(n515), .A4(n516), .ZN(n254) );
  NOR4_X1 U460 ( .A1(IR_IN_31), .A2(IR_IN[9]), .A3(IR_IN[8]), .A4(IR_IN[7]), 
        .ZN(n516) );
  NOR2_X1 U461 ( .A1(IR_IN[6]), .A2(IR_IN[10]), .ZN(n515) );
  NOR2_X1 U462 ( .A1(IR_IN_26), .A2(IR_IN_27), .ZN(n457) );
  NOR3_X1 U463 ( .A1(IR_IN_29), .A2(IR_IN_30), .A3(IR_IN_28), .ZN(n494) );
  INV_X1 U464 ( .A(n356), .ZN(n484) );
  NOR3_X1 U465 ( .A1(IR_IN_30), .A2(IR_IN_31), .A3(n498), .ZN(n356) );
  NAND2_X1 U466 ( .A1(IR_IN_29), .A2(n244), .ZN(n498) );
  NAND3_X1 U467 ( .A1(n244), .A2(n242), .A3(n449), .ZN(n483) );
  NAND2_X1 U468 ( .A1(n462), .A2(n495), .ZN(n449) );
  INV_X1 U469 ( .A(n489), .ZN(n462) );
  NOR2_X1 U470 ( .A1(n502), .A2(IR_IN_26), .ZN(n489) );
  INV_X1 U471 ( .A(IR_IN_27), .ZN(n502) );
endmodule


module regFFD_NBIT32_0 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;

  DFFR_X1 \Q_reg[31]  ( .D(n96), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n64) );
  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n63) );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n62) );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n61) );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n60) );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n59) );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n58) );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n57) );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n56) );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n55) );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n54) );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n53) );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n52) );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n51) );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n50) );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n49) );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n48) );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n47) );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n46) );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n45) );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n44) );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n43) );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n42) );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n41) );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n40) );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n39) );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n38) );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n37) );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n36) );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n35) );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n34) );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n33) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n33), .B2(ENABLE), .A(n1), .ZN(n65) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n1) );
  OAI21_X1 U7 ( .B1(n34), .B2(ENABLE), .A(n2), .ZN(n66) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n2) );
  OAI21_X1 U9 ( .B1(n35), .B2(ENABLE), .A(n3), .ZN(n67) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n3) );
  OAI21_X1 U11 ( .B1(n36), .B2(ENABLE), .A(n4), .ZN(n68) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n4) );
  OAI21_X1 U13 ( .B1(n37), .B2(ENABLE), .A(n5), .ZN(n69) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n5) );
  OAI21_X1 U15 ( .B1(n38), .B2(ENABLE), .A(n6), .ZN(n70) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n6) );
  OAI21_X1 U17 ( .B1(n39), .B2(ENABLE), .A(n7), .ZN(n71) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n7) );
  OAI21_X1 U19 ( .B1(n40), .B2(ENABLE), .A(n8), .ZN(n72) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n8) );
  OAI21_X1 U21 ( .B1(n41), .B2(ENABLE), .A(n9), .ZN(n73) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n9) );
  OAI21_X1 U23 ( .B1(n42), .B2(ENABLE), .A(n10), .ZN(n74) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n10) );
  OAI21_X1 U25 ( .B1(n43), .B2(ENABLE), .A(n11), .ZN(n75) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n11) );
  OAI21_X1 U27 ( .B1(n44), .B2(ENABLE), .A(n12), .ZN(n76) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n12) );
  OAI21_X1 U29 ( .B1(n45), .B2(ENABLE), .A(n13), .ZN(n77) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n13) );
  OAI21_X1 U31 ( .B1(n46), .B2(ENABLE), .A(n14), .ZN(n78) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n14) );
  OAI21_X1 U33 ( .B1(n47), .B2(ENABLE), .A(n15), .ZN(n79) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n15) );
  OAI21_X1 U35 ( .B1(n48), .B2(ENABLE), .A(n16), .ZN(n80) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n16) );
  OAI21_X1 U37 ( .B1(n49), .B2(ENABLE), .A(n17), .ZN(n81) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n17) );
  OAI21_X1 U39 ( .B1(n50), .B2(ENABLE), .A(n18), .ZN(n82) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n18) );
  OAI21_X1 U41 ( .B1(n51), .B2(ENABLE), .A(n19), .ZN(n83) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n19) );
  OAI21_X1 U43 ( .B1(n52), .B2(ENABLE), .A(n20), .ZN(n84) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n20) );
  OAI21_X1 U45 ( .B1(n53), .B2(ENABLE), .A(n21), .ZN(n85) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n21) );
  OAI21_X1 U47 ( .B1(n54), .B2(ENABLE), .A(n22), .ZN(n86) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n22) );
  OAI21_X1 U49 ( .B1(n55), .B2(ENABLE), .A(n23), .ZN(n87) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n23) );
  OAI21_X1 U51 ( .B1(n56), .B2(ENABLE), .A(n24), .ZN(n88) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n24) );
  OAI21_X1 U53 ( .B1(n57), .B2(ENABLE), .A(n25), .ZN(n89) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n25) );
  OAI21_X1 U55 ( .B1(n58), .B2(ENABLE), .A(n26), .ZN(n90) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n26) );
  OAI21_X1 U57 ( .B1(n59), .B2(ENABLE), .A(n27), .ZN(n91) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n27) );
  OAI21_X1 U59 ( .B1(n60), .B2(ENABLE), .A(n28), .ZN(n92) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n28) );
  OAI21_X1 U61 ( .B1(n61), .B2(ENABLE), .A(n29), .ZN(n93) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n29) );
  OAI21_X1 U63 ( .B1(n62), .B2(ENABLE), .A(n30), .ZN(n94) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n30) );
  OAI21_X1 U65 ( .B1(n63), .B2(ENABLE), .A(n31), .ZN(n95) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n31) );
  OAI21_X1 U67 ( .B1(n64), .B2(ENABLE), .A(n32), .ZN(n96) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n32) );
endmodule


module regFFD_NBIT32_18 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_17 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_767 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_766 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0 UIV ( .A(S), .Y(SB) );
  ND2_0 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_767 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_766 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_255 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_765 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_764 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_763 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_255 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_255 UIV ( .A(S), .Y(SB) );
  ND2_765 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_764 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_763 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_254 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_762 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_761 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_760 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_254 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_254 UIV ( .A(S), .Y(SB) );
  ND2_762 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_761 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_760 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_253 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_759 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_758 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_757 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_253 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_253 UIV ( .A(S), .Y(SB) );
  ND2_759 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_758 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_757 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_252 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_756 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_755 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_754 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_252 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_252 UIV ( .A(S), .Y(SB) );
  ND2_756 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_755 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_754 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_251 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_753 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_752 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_751 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_251 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_251 UIV ( .A(S), .Y(SB) );
  ND2_753 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_752 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_751 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_250 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_750 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_749 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_748 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_250 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_250 UIV ( .A(S), .Y(SB) );
  ND2_750 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_749 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_748 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_249 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_747 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_746 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_745 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_249 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_249 UIV ( .A(S), .Y(SB) );
  ND2_747 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_746 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_745 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_248 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_744 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_743 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_742 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_248 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_248 UIV ( .A(S), .Y(SB) );
  ND2_744 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_743 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_742 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_247 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_741 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_740 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_739 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_247 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_247 UIV ( .A(S), .Y(SB) );
  ND2_741 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_740 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_739 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_246 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_738 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_737 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_736 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_246 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_246 UIV ( .A(S), .Y(SB) );
  ND2_738 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_737 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_736 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_245 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_735 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_734 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_733 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_245 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_245 UIV ( .A(S), .Y(SB) );
  ND2_735 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_734 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_733 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_244 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_732 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_731 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_730 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_244 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_244 UIV ( .A(S), .Y(SB) );
  ND2_732 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_731 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_730 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_243 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_729 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_728 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_727 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_243 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_243 UIV ( .A(S), .Y(SB) );
  ND2_729 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_728 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_727 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_242 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_726 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_725 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_724 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_242 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_242 UIV ( .A(S), .Y(SB) );
  ND2_726 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_725 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_724 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_241 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_723 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_722 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_721 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_241 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_241 UIV ( .A(S), .Y(SB) );
  ND2_723 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_722 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_721 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_240 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_720 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_719 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_718 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_240 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_240 UIV ( .A(S), .Y(SB) );
  ND2_720 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_719 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_718 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_239 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_717 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_716 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_715 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_239 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_239 UIV ( .A(S), .Y(SB) );
  ND2_717 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_716 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_715 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_238 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_714 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_713 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_712 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_238 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_238 UIV ( .A(S), .Y(SB) );
  ND2_714 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_713 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_712 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_237 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_711 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_710 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_709 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_237 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_237 UIV ( .A(S), .Y(SB) );
  ND2_711 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_710 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_709 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_236 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_708 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_707 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_706 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_236 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_236 UIV ( .A(S), .Y(SB) );
  ND2_708 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_707 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_706 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_235 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_705 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_704 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_703 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_235 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_235 UIV ( .A(S), .Y(SB) );
  ND2_705 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_704 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_703 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_234 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_702 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_701 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_700 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_234 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_234 UIV ( .A(S), .Y(SB) );
  ND2_702 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_701 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_700 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_233 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_699 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_698 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_697 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_233 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_233 UIV ( .A(S), .Y(SB) );
  ND2_699 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_698 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_697 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_232 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_696 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_695 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_694 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_232 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_232 UIV ( .A(S), .Y(SB) );
  ND2_696 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_695 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_694 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_231 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_693 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_692 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_691 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_231 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_231 UIV ( .A(S), .Y(SB) );
  ND2_693 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_692 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_691 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_230 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_690 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_689 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_688 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_230 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_230 UIV ( .A(S), .Y(SB) );
  ND2_690 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_689 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_688 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_229 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_687 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_686 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_685 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_229 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_229 UIV ( .A(S), .Y(SB) );
  ND2_687 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_686 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_685 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_228 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_684 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_683 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_682 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_228 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_228 UIV ( .A(S), .Y(SB) );
  ND2_684 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_683 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_682 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_227 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_681 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_680 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_679 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_227 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_227 UIV ( .A(S), .Y(SB) );
  ND2_681 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_680 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_679 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_226 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_678 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_677 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_676 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_226 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_226 UIV ( .A(S), .Y(SB) );
  ND2_678 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_677 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_676 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_225 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_675 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_674 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_673 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_225 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_225 UIV ( .A(S), .Y(SB) );
  ND2_675 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_674 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_673 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_0 gen1_0 ( .A(A[0]), .B(B[0]), .S(n3), .Y(Y[0]) );
  MUX21_255 gen1_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_254 gen1_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_253 gen1_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_252 gen1_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_251 gen1_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_250 gen1_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_249 gen1_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_248 gen1_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_247 gen1_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_246 gen1_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_245 gen1_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_244 gen1_12 ( .A(A[12]), .B(B[12]), .S(n1), .Y(Y[12]) );
  MUX21_243 gen1_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_242 gen1_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_241 gen1_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_240 gen1_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_239 gen1_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_238 gen1_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_237 gen1_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_236 gen1_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_235 gen1_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_234 gen1_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_233 gen1_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_232 gen1_24 ( .A(A[24]), .B(B[24]), .S(n2), .Y(Y[24]) );
  MUX21_231 gen1_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_230 gen1_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_229 gen1_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_228 gen1_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_227 gen1_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_226 gen1_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_225 gen1_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module regFFD_NBIT32_16 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_15 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_14 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_13 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_12 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_11 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module sign_eval_N_in5_N_out32 ( IR_out, signed_val, Immediate );
  input [4:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   N0, n1;
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];
  assign Immediate[5] = N0;
  assign Immediate[6] = N0;
  assign Immediate[7] = N0;
  assign Immediate[8] = N0;
  assign Immediate[9] = N0;
  assign Immediate[10] = N0;
  assign Immediate[11] = N0;
  assign Immediate[12] = N0;
  assign Immediate[13] = N0;
  assign Immediate[14] = N0;
  assign Immediate[15] = N0;
  assign Immediate[16] = N0;
  assign Immediate[17] = N0;
  assign Immediate[18] = N0;
  assign Immediate[19] = N0;
  assign Immediate[20] = N0;
  assign Immediate[21] = N0;
  assign Immediate[22] = N0;
  assign Immediate[23] = N0;
  assign Immediate[24] = N0;
  assign Immediate[25] = N0;
  assign Immediate[26] = N0;
  assign Immediate[27] = N0;
  assign Immediate[28] = N0;
  assign Immediate[29] = N0;
  assign Immediate[30] = N0;
  assign Immediate[31] = N0;

  NOR2_X1 U1 ( .A1(signed_val), .A2(n1), .ZN(N0) );
  INV_X1 U2 ( .A(IR_out[4]), .ZN(n1) );
endmodule


module sign_eval_N_in16_N_out32 ( IR_out, signed_val, Immediate );
  input [15:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   N0, n1;
  assign Immediate[15] = IR_out[15];
  assign Immediate[14] = IR_out[14];
  assign Immediate[13] = IR_out[13];
  assign Immediate[12] = IR_out[12];
  assign Immediate[11] = IR_out[11];
  assign Immediate[10] = IR_out[10];
  assign Immediate[9] = IR_out[9];
  assign Immediate[8] = IR_out[8];
  assign Immediate[7] = IR_out[7];
  assign Immediate[6] = IR_out[6];
  assign Immediate[5] = IR_out[5];
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];
  assign Immediate[16] = N0;
  assign Immediate[17] = N0;
  assign Immediate[18] = N0;
  assign Immediate[19] = N0;
  assign Immediate[20] = N0;
  assign Immediate[21] = N0;
  assign Immediate[22] = N0;
  assign Immediate[23] = N0;
  assign Immediate[24] = N0;
  assign Immediate[25] = N0;
  assign Immediate[26] = N0;
  assign Immediate[27] = N0;
  assign Immediate[28] = N0;
  assign Immediate[29] = N0;
  assign Immediate[30] = N0;
  assign Immediate[31] = N0;

  NOR2_X1 U1 ( .A1(signed_val), .A2(n1), .ZN(N0) );
  INV_X1 U2 ( .A(IR_out[15]), .ZN(n1) );
endmodule


module sign_eval_N_in26_N_out32 ( IR_out, signed_val, Immediate );
  input [25:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   N0, n1;
  assign Immediate[25] = IR_out[25];
  assign Immediate[24] = IR_out[24];
  assign Immediate[23] = IR_out[23];
  assign Immediate[22] = IR_out[22];
  assign Immediate[21] = IR_out[21];
  assign Immediate[20] = IR_out[20];
  assign Immediate[19] = IR_out[19];
  assign Immediate[18] = IR_out[18];
  assign Immediate[17] = IR_out[17];
  assign Immediate[16] = IR_out[16];
  assign Immediate[15] = IR_out[15];
  assign Immediate[14] = IR_out[14];
  assign Immediate[13] = IR_out[13];
  assign Immediate[12] = IR_out[12];
  assign Immediate[11] = IR_out[11];
  assign Immediate[10] = IR_out[10];
  assign Immediate[9] = IR_out[9];
  assign Immediate[8] = IR_out[8];
  assign Immediate[7] = IR_out[7];
  assign Immediate[6] = IR_out[6];
  assign Immediate[5] = IR_out[5];
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];
  assign Immediate[26] = N0;
  assign Immediate[27] = N0;
  assign Immediate[28] = N0;
  assign Immediate[29] = N0;
  assign Immediate[30] = N0;
  assign Immediate[31] = N0;

  NOR2_X1 U1 ( .A1(signed_val), .A2(n1), .ZN(N0) );
  INV_X1 U2 ( .A(IR_out[25]), .ZN(n1) );
endmodule


module IR_DECODE_NBIT32_opBIT6_regBIT5 ( CLK, IR_26, OPCODE, is_signed, RS1, 
        RS2, RD, IMMEDIATE );
  input [25:0] IR_26;
  input [5:0] OPCODE;
  output [4:0] RS1;
  output [4:0] RS2;
  output [4:0] RD;
  output [31:0] IMMEDIATE;
  input CLK, is_signed;
  wire   N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, net105089, net137935, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23;
  wire   [31:0] IMMEDIATE_16;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;
  assign N133 = IR_26[21];
  assign N134 = IR_26[22];
  assign N135 = IR_26[23];
  assign N136 = IR_26[24];
  assign N137 = IR_26[25];
  assign N138 = IR_26[16];
  assign N139 = IR_26[17];
  assign N140 = IR_26[18];
  assign N141 = IR_26[19];
  assign N142 = IR_26[20];

  DLH_X1 \RD_reg[4]  ( .G(CLK), .D(N147), .Q(RD[4]) );
  DLH_X1 \RD_reg[3]  ( .G(CLK), .D(N146), .Q(RD[3]) );
  DLH_X1 \RD_reg[2]  ( .G(CLK), .D(N145), .Q(RD[2]) );
  DLH_X1 \RD_reg[1]  ( .G(CLK), .D(N144), .Q(RD[1]) );
  DLH_X1 \RD_reg[0]  ( .G(CLK), .D(N143), .Q(RD[0]) );
  DLH_X1 \IMMEDIATE_reg[31]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[31]) );
  DLH_X1 \IMMEDIATE_reg[30]  ( .G(CLK), .D(n23), .Q(IMMEDIATE[30]) );
  DLH_X1 \IMMEDIATE_reg[29]  ( .G(CLK), .D(n23), .Q(IMMEDIATE[29]) );
  DLH_X1 \IMMEDIATE_reg[28]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[28]) );
  DLH_X1 \IMMEDIATE_reg[27]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[27]) );
  DLH_X1 \IMMEDIATE_reg[26]  ( .G(CLK), .D(n23), .Q(IMMEDIATE[26]) );
  DLH_X1 \IMMEDIATE_reg[25]  ( .G(CLK), .D(n23), .Q(IMMEDIATE[25]) );
  DLH_X1 \IMMEDIATE_reg[24]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[24]) );
  DLH_X1 \IMMEDIATE_reg[23]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[23]) );
  DLH_X1 \IMMEDIATE_reg[22]  ( .G(CLK), .D(n23), .Q(IMMEDIATE[22]) );
  DLH_X1 \IMMEDIATE_reg[21]  ( .G(CLK), .D(n23), .Q(IMMEDIATE[21]) );
  DLH_X1 \IMMEDIATE_reg[20]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[20]) );
  DLH_X1 \IMMEDIATE_reg[19]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[19]) );
  DLH_X1 \IMMEDIATE_reg[18]  ( .G(CLK), .D(n23), .Q(IMMEDIATE[18]) );
  DLH_X1 \IMMEDIATE_reg[17]  ( .G(CLK), .D(n23), .Q(IMMEDIATE[17]) );
  DLH_X1 \IMMEDIATE_reg[16]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[16]) );
  DLH_X1 \IMMEDIATE_reg[15]  ( .G(CLK), .D(n22), .Q(IMMEDIATE[15]) );
  DLH_X1 \IMMEDIATE_reg[14]  ( .G(CLK), .D(n21), .Q(IMMEDIATE[14]) );
  DLH_X1 \IMMEDIATE_reg[13]  ( .G(CLK), .D(n20), .Q(IMMEDIATE[13]) );
  DLH_X1 \IMMEDIATE_reg[12]  ( .G(CLK), .D(net105089), .Q(IMMEDIATE[12]) );
  DLH_X1 \IMMEDIATE_reg[11]  ( .G(CLK), .D(n19), .Q(IMMEDIATE[11]) );
  DLH_X1 \IMMEDIATE_reg[10]  ( .G(CLK), .D(n18), .Q(IMMEDIATE[10]) );
  DLH_X1 \IMMEDIATE_reg[9]  ( .G(CLK), .D(n17), .Q(IMMEDIATE[9]) );
  DLH_X1 \IMMEDIATE_reg[8]  ( .G(CLK), .D(n16), .Q(IMMEDIATE[8]) );
  DLH_X1 \IMMEDIATE_reg[7]  ( .G(CLK), .D(n15), .Q(IMMEDIATE[7]) );
  DLH_X1 \IMMEDIATE_reg[6]  ( .G(CLK), .D(n14), .Q(IMMEDIATE[6]) );
  DLH_X1 \IMMEDIATE_reg[5]  ( .G(CLK), .D(n13), .Q(IMMEDIATE[5]) );
  DLH_X1 \IMMEDIATE_reg[4]  ( .G(CLK), .D(n12), .Q(IMMEDIATE[4]) );
  DLH_X1 \IMMEDIATE_reg[3]  ( .G(CLK), .D(n11), .Q(IMMEDIATE[3]) );
  DLH_X1 \IMMEDIATE_reg[2]  ( .G(CLK), .D(n10), .Q(IMMEDIATE[2]) );
  DLH_X1 \IMMEDIATE_reg[1]  ( .G(CLK), .D(n9), .Q(IMMEDIATE[1]) );
  DLH_X1 \IMMEDIATE_reg[0]  ( .G(CLK), .D(n8), .Q(IMMEDIATE[0]) );
  DLH_X1 \RS1_reg[4]  ( .G(CLK), .D(N137), .Q(RS1[4]) );
  DLH_X1 \RS1_reg[3]  ( .G(CLK), .D(N136), .Q(RS1[3]) );
  DLH_X1 \RS1_reg[2]  ( .G(CLK), .D(N135), .Q(RS1[2]) );
  DLH_X1 \RS1_reg[1]  ( .G(CLK), .D(N134), .Q(RS1[1]) );
  DLH_X1 \RS1_reg[0]  ( .G(CLK), .D(N133), .Q(RS1[0]) );
  DLH_X1 \RS2_reg[4]  ( .G(CLK), .D(N142), .Q(RS2[4]) );
  DLH_X1 \RS2_reg[3]  ( .G(CLK), .D(N141), .Q(RS2[3]) );
  DLH_X1 \RS2_reg[2]  ( .G(CLK), .D(N140), .Q(RS2[2]) );
  DLH_X1 \RS2_reg[1]  ( .G(CLK), .D(N139), .Q(RS2[1]) );
  DLH_X1 \RS2_reg[0]  ( .G(CLK), .D(N138), .Q(RS2[0]) );
  sign_eval_N_in5_N_out32 SIGN_EXTENSION_imm5 ( .IR_out(IR_26[15:11]), 
        .signed_val(is_signed) );
  sign_eval_N_in16_N_out32 SIGN_EXTENSION_imm16 ( .IR_out(IR_26[15:0]), 
        .signed_val(is_signed), .Immediate({IMMEDIATE_16[31], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, IMMEDIATE_16[15:0]}) );
  sign_eval_N_in26_N_out32 SIGN_EXTENSION_imm26 ( .IR_out({N137, N136, N135, 
        N134, N133, N142, N141, N140, N139, N138, IR_26[15:0]}), .signed_val(
        1'b0) );
  NOR2_X1 U3 ( .A1(n1), .A2(n5), .ZN(net105089) );
  INV_X1 U4 ( .A(IMMEDIATE_16[12]), .ZN(n5) );
  AND2_X1 U5 ( .A1(n3), .A2(n2), .ZN(n1) );
  NOR3_X1 U6 ( .A1(OPCODE[2]), .A2(OPCODE[1]), .A3(OPCODE[0]), .ZN(n2) );
  NOR3_X1 U7 ( .A1(OPCODE[2]), .A2(OPCODE[1]), .A3(OPCODE[0]), .ZN(n4) );
  MUX2_X1 U8 ( .A(N141), .B(IR_26[14]), .S(n1), .Z(N146) );
  MUX2_X1 U9 ( .A(N138), .B(IR_26[11]), .S(n1), .Z(N143) );
  NOR3_X2 U10 ( .A1(OPCODE[5]), .A2(OPCODE[4]), .A3(OPCODE[3]), .ZN(n3) );
  NAND2_X1 U11 ( .A1(n3), .A2(n4), .ZN(net137935) );
  NAND2_X1 U12 ( .A1(n3), .A2(n4), .ZN(n6) );
  AND2_X1 U13 ( .A1(IMMEDIATE_16[31]), .A2(net137935), .ZN(n7) );
  AND2_X1 U14 ( .A1(IMMEDIATE_16[0]), .A2(n6), .ZN(n8) );
  AND2_X1 U15 ( .A1(IMMEDIATE_16[1]), .A2(n6), .ZN(n9) );
  AND2_X1 U16 ( .A1(IMMEDIATE_16[2]), .A2(net137935), .ZN(n10) );
  AND2_X1 U17 ( .A1(IMMEDIATE_16[3]), .A2(net137935), .ZN(n11) );
  AND2_X1 U18 ( .A1(IMMEDIATE_16[4]), .A2(n6), .ZN(n12) );
  AND2_X1 U19 ( .A1(IMMEDIATE_16[5]), .A2(n6), .ZN(n13) );
  AND2_X1 U20 ( .A1(IMMEDIATE_16[6]), .A2(n6), .ZN(n14) );
  AND2_X1 U21 ( .A1(IMMEDIATE_16[7]), .A2(n6), .ZN(n15) );
  AND2_X1 U22 ( .A1(IMMEDIATE_16[8]), .A2(net137935), .ZN(n16) );
  AND2_X1 U23 ( .A1(IMMEDIATE_16[9]), .A2(net137935), .ZN(n17) );
  AND2_X1 U24 ( .A1(IMMEDIATE_16[10]), .A2(net137935), .ZN(n18) );
  AND2_X1 U25 ( .A1(IMMEDIATE_16[11]), .A2(n6), .ZN(n19) );
  AND2_X1 U26 ( .A1(IMMEDIATE_16[13]), .A2(net137935), .ZN(n20) );
  AND2_X1 U27 ( .A1(IMMEDIATE_16[14]), .A2(n6), .ZN(n21) );
  AND2_X1 U28 ( .A1(IMMEDIATE_16[15]), .A2(n6), .ZN(n22) );
  AND2_X1 U29 ( .A1(IMMEDIATE_16[31]), .A2(net137935), .ZN(n23) );
  MUX2_X1 U30 ( .A(IR_26[15]), .B(N142), .S(n6), .Z(N147) );
  MUX2_X1 U31 ( .A(IR_26[13]), .B(N140), .S(net137935), .Z(N145) );
  MUX2_X1 U32 ( .A(IR_26[12]), .B(N139), .S(n6), .Z(N144) );
endmodule


module windRF_M8_N8_F5_NBIT32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n4, n5;
  wire   [6:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n4), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(A[5]), .B(carry[5]), .Z(SUM[5]) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XNOR2_X1 U3 ( .A(A[6]), .B(n5), .ZN(SUM[6]) );
  NAND2_X1 U4 ( .A1(A[5]), .A2(carry[5]), .ZN(n5) );
  AND2_X1 U5 ( .A1(B[0]), .A2(A[0]), .ZN(n4) );
endmodule


module windRF_M8_N8_F5_NBIT32_DW01_add_3 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n4, n5;
  wire   [6:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n4), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(A[5]), .B(carry[5]), .Z(SUM[5]) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XNOR2_X1 U3 ( .A(A[6]), .B(n5), .ZN(SUM[6]) );
  NAND2_X1 U4 ( .A1(A[5]), .A2(carry[5]), .ZN(n5) );
  AND2_X1 U5 ( .A1(B[0]), .A2(A[0]), .ZN(n4) );
endmodule


module windRF_M8_N8_F5_NBIT32_DW01_add_5 ( A, B, CI, SUM, CO );
  input [6:0] A;
  input [6:0] B;
  output [6:0] SUM;
  input CI;
  output CO;
  wire   n4, n5;
  wire   [6:1] carry;

  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n4), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XNOR2_X1 U2 ( .A(A[6]), .B(n5), .ZN(SUM[6]) );
  XOR2_X1 U3 ( .A(A[5]), .B(carry[5]), .Z(SUM[5]) );
  NAND2_X1 U4 ( .A1(A[5]), .A2(carry[5]), .ZN(n5) );
  AND2_X1 U5 ( .A1(B[0]), .A2(A[0]), .ZN(n4) );
endmodule


module windRF_M8_N8_F5_NBIT32 ( CLK, RESET, ENABLE, CALL, RETRN, FILL, SPILL, 
        BUSin, BUSout, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, 
        OUT2, wr_signal );
  input [31:0] BUSin;
  output [31:0] BUSout;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, CALL, RETRN, RD1, RD2, WR, wr_signal;
  output FILL, SPILL;
  wire   \REGISTERS[11][31] , \REGISTERS[11][30] , \REGISTERS[11][29] ,
         \REGISTERS[11][28] , \REGISTERS[11][27] , \REGISTERS[11][26] ,
         \REGISTERS[11][25] , \REGISTERS[11][24] , \REGISTERS[11][23] ,
         \REGISTERS[11][22] , \REGISTERS[11][21] , \REGISTERS[11][20] ,
         \REGISTERS[11][19] , \REGISTERS[11][18] , \REGISTERS[11][17] ,
         \REGISTERS[11][16] , \REGISTERS[11][15] , \REGISTERS[11][14] ,
         \REGISTERS[11][13] , \REGISTERS[11][12] , \REGISTERS[11][11] ,
         \REGISTERS[11][10] , \REGISTERS[11][9] , \REGISTERS[11][8] ,
         \REGISTERS[11][7] , \REGISTERS[11][6] , \REGISTERS[11][5] ,
         \REGISTERS[11][4] , \REGISTERS[11][3] , \REGISTERS[11][2] ,
         \REGISTERS[11][1] , \REGISTERS[11][0] , \REGISTERS[12][31] ,
         \REGISTERS[12][30] , \REGISTERS[12][29] , \REGISTERS[12][28] ,
         \REGISTERS[12][27] , \REGISTERS[12][26] , \REGISTERS[12][25] ,
         \REGISTERS[12][24] , \REGISTERS[12][23] , \REGISTERS[12][22] ,
         \REGISTERS[12][21] , \REGISTERS[12][20] , \REGISTERS[12][19] ,
         \REGISTERS[12][18] , \REGISTERS[12][17] , \REGISTERS[12][16] ,
         \REGISTERS[12][15] , \REGISTERS[12][14] , \REGISTERS[12][13] ,
         \REGISTERS[12][12] , \REGISTERS[12][11] , \REGISTERS[12][10] ,
         \REGISTERS[12][9] , \REGISTERS[12][8] , \REGISTERS[12][7] ,
         \REGISTERS[12][6] , \REGISTERS[12][5] , \REGISTERS[12][4] ,
         \REGISTERS[12][3] , \REGISTERS[12][2] , \REGISTERS[12][1] ,
         \REGISTERS[12][0] , \REGISTERS[16][31] , \REGISTERS[16][30] ,
         \REGISTERS[16][29] , \REGISTERS[16][28] , \REGISTERS[16][27] ,
         \REGISTERS[16][26] , \REGISTERS[16][25] , \REGISTERS[16][24] ,
         \REGISTERS[16][23] , \REGISTERS[16][22] , \REGISTERS[16][21] ,
         \REGISTERS[16][20] , \REGISTERS[16][19] , \REGISTERS[16][18] ,
         \REGISTERS[16][17] , \REGISTERS[16][16] , \REGISTERS[16][15] ,
         \REGISTERS[16][14] , \REGISTERS[16][13] , \REGISTERS[16][12] ,
         \REGISTERS[16][11] , \REGISTERS[16][10] , \REGISTERS[16][9] ,
         \REGISTERS[16][8] , \REGISTERS[16][7] , \REGISTERS[16][6] ,
         \REGISTERS[16][5] , \REGISTERS[16][4] , \REGISTERS[16][3] ,
         \REGISTERS[16][2] , \REGISTERS[16][1] , \REGISTERS[16][0] ,
         \REGISTERS[17][31] , \REGISTERS[17][30] , \REGISTERS[17][29] ,
         \REGISTERS[17][28] , \REGISTERS[17][27] , \REGISTERS[17][26] ,
         \REGISTERS[17][25] , \REGISTERS[17][24] , \REGISTERS[17][23] ,
         \REGISTERS[17][22] , \REGISTERS[17][21] , \REGISTERS[17][20] ,
         \REGISTERS[17][19] , \REGISTERS[17][18] , \REGISTERS[17][17] ,
         \REGISTERS[17][16] , \REGISTERS[17][15] , \REGISTERS[17][14] ,
         \REGISTERS[17][13] , \REGISTERS[17][12] , \REGISTERS[17][11] ,
         \REGISTERS[17][10] , \REGISTERS[17][9] , \REGISTERS[17][8] ,
         \REGISTERS[17][7] , \REGISTERS[17][6] , \REGISTERS[17][5] ,
         \REGISTERS[17][4] , \REGISTERS[17][3] , \REGISTERS[17][2] ,
         \REGISTERS[17][1] , \REGISTERS[17][0] , \REGISTERS[18][31] ,
         \REGISTERS[18][30] , \REGISTERS[18][29] , \REGISTERS[18][28] ,
         \REGISTERS[18][27] , \REGISTERS[18][26] , \REGISTERS[18][25] ,
         \REGISTERS[18][24] , \REGISTERS[18][23] , \REGISTERS[18][22] ,
         \REGISTERS[18][21] , \REGISTERS[18][20] , \REGISTERS[18][19] ,
         \REGISTERS[18][18] , \REGISTERS[18][17] , \REGISTERS[18][16] ,
         \REGISTERS[18][15] , \REGISTERS[18][14] , \REGISTERS[18][13] ,
         \REGISTERS[18][12] , \REGISTERS[18][11] , \REGISTERS[18][10] ,
         \REGISTERS[18][9] , \REGISTERS[18][8] , \REGISTERS[18][7] ,
         \REGISTERS[18][6] , \REGISTERS[18][5] , \REGISTERS[18][4] ,
         \REGISTERS[18][3] , \REGISTERS[18][2] , \REGISTERS[18][1] ,
         \REGISTERS[18][0] , \REGISTERS[19][31] , \REGISTERS[19][30] ,
         \REGISTERS[19][29] , \REGISTERS[19][28] , \REGISTERS[19][27] ,
         \REGISTERS[19][26] , \REGISTERS[19][25] , \REGISTERS[19][24] ,
         \REGISTERS[19][23] , \REGISTERS[19][22] , \REGISTERS[19][21] ,
         \REGISTERS[19][20] , \REGISTERS[19][19] , \REGISTERS[19][18] ,
         \REGISTERS[19][17] , \REGISTERS[19][16] , \REGISTERS[19][15] ,
         \REGISTERS[19][14] , \REGISTERS[19][13] , \REGISTERS[19][12] ,
         \REGISTERS[19][11] , \REGISTERS[19][10] , \REGISTERS[19][9] ,
         \REGISTERS[19][8] , \REGISTERS[19][7] , \REGISTERS[19][6] ,
         \REGISTERS[19][5] , \REGISTERS[19][4] , \REGISTERS[19][3] ,
         \REGISTERS[19][2] , \REGISTERS[19][1] , \REGISTERS[19][0] ,
         \REGISTERS[20][31] , \REGISTERS[20][30] , \REGISTERS[20][29] ,
         \REGISTERS[20][28] , \REGISTERS[20][27] , \REGISTERS[20][26] ,
         \REGISTERS[20][25] , \REGISTERS[20][24] , \REGISTERS[20][23] ,
         \REGISTERS[20][22] , \REGISTERS[20][21] , \REGISTERS[20][20] ,
         \REGISTERS[20][19] , \REGISTERS[20][18] , \REGISTERS[20][17] ,
         \REGISTERS[20][16] , \REGISTERS[20][15] , \REGISTERS[20][14] ,
         \REGISTERS[20][13] , \REGISTERS[20][12] , \REGISTERS[20][11] ,
         \REGISTERS[20][10] , \REGISTERS[20][9] , \REGISTERS[20][8] ,
         \REGISTERS[20][7] , \REGISTERS[20][6] , \REGISTERS[20][5] ,
         \REGISTERS[20][4] , \REGISTERS[20][3] , \REGISTERS[20][2] ,
         \REGISTERS[20][1] , \REGISTERS[20][0] , \REGISTERS[21][31] ,
         \REGISTERS[21][30] , \REGISTERS[21][29] , \REGISTERS[21][28] ,
         \REGISTERS[21][27] , \REGISTERS[21][26] , \REGISTERS[21][25] ,
         \REGISTERS[21][24] , \REGISTERS[21][23] , \REGISTERS[21][22] ,
         \REGISTERS[21][21] , \REGISTERS[21][20] , \REGISTERS[21][19] ,
         \REGISTERS[21][18] , \REGISTERS[21][17] , \REGISTERS[21][16] ,
         \REGISTERS[21][15] , \REGISTERS[21][14] , \REGISTERS[21][13] ,
         \REGISTERS[21][12] , \REGISTERS[21][11] , \REGISTERS[21][10] ,
         \REGISTERS[21][9] , \REGISTERS[21][8] , \REGISTERS[21][7] ,
         \REGISTERS[21][6] , \REGISTERS[21][5] , \REGISTERS[21][4] ,
         \REGISTERS[21][3] , \REGISTERS[21][2] , \REGISTERS[21][1] ,
         \REGISTERS[21][0] , \REGISTERS[33][31] , \REGISTERS[33][30] ,
         \REGISTERS[33][29] , \REGISTERS[33][28] , \REGISTERS[33][27] ,
         \REGISTERS[33][26] , \REGISTERS[33][25] , \REGISTERS[33][24] ,
         \REGISTERS[33][23] , \REGISTERS[33][22] , \REGISTERS[33][21] ,
         \REGISTERS[33][20] , \REGISTERS[33][19] , \REGISTERS[33][18] ,
         \REGISTERS[33][17] , \REGISTERS[33][16] , \REGISTERS[33][15] ,
         \REGISTERS[33][14] , \REGISTERS[33][13] , \REGISTERS[33][12] ,
         \REGISTERS[33][11] , \REGISTERS[33][10] , \REGISTERS[33][9] ,
         \REGISTERS[33][8] , \REGISTERS[33][7] , \REGISTERS[33][6] ,
         \REGISTERS[33][5] , \REGISTERS[33][4] , \REGISTERS[33][3] ,
         \REGISTERS[33][2] , \REGISTERS[33][1] , \REGISTERS[33][0] ,
         \REGISTERS[34][31] , \REGISTERS[34][30] , \REGISTERS[34][29] ,
         \REGISTERS[34][28] , \REGISTERS[34][27] , \REGISTERS[34][26] ,
         \REGISTERS[34][25] , \REGISTERS[34][24] , \REGISTERS[34][23] ,
         \REGISTERS[34][22] , \REGISTERS[34][21] , \REGISTERS[34][20] ,
         \REGISTERS[34][19] , \REGISTERS[34][18] , \REGISTERS[34][17] ,
         \REGISTERS[34][16] , \REGISTERS[34][15] , \REGISTERS[34][14] ,
         \REGISTERS[34][13] , \REGISTERS[34][12] , \REGISTERS[34][11] ,
         \REGISTERS[34][10] , \REGISTERS[34][9] , \REGISTERS[34][8] ,
         \REGISTERS[34][7] , \REGISTERS[34][6] , \REGISTERS[34][5] ,
         \REGISTERS[34][4] , \REGISTERS[34][3] , \REGISTERS[34][2] ,
         \REGISTERS[34][1] , \REGISTERS[34][0] , \REGISTERS[38][31] ,
         \REGISTERS[38][30] , \REGISTERS[38][29] , \REGISTERS[38][28] ,
         \REGISTERS[38][27] , \REGISTERS[38][26] , \REGISTERS[38][25] ,
         \REGISTERS[38][24] , \REGISTERS[38][23] , \REGISTERS[38][22] ,
         \REGISTERS[38][21] , \REGISTERS[38][20] , \REGISTERS[38][19] ,
         \REGISTERS[38][18] , \REGISTERS[38][17] , \REGISTERS[38][16] ,
         \REGISTERS[38][15] , \REGISTERS[38][14] , \REGISTERS[38][13] ,
         \REGISTERS[38][12] , \REGISTERS[38][11] , \REGISTERS[38][10] ,
         \REGISTERS[38][9] , \REGISTERS[38][8] , \REGISTERS[38][7] ,
         \REGISTERS[38][6] , \REGISTERS[38][5] , \REGISTERS[38][4] ,
         \REGISTERS[38][3] , \REGISTERS[38][2] , \REGISTERS[38][1] ,
         \REGISTERS[38][0] , \REGISTERS[39][31] , \REGISTERS[39][30] ,
         \REGISTERS[39][29] , \REGISTERS[39][28] , \REGISTERS[39][27] ,
         \REGISTERS[39][26] , \REGISTERS[39][25] , \REGISTERS[39][24] ,
         \REGISTERS[39][23] , \REGISTERS[39][22] , \REGISTERS[39][21] ,
         \REGISTERS[39][20] , \REGISTERS[39][19] , \REGISTERS[39][18] ,
         \REGISTERS[39][17] , \REGISTERS[39][16] , \REGISTERS[39][15] ,
         \REGISTERS[39][14] , \REGISTERS[39][13] , \REGISTERS[39][12] ,
         \REGISTERS[39][11] , \REGISTERS[39][10] , \REGISTERS[39][9] ,
         \REGISTERS[39][8] , \REGISTERS[39][7] , \REGISTERS[39][6] ,
         \REGISTERS[39][5] , \REGISTERS[39][4] , \REGISTERS[39][3] ,
         \REGISTERS[39][2] , \REGISTERS[39][1] , \REGISTERS[39][0] ,
         \REGISTERS[40][31] , \REGISTERS[40][30] , \REGISTERS[40][29] ,
         \REGISTERS[40][28] , \REGISTERS[40][27] , \REGISTERS[40][26] ,
         \REGISTERS[40][25] , \REGISTERS[40][24] , \REGISTERS[40][23] ,
         \REGISTERS[40][22] , \REGISTERS[40][21] , \REGISTERS[40][20] ,
         \REGISTERS[40][19] , \REGISTERS[40][18] , \REGISTERS[40][17] ,
         \REGISTERS[40][16] , \REGISTERS[40][15] , \REGISTERS[40][14] ,
         \REGISTERS[40][13] , \REGISTERS[40][12] , \REGISTERS[40][11] ,
         \REGISTERS[40][10] , \REGISTERS[40][9] , \REGISTERS[40][8] ,
         \REGISTERS[40][7] , \REGISTERS[40][6] , \REGISTERS[40][5] ,
         \REGISTERS[40][4] , \REGISTERS[40][3] , \REGISTERS[40][2] ,
         \REGISTERS[40][1] , \REGISTERS[40][0] , \REGISTERS[41][31] ,
         \REGISTERS[41][30] , \REGISTERS[41][29] , \REGISTERS[41][28] ,
         \REGISTERS[41][27] , \REGISTERS[41][26] , \REGISTERS[41][25] ,
         \REGISTERS[41][24] , \REGISTERS[41][23] , \REGISTERS[41][22] ,
         \REGISTERS[41][21] , \REGISTERS[41][20] , \REGISTERS[41][19] ,
         \REGISTERS[41][18] , \REGISTERS[41][17] , \REGISTERS[41][16] ,
         \REGISTERS[41][15] , \REGISTERS[41][14] , \REGISTERS[41][13] ,
         \REGISTERS[41][12] , \REGISTERS[41][11] , \REGISTERS[41][10] ,
         \REGISTERS[41][9] , \REGISTERS[41][8] , \REGISTERS[41][7] ,
         \REGISTERS[41][6] , \REGISTERS[41][5] , \REGISTERS[41][4] ,
         \REGISTERS[41][3] , \REGISTERS[41][2] , \REGISTERS[41][1] ,
         \REGISTERS[41][0] , \REGISTERS[42][31] , \REGISTERS[42][30] ,
         \REGISTERS[42][29] , \REGISTERS[42][28] , \REGISTERS[42][27] ,
         \REGISTERS[42][26] , \REGISTERS[42][25] , \REGISTERS[42][24] ,
         \REGISTERS[42][23] , \REGISTERS[42][22] , \REGISTERS[42][21] ,
         \REGISTERS[42][20] , \REGISTERS[42][19] , \REGISTERS[42][18] ,
         \REGISTERS[42][17] , \REGISTERS[42][16] , \REGISTERS[42][15] ,
         \REGISTERS[42][14] , \REGISTERS[42][13] , \REGISTERS[42][12] ,
         \REGISTERS[42][11] , \REGISTERS[42][10] , \REGISTERS[42][9] ,
         \REGISTERS[42][8] , \REGISTERS[42][7] , \REGISTERS[42][6] ,
         \REGISTERS[42][5] , \REGISTERS[42][4] , \REGISTERS[42][3] ,
         \REGISTERS[42][2] , \REGISTERS[42][1] , \REGISTERS[42][0] ,
         \REGISTERS[43][31] , \REGISTERS[43][30] , \REGISTERS[43][29] ,
         \REGISTERS[43][28] , \REGISTERS[43][27] , \REGISTERS[43][26] ,
         \REGISTERS[43][25] , \REGISTERS[43][24] , \REGISTERS[43][23] ,
         \REGISTERS[43][22] , \REGISTERS[43][21] , \REGISTERS[43][20] ,
         \REGISTERS[43][19] , \REGISTERS[43][18] , \REGISTERS[43][17] ,
         \REGISTERS[43][16] , \REGISTERS[43][15] , \REGISTERS[43][14] ,
         \REGISTERS[43][13] , \REGISTERS[43][12] , \REGISTERS[43][11] ,
         \REGISTERS[43][10] , \REGISTERS[43][9] , \REGISTERS[43][8] ,
         \REGISTERS[43][7] , \REGISTERS[43][6] , \REGISTERS[43][5] ,
         \REGISTERS[43][4] , \REGISTERS[43][3] , \REGISTERS[43][2] ,
         \REGISTERS[43][1] , \REGISTERS[43][0] , \REGISTERS[44][31] ,
         \REGISTERS[44][30] , \REGISTERS[44][29] , \REGISTERS[44][28] ,
         \REGISTERS[44][27] , \REGISTERS[44][26] , \REGISTERS[44][25] ,
         \REGISTERS[44][24] , \REGISTERS[44][23] , \REGISTERS[44][22] ,
         \REGISTERS[44][21] , \REGISTERS[44][20] , \REGISTERS[44][19] ,
         \REGISTERS[44][18] , \REGISTERS[44][17] , \REGISTERS[44][16] ,
         \REGISTERS[44][15] , \REGISTERS[44][14] , \REGISTERS[44][13] ,
         \REGISTERS[44][12] , \REGISTERS[44][11] , \REGISTERS[44][10] ,
         \REGISTERS[44][9] , \REGISTERS[44][8] , \REGISTERS[44][7] ,
         \REGISTERS[44][6] , \REGISTERS[44][5] , \REGISTERS[44][4] ,
         \REGISTERS[44][3] , \REGISTERS[44][2] , \REGISTERS[44][1] ,
         \REGISTERS[44][0] , \REGISTERS[45][31] , \REGISTERS[45][30] ,
         \REGISTERS[45][29] , \REGISTERS[45][28] , \REGISTERS[45][27] ,
         \REGISTERS[45][26] , \REGISTERS[45][25] , \REGISTERS[45][24] ,
         \REGISTERS[45][23] , \REGISTERS[45][22] , \REGISTERS[45][21] ,
         \REGISTERS[45][20] , \REGISTERS[45][19] , \REGISTERS[45][18] ,
         \REGISTERS[45][17] , \REGISTERS[45][16] , \REGISTERS[45][15] ,
         \REGISTERS[45][14] , \REGISTERS[45][13] , \REGISTERS[45][12] ,
         \REGISTERS[45][11] , \REGISTERS[45][10] , \REGISTERS[45][9] ,
         \REGISTERS[45][8] , \REGISTERS[45][7] , \REGISTERS[45][6] ,
         \REGISTERS[45][5] , \REGISTERS[45][4] , \REGISTERS[45][3] ,
         \REGISTERS[45][2] , \REGISTERS[45][1] , \REGISTERS[45][0] ,
         \REGISTERS[49][31] , \REGISTERS[49][30] , \REGISTERS[49][29] ,
         \REGISTERS[49][28] , \REGISTERS[49][27] , \REGISTERS[49][26] ,
         \REGISTERS[49][25] , \REGISTERS[49][24] , \REGISTERS[49][23] ,
         \REGISTERS[49][22] , \REGISTERS[49][21] , \REGISTERS[49][20] ,
         \REGISTERS[49][19] , \REGISTERS[49][18] , \REGISTERS[49][17] ,
         \REGISTERS[49][16] , \REGISTERS[49][15] , \REGISTERS[49][14] ,
         \REGISTERS[49][13] , \REGISTERS[49][12] , \REGISTERS[49][11] ,
         \REGISTERS[49][10] , \REGISTERS[49][9] , \REGISTERS[49][8] ,
         \REGISTERS[49][7] , \REGISTERS[49][6] , \REGISTERS[49][5] ,
         \REGISTERS[49][4] , \REGISTERS[49][3] , \REGISTERS[49][2] ,
         \REGISTERS[49][1] , \REGISTERS[49][0] , \REGISTERS[50][31] ,
         \REGISTERS[50][30] , \REGISTERS[50][29] , \REGISTERS[50][28] ,
         \REGISTERS[50][27] , \REGISTERS[50][26] , \REGISTERS[50][25] ,
         \REGISTERS[50][24] , \REGISTERS[50][23] , \REGISTERS[50][22] ,
         \REGISTERS[50][21] , \REGISTERS[50][20] , \REGISTERS[50][19] ,
         \REGISTERS[50][18] , \REGISTERS[50][17] , \REGISTERS[50][16] ,
         \REGISTERS[50][15] , \REGISTERS[50][14] , \REGISTERS[50][13] ,
         \REGISTERS[50][12] , \REGISTERS[50][11] , \REGISTERS[50][10] ,
         \REGISTERS[50][9] , \REGISTERS[50][8] , \REGISTERS[50][7] ,
         \REGISTERS[50][6] , \REGISTERS[50][5] , \REGISTERS[50][4] ,
         \REGISTERS[50][3] , \REGISTERS[50][2] , \REGISTERS[50][1] ,
         \REGISTERS[50][0] , \REGISTERS[51][31] , \REGISTERS[51][30] ,
         \REGISTERS[51][29] , \REGISTERS[51][28] , \REGISTERS[51][27] ,
         \REGISTERS[51][26] , \REGISTERS[51][25] , \REGISTERS[51][24] ,
         \REGISTERS[51][23] , \REGISTERS[51][22] , \REGISTERS[51][21] ,
         \REGISTERS[51][20] , \REGISTERS[51][19] , \REGISTERS[51][18] ,
         \REGISTERS[51][17] , \REGISTERS[51][16] , \REGISTERS[51][15] ,
         \REGISTERS[51][14] , \REGISTERS[51][13] , \REGISTERS[51][12] ,
         \REGISTERS[51][11] , \REGISTERS[51][10] , \REGISTERS[51][9] ,
         \REGISTERS[51][8] , \REGISTERS[51][7] , \REGISTERS[51][6] ,
         \REGISTERS[51][5] , \REGISTERS[51][4] , \REGISTERS[51][3] ,
         \REGISTERS[51][2] , \REGISTERS[51][1] , \REGISTERS[51][0] ,
         \REGISTERS[52][31] , \REGISTERS[52][30] , \REGISTERS[52][29] ,
         \REGISTERS[52][28] , \REGISTERS[52][27] , \REGISTERS[52][26] ,
         \REGISTERS[52][25] , \REGISTERS[52][24] , \REGISTERS[52][23] ,
         \REGISTERS[52][22] , \REGISTERS[52][21] , \REGISTERS[52][20] ,
         \REGISTERS[52][19] , \REGISTERS[52][18] , \REGISTERS[52][17] ,
         \REGISTERS[52][16] , \REGISTERS[52][15] , \REGISTERS[52][14] ,
         \REGISTERS[52][13] , \REGISTERS[52][12] , \REGISTERS[52][11] ,
         \REGISTERS[52][10] , \REGISTERS[52][9] , \REGISTERS[52][8] ,
         \REGISTERS[52][7] , \REGISTERS[52][6] , \REGISTERS[52][5] ,
         \REGISTERS[52][4] , \REGISTERS[52][3] , \REGISTERS[52][2] ,
         \REGISTERS[52][1] , \REGISTERS[52][0] , \REGISTERS[53][31] ,
         \REGISTERS[53][30] , \REGISTERS[53][29] , \REGISTERS[53][28] ,
         \REGISTERS[53][27] , \REGISTERS[53][26] , \REGISTERS[53][25] ,
         \REGISTERS[53][24] , \REGISTERS[53][23] , \REGISTERS[53][22] ,
         \REGISTERS[53][21] , \REGISTERS[53][20] , \REGISTERS[53][19] ,
         \REGISTERS[53][18] , \REGISTERS[53][17] , \REGISTERS[53][16] ,
         \REGISTERS[53][15] , \REGISTERS[53][14] , \REGISTERS[53][13] ,
         \REGISTERS[53][12] , \REGISTERS[53][11] , \REGISTERS[53][10] ,
         \REGISTERS[53][9] , \REGISTERS[53][8] , \REGISTERS[53][7] ,
         \REGISTERS[53][6] , \REGISTERS[53][5] , \REGISTERS[53][4] ,
         \REGISTERS[53][3] , \REGISTERS[53][2] , \REGISTERS[53][1] ,
         \REGISTERS[53][0] , \REGISTERS[54][31] , \REGISTERS[54][30] ,
         \REGISTERS[54][29] , \REGISTERS[54][28] , \REGISTERS[54][27] ,
         \REGISTERS[54][26] , \REGISTERS[54][25] , \REGISTERS[54][24] ,
         \REGISTERS[54][23] , \REGISTERS[54][22] , \REGISTERS[54][21] ,
         \REGISTERS[54][20] , \REGISTERS[54][19] , \REGISTERS[54][18] ,
         \REGISTERS[54][17] , \REGISTERS[54][16] , \REGISTERS[54][15] ,
         \REGISTERS[54][14] , \REGISTERS[54][13] , \REGISTERS[54][12] ,
         \REGISTERS[54][11] , \REGISTERS[54][10] , \REGISTERS[54][9] ,
         \REGISTERS[54][8] , \REGISTERS[54][7] , \REGISTERS[54][6] ,
         \REGISTERS[54][5] , \REGISTERS[54][4] , \REGISTERS[54][3] ,
         \REGISTERS[54][2] , \REGISTERS[54][1] , \REGISTERS[54][0] ,
         \REGISTERS[77][31] , \REGISTERS[77][30] , \REGISTERS[77][29] ,
         \REGISTERS[77][28] , \REGISTERS[77][27] , \REGISTERS[77][26] ,
         \REGISTERS[77][25] , \REGISTERS[77][24] , \REGISTERS[77][23] ,
         \REGISTERS[77][22] , \REGISTERS[77][21] , \REGISTERS[77][20] ,
         \REGISTERS[77][19] , \REGISTERS[77][18] , \REGISTERS[77][17] ,
         \REGISTERS[77][16] , \REGISTERS[77][15] , \REGISTERS[77][14] ,
         \REGISTERS[77][13] , \REGISTERS[77][12] , \REGISTERS[77][11] ,
         \REGISTERS[77][10] , \REGISTERS[77][9] , \REGISTERS[77][8] ,
         \REGISTERS[77][7] , \REGISTERS[77][6] , \REGISTERS[77][5] ,
         \REGISTERS[77][4] , \REGISTERS[77][3] , \REGISTERS[77][2] ,
         \REGISTERS[77][1] , \REGISTERS[77][0] , \REGISTERS[78][31] ,
         \REGISTERS[78][30] , \REGISTERS[78][29] , \REGISTERS[78][28] ,
         \REGISTERS[78][27] , \REGISTERS[78][26] , \REGISTERS[78][25] ,
         \REGISTERS[78][24] , \REGISTERS[78][23] , \REGISTERS[78][22] ,
         \REGISTERS[78][21] , \REGISTERS[78][20] , \REGISTERS[78][19] ,
         \REGISTERS[78][18] , \REGISTERS[78][17] , \REGISTERS[78][16] ,
         \REGISTERS[78][15] , \REGISTERS[78][14] , \REGISTERS[78][13] ,
         \REGISTERS[78][12] , \REGISTERS[78][11] , \REGISTERS[78][10] ,
         \REGISTERS[78][9] , \REGISTERS[78][8] , \REGISTERS[78][7] ,
         \REGISTERS[78][6] , \REGISTERS[78][5] , \REGISTERS[78][4] ,
         \REGISTERS[78][3] , \REGISTERS[78][2] , \REGISTERS[78][1] ,
         \REGISTERS[78][0] , \REGISTERS[82][31] , \REGISTERS[82][30] ,
         \REGISTERS[82][29] , \REGISTERS[82][28] , \REGISTERS[82][27] ,
         \REGISTERS[82][26] , \REGISTERS[82][25] , \REGISTERS[82][24] ,
         \REGISTERS[82][23] , \REGISTERS[82][22] , \REGISTERS[82][21] ,
         \REGISTERS[82][20] , \REGISTERS[82][19] , \REGISTERS[82][18] ,
         \REGISTERS[82][17] , \REGISTERS[82][16] , \REGISTERS[82][15] ,
         \REGISTERS[82][14] , \REGISTERS[82][13] , \REGISTERS[82][12] ,
         \REGISTERS[82][11] , \REGISTERS[82][10] , \REGISTERS[82][9] ,
         \REGISTERS[82][8] , \REGISTERS[82][7] , \REGISTERS[82][6] ,
         \REGISTERS[82][5] , \REGISTERS[82][4] , \REGISTERS[82][3] ,
         \REGISTERS[82][2] , \REGISTERS[82][1] , \REGISTERS[82][0] ,
         \REGISTERS[83][31] , \REGISTERS[83][30] , \REGISTERS[83][29] ,
         \REGISTERS[83][28] , \REGISTERS[83][27] , \REGISTERS[83][26] ,
         \REGISTERS[83][25] , \REGISTERS[83][24] , \REGISTERS[83][23] ,
         \REGISTERS[83][22] , \REGISTERS[83][21] , \REGISTERS[83][20] ,
         \REGISTERS[83][19] , \REGISTERS[83][18] , \REGISTERS[83][17] ,
         \REGISTERS[83][16] , \REGISTERS[83][15] , \REGISTERS[83][14] ,
         \REGISTERS[83][13] , \REGISTERS[83][12] , \REGISTERS[83][11] ,
         \REGISTERS[83][10] , \REGISTERS[83][9] , \REGISTERS[83][8] ,
         \REGISTERS[83][7] , \REGISTERS[83][6] , \REGISTERS[83][5] ,
         \REGISTERS[83][4] , \REGISTERS[83][3] , \REGISTERS[83][2] ,
         \REGISTERS[83][1] , \REGISTERS[83][0] , \REGISTERS[84][31] ,
         \REGISTERS[84][30] , \REGISTERS[84][29] , \REGISTERS[84][28] ,
         \REGISTERS[84][27] , \REGISTERS[84][26] , \REGISTERS[84][25] ,
         \REGISTERS[84][24] , \REGISTERS[84][23] , \REGISTERS[84][22] ,
         \REGISTERS[84][21] , \REGISTERS[84][20] , \REGISTERS[84][19] ,
         \REGISTERS[84][18] , \REGISTERS[84][17] , \REGISTERS[84][16] ,
         \REGISTERS[84][15] , \REGISTERS[84][14] , \REGISTERS[84][13] ,
         \REGISTERS[84][12] , \REGISTERS[84][11] , \REGISTERS[84][10] ,
         \REGISTERS[84][9] , \REGISTERS[84][8] , \REGISTERS[84][7] ,
         \REGISTERS[84][6] , \REGISTERS[84][5] , \REGISTERS[84][4] ,
         \REGISTERS[84][3] , \REGISTERS[84][2] , \REGISTERS[84][1] ,
         \REGISTERS[84][0] , \REGISTERS[85][31] , \REGISTERS[85][30] ,
         \REGISTERS[85][29] , \REGISTERS[85][28] , \REGISTERS[85][27] ,
         \REGISTERS[85][26] , \REGISTERS[85][25] , \REGISTERS[85][24] ,
         \REGISTERS[85][23] , \REGISTERS[85][22] , \REGISTERS[85][21] ,
         \REGISTERS[85][20] , \REGISTERS[85][19] , \REGISTERS[85][18] ,
         \REGISTERS[85][17] , \REGISTERS[85][16] , \REGISTERS[85][15] ,
         \REGISTERS[85][14] , \REGISTERS[85][13] , \REGISTERS[85][12] ,
         \REGISTERS[85][11] , \REGISTERS[85][10] , \REGISTERS[85][9] ,
         \REGISTERS[85][8] , \REGISTERS[85][7] , \REGISTERS[85][6] ,
         \REGISTERS[85][5] , \REGISTERS[85][4] , \REGISTERS[85][3] ,
         \REGISTERS[85][2] , \REGISTERS[85][1] , \REGISTERS[85][0] ,
         \REGISTERS[86][31] , \REGISTERS[86][30] , \REGISTERS[86][29] ,
         \REGISTERS[86][28] , \REGISTERS[86][27] , \REGISTERS[86][26] ,
         \REGISTERS[86][25] , \REGISTERS[86][24] , \REGISTERS[86][23] ,
         \REGISTERS[86][22] , \REGISTERS[86][21] , \REGISTERS[86][20] ,
         \REGISTERS[86][19] , \REGISTERS[86][18] , \REGISTERS[86][17] ,
         \REGISTERS[86][16] , \REGISTERS[86][15] , \REGISTERS[86][14] ,
         \REGISTERS[86][13] , \REGISTERS[86][12] , \REGISTERS[86][11] ,
         \REGISTERS[86][10] , \REGISTERS[86][9] , \REGISTERS[86][8] ,
         \REGISTERS[86][7] , \REGISTERS[86][6] , \REGISTERS[86][5] ,
         \REGISTERS[86][4] , \REGISTERS[86][3] , \REGISTERS[86][2] ,
         \REGISTERS[86][1] , \REGISTERS[86][0] , \REGISTERS[87][31] ,
         \REGISTERS[87][30] , \REGISTERS[87][29] , \REGISTERS[87][28] ,
         \REGISTERS[87][27] , \REGISTERS[87][26] , \REGISTERS[87][25] ,
         \REGISTERS[87][24] , \REGISTERS[87][23] , \REGISTERS[87][22] ,
         \REGISTERS[87][21] , \REGISTERS[87][20] , \REGISTERS[87][19] ,
         \REGISTERS[87][18] , \REGISTERS[87][17] , \REGISTERS[87][16] ,
         \REGISTERS[87][15] , \REGISTERS[87][14] , \REGISTERS[87][13] ,
         \REGISTERS[87][12] , \REGISTERS[87][11] , \REGISTERS[87][10] ,
         \REGISTERS[87][9] , \REGISTERS[87][8] , \REGISTERS[87][7] ,
         \REGISTERS[87][6] , \REGISTERS[87][5] , \REGISTERS[87][4] ,
         \REGISTERS[87][3] , \REGISTERS[87][2] , \REGISTERS[87][1] ,
         \REGISTERS[87][0] , N2151, N2153, N2154, N2155, N2156, N2157, N2158,
         N2159, N2160, N2161, N2162, N2163, N2164, N2165, N2166, N8415, N8417,
         N8418, N8419, N8420, N8421, N8422, N8423, N8424, N8425, N8426, N8427,
         N8428, N8429, N8430, N8559, N8561, N8562, N8563, N8564, N8565, N8566,
         N8567, N8568, N8569, N8570, N8571, N8572, N8573, N8574, N8702, N8703,
         N8704, N8705, N8706, N8707, N8708, N8709, N8710, N8711, N8712, N8713,
         N8714, N8715, N8716, N8717, N8718, N8719, N8720, N8721, N8722, N8723,
         N8724, N8725, N8726, N8727, N8728, N8729, N8730, N8731, N8732, N8733,
         N8734, N8735, N8736, N8737, N8738, N8739, N8740, N8741, N8742, N8743,
         N8744, N8745, N8746, N8747, N8748, N8749, N8750, N8751, N8752, N8753,
         N8754, N8755, N8756, N8757, N8758, N8759, N8760, N8761, N8762, N8763,
         N8764, N8765, N8766, N8767, N8787, N8788, N8789, N8790, N8791, N8833,
         N8834, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2898,
         n2916, n2918, n2919, n2920, n2921, n2996, n3029, n3030, n3033, n3035,
         n3038, n3040, n3043, n3045, n3048, n3050, n3053, n3055, n3058, n3060,
         n3063, n3065, n3068, n3070, n3073, n3075, n3078, n3080, n3083, n3085,
         n3088, n3090, n3093, n3095, n3098, n3100, n3103, n3105, n3106, n3107,
         n3108, n3109, n3112, n3114, n3117, n3121, n3125, n3129, n3133, n3137,
         n3141, n3145, n3149, n3153, n3157, n3161, n3165, n3169, n3173, n3177,
         n3179, n3182, n3186, n3190, n3194, n3198, n3202, n3206, n3210, n3214,
         n3218, n3222, n3226, n3230, n3234, n3238, n3242, n3244, n3247, n3251,
         n3255, n3259, n3263, n3267, n3271, n3275, n3279, n3283, n3287, n3291,
         n3295, n3299, n3303, n3307, n3309, n3312, n3316, n3320, n3324, n3328,
         n3332, n3336, n3340, n3342, n3343, n3346, n3348, n3351, n3353, n3356,
         n3358, n3359, n3362, n3364, n3367, n3371, n3375, n3377, n3380, n3382,
         n3383, n3386, n3390, n3394, n3398, n3400, n3403, n3405, n3406, n3409,
         n3413, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, \sub_189/carry[6] , n1, n2,
         n3, n4, n5, n6, n8, n9, n10, n12, n13, n14, n15, n16, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2917, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3031,
         n3032, n3034, n3036, n3037, n3039, n3041, n3042, n3044, n3046, n3047,
         n3049, n3051, n3052, n3054, n3056, n3057, n3059, n3061, n3062, n3064,
         n3066, n3067, n3069, n3071, n3072, n3074, n3076, n3077, n3079, n3081,
         n3082, n3084, n3086, n3087, n3089, n3091, n3092, n3094, n3096, n3097,
         n3099, n3101, n3102, n3104, n3110, n3111, n3113, n3115, n3116, n3118,
         n3119, n3120, n3122, n3123, n3124, n3126, n3127, n3128, n3130, n3131,
         n3132, n3134, n3135, n3136, n3138, n3139, n3140, n3142, n3143, n3144,
         n3146, n3147, n3148, n3150, n3151, n3152, n3154, n3155, n3156, n3158,
         n3159, n3160, n3162, n3163, n3164, n3166, n3167, n3168, n3170, n3171,
         n3172, n3174, n3175, n3176, n3178, n3180, n3181, n3183, n3184, n3185,
         n3187, n3188, n3189, n3191, n3192, n3193, n3195, n3196, n3197, n3199,
         n3200, n3201, n3203, n3204, n3205, n3207, n3208, n3209, n3211, n3212,
         n3213, n3215, n3216, n3217, n3219, n3220, n3221, n3223, n3224, n3225,
         n3227, n3228, n3229, n3231, n3232, n3233, n3235, n3236, n3237, n3239,
         n3240, n3241, n3243, n3245, n3246, n3248, n3249, n3250, n3252, n3253,
         n3254, n3256, n3257, n3258, n3260, n3261, n3262, n3264, n3265, n3266,
         n3268, n3269, n3270, n3272, n3273, n3274, n3276, n3277, n3278, n3280,
         n3281, n3282, n3284, n3285, n3286, n3288, n3289, n3290, n3292, n3293,
         n3294, n3296, n3297, n3298, n3300, n3301, n3302, n3304, n3305, n3306,
         n3308, n3310, n3311, n3313, n3314, n3315, n3317, n3318, n3319, n3321,
         n3322, n3323, n3325, n3326, n3327, n3329, n3330, n3331, n3333, n3334,
         n3335, n3337, n3338, n3339, n3341, n3344, n3345, n3347, n3349, n3350,
         n3352, n3354, n3355, n3357, n3360, n3361, n3363, n3365, n3366, n3368,
         n3369, n3370, n3372, n3373, n3374, n3376, n3378, n3379, n3381, n3384,
         n3385, n3387, n3388, n3389, n3391, n3392, n3393, n3395, n3396, n3397,
         n3399, n3401, n3402, n3404, n3407, n3408, n3410, n3411, n3412, n3414,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921;
  wire   [6:0] CWP;
  assign SPILL = 1'b0;
  assign BUSout[31] = 1'b0;
  assign BUSout[30] = 1'b0;
  assign BUSout[29] = 1'b0;
  assign BUSout[28] = 1'b0;
  assign BUSout[27] = 1'b0;
  assign BUSout[26] = 1'b0;
  assign BUSout[25] = 1'b0;
  assign BUSout[24] = 1'b0;
  assign BUSout[23] = 1'b0;
  assign BUSout[22] = 1'b0;
  assign BUSout[21] = 1'b0;
  assign BUSout[20] = 1'b0;
  assign BUSout[19] = 1'b0;
  assign BUSout[18] = 1'b0;
  assign BUSout[17] = 1'b0;
  assign BUSout[16] = 1'b0;
  assign BUSout[15] = 1'b0;
  assign BUSout[14] = 1'b0;
  assign BUSout[13] = 1'b0;
  assign BUSout[12] = 1'b0;
  assign BUSout[11] = 1'b0;
  assign BUSout[10] = 1'b0;
  assign BUSout[9] = 1'b0;
  assign BUSout[8] = 1'b0;
  assign BUSout[7] = 1'b0;
  assign BUSout[6] = 1'b0;
  assign BUSout[5] = 1'b0;
  assign BUSout[4] = 1'b0;
  assign BUSout[3] = 1'b0;
  assign BUSout[2] = 1'b0;
  assign BUSout[1] = 1'b0;
  assign BUSout[0] = 1'b0;
  assign N2160 = ADD_WR[0];
  assign N2161 = ADD_WR[1];
  assign N2162 = ADD_WR[2];
  assign N8424 = ADD_RD1[0];
  assign N8425 = ADD_RD1[1];
  assign N8426 = ADD_RD1[2];
  assign N8568 = ADD_RD2[0];
  assign N8569 = ADD_RD2[1];
  assign N8570 = ADD_RD2[2];
  assign FILL = 1'b0;

  DFFR_X1 \REGISTERS_reg[0][31]  ( .D(n6317), .CK(CLK), .RN(n2974), .Q(n3393), 
        .QN(n80) );
  DFFR_X1 \REGISTERS_reg[0][30]  ( .D(n6318), .CK(CLK), .RN(n2973), .Q(n3395), 
        .QN(n81) );
  DFFR_X1 \REGISTERS_reg[0][29]  ( .D(n6319), .CK(CLK), .RN(n2971), .Q(n3396), 
        .QN(n82) );
  DFFR_X1 \REGISTERS_reg[0][28]  ( .D(n6320), .CK(CLK), .RN(n2972), .Q(n3397), 
        .QN(n83) );
  DFFR_X1 \REGISTERS_reg[0][27]  ( .D(n6321), .CK(CLK), .RN(n3264), .Q(n3399), 
        .QN(n84) );
  DFFR_X1 \REGISTERS_reg[0][26]  ( .D(n6322), .CK(CLK), .RN(n3264), .Q(n3401), 
        .QN(n85) );
  DFFR_X1 \REGISTERS_reg[0][25]  ( .D(n6323), .CK(CLK), .RN(n3264), .Q(n3402), 
        .QN(n86) );
  DFFR_X1 \REGISTERS_reg[0][24]  ( .D(n6324), .CK(CLK), .RN(n3264), .Q(n3404), 
        .QN(n87) );
  DFFR_X1 \REGISTERS_reg[0][23]  ( .D(n6325), .CK(CLK), .RN(n3264), .Q(n3407), 
        .QN(n88) );
  DFFR_X1 \REGISTERS_reg[0][22]  ( .D(n6326), .CK(CLK), .RN(n3264), .Q(n3408), 
        .QN(n89) );
  DFFR_X1 \REGISTERS_reg[0][21]  ( .D(n6327), .CK(CLK), .RN(n3264), .Q(n3410), 
        .QN(n90) );
  DFFR_X1 \REGISTERS_reg[0][20]  ( .D(n6328), .CK(CLK), .RN(n3264), .Q(n3411), 
        .QN(n91) );
  DFFR_X1 \REGISTERS_reg[0][19]  ( .D(n6329), .CK(CLK), .RN(n3264), .Q(n3412), 
        .QN(n92) );
  DFFR_X1 \REGISTERS_reg[0][18]  ( .D(n6330), .CK(CLK), .RN(n3264), .Q(n3414), 
        .QN(n93) );
  DFFR_X1 \REGISTERS_reg[0][17]  ( .D(n6331), .CK(CLK), .RN(n3264), .Q(n9140), 
        .QN(n94) );
  DFFR_X1 \REGISTERS_reg[0][16]  ( .D(n6332), .CK(CLK), .RN(n3264), .Q(n9141), 
        .QN(n95) );
  DFFR_X1 \REGISTERS_reg[0][15]  ( .D(n6333), .CK(CLK), .RN(n3262), .Q(n9142), 
        .QN(n96) );
  DFFR_X1 \REGISTERS_reg[0][14]  ( .D(n6334), .CK(CLK), .RN(n3262), .Q(n9143), 
        .QN(n97) );
  DFFR_X1 \REGISTERS_reg[0][13]  ( .D(n6335), .CK(CLK), .RN(n3262), .Q(n9144), 
        .QN(n98) );
  DFFR_X1 \REGISTERS_reg[0][12]  ( .D(n6336), .CK(CLK), .RN(n3262), .Q(n9145), 
        .QN(n99) );
  DFFR_X1 \REGISTERS_reg[0][11]  ( .D(n6337), .CK(CLK), .RN(n3262), .Q(n9146), 
        .QN(n100) );
  DFFR_X1 \REGISTERS_reg[0][10]  ( .D(n6338), .CK(CLK), .RN(n3262), .Q(n9147), 
        .QN(n101) );
  DFFR_X1 \REGISTERS_reg[0][9]  ( .D(n6339), .CK(CLK), .RN(n3262), .Q(n9148), 
        .QN(n102) );
  DFFR_X1 \REGISTERS_reg[0][8]  ( .D(n6340), .CK(CLK), .RN(n3262), .Q(n9149), 
        .QN(n103) );
  DFFR_X1 \REGISTERS_reg[0][7]  ( .D(n6341), .CK(CLK), .RN(n3262), .Q(n9150), 
        .QN(n104) );
  DFFR_X1 \REGISTERS_reg[0][6]  ( .D(n6342), .CK(CLK), .RN(n3262), .Q(n9151), 
        .QN(n105) );
  DFFR_X1 \REGISTERS_reg[0][5]  ( .D(n6343), .CK(CLK), .RN(n3262), .Q(n9152), 
        .QN(n106) );
  DFFR_X1 \REGISTERS_reg[0][4]  ( .D(n6344), .CK(CLK), .RN(n3262), .Q(n9153), 
        .QN(n107) );
  DFFR_X1 \REGISTERS_reg[0][3]  ( .D(n6345), .CK(CLK), .RN(n2977), .Q(n9154), 
        .QN(n108) );
  DFFR_X1 \REGISTERS_reg[0][2]  ( .D(n6346), .CK(CLK), .RN(n2975), .Q(n9155), 
        .QN(n109) );
  DFFR_X1 \REGISTERS_reg[0][1]  ( .D(n6347), .CK(CLK), .RN(n2976), .Q(n9156), 
        .QN(n110) );
  DFFR_X1 \REGISTERS_reg[0][0]  ( .D(n6348), .CK(CLK), .RN(n3006), .Q(n9157), 
        .QN(n111) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n6349), .CK(CLK), .RN(n3007), .Q(n9158), 
        .QN(n112) );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n6350), .CK(CLK), .RN(n2983), .Q(n9159), 
        .QN(n113) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n6351), .CK(CLK), .RN(n2981), .Q(n9160), 
        .QN(n114) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n6352), .CK(CLK), .RN(n2982), .Q(n9161), 
        .QN(n115) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n6353), .CK(CLK), .RN(n2984), .Q(n9162), 
        .QN(n116) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n6354), .CK(CLK), .RN(n2979), .Q(n9163), 
        .QN(n117) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n6355), .CK(CLK), .RN(n2980), .Q(n9164), 
        .QN(n118) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n6356), .CK(CLK), .RN(n2978), .Q(n9165), 
        .QN(n119) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n6357), .CK(CLK), .RN(n3018), .Q(n9166), 
        .QN(n120) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n6358), .CK(CLK), .RN(n3016), .Q(n9167), 
        .QN(n121) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n6359), .CK(CLK), .RN(n3014), .Q(n9168), 
        .QN(n122) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n6360), .CK(CLK), .RN(n3010), .Q(n9169), 
        .QN(n123) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n6361), .CK(CLK), .RN(n3017), .Q(n9170), 
        .QN(n124) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n6362), .CK(CLK), .RN(n3015), .Q(n9171), 
        .QN(n125) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n6363), .CK(CLK), .RN(n3011), .Q(n9172), 
        .QN(n126) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n6364), .CK(CLK), .RN(n3008), .Q(n9173), 
        .QN(n127) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n6365), .CK(CLK), .RN(n3019), .Q(n9174), 
        .QN(n128) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n6366), .CK(CLK), .RN(n3012), .Q(n9175), 
        .QN(n129) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n6367), .CK(CLK), .RN(n3013), .Q(n9176), 
        .QN(n130) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n6368), .CK(CLK), .RN(n3009), .Q(n9177), 
        .QN(n131) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n6369), .CK(CLK), .RN(n2990), .Q(n9178), 
        .QN(n132) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n6370), .CK(CLK), .RN(n2985), .Q(n9179), 
        .QN(n133) );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n6371), .CK(CLK), .RN(n2986), .Q(n9180), 
        .QN(n134) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n6372), .CK(CLK), .RN(n3025), .Q(n9181), 
        .QN(n135) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n6373), .CK(CLK), .RN(n2989), .Q(n9182), 
        .QN(n136) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n6374), .CK(CLK), .RN(n2987), .Q(n9183), 
        .QN(n137) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n6375), .CK(CLK), .RN(n3023), .Q(n9184), 
        .QN(n138) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n6376), .CK(CLK), .RN(n3024), .Q(n9185), 
        .QN(n139) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n6377), .CK(CLK), .RN(n3022), .Q(n9186), 
        .QN(n140) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n6378), .CK(CLK), .RN(n3020), .Q(n9187), 
        .QN(n141) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n6379), .CK(CLK), .RN(n3021), .Q(n9188), 
        .QN(n142) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n6380), .CK(CLK), .RN(n2988), .Q(n9189), 
        .QN(n143) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n6381), .CK(CLK), .RN(n3261), .Q(n9190), 
        .QN(n144) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n6382), .CK(CLK), .RN(n3261), .Q(n9191), 
        .QN(n145) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n6383), .CK(CLK), .RN(n3261), .Q(n9192), 
        .QN(n146) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n6384), .CK(CLK), .RN(n3261), .Q(n9193), 
        .QN(n147) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n6385), .CK(CLK), .RN(n3261), .Q(n9194), 
        .QN(n148) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n6386), .CK(CLK), .RN(n3261), .Q(n9195), 
        .QN(n149) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n6387), .CK(CLK), .RN(n3261), .Q(n9196), 
        .QN(n150) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n6388), .CK(CLK), .RN(n3261), .Q(n9197), 
        .QN(n151) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n6389), .CK(CLK), .RN(n3261), .Q(n9198), 
        .QN(n152) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n6390), .CK(CLK), .RN(n3261), .Q(n9199), 
        .QN(n153) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n6391), .CK(CLK), .RN(n3261), .Q(n9200), 
        .QN(n154) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n6392), .CK(CLK), .RN(n3261), .Q(n9201), 
        .QN(n155) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n6393), .CK(CLK), .RN(n3260), .Q(n9202), 
        .QN(n156) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n6394), .CK(CLK), .RN(n3260), .Q(n9203), 
        .QN(n157) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n6395), .CK(CLK), .RN(n3260), .Q(n9204), 
        .QN(n158) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n6396), .CK(CLK), .RN(n3260), .Q(n9205), 
        .QN(n159) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n6397), .CK(CLK), .RN(n3260), .Q(n9206), 
        .QN(n160) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n6398), .CK(CLK), .RN(n3260), .Q(n9207), 
        .QN(n161) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n6399), .CK(CLK), .RN(n3260), .Q(n9208), 
        .QN(n162) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n6400), .CK(CLK), .RN(n3260), .Q(n9209), 
        .QN(n163) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n6401), .CK(CLK), .RN(n3260), .Q(n9210), 
        .QN(n164) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n6402), .CK(CLK), .RN(n3260), .Q(n9211), 
        .QN(n165) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n6403), .CK(CLK), .RN(n3260), .Q(n9212), 
        .QN(n166) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n6404), .CK(CLK), .RN(n3260), .Q(n9213), 
        .QN(n167) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n6405), .CK(CLK), .RN(n3258), .Q(n9214), 
        .QN(n168) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n6406), .CK(CLK), .RN(n3258), .Q(n9215), 
        .QN(n169) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n6407), .CK(CLK), .RN(n3258), .Q(n9216), 
        .QN(n170) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n6408), .CK(CLK), .RN(n3258), .Q(n9217), 
        .QN(n171) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n6409), .CK(CLK), .RN(n3258), .Q(n9218), 
        .QN(n172) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n6410), .CK(CLK), .RN(n3258), .Q(n9219), 
        .QN(n173) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n6411), .CK(CLK), .RN(n3258), .Q(n9220), 
        .QN(n174) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n6412), .CK(CLK), .RN(n3258), .Q(n9221), 
        .QN(n175) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n6413), .CK(CLK), .RN(n3258), .Q(n9222), 
        .QN(n176) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n6414), .CK(CLK), .RN(n3258), .Q(n9223), 
        .QN(n177) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n6415), .CK(CLK), .RN(n3258), .Q(n9224), 
        .QN(n178) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n6416), .CK(CLK), .RN(n3258), .Q(n9225), 
        .QN(n179) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n6417), .CK(CLK), .RN(n3257), .Q(n9226), 
        .QN(n180) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n6418), .CK(CLK), .RN(n3257), .Q(n9227), 
        .QN(n181) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n6419), .CK(CLK), .RN(n3257), .Q(n9228), 
        .QN(n182) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n6420), .CK(CLK), .RN(n3257), .Q(n9229), 
        .QN(n183) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n6421), .CK(CLK), .RN(n3257), .Q(n9230), 
        .QN(n184) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n6422), .CK(CLK), .RN(n3257), .Q(n9231), 
        .QN(n185) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n6423), .CK(CLK), .RN(n3257), .Q(n9232), 
        .QN(n186) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n6424), .CK(CLK), .RN(n3257), .Q(n9233), 
        .QN(n187) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n6425), .CK(CLK), .RN(n3257), .Q(n9234), 
        .QN(n188) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n6426), .CK(CLK), .RN(n3257), .Q(n9235), 
        .QN(n189) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n6427), .CK(CLK), .RN(n3257), .Q(n9236), 
        .QN(n190) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n6428), .CK(CLK), .RN(n3257), .Q(n9237), 
        .QN(n191) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n6429), .CK(CLK), .RN(n3256), .Q(n9238), 
        .QN(n192) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n6430), .CK(CLK), .RN(n3256), .Q(n9239), 
        .QN(n193) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n6431), .CK(CLK), .RN(n3256), .Q(n9240), 
        .QN(n194) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n6432), .CK(CLK), .RN(n3256), .Q(n9241), 
        .QN(n195) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n6433), .CK(CLK), .RN(n3256), .Q(n9242), 
        .QN(n196) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n6434), .CK(CLK), .RN(n3256), .Q(n9243), 
        .QN(n197) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n6435), .CK(CLK), .RN(n3256), .Q(n9244), 
        .QN(n198) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n6436), .CK(CLK), .RN(n3256), .Q(n9245), 
        .QN(n199) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n6437), .CK(CLK), .RN(n3256), .Q(n9246), 
        .QN(n200) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n6438), .CK(CLK), .RN(n3256), .Q(n9247), 
        .QN(n201) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n6439), .CK(CLK), .RN(n3256), .Q(n9248), 
        .QN(n202) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n6440), .CK(CLK), .RN(n3256), .Q(n9249), 
        .QN(n203) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n6441), .CK(CLK), .RN(n3254), .Q(n9250), 
        .QN(n204) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n6442), .CK(CLK), .RN(n3254), .Q(n9251), 
        .QN(n205) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n6443), .CK(CLK), .RN(n3254), .Q(n9252), 
        .QN(n206) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n6444), .CK(CLK), .RN(n3254), .Q(n9253), 
        .QN(n207) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n6445), .CK(CLK), .RN(n3254), .Q(n9254), 
        .QN(n208) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n6446), .CK(CLK), .RN(n3254), .Q(n9255), 
        .QN(n209) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n6447), .CK(CLK), .RN(n3254), .Q(n9256), 
        .QN(n210) );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n6448), .CK(CLK), .RN(n3254), .Q(n9257), 
        .QN(n211) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n6449), .CK(CLK), .RN(n3254), .Q(n9258), 
        .QN(n212) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n6450), .CK(CLK), .RN(n3254), .Q(n9259), 
        .QN(n213) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n6451), .CK(CLK), .RN(n3254), .Q(n9260), 
        .QN(n214) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n6452), .CK(CLK), .RN(n3254), .Q(n9261), 
        .QN(n215) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n6453), .CK(CLK), .RN(n3253), .Q(n9262), 
        .QN(n216) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n6454), .CK(CLK), .RN(n3253), .Q(n9263), 
        .QN(n217) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n6455), .CK(CLK), .RN(n3253), .Q(n9264), 
        .QN(n218) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n6456), .CK(CLK), .RN(n3253), .Q(n9265), 
        .QN(n219) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n6457), .CK(CLK), .RN(n3253), .Q(n9266), 
        .QN(n220) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n6458), .CK(CLK), .RN(n3253), .Q(n9267), 
        .QN(n221) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n6459), .CK(CLK), .RN(n3253), .Q(n9268), 
        .QN(n222) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n6460), .CK(CLK), .RN(n3253), .Q(n9269), 
        .QN(n223) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n6461), .CK(CLK), .RN(n3253), .Q(n9270), 
        .QN(n224) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n6462), .CK(CLK), .RN(n3253), .Q(n9271), 
        .QN(n225) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n6463), .CK(CLK), .RN(n3253), .Q(n9272), 
        .QN(n226) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n6464), .CK(CLK), .RN(n3253), .Q(n9273), 
        .QN(n227) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n6465), .CK(CLK), .RN(n3252), .Q(n9274), 
        .QN(n228) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n6466), .CK(CLK), .RN(n3252), .Q(n9275), 
        .QN(n229) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n6467), .CK(CLK), .RN(n3252), .Q(n9276), 
        .QN(n230) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n6468), .CK(CLK), .RN(n3252), .Q(n9277), 
        .QN(n231) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n6469), .CK(CLK), .RN(n3252), .Q(n9278), 
        .QN(n232) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n6470), .CK(CLK), .RN(n3252), .Q(n9279), 
        .QN(n233) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n6471), .CK(CLK), .RN(n3252), .Q(n9280), 
        .QN(n234) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n6472), .CK(CLK), .RN(n3252), .Q(n9281), 
        .QN(n235) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n6473), .CK(CLK), .RN(n3252), .Q(n9282), 
        .QN(n236) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n6474), .CK(CLK), .RN(n3252), .Q(n9283), 
        .QN(n237) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n6475), .CK(CLK), .RN(n3252), .Q(n9284), 
        .QN(n238) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n6476), .CK(CLK), .RN(n3252), .Q(n9285), 
        .QN(n239) );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n6477), .CK(CLK), .RN(n3250), .Q(n9286), 
        .QN(n240) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n6478), .CK(CLK), .RN(n3250), .Q(n9287), 
        .QN(n241) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n6479), .CK(CLK), .RN(n3250), .Q(n9288), 
        .QN(n242) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n6480), .CK(CLK), .RN(n3250), .Q(n9289), 
        .QN(n243) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n6481), .CK(CLK), .RN(n3250), .Q(n9290), 
        .QN(n244) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n6482), .CK(CLK), .RN(n3250), .Q(n9291), 
        .QN(n245) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n6483), .CK(CLK), .RN(n3250), .Q(n9292), 
        .QN(n246) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n6484), .CK(CLK), .RN(n3250), .Q(n9293), 
        .QN(n247) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n6485), .CK(CLK), .RN(n3250), .Q(n9294), 
        .QN(n248) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n6486), .CK(CLK), .RN(n3250), .Q(n9295), 
        .QN(n249) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n6487), .CK(CLK), .RN(n3250), .Q(n9296), 
        .QN(n250) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n6488), .CK(CLK), .RN(n3250), .Q(n9297), 
        .QN(n251) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n6489), .CK(CLK), .RN(n3249), .Q(n9298), 
        .QN(n252) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n6490), .CK(CLK), .RN(n3249), .Q(n9299), 
        .QN(n253) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n6491), .CK(CLK), .RN(n3249), .Q(n9300), 
        .QN(n254) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n6492), .CK(CLK), .RN(n3249), .Q(n9301), 
        .QN(n255) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n6493), .CK(CLK), .RN(n3249), .Q(n9302), 
        .QN(n256) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n6494), .CK(CLK), .RN(n3249), .Q(n9303), 
        .QN(n257) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n6495), .CK(CLK), .RN(n3249), .Q(n9304), 
        .QN(n258) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n6496), .CK(CLK), .RN(n3249), .Q(n9305), 
        .QN(n259) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n6497), .CK(CLK), .RN(n3249), .Q(n9306), 
        .QN(n260) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n6498), .CK(CLK), .RN(n3249), .Q(n9307), 
        .QN(n261) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n6499), .CK(CLK), .RN(n3249), .Q(n9308), 
        .QN(n262) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n6500), .CK(CLK), .RN(n3249), .Q(n9309), 
        .QN(n263) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n6501), .CK(CLK), .RN(n3248), .Q(n9310), 
        .QN(n264) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n6502), .CK(CLK), .RN(n3248), .Q(n9311), 
        .QN(n265) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n6503), .CK(CLK), .RN(n3248), .Q(n9312), 
        .QN(n266) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n6504), .CK(CLK), .RN(n3248), .Q(n9313), 
        .QN(n267) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n6505), .CK(CLK), .RN(n3248), .Q(n9314), 
        .QN(n268) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n6506), .CK(CLK), .RN(n3248), .Q(n9315), 
        .QN(n269) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n6507), .CK(CLK), .RN(n3248), .Q(n9316), 
        .QN(n270) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n6508), .CK(CLK), .RN(n3248), .Q(n9317), 
        .QN(n271) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n6509), .CK(CLK), .RN(n3248), .Q(n9318), 
        .QN(n272) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n6510), .CK(CLK), .RN(n3248), .Q(n9319), 
        .QN(n273) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n6511), .CK(CLK), .RN(n3248), .Q(n9320), 
        .QN(n274) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n6512), .CK(CLK), .RN(n3248), .Q(n9321), 
        .QN(n275) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n6513), .CK(CLK), .RN(n3246), .Q(n9322), 
        .QN(n276) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n6514), .CK(CLK), .RN(n3246), .Q(n9323), 
        .QN(n277) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n6515), .CK(CLK), .RN(n3246), .Q(n9324), 
        .QN(n278) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n6516), .CK(CLK), .RN(n3246), .Q(n9325), 
        .QN(n279) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n6517), .CK(CLK), .RN(n3246), .Q(n9326), 
        .QN(n280) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n6518), .CK(CLK), .RN(n3246), .Q(n9327), 
        .QN(n281) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n6519), .CK(CLK), .RN(n3246), .Q(n9328), 
        .QN(n282) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n6520), .CK(CLK), .RN(n3246), .Q(n9329), 
        .QN(n283) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n6521), .CK(CLK), .RN(n3246), .Q(n9330), 
        .QN(n284) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n6522), .CK(CLK), .RN(n3246), .Q(n9331), 
        .QN(n285) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n6523), .CK(CLK), .RN(n3246), .Q(n9332), 
        .QN(n286) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n6524), .CK(CLK), .RN(n3246), .Q(n9333), 
        .QN(n287) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n6525), .CK(CLK), .RN(n3245), .Q(n9334), 
        .QN(n288) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n6526), .CK(CLK), .RN(n3245), .Q(n9335), 
        .QN(n289) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n6527), .CK(CLK), .RN(n3245), .Q(n9336), 
        .QN(n290) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n6528), .CK(CLK), .RN(n3245), .Q(n9337), 
        .QN(n291) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n6529), .CK(CLK), .RN(n3245), .Q(n9338), 
        .QN(n292) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n6530), .CK(CLK), .RN(n3245), .Q(n9339), 
        .QN(n293) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n6531), .CK(CLK), .RN(n3245), .Q(n9340), 
        .QN(n294) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n6532), .CK(CLK), .RN(n3245), .Q(n9341), 
        .QN(n295) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n6533), .CK(CLK), .RN(n3245), .Q(n9342), 
        .QN(n296) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n6534), .CK(CLK), .RN(n3245), .Q(n9343), 
        .QN(n297) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n6535), .CK(CLK), .RN(n3245), .Q(n9344), 
        .QN(n298) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n6536), .CK(CLK), .RN(n3245), .Q(n9345), 
        .QN(n299) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n6537), .CK(CLK), .RN(n3243), .Q(n9346), 
        .QN(n300) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n6538), .CK(CLK), .RN(n3243), .Q(n9347), 
        .QN(n301) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n6539), .CK(CLK), .RN(n3243), .Q(n9348), 
        .QN(n302) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n6540), .CK(CLK), .RN(n3243), .Q(n9349), 
        .QN(n303) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n6541), .CK(CLK), .RN(n3243), .Q(n9350), 
        .QN(n304) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n6542), .CK(CLK), .RN(n3243), .Q(n9351), 
        .QN(n305) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n6543), .CK(CLK), .RN(n3243), .Q(n9352), 
        .QN(n306) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n6544), .CK(CLK), .RN(n3243), .Q(n9353), 
        .QN(n307) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n6545), .CK(CLK), .RN(n3243), .Q(n9354), 
        .QN(n308) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n6546), .CK(CLK), .RN(n3243), .Q(n9355), 
        .QN(n309) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n6547), .CK(CLK), .RN(n3243), .Q(n9356), 
        .QN(n310) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n6548), .CK(CLK), .RN(n3243), .Q(n9357), 
        .QN(n311) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n6549), .CK(CLK), .RN(n3241), .Q(n9358), 
        .QN(n312) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n6550), .CK(CLK), .RN(n3241), .Q(n9359), 
        .QN(n313) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n6551), .CK(CLK), .RN(n3241), .Q(n9360), 
        .QN(n314) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n6552), .CK(CLK), .RN(n3241), .Q(n9361), 
        .QN(n315) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n6553), .CK(CLK), .RN(n3241), .Q(n9362), 
        .QN(n316) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n6554), .CK(CLK), .RN(n3241), .Q(n9363), 
        .QN(n317) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n6555), .CK(CLK), .RN(n3241), .Q(n9364), 
        .QN(n318) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n6556), .CK(CLK), .RN(n3241), .Q(n9365), 
        .QN(n319) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n6557), .CK(CLK), .RN(n3241), .Q(n9366), 
        .QN(n320) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n6558), .CK(CLK), .RN(n3241), .Q(n9367), 
        .QN(n321) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n6559), .CK(CLK), .RN(n3241), .Q(n9368), 
        .QN(n322) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n6560), .CK(CLK), .RN(n3241), .Q(n9369), 
        .QN(n323) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n6561), .CK(CLK), .RN(n3240), .Q(n9370), 
        .QN(n324) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n6562), .CK(CLK), .RN(n3240), .Q(n9371), 
        .QN(n325) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n6563), .CK(CLK), .RN(n3240), .Q(n9372), 
        .QN(n326) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n6564), .CK(CLK), .RN(n3240), .Q(n9373), 
        .QN(n327) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n6565), .CK(CLK), .RN(n3240), .Q(n9374), 
        .QN(n328) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n6566), .CK(CLK), .RN(n3240), .Q(n9375), 
        .QN(n329) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n6567), .CK(CLK), .RN(n3240), .Q(n9376), 
        .QN(n330) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n6568), .CK(CLK), .RN(n3240), .Q(n9377), 
        .QN(n331) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n6569), .CK(CLK), .RN(n3240), .Q(n9378), 
        .QN(n332) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n6570), .CK(CLK), .RN(n3240), .Q(n9379), 
        .QN(n333) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n6571), .CK(CLK), .RN(n3240), .Q(n9380), 
        .QN(n334) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n6572), .CK(CLK), .RN(n3240), .Q(n9381), 
        .QN(n335) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n6573), .CK(CLK), .RN(n3239), .Q(n9382), 
        .QN(n336) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n6574), .CK(CLK), .RN(n3239), .Q(n9383), 
        .QN(n337) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n6575), .CK(CLK), .RN(n3239), .Q(n9384), 
        .QN(n338) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n6576), .CK(CLK), .RN(n3239), .Q(n9385), 
        .QN(n339) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n6577), .CK(CLK), .RN(n3239), .Q(n9386), 
        .QN(n340) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n6578), .CK(CLK), .RN(n3239), .Q(n9387), 
        .QN(n341) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n6579), .CK(CLK), .RN(n3239), .Q(n9388), 
        .QN(n342) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n6580), .CK(CLK), .RN(n3239), .Q(n9389), 
        .QN(n343) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n6581), .CK(CLK), .RN(n3239), .Q(n9390), 
        .QN(n344) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n6582), .CK(CLK), .RN(n3239), .Q(n9391), 
        .QN(n345) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n6583), .CK(CLK), .RN(n3239), .Q(n9392), 
        .QN(n346) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n6584), .CK(CLK), .RN(n3239), .Q(n9393), 
        .QN(n347) );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n6585), .CK(CLK), .RN(n3237), .Q(n9394), 
        .QN(n348) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n6586), .CK(CLK), .RN(n3237), .Q(n9395), 
        .QN(n349) );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n6587), .CK(CLK), .RN(n3237), .Q(n9396), 
        .QN(n350) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n6588), .CK(CLK), .RN(n3237), .Q(n9397), 
        .QN(n351) );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n6589), .CK(CLK), .RN(n3237), .Q(n9398), 
        .QN(n352) );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n6590), .CK(CLK), .RN(n3237), .Q(n9399), 
        .QN(n353) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n6591), .CK(CLK), .RN(n3237), .Q(n9400), 
        .QN(n354) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n6592), .CK(CLK), .RN(n3237), .Q(n9401), 
        .QN(n355) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n6593), .CK(CLK), .RN(n3237), .Q(n9402), 
        .QN(n356) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n6594), .CK(CLK), .RN(n3237), .Q(n9403), 
        .QN(n357) );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n6595), .CK(CLK), .RN(n3237), .Q(n9404), 
        .QN(n358) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n6596), .CK(CLK), .RN(n3237), .Q(n9405), 
        .QN(n359) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n6597), .CK(CLK), .RN(n3236), .Q(n9406), 
        .QN(n360) );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n6598), .CK(CLK), .RN(n3236), .Q(n9407), 
        .QN(n361) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n6599), .CK(CLK), .RN(n3236), .Q(n9408), 
        .QN(n362) );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n6600), .CK(CLK), .RN(n3236), .Q(n9409), 
        .QN(n363) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n6601), .CK(CLK), .RN(n3236), .Q(n9410), 
        .QN(n364) );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n6602), .CK(CLK), .RN(n3236), .Q(n9411), 
        .QN(n365) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n6603), .CK(CLK), .RN(n3236), .Q(n9412), 
        .QN(n366) );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n6604), .CK(CLK), .RN(n3236), .Q(n9413), 
        .QN(n367) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n6605), .CK(CLK), .RN(n3236), .Q(n9414), 
        .QN(n368) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n6606), .CK(CLK), .RN(n3236), .Q(n9415), 
        .QN(n369) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n6607), .CK(CLK), .RN(n3236), .Q(n9416), 
        .QN(n370) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n6608), .CK(CLK), .RN(n3236), .Q(n9417), 
        .QN(n371) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n6609), .CK(CLK), .RN(n3235), .Q(n9418), 
        .QN(n372) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n6610), .CK(CLK), .RN(n3235), .Q(n9419), 
        .QN(n373) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n6611), .CK(CLK), .RN(n3235), .Q(n9420), 
        .QN(n374) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n6612), .CK(CLK), .RN(n3235), .Q(n9421), 
        .QN(n375) );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n6613), .CK(CLK), .RN(n3235), .Q(n9422), 
        .QN(n376) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n6614), .CK(CLK), .RN(n3235), .Q(n9423), 
        .QN(n377) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n6615), .CK(CLK), .RN(n3235), .Q(n9424), 
        .QN(n378) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n6616), .CK(CLK), .RN(n3235), .Q(n9425), 
        .QN(n379) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n6617), .CK(CLK), .RN(n3235), .Q(n9426), 
        .QN(n380) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n6618), .CK(CLK), .RN(n3235), .Q(n9427), 
        .QN(n381) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n6619), .CK(CLK), .RN(n3235), .Q(n9428), 
        .QN(n382) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n6620), .CK(CLK), .RN(n3235), .Q(n9429), 
        .QN(n383) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n6621), .CK(CLK), .RN(n3233), .Q(n9430), 
        .QN(n384) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n6622), .CK(CLK), .RN(n3233), .Q(n9431), 
        .QN(n385) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n6623), .CK(CLK), .RN(n3233), .Q(n9432), 
        .QN(n386) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n6624), .CK(CLK), .RN(n3233), .Q(n9433), 
        .QN(n387) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n6625), .CK(CLK), .RN(n3233), .Q(n9434), 
        .QN(n388) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n6626), .CK(CLK), .RN(n3233), .Q(n9435), 
        .QN(n389) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n6627), .CK(CLK), .RN(n3233), .Q(n9436), 
        .QN(n390) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n6628), .CK(CLK), .RN(n3233), .Q(n9437), 
        .QN(n391) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n6629), .CK(CLK), .RN(n3233), .Q(n9438), 
        .QN(n392) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n6630), .CK(CLK), .RN(n3233), .Q(n9439), 
        .QN(n393) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n6631), .CK(CLK), .RN(n3233), .Q(n9440), 
        .QN(n394) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n6632), .CK(CLK), .RN(n3233), .Q(n9441), 
        .QN(n395) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n6633), .CK(CLK), .RN(n3232), .Q(n9442), 
        .QN(n396) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n6634), .CK(CLK), .RN(n3232), .Q(n9443), 
        .QN(n397) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n6635), .CK(CLK), .RN(n3232), .Q(n9444), 
        .QN(n398) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n6636), .CK(CLK), .RN(n3232), .Q(n9445), 
        .QN(n399) );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n6637), .CK(CLK), .RN(n3232), .Q(n9446), 
        .QN(n400) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n6638), .CK(CLK), .RN(n3232), .Q(n9447), 
        .QN(n401) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n6639), .CK(CLK), .RN(n3232), .Q(n9448), 
        .QN(n402) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n6640), .CK(CLK), .RN(n3232), .Q(n9449), 
        .QN(n403) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n6641), .CK(CLK), .RN(n3232), .Q(n9450), 
        .QN(n404) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n6642), .CK(CLK), .RN(n3232), .Q(n9451), 
        .QN(n405) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n6643), .CK(CLK), .RN(n3232), .Q(n9452), 
        .QN(n406) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n6644), .CK(CLK), .RN(n3232), .Q(n9453), 
        .QN(n407) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n6645), .CK(CLK), .RN(n3231), .Q(n9454), 
        .QN(n408) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n6646), .CK(CLK), .RN(n3231), .Q(n9455), 
        .QN(n409) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n6647), .CK(CLK), .RN(n3231), .Q(n9456), 
        .QN(n410) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n6648), .CK(CLK), .RN(n3231), .Q(n9457), 
        .QN(n411) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n6649), .CK(CLK), .RN(n3231), .Q(n9458), 
        .QN(n412) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n6650), .CK(CLK), .RN(n3231), .Q(n9459), 
        .QN(n413) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n6651), .CK(CLK), .RN(n3231), .Q(n9460), 
        .QN(n414) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n6652), .CK(CLK), .RN(n3231), .Q(n9461), 
        .QN(n415) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n6653), .CK(CLK), .RN(n3231), .Q(n9462), 
        .QN(n416) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n6654), .CK(CLK), .RN(n3231), .Q(n9463), 
        .QN(n417) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n6655), .CK(CLK), .RN(n3231), .Q(n9464), 
        .QN(n418) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n6656), .CK(CLK), .RN(n3231), .Q(n9465), 
        .QN(n419) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n6657), .CK(CLK), .RN(n3229), .Q(n9466), 
        .QN(n420) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n6658), .CK(CLK), .RN(n3229), .Q(n9467), 
        .QN(n421) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n6659), .CK(CLK), .RN(n3229), .Q(n9468), 
        .QN(n422) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n6660), .CK(CLK), .RN(n3229), .Q(n9469), 
        .QN(n423) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n6661), .CK(CLK), .RN(n3229), .Q(n9470), 
        .QN(n424) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n6662), .CK(CLK), .RN(n3229), .Q(n9471), 
        .QN(n425) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n6663), .CK(CLK), .RN(n3229), .Q(n9472), 
        .QN(n426) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n6664), .CK(CLK), .RN(n3229), .Q(n9473), 
        .QN(n427) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n6665), .CK(CLK), .RN(n3229), .Q(n9474), 
        .QN(n428) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n6666), .CK(CLK), .RN(n3229), .Q(n9475), 
        .QN(n429) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n6667), .CK(CLK), .RN(n3229), .Q(n9476), 
        .QN(n430) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n6668), .CK(CLK), .RN(n3229), .Q(n9477), 
        .QN(n431) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n6733), .CK(CLK), .RN(n3221), .Q(n9478), 
        .QN(n496) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n6734), .CK(CLK), .RN(n3221), .Q(n9479), 
        .QN(n497) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n6735), .CK(CLK), .RN(n3221), .Q(n9480), 
        .QN(n498) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n6736), .CK(CLK), .RN(n3221), .Q(n9481), 
        .QN(n499) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n6737), .CK(CLK), .RN(n3221), .Q(n9482), 
        .QN(n500) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n6738), .CK(CLK), .RN(n3221), .Q(n9483), 
        .QN(n501) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n6739), .CK(CLK), .RN(n3221), .Q(n9484), 
        .QN(n502) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n6740), .CK(CLK), .RN(n3221), .Q(n9485), 
        .QN(n503) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n6741), .CK(CLK), .RN(n3220), .Q(n9486), 
        .QN(n504) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n6742), .CK(CLK), .RN(n3220), .Q(n9487), 
        .QN(n505) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n6743), .CK(CLK), .RN(n3220), .Q(n9488), 
        .QN(n506) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n6744), .CK(CLK), .RN(n3220), .Q(n9489), 
        .QN(n507) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n6745), .CK(CLK), .RN(n3220), .Q(n9490), 
        .QN(n508) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n6746), .CK(CLK), .RN(n3220), .Q(n9491), 
        .QN(n509) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n6747), .CK(CLK), .RN(n3220), .Q(n9492), 
        .QN(n510) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n6748), .CK(CLK), .RN(n3220), .Q(n9493), 
        .QN(n511) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n6749), .CK(CLK), .RN(n3220), .Q(n9494), 
        .QN(n512) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n6750), .CK(CLK), .RN(n3220), .Q(n9495), 
        .QN(n513) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n6751), .CK(CLK), .RN(n3220), .Q(n9496), 
        .QN(n514) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n6752), .CK(CLK), .RN(n3220), .Q(n9497), 
        .QN(n515) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n6753), .CK(CLK), .RN(n3219), .Q(n9498), 
        .QN(n516) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n6754), .CK(CLK), .RN(n3219), .Q(n9499), 
        .QN(n517) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n6755), .CK(CLK), .RN(n3219), .Q(n9500), 
        .QN(n518) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n6756), .CK(CLK), .RN(n3219), .Q(n9501), 
        .QN(n519) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n6757), .CK(CLK), .RN(n3219), .Q(n9502), 
        .QN(n520) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n6758), .CK(CLK), .RN(n3219), .Q(n9503), 
        .QN(n521) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n6759), .CK(CLK), .RN(n3219), .Q(n9504), 
        .QN(n522) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n6760), .CK(CLK), .RN(n3219), .Q(n9505), 
        .QN(n523) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n6761), .CK(CLK), .RN(n3219), .Q(n9506), 
        .QN(n524) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n6762), .CK(CLK), .RN(n3219), .Q(n9507), 
        .QN(n525) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n6763), .CK(CLK), .RN(n3219), .Q(n9508), 
        .QN(n526) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n6764), .CK(CLK), .RN(n3219), .Q(n9509), 
        .QN(n527) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n6765), .CK(CLK), .RN(n3217), .Q(n9510), 
        .QN(n528) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n6766), .CK(CLK), .RN(n3217), .Q(n9511), 
        .QN(n529) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n6767), .CK(CLK), .RN(n3217), .Q(n9512), 
        .QN(n530) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n6768), .CK(CLK), .RN(n3217), .Q(n9513), 
        .QN(n531) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n6769), .CK(CLK), .RN(n3217), .Q(n9514), 
        .QN(n532) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n6770), .CK(CLK), .RN(n3217), .Q(n9515), 
        .QN(n533) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n6771), .CK(CLK), .RN(n3217), .Q(n9516), 
        .QN(n534) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n6772), .CK(CLK), .RN(n3217), .Q(n9517), 
        .QN(n535) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n6773), .CK(CLK), .RN(n3217), .Q(n9518), 
        .QN(n536) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n6774), .CK(CLK), .RN(n3217), .Q(n9519), 
        .QN(n537) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n6775), .CK(CLK), .RN(n3217), .Q(n9520), 
        .QN(n538) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n6776), .CK(CLK), .RN(n3217), .Q(n9521), 
        .QN(n539) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n6777), .CK(CLK), .RN(n3216), .Q(n9522), 
        .QN(n540) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n6778), .CK(CLK), .RN(n3216), .Q(n9523), 
        .QN(n541) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n6779), .CK(CLK), .RN(n3216), .Q(n9524), 
        .QN(n542) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n6780), .CK(CLK), .RN(n3216), .Q(n9525), 
        .QN(n543) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n6781), .CK(CLK), .RN(n3216), .Q(n9526), 
        .QN(n544) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n6782), .CK(CLK), .RN(n3216), .Q(n9527), 
        .QN(n545) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n6783), .CK(CLK), .RN(n3216), .Q(n9528), 
        .QN(n546) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n6784), .CK(CLK), .RN(n3216), .Q(n9529), 
        .QN(n547) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n6785), .CK(CLK), .RN(n3216), .Q(n9530), 
        .QN(n548) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n6786), .CK(CLK), .RN(n3216), .Q(n9531), 
        .QN(n549) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n6787), .CK(CLK), .RN(n3216), .Q(n9532), 
        .QN(n550) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n6788), .CK(CLK), .RN(n3216), .Q(n9533), 
        .QN(n551) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n6789), .CK(CLK), .RN(n3215), .Q(n9534), 
        .QN(n552) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n6790), .CK(CLK), .RN(n3215), .Q(n9535), 
        .QN(n553) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n6791), .CK(CLK), .RN(n3215), .Q(n9536), 
        .QN(n554) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n6792), .CK(CLK), .RN(n3215), .Q(n9537), 
        .QN(n555) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n6793), .CK(CLK), .RN(n3215), .Q(n9538), 
        .QN(n556) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n6794), .CK(CLK), .RN(n3215), .Q(n9539), 
        .QN(n557) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n6795), .CK(CLK), .RN(n3215), .Q(n9540), 
        .QN(n558) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n6796), .CK(CLK), .RN(n3215), .Q(n9541), 
        .QN(n559) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n6797), .CK(CLK), .RN(n3215), .Q(n9542), 
        .QN(n560) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n6798), .CK(CLK), .RN(n3215), .Q(n9543), 
        .QN(n561) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n6799), .CK(CLK), .RN(n3215), .Q(n9544), 
        .QN(n562) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n6800), .CK(CLK), .RN(n3215), .Q(n9545), 
        .QN(n563) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n6801), .CK(CLK), .RN(n3213), .Q(n9546), 
        .QN(n564) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n6802), .CK(CLK), .RN(n3213), .Q(n9547), 
        .QN(n565) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n6803), .CK(CLK), .RN(n3213), .Q(n9548), 
        .QN(n566) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n6804), .CK(CLK), .RN(n3213), .Q(n9549), 
        .QN(n567) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n6805), .CK(CLK), .RN(n3213), .Q(n9550), 
        .QN(n568) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n6806), .CK(CLK), .RN(n3213), .Q(n9551), 
        .QN(n569) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n6807), .CK(CLK), .RN(n3213), .Q(n9552), 
        .QN(n570) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n6808), .CK(CLK), .RN(n3213), .Q(n9553), 
        .QN(n571) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n6809), .CK(CLK), .RN(n3213), .Q(n9554), 
        .QN(n572) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n6810), .CK(CLK), .RN(n3213), .Q(n9555), 
        .QN(n573) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n6811), .CK(CLK), .RN(n3213), .Q(n9556), 
        .QN(n574) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n6812), .CK(CLK), .RN(n3213), .Q(n9557), 
        .QN(n575) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n6813), .CK(CLK), .RN(n3212), .Q(n9558), 
        .QN(n576) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n6814), .CK(CLK), .RN(n3212), .Q(n9559), 
        .QN(n577) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n6815), .CK(CLK), .RN(n3212), .Q(n9560), 
        .QN(n578) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n6816), .CK(CLK), .RN(n3212), .Q(n9561), 
        .QN(n579) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n6817), .CK(CLK), .RN(n3212), .Q(n9562), 
        .QN(n580) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n6818), .CK(CLK), .RN(n3212), .Q(n9563), 
        .QN(n581) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n6819), .CK(CLK), .RN(n3212), .Q(n9564), 
        .QN(n582) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n6820), .CK(CLK), .RN(n3212), .Q(n9565), 
        .QN(n583) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n6821), .CK(CLK), .RN(n3212), .Q(n9566), 
        .QN(n584) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n6822), .CK(CLK), .RN(n3212), .Q(n9567), 
        .QN(n585) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n6823), .CK(CLK), .RN(n3212), .Q(n9568), 
        .QN(n586) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n6824), .CK(CLK), .RN(n3212), .Q(n9569), 
        .QN(n587) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n6825), .CK(CLK), .RN(n3211), .Q(n9570), 
        .QN(n588) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n6826), .CK(CLK), .RN(n3211), .Q(n9571), 
        .QN(n589) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n6827), .CK(CLK), .RN(n3211), .Q(n9572), 
        .QN(n590) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n6828), .CK(CLK), .RN(n3211), .Q(n9573), 
        .QN(n591) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n7021), .CK(CLK), .RN(n3189), .Q(n9574), 
        .QN(n784) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n7022), .CK(CLK), .RN(n3189), .Q(n9575), 
        .QN(n785) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n7023), .CK(CLK), .RN(n3189), .Q(n9576), 
        .QN(n786) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n7024), .CK(CLK), .RN(n3189), .Q(n9577), 
        .QN(n787) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n7025), .CK(CLK), .RN(n3189), .Q(n9578), 
        .QN(n788) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n7026), .CK(CLK), .RN(n3189), .Q(n9579), 
        .QN(n789) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n7027), .CK(CLK), .RN(n3189), .Q(n9580), 
        .QN(n790) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n7028), .CK(CLK), .RN(n3189), .Q(n9581), 
        .QN(n791) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n7029), .CK(CLK), .RN(n3188), .Q(n9582), 
        .QN(n792) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n7030), .CK(CLK), .RN(n3188), .Q(n9583), 
        .QN(n793) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n7031), .CK(CLK), .RN(n3188), .Q(n9584), 
        .QN(n794) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n7032), .CK(CLK), .RN(n3188), .Q(n9585), 
        .QN(n795) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n7033), .CK(CLK), .RN(n3188), .Q(n9586), 
        .QN(n796) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n7034), .CK(CLK), .RN(n3188), .Q(n9587), 
        .QN(n797) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n7035), .CK(CLK), .RN(n3188), .Q(n9588), 
        .QN(n798) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n7036), .CK(CLK), .RN(n3188), .Q(n9589), 
        .QN(n799) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n7037), .CK(CLK), .RN(n3188), .Q(n9590), 
        .QN(n800) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n7038), .CK(CLK), .RN(n3188), .Q(n9591), 
        .QN(n801) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n7039), .CK(CLK), .RN(n3188), .Q(n9592), 
        .QN(n802) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n7040), .CK(CLK), .RN(n3188), .Q(n9593), 
        .QN(n803) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n7041), .CK(CLK), .RN(n3187), .Q(n9594), 
        .QN(n804) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n7042), .CK(CLK), .RN(n3187), .Q(n9595), 
        .QN(n805) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n7043), .CK(CLK), .RN(n3187), .Q(n9596), 
        .QN(n806) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n7044), .CK(CLK), .RN(n3187), .Q(n9597), 
        .QN(n807) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n7045), .CK(CLK), .RN(n3187), .Q(n9598), 
        .QN(n808) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n7046), .CK(CLK), .RN(n3187), .Q(n9599), 
        .QN(n809) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n7047), .CK(CLK), .RN(n3187), .Q(n9600), 
        .QN(n810) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n7048), .CK(CLK), .RN(n3187), .Q(n9601), 
        .QN(n811) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n7049), .CK(CLK), .RN(n3187), .Q(n9602), 
        .QN(n812) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n7050), .CK(CLK), .RN(n3187), .Q(n9603), 
        .QN(n813) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n7051), .CK(CLK), .RN(n3187), .Q(n9604), 
        .QN(n814) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n7052), .CK(CLK), .RN(n3187), .Q(n9605), 
        .QN(n815) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n7053), .CK(CLK), .RN(n3185), .Q(n9606), 
        .QN(n816) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n7054), .CK(CLK), .RN(n3185), .Q(n9607), 
        .QN(n817) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n7055), .CK(CLK), .RN(n3185), .Q(n9608), 
        .QN(n818) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n7056), .CK(CLK), .RN(n3185), .Q(n9609), 
        .QN(n819) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n7057), .CK(CLK), .RN(n3185), .Q(n9610), 
        .QN(n820) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n7058), .CK(CLK), .RN(n3185), .Q(n9611), 
        .QN(n821) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n7059), .CK(CLK), .RN(n3185), .Q(n9612), 
        .QN(n822) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n7060), .CK(CLK), .RN(n3185), .Q(n9613), 
        .QN(n823) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n7061), .CK(CLK), .RN(n3185), .Q(n9614), 
        .QN(n824) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n7062), .CK(CLK), .RN(n3185), .Q(n9615), 
        .QN(n825) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n7063), .CK(CLK), .RN(n3185), .Q(n9616), 
        .QN(n826) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n7064), .CK(CLK), .RN(n3185), .Q(n9617), 
        .QN(n827) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n7065), .CK(CLK), .RN(n3184), .Q(n9618), 
        .QN(n828) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n7066), .CK(CLK), .RN(n3184), .Q(n9619), 
        .QN(n829) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n7067), .CK(CLK), .RN(n3184), .Q(n9620), 
        .QN(n830) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n7068), .CK(CLK), .RN(n3184), .Q(n9621), 
        .QN(n831) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n7069), .CK(CLK), .RN(n3184), .Q(n9622), 
        .QN(n832) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n7070), .CK(CLK), .RN(n3184), .Q(n9623), 
        .QN(n833) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n7071), .CK(CLK), .RN(n3184), .Q(n9624), 
        .QN(n834) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n7072), .CK(CLK), .RN(n3184), .Q(n9625), 
        .QN(n835) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n7073), .CK(CLK), .RN(n3184), .Q(n9626), 
        .QN(n836) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n7074), .CK(CLK), .RN(n3184), .Q(n9627), 
        .QN(n837) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n7075), .CK(CLK), .RN(n3184), .Q(n9628), 
        .QN(n838) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n7076), .CK(CLK), .RN(n3184), .Q(n9629), 
        .QN(n839) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n7077), .CK(CLK), .RN(n3183), .Q(n9630), 
        .QN(n840) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n7078), .CK(CLK), .RN(n3183), .Q(n9631), 
        .QN(n841) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n7079), .CK(CLK), .RN(n3183), .Q(n9632), 
        .QN(n842) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n7080), .CK(CLK), .RN(n3183), .Q(n9633), 
        .QN(n843) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n7081), .CK(CLK), .RN(n3183), .Q(n9634), 
        .QN(n844) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n7082), .CK(CLK), .RN(n3183), .Q(n9635), 
        .QN(n845) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n7083), .CK(CLK), .RN(n3183), .Q(n9636), 
        .QN(n846) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n7084), .CK(CLK), .RN(n3183), .Q(n9637), 
        .QN(n847) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n7085), .CK(CLK), .RN(n3183), .Q(n9638), 
        .QN(n848) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n7086), .CK(CLK), .RN(n3183), .Q(n9639), 
        .QN(n849) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n7087), .CK(CLK), .RN(n3183), .Q(n9640), 
        .QN(n850) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n7088), .CK(CLK), .RN(n3183), .Q(n9641), 
        .QN(n851) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n7089), .CK(CLK), .RN(n3181), .Q(n9642), 
        .QN(n852) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n7090), .CK(CLK), .RN(n3181), .Q(n9643), 
        .QN(n853) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n7091), .CK(CLK), .RN(n3181), .Q(n9644), 
        .QN(n854) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n7092), .CK(CLK), .RN(n3181), .Q(n9645), 
        .QN(n855) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n7093), .CK(CLK), .RN(n3181), .Q(n9646), 
        .QN(n856) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n7094), .CK(CLK), .RN(n3181), .Q(n9647), 
        .QN(n857) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n7095), .CK(CLK), .RN(n3181), .Q(n9648), 
        .QN(n858) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n7096), .CK(CLK), .RN(n3181), .Q(n9649), 
        .QN(n859) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n7097), .CK(CLK), .RN(n3181), .Q(n9650), 
        .QN(n860) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n7098), .CK(CLK), .RN(n3181), .Q(n9651), 
        .QN(n861) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n7099), .CK(CLK), .RN(n3181), .Q(n9652), 
        .QN(n862) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n7100), .CK(CLK), .RN(n3181), .Q(n9653), 
        .QN(n863) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n7101), .CK(CLK), .RN(n3180), .Q(n9654), 
        .QN(n864) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n7102), .CK(CLK), .RN(n3180), .Q(n9655), 
        .QN(n865) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n7103), .CK(CLK), .RN(n3180), .Q(n9656), 
        .QN(n866) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n7104), .CK(CLK), .RN(n3180), .Q(n9657), 
        .QN(n867) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n7105), .CK(CLK), .RN(n3180), .Q(n9658), 
        .QN(n868) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n7106), .CK(CLK), .RN(n3180), .Q(n9659), 
        .QN(n869) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n7107), .CK(CLK), .RN(n3180), .Q(n9660), 
        .QN(n870) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n7108), .CK(CLK), .RN(n3180), .Q(n9661), 
        .QN(n871) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n7109), .CK(CLK), .RN(n3180), .Q(n9662), 
        .QN(n872) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n7110), .CK(CLK), .RN(n3180), .Q(n9663), 
        .QN(n873) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n7111), .CK(CLK), .RN(n3180), .Q(n9664), 
        .QN(n874) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n7112), .CK(CLK), .RN(n3180), .Q(n9665), 
        .QN(n875) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n7113), .CK(CLK), .RN(n3178), .Q(n9666), 
        .QN(n876) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n7114), .CK(CLK), .RN(n3178), .Q(n9667), 
        .QN(n877) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n7115), .CK(CLK), .RN(n3178), .Q(n9668), 
        .QN(n878) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n7116), .CK(CLK), .RN(n3178), .Q(n9669), 
        .QN(n879) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n7117), .CK(CLK), .RN(n3178), .Q(n9670), 
        .QN(n880) );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n7118), .CK(CLK), .RN(n3178), .Q(n9671), 
        .QN(n881) );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n7119), .CK(CLK), .RN(n3178), .Q(n9672), 
        .QN(n882) );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n7120), .CK(CLK), .RN(n3178), .Q(n9673), 
        .QN(n883) );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n7121), .CK(CLK), .RN(n3178), .Q(n9674), 
        .QN(n884) );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n7122), .CK(CLK), .RN(n3178), .Q(n9675), 
        .QN(n885) );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n7123), .CK(CLK), .RN(n3178), .Q(n9676), 
        .QN(n886) );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n7124), .CK(CLK), .RN(n3178), .Q(n9677), 
        .QN(n887) );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n7125), .CK(CLK), .RN(n3176), .Q(n9678), 
        .QN(n888) );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n7126), .CK(CLK), .RN(n3176), .Q(n9679), 
        .QN(n889) );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n7127), .CK(CLK), .RN(n3176), .Q(n9680), 
        .QN(n890) );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n7128), .CK(CLK), .RN(n3176), .Q(n9681), 
        .QN(n891) );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n7129), .CK(CLK), .RN(n3176), .Q(n9682), 
        .QN(n892) );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n7130), .CK(CLK), .RN(n3176), .Q(n9683), 
        .QN(n893) );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n7131), .CK(CLK), .RN(n3176), .Q(n9684), 
        .QN(n894) );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n7132), .CK(CLK), .RN(n3176), .Q(n9685), 
        .QN(n895) );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n7133), .CK(CLK), .RN(n3176), .Q(n9686), 
        .QN(n896) );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n7134), .CK(CLK), .RN(n3176), .Q(n9687), 
        .QN(n897) );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n7135), .CK(CLK), .RN(n3176), .Q(n9688), 
        .QN(n898) );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n7136), .CK(CLK), .RN(n3176), .Q(n9689), 
        .QN(n899) );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n7137), .CK(CLK), .RN(n3175), .Q(n9690), 
        .QN(n900) );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n7138), .CK(CLK), .RN(n3175), .Q(n9691), 
        .QN(n901) );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n7139), .CK(CLK), .RN(n3175), .Q(n9692), 
        .QN(n902) );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n7140), .CK(CLK), .RN(n3175), .Q(n9693), 
        .QN(n903) );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n7141), .CK(CLK), .RN(n3175), .Q(n9694), 
        .QN(n904) );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n7142), .CK(CLK), .RN(n3175), .Q(n9695), 
        .QN(n905) );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n7143), .CK(CLK), .RN(n3175), .Q(n9696), 
        .QN(n906) );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n7144), .CK(CLK), .RN(n3175), .Q(n9697), 
        .QN(n907) );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n7145), .CK(CLK), .RN(n3175), .Q(n9698), 
        .QN(n908) );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n7146), .CK(CLK), .RN(n3175), .Q(n9699), 
        .QN(n909) );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n7147), .CK(CLK), .RN(n3175), .Q(n9700), 
        .QN(n910) );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n7148), .CK(CLK), .RN(n3175), .Q(n9701), 
        .QN(n911) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n7149), .CK(CLK), .RN(n3174), .Q(n9702), 
        .QN(n912) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n7150), .CK(CLK), .RN(n3174), .Q(n9703), 
        .QN(n913) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n7151), .CK(CLK), .RN(n3174), .Q(n9704), 
        .QN(n914) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n7152), .CK(CLK), .RN(n3174), .Q(n9705), 
        .QN(n915) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n7153), .CK(CLK), .RN(n3174), .Q(n9706), 
        .QN(n916) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n7154), .CK(CLK), .RN(n3174), .Q(n9707), 
        .QN(n917) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n7155), .CK(CLK), .RN(n3174), .Q(n9708), 
        .QN(n918) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n7156), .CK(CLK), .RN(n3174), .Q(n9709), 
        .QN(n919) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n7157), .CK(CLK), .RN(n3174), .Q(n9710), 
        .QN(n920) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n7158), .CK(CLK), .RN(n3174), .Q(n9711), 
        .QN(n921) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n7159), .CK(CLK), .RN(n3174), .Q(n9712), 
        .QN(n922) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n7160), .CK(CLK), .RN(n3174), .Q(n9713), 
        .QN(n923) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n7161), .CK(CLK), .RN(n3172), .Q(n9714), 
        .QN(n924) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n7162), .CK(CLK), .RN(n3172), .Q(n9715), 
        .QN(n925) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n7163), .CK(CLK), .RN(n3172), .Q(n9716), 
        .QN(n926) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n7164), .CK(CLK), .RN(n3172), .Q(n9717), 
        .QN(n927) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n7165), .CK(CLK), .RN(n3172), .Q(n9718), 
        .QN(n928) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n7166), .CK(CLK), .RN(n3172), .Q(n9719), 
        .QN(n929) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n7167), .CK(CLK), .RN(n3172), .Q(n9720), 
        .QN(n930) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n7168), .CK(CLK), .RN(n3172), .Q(n9721), 
        .QN(n931) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n7169), .CK(CLK), .RN(n3172), .Q(n9722), 
        .QN(n932) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n7170), .CK(CLK), .RN(n3172), .Q(n9723), 
        .QN(n933) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n7171), .CK(CLK), .RN(n3172), .Q(n9724), 
        .QN(n934) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n7172), .CK(CLK), .RN(n3172), .Q(n9725), 
        .QN(n935) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n7173), .CK(CLK), .RN(n3171), .Q(n9726), 
        .QN(n936) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n7174), .CK(CLK), .RN(n3171), .Q(n9727), 
        .QN(n937) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n7175), .CK(CLK), .RN(n3171), .Q(n9728), 
        .QN(n938) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n7176), .CK(CLK), .RN(n3171), .Q(n9729), 
        .QN(n939) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n7177), .CK(CLK), .RN(n3171), .Q(n9730), 
        .QN(n940) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n7178), .CK(CLK), .RN(n3171), .Q(n9731), 
        .QN(n941) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n7179), .CK(CLK), .RN(n3171), .Q(n9732), 
        .QN(n942) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n7180), .CK(CLK), .RN(n3171), .Q(n9733), 
        .QN(n943) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n7181), .CK(CLK), .RN(n3171), .Q(n9734), 
        .QN(n944) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n7182), .CK(CLK), .RN(n3171), .Q(n9735), 
        .QN(n945) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n7183), .CK(CLK), .RN(n3171), .Q(n9736), 
        .QN(n946) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n7184), .CK(CLK), .RN(n3171), .Q(n9737), 
        .QN(n947) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n7185), .CK(CLK), .RN(n3170), .Q(n9738), 
        .QN(n948) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n7186), .CK(CLK), .RN(n3170), .Q(n9739), 
        .QN(n949) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n7187), .CK(CLK), .RN(n3170), .Q(n9740), 
        .QN(n950) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n7188), .CK(CLK), .RN(n3170), .Q(n9741), 
        .QN(n951) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n7189), .CK(CLK), .RN(n3170), .Q(n9742), 
        .QN(n952) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n7190), .CK(CLK), .RN(n3170), .Q(n9743), 
        .QN(n953) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n7191), .CK(CLK), .RN(n3170), .Q(n9744), 
        .QN(n954) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n7192), .CK(CLK), .RN(n3170), .Q(n9745), 
        .QN(n955) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n7193), .CK(CLK), .RN(n3170), .Q(n9746), 
        .QN(n956) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n7194), .CK(CLK), .RN(n3170), .Q(n9747), 
        .QN(n957) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n7195), .CK(CLK), .RN(n3170), .Q(n9748), 
        .QN(n958) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n7196), .CK(CLK), .RN(n3170), .Q(n9749), 
        .QN(n959) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n7197), .CK(CLK), .RN(n3168), .Q(n9750), 
        .QN(n960) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n7198), .CK(CLK), .RN(n3168), .Q(n9751), 
        .QN(n961) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n7199), .CK(CLK), .RN(n3168), .Q(n9752), 
        .QN(n962) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n7200), .CK(CLK), .RN(n3168), .Q(n9753), 
        .QN(n963) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n7201), .CK(CLK), .RN(n3168), .Q(n9754), 
        .QN(n964) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n7202), .CK(CLK), .RN(n3168), .Q(n9755), 
        .QN(n965) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n7203), .CK(CLK), .RN(n3168), .Q(n9756), 
        .QN(n966) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n7204), .CK(CLK), .RN(n3168), .Q(n9757), 
        .QN(n967) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n7205), .CK(CLK), .RN(n3168), .Q(n9758), 
        .QN(n968) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n7206), .CK(CLK), .RN(n3168), .Q(n9759), 
        .QN(n969) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n7207), .CK(CLK), .RN(n3168), .Q(n9760), 
        .QN(n970) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n7208), .CK(CLK), .RN(n3168), .Q(n9761), 
        .QN(n971) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n7209), .CK(CLK), .RN(n3167), .Q(n9762), 
        .QN(n972) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n7210), .CK(CLK), .RN(n3167), .Q(n9763), 
        .QN(n973) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n7211), .CK(CLK), .RN(n3167), .Q(n9764), 
        .QN(n974) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n7212), .CK(CLK), .RN(n3167), .Q(n9765), 
        .QN(n975) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n7213), .CK(CLK), .RN(n3167), .Q(n9766), 
        .QN(n976) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n7214), .CK(CLK), .RN(n3167), .Q(n9767), 
        .QN(n977) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n7215), .CK(CLK), .RN(n3167), .Q(n9768), 
        .QN(n978) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n7216), .CK(CLK), .RN(n3167), .Q(n9769), 
        .QN(n979) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n7217), .CK(CLK), .RN(n3167), .Q(n9770), 
        .QN(n980) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n7218), .CK(CLK), .RN(n3167), .Q(n9771), 
        .QN(n981) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n7219), .CK(CLK), .RN(n3167), .Q(n9772), 
        .QN(n982) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n7220), .CK(CLK), .RN(n3167), .Q(n9773), 
        .QN(n983) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n7221), .CK(CLK), .RN(n3166), .Q(n9774), 
        .QN(n984) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n7222), .CK(CLK), .RN(n3166), .Q(n9775), 
        .QN(n985) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n7223), .CK(CLK), .RN(n3166), .Q(n9776), 
        .QN(n986) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n7224), .CK(CLK), .RN(n3166), .Q(n9777), 
        .QN(n987) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n7225), .CK(CLK), .RN(n3166), .Q(n9778), 
        .QN(n988) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n7226), .CK(CLK), .RN(n3166), .Q(n9779), 
        .QN(n989) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n7227), .CK(CLK), .RN(n3166), .Q(n9780), 
        .QN(n990) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n7228), .CK(CLK), .RN(n3166), .Q(n9781), 
        .QN(n991) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n7229), .CK(CLK), .RN(n3166), .Q(n9782), 
        .QN(n992) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n7230), .CK(CLK), .RN(n3166), .Q(n9783), 
        .QN(n993) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n7231), .CK(CLK), .RN(n3166), .Q(n9784), 
        .QN(n994) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n7232), .CK(CLK), .RN(n3166), .Q(n9785), 
        .QN(n995) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n7233), .CK(CLK), .RN(n3164), .Q(n9786), 
        .QN(n996) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n7234), .CK(CLK), .RN(n3164), .Q(n9787), 
        .QN(n997) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n7235), .CK(CLK), .RN(n3164), .Q(n9788), 
        .QN(n998) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n7236), .CK(CLK), .RN(n3164), .Q(n9789), 
        .QN(n999) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n7237), .CK(CLK), .RN(n3164), .Q(n9790), 
        .QN(n1000) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n7238), .CK(CLK), .RN(n3164), .Q(n9791), 
        .QN(n1001) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n7239), .CK(CLK), .RN(n3164), .Q(n9792), 
        .QN(n1002) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n7240), .CK(CLK), .RN(n3164), .Q(n9793), 
        .QN(n1003) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n7241), .CK(CLK), .RN(n3164), .Q(n9794), 
        .QN(n1004) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n7242), .CK(CLK), .RN(n3164), .Q(n9795), 
        .QN(n1005) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n7243), .CK(CLK), .RN(n3164), .Q(n9796), 
        .QN(n1006) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n7244), .CK(CLK), .RN(n3164), .Q(n9797), 
        .QN(n1007) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n7245), .CK(CLK), .RN(n3163), .Q(n9798), 
        .QN(n1008) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n7246), .CK(CLK), .RN(n3163), .Q(n9799), 
        .QN(n1009) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n7247), .CK(CLK), .RN(n3163), .Q(n9800), 
        .QN(n1010) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n7248), .CK(CLK), .RN(n3163), .Q(n9801), 
        .QN(n1011) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n7249), .CK(CLK), .RN(n3163), .Q(n9802), 
        .QN(n1012) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n7250), .CK(CLK), .RN(n3163), .Q(n9803), 
        .QN(n1013) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n7251), .CK(CLK), .RN(n3163), .Q(n9804), 
        .QN(n1014) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n7252), .CK(CLK), .RN(n3163), .Q(n9805), 
        .QN(n1015) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n7253), .CK(CLK), .RN(n3163), .Q(n9806), 
        .QN(n1016) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n7254), .CK(CLK), .RN(n3163), .Q(n9807), 
        .QN(n1017) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n7255), .CK(CLK), .RN(n3163), .Q(n9808), 
        .QN(n1018) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n7256), .CK(CLK), .RN(n3163), .Q(n9809), 
        .QN(n1019) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n7257), .CK(CLK), .RN(n3162), .Q(n9810), 
        .QN(n1020) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n7258), .CK(CLK), .RN(n3162), .Q(n9811), 
        .QN(n1021) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n7259), .CK(CLK), .RN(n3162), .Q(n9812), 
        .QN(n1022) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n7260), .CK(CLK), .RN(n3162), .Q(n9813), 
        .QN(n1023) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n7261), .CK(CLK), .RN(n3162), .Q(n9814), 
        .QN(n1024) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n7262), .CK(CLK), .RN(n3162), .Q(n9815), 
        .QN(n1025) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n7263), .CK(CLK), .RN(n3162), .Q(n9816), 
        .QN(n1026) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n7264), .CK(CLK), .RN(n3162), .Q(n9817), 
        .QN(n1027) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n7265), .CK(CLK), .RN(n3162), .Q(n9818), 
        .QN(n1028) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n7266), .CK(CLK), .RN(n3162), .Q(n9819), 
        .QN(n1029) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n7267), .CK(CLK), .RN(n3162), .Q(n9820), 
        .QN(n1030) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n7268), .CK(CLK), .RN(n3162), .Q(n9821), 
        .QN(n1031) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n7269), .CK(CLK), .RN(n3160), .Q(n9822), 
        .QN(n1032) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n7270), .CK(CLK), .RN(n3160), .Q(n9823), 
        .QN(n1033) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n7271), .CK(CLK), .RN(n3160), .Q(n9824), 
        .QN(n1034) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n7272), .CK(CLK), .RN(n3160), .Q(n9825), 
        .QN(n1035) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n7273), .CK(CLK), .RN(n3160), .Q(n9826), 
        .QN(n1036) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n7274), .CK(CLK), .RN(n3160), .Q(n9827), 
        .QN(n1037) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n7275), .CK(CLK), .RN(n3160), .Q(n9828), 
        .QN(n1038) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n7276), .CK(CLK), .RN(n3160), .Q(n9829), 
        .QN(n1039) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n7277), .CK(CLK), .RN(n3160), .Q(n9830), 
        .QN(n1040) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n7278), .CK(CLK), .RN(n3160), .Q(n9831), 
        .QN(n1041) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n7279), .CK(CLK), .RN(n3160), .Q(n9832), 
        .QN(n1042) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n7280), .CK(CLK), .RN(n3160), .Q(n9833), 
        .QN(n1043) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n7281), .CK(CLK), .RN(n3159), .Q(n9834), 
        .QN(n1044) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n7282), .CK(CLK), .RN(n3159), .Q(n9835), 
        .QN(n1045) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n7283), .CK(CLK), .RN(n3159), .Q(n9836), 
        .QN(n1046) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n7284), .CK(CLK), .RN(n3159), .Q(n9837), 
        .QN(n1047) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n7285), .CK(CLK), .RN(n3159), .Q(n9838), 
        .QN(n1048) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n7286), .CK(CLK), .RN(n3159), .Q(n9839), 
        .QN(n1049) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n7287), .CK(CLK), .RN(n3159), .Q(n9840), 
        .QN(n1050) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n7288), .CK(CLK), .RN(n3159), .Q(n9841), 
        .QN(n1051) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n7289), .CK(CLK), .RN(n3159), .Q(n9842), 
        .QN(n1052) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n7290), .CK(CLK), .RN(n3159), .Q(n9843), 
        .QN(n1053) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n7291), .CK(CLK), .RN(n3159), .Q(n9844), 
        .QN(n1054) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n7292), .CK(CLK), .RN(n3159), .Q(n9845), 
        .QN(n1055) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n7293), .CK(CLK), .RN(n3158), .Q(n9846), 
        .QN(n1056) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n7294), .CK(CLK), .RN(n3158), .Q(n9847), 
        .QN(n1057) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n7295), .CK(CLK), .RN(n3158), .Q(n9848), 
        .QN(n1058) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n7296), .CK(CLK), .RN(n3158), .Q(n9849), 
        .QN(n1059) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n7297), .CK(CLK), .RN(n3158), .Q(n9850), 
        .QN(n1060) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n7298), .CK(CLK), .RN(n3158), .Q(n9851), 
        .QN(n1061) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n7299), .CK(CLK), .RN(n3158), .Q(n9852), 
        .QN(n1062) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n7300), .CK(CLK), .RN(n3158), .Q(n9853), 
        .QN(n1063) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n7301), .CK(CLK), .RN(n3158), .Q(n9854), 
        .QN(n1064) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n7302), .CK(CLK), .RN(n3158), .Q(n9855), 
        .QN(n1065) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n7303), .CK(CLK), .RN(n3158), .Q(n9856), 
        .QN(n1066) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n7304), .CK(CLK), .RN(n3158), .Q(n9857), 
        .QN(n1067) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n7305), .CK(CLK), .RN(n3156), .Q(n9858), 
        .QN(n1068) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n7306), .CK(CLK), .RN(n3156), .Q(n9859), 
        .QN(n1069) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n7307), .CK(CLK), .RN(n3156), .Q(n9860), 
        .QN(n1070) );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n7308), .CK(CLK), .RN(n3156), .Q(n9861), 
        .QN(n1071) );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n7309), .CK(CLK), .RN(n3156), .Q(n9862), 
        .QN(n1072) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n7310), .CK(CLK), .RN(n3156), .Q(n9863), 
        .QN(n1073) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n7311), .CK(CLK), .RN(n3156), .Q(n9864), 
        .QN(n1074) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n7312), .CK(CLK), .RN(n3156), .Q(n9865), 
        .QN(n1075) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n7313), .CK(CLK), .RN(n3156), .Q(n9866), 
        .QN(n1076) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n7314), .CK(CLK), .RN(n3156), .Q(n9867), 
        .QN(n1077) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n7315), .CK(CLK), .RN(n3156), .Q(n9868), 
        .QN(n1078) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n7316), .CK(CLK), .RN(n3156), .Q(n9869), 
        .QN(n1079) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n7317), .CK(CLK), .RN(n3155), .Q(n9870), 
        .QN(n1080) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n7318), .CK(CLK), .RN(n3155), .Q(n9871), 
        .QN(n1081) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n7319), .CK(CLK), .RN(n3155), .Q(n9872), 
        .QN(n1082) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n7320), .CK(CLK), .RN(n3155), .Q(n9873), 
        .QN(n1083) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n7321), .CK(CLK), .RN(n3155), .Q(n9874), 
        .QN(n1084) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n7322), .CK(CLK), .RN(n3155), .Q(n9875), 
        .QN(n1085) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n7323), .CK(CLK), .RN(n3155), .Q(n9876), 
        .QN(n1086) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n7324), .CK(CLK), .RN(n3155), .Q(n9877), 
        .QN(n1087) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n7325), .CK(CLK), .RN(n3155), .Q(n9878), 
        .QN(n1088) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n7326), .CK(CLK), .RN(n3155), .Q(n9879), 
        .QN(n1089) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n7327), .CK(CLK), .RN(n3155), .Q(n9880), 
        .QN(n1090) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n7328), .CK(CLK), .RN(n3155), .Q(n9881), 
        .QN(n1091) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n7329), .CK(CLK), .RN(n3154), .Q(n9882), 
        .QN(n1092) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n7330), .CK(CLK), .RN(n3154), .Q(n9883), 
        .QN(n1093) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n7331), .CK(CLK), .RN(n3154), .Q(n9884), 
        .QN(n1094) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n7332), .CK(CLK), .RN(n3154), .Q(n9885), 
        .QN(n1095) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n7333), .CK(CLK), .RN(n3154), .Q(n9886), 
        .QN(n1096) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n7334), .CK(CLK), .RN(n3154), .Q(n9887), 
        .QN(n1097) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n7335), .CK(CLK), .RN(n3154), .Q(n9888), 
        .QN(n1098) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n7336), .CK(CLK), .RN(n3154), .Q(n9889), 
        .QN(n1099) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n7337), .CK(CLK), .RN(n3154), .Q(n9890), 
        .QN(n1100) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n7338), .CK(CLK), .RN(n3154), .Q(n9891), 
        .QN(n1101) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n7339), .CK(CLK), .RN(n3154), .Q(n9892), 
        .QN(n1102) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n7340), .CK(CLK), .RN(n3154), .Q(n9893), 
        .QN(n1103) );
  DFFR_X1 \REGISTERS_reg[32][31]  ( .D(n7341), .CK(CLK), .RN(n3152), .Q(n9894), 
        .QN(n1104) );
  DFFR_X1 \REGISTERS_reg[32][30]  ( .D(n7342), .CK(CLK), .RN(n3152), .Q(n9895), 
        .QN(n1105) );
  DFFR_X1 \REGISTERS_reg[32][29]  ( .D(n7343), .CK(CLK), .RN(n3152), .Q(n9896), 
        .QN(n1106) );
  DFFR_X1 \REGISTERS_reg[32][28]  ( .D(n7344), .CK(CLK), .RN(n3152), .Q(n9897), 
        .QN(n1107) );
  DFFR_X1 \REGISTERS_reg[32][27]  ( .D(n7345), .CK(CLK), .RN(n3152), .Q(n9898), 
        .QN(n1108) );
  DFFR_X1 \REGISTERS_reg[32][26]  ( .D(n7346), .CK(CLK), .RN(n3152), .Q(n9899), 
        .QN(n1109) );
  DFFR_X1 \REGISTERS_reg[32][25]  ( .D(n7347), .CK(CLK), .RN(n3152), .Q(n9900), 
        .QN(n1110) );
  DFFR_X1 \REGISTERS_reg[32][24]  ( .D(n7348), .CK(CLK), .RN(n3152), .Q(n9901), 
        .QN(n1111) );
  DFFR_X1 \REGISTERS_reg[32][23]  ( .D(n7349), .CK(CLK), .RN(n3152), .Q(n9902), 
        .QN(n1112) );
  DFFR_X1 \REGISTERS_reg[32][22]  ( .D(n7350), .CK(CLK), .RN(n3152), .Q(n9903), 
        .QN(n1113) );
  DFFR_X1 \REGISTERS_reg[32][21]  ( .D(n7351), .CK(CLK), .RN(n3152), .Q(n9904), 
        .QN(n1114) );
  DFFR_X1 \REGISTERS_reg[32][20]  ( .D(n7352), .CK(CLK), .RN(n3152), .Q(n9905), 
        .QN(n1115) );
  DFFR_X1 \REGISTERS_reg[32][19]  ( .D(n7353), .CK(CLK), .RN(n3151), .Q(n9906), 
        .QN(n1116) );
  DFFR_X1 \REGISTERS_reg[32][18]  ( .D(n7354), .CK(CLK), .RN(n3151), .Q(n9907), 
        .QN(n1117) );
  DFFR_X1 \REGISTERS_reg[32][17]  ( .D(n7355), .CK(CLK), .RN(n3151), .Q(n9908), 
        .QN(n1118) );
  DFFR_X1 \REGISTERS_reg[32][16]  ( .D(n7356), .CK(CLK), .RN(n3151), .Q(n9909), 
        .QN(n1119) );
  DFFR_X1 \REGISTERS_reg[32][15]  ( .D(n7357), .CK(CLK), .RN(n3151), .Q(n9910), 
        .QN(n1120) );
  DFFR_X1 \REGISTERS_reg[32][14]  ( .D(n7358), .CK(CLK), .RN(n3151), .Q(n9911), 
        .QN(n1121) );
  DFFR_X1 \REGISTERS_reg[32][13]  ( .D(n7359), .CK(CLK), .RN(n3151), .Q(n9912), 
        .QN(n1122) );
  DFFR_X1 \REGISTERS_reg[32][12]  ( .D(n7360), .CK(CLK), .RN(n3151), .Q(n9913), 
        .QN(n1123) );
  DFFR_X1 \REGISTERS_reg[32][11]  ( .D(n7361), .CK(CLK), .RN(n3151), .Q(n9914), 
        .QN(n1124) );
  DFFR_X1 \REGISTERS_reg[32][10]  ( .D(n7362), .CK(CLK), .RN(n3151), .Q(n9915), 
        .QN(n1125) );
  DFFR_X1 \REGISTERS_reg[32][9]  ( .D(n7363), .CK(CLK), .RN(n3151), .Q(n9916), 
        .QN(n1126) );
  DFFR_X1 \REGISTERS_reg[32][8]  ( .D(n7364), .CK(CLK), .RN(n3151), .Q(n9917), 
        .QN(n1127) );
  DFFR_X1 \REGISTERS_reg[32][7]  ( .D(n7365), .CK(CLK), .RN(n3150), .Q(n9918), 
        .QN(n1128) );
  DFFR_X1 \REGISTERS_reg[32][6]  ( .D(n7366), .CK(CLK), .RN(n3150), .Q(n9919), 
        .QN(n1129) );
  DFFR_X1 \REGISTERS_reg[32][5]  ( .D(n7367), .CK(CLK), .RN(n3150), .Q(n9920), 
        .QN(n1130) );
  DFFR_X1 \REGISTERS_reg[32][4]  ( .D(n7368), .CK(CLK), .RN(n3150), .Q(n9921), 
        .QN(n1131) );
  DFFR_X1 \REGISTERS_reg[32][3]  ( .D(n7369), .CK(CLK), .RN(n3150), .Q(n9922), 
        .QN(n1132) );
  DFFR_X1 \REGISTERS_reg[32][2]  ( .D(n7370), .CK(CLK), .RN(n3150), .Q(n9923), 
        .QN(n1133) );
  DFFR_X1 \REGISTERS_reg[32][1]  ( .D(n7371), .CK(CLK), .RN(n3150), .Q(n9924), 
        .QN(n1134) );
  DFFR_X1 \REGISTERS_reg[32][0]  ( .D(n7372), .CK(CLK), .RN(n3150), .Q(n9925), 
        .QN(n1135) );
  DFFR_X1 \REGISTERS_reg[35][31]  ( .D(n7437), .CK(CLK), .RN(n3142), .Q(n9926), 
        .QN(n1200) );
  DFFR_X1 \REGISTERS_reg[35][30]  ( .D(n7438), .CK(CLK), .RN(n3142), .Q(n9927), 
        .QN(n1201) );
  DFFR_X1 \REGISTERS_reg[35][29]  ( .D(n7439), .CK(CLK), .RN(n3142), .Q(n9928), 
        .QN(n1202) );
  DFFR_X1 \REGISTERS_reg[35][28]  ( .D(n7440), .CK(CLK), .RN(n3142), .Q(n9929), 
        .QN(n1203) );
  DFFR_X1 \REGISTERS_reg[35][27]  ( .D(n7441), .CK(CLK), .RN(n3142), .Q(n9930), 
        .QN(n1204) );
  DFFR_X1 \REGISTERS_reg[35][26]  ( .D(n7442), .CK(CLK), .RN(n3142), .Q(n9931), 
        .QN(n1205) );
  DFFR_X1 \REGISTERS_reg[35][25]  ( .D(n7443), .CK(CLK), .RN(n3142), .Q(n9932), 
        .QN(n1206) );
  DFFR_X1 \REGISTERS_reg[35][24]  ( .D(n7444), .CK(CLK), .RN(n3142), .Q(n9933), 
        .QN(n1207) );
  DFFR_X1 \REGISTERS_reg[35][23]  ( .D(n7445), .CK(CLK), .RN(n3142), .Q(n9934), 
        .QN(n1208) );
  DFFR_X1 \REGISTERS_reg[35][22]  ( .D(n7446), .CK(CLK), .RN(n3142), .Q(n9935), 
        .QN(n1209) );
  DFFR_X1 \REGISTERS_reg[35][21]  ( .D(n7447), .CK(CLK), .RN(n3142), .Q(n9936), 
        .QN(n1210) );
  DFFR_X1 \REGISTERS_reg[35][20]  ( .D(n7448), .CK(CLK), .RN(n3142), .Q(n9937), 
        .QN(n1211) );
  DFFR_X1 \REGISTERS_reg[35][19]  ( .D(n7449), .CK(CLK), .RN(n3140), .Q(n9938), 
        .QN(n1212) );
  DFFR_X1 \REGISTERS_reg[35][18]  ( .D(n7450), .CK(CLK), .RN(n3140), .Q(n9939), 
        .QN(n1213) );
  DFFR_X1 \REGISTERS_reg[35][17]  ( .D(n7451), .CK(CLK), .RN(n3140), .Q(n9940), 
        .QN(n1214) );
  DFFR_X1 \REGISTERS_reg[35][16]  ( .D(n7452), .CK(CLK), .RN(n3140), .Q(n9941), 
        .QN(n1215) );
  DFFR_X1 \REGISTERS_reg[35][15]  ( .D(n7453), .CK(CLK), .RN(n3140), .Q(n9942), 
        .QN(n1216) );
  DFFR_X1 \REGISTERS_reg[35][14]  ( .D(n7454), .CK(CLK), .RN(n3140), .Q(n9943), 
        .QN(n1217) );
  DFFR_X1 \REGISTERS_reg[35][13]  ( .D(n7455), .CK(CLK), .RN(n3140), .Q(n9944), 
        .QN(n1218) );
  DFFR_X1 \REGISTERS_reg[35][12]  ( .D(n7456), .CK(CLK), .RN(n3140), .Q(n9945), 
        .QN(n1219) );
  DFFR_X1 \REGISTERS_reg[35][11]  ( .D(n7457), .CK(CLK), .RN(n3140), .Q(n9946), 
        .QN(n1220) );
  DFFR_X1 \REGISTERS_reg[35][10]  ( .D(n7458), .CK(CLK), .RN(n3140), .Q(n9947), 
        .QN(n1221) );
  DFFR_X1 \REGISTERS_reg[35][9]  ( .D(n7459), .CK(CLK), .RN(n3140), .Q(n9948), 
        .QN(n1222) );
  DFFR_X1 \REGISTERS_reg[35][8]  ( .D(n7460), .CK(CLK), .RN(n3140), .Q(n9949), 
        .QN(n1223) );
  DFFR_X1 \REGISTERS_reg[35][7]  ( .D(n7461), .CK(CLK), .RN(n3139), .Q(n9950), 
        .QN(n1224) );
  DFFR_X1 \REGISTERS_reg[35][6]  ( .D(n7462), .CK(CLK), .RN(n3139), .Q(n9951), 
        .QN(n1225) );
  DFFR_X1 \REGISTERS_reg[35][5]  ( .D(n7463), .CK(CLK), .RN(n3139), .Q(n9952), 
        .QN(n1226) );
  DFFR_X1 \REGISTERS_reg[35][4]  ( .D(n7464), .CK(CLK), .RN(n3139), .Q(n9953), 
        .QN(n1227) );
  DFFR_X1 \REGISTERS_reg[35][3]  ( .D(n7465), .CK(CLK), .RN(n3139), .Q(n9954), 
        .QN(n1228) );
  DFFR_X1 \REGISTERS_reg[35][2]  ( .D(n7466), .CK(CLK), .RN(n3139), .Q(n9955), 
        .QN(n1229) );
  DFFR_X1 \REGISTERS_reg[35][1]  ( .D(n7467), .CK(CLK), .RN(n3139), .Q(n9956), 
        .QN(n1230) );
  DFFR_X1 \REGISTERS_reg[35][0]  ( .D(n7468), .CK(CLK), .RN(n3139), .Q(n9957), 
        .QN(n1231) );
  DFFR_X1 \REGISTERS_reg[36][31]  ( .D(n7469), .CK(CLK), .RN(n3139), .Q(n9958), 
        .QN(n1232) );
  DFFR_X1 \REGISTERS_reg[36][30]  ( .D(n7470), .CK(CLK), .RN(n3139), .Q(n9959), 
        .QN(n1233) );
  DFFR_X1 \REGISTERS_reg[36][29]  ( .D(n7471), .CK(CLK), .RN(n3139), .Q(n9960), 
        .QN(n1234) );
  DFFR_X1 \REGISTERS_reg[36][28]  ( .D(n7472), .CK(CLK), .RN(n3139), .Q(n9961), 
        .QN(n1235) );
  DFFR_X1 \REGISTERS_reg[36][27]  ( .D(n7473), .CK(CLK), .RN(n3138), .Q(n9962), 
        .QN(n1236) );
  DFFR_X1 \REGISTERS_reg[36][26]  ( .D(n7474), .CK(CLK), .RN(n3138), .Q(n9963), 
        .QN(n1237) );
  DFFR_X1 \REGISTERS_reg[36][25]  ( .D(n7475), .CK(CLK), .RN(n3138), .Q(n9964), 
        .QN(n1238) );
  DFFR_X1 \REGISTERS_reg[36][24]  ( .D(n7476), .CK(CLK), .RN(n3138), .Q(n9965), 
        .QN(n1239) );
  DFFR_X1 \REGISTERS_reg[36][23]  ( .D(n7477), .CK(CLK), .RN(n3138), .Q(n9966), 
        .QN(n1240) );
  DFFR_X1 \REGISTERS_reg[36][22]  ( .D(n7478), .CK(CLK), .RN(n3138), .Q(n9967), 
        .QN(n1241) );
  DFFR_X1 \REGISTERS_reg[36][21]  ( .D(n7479), .CK(CLK), .RN(n3138), .Q(n9968), 
        .QN(n1242) );
  DFFR_X1 \REGISTERS_reg[36][20]  ( .D(n7480), .CK(CLK), .RN(n3138), .Q(n9969), 
        .QN(n1243) );
  DFFR_X1 \REGISTERS_reg[36][19]  ( .D(n7481), .CK(CLK), .RN(n3138), .Q(n9970), 
        .QN(n1244) );
  DFFR_X1 \REGISTERS_reg[36][18]  ( .D(n7482), .CK(CLK), .RN(n3138), .Q(n9971), 
        .QN(n1245) );
  DFFR_X1 \REGISTERS_reg[36][17]  ( .D(n7483), .CK(CLK), .RN(n3138), .Q(n9972), 
        .QN(n1246) );
  DFFR_X1 \REGISTERS_reg[36][16]  ( .D(n7484), .CK(CLK), .RN(n3138), .Q(n9973), 
        .QN(n1247) );
  DFFR_X1 \REGISTERS_reg[36][15]  ( .D(n7485), .CK(CLK), .RN(n3136), .Q(n9974), 
        .QN(n1248) );
  DFFR_X1 \REGISTERS_reg[36][14]  ( .D(n7486), .CK(CLK), .RN(n3136), .Q(n9975), 
        .QN(n1249) );
  DFFR_X1 \REGISTERS_reg[36][13]  ( .D(n7487), .CK(CLK), .RN(n3136), .Q(n9976), 
        .QN(n1250) );
  DFFR_X1 \REGISTERS_reg[36][12]  ( .D(n7488), .CK(CLK), .RN(n3136), .Q(n9977), 
        .QN(n1251) );
  DFFR_X1 \REGISTERS_reg[36][11]  ( .D(n7489), .CK(CLK), .RN(n3136), .Q(n9978), 
        .QN(n1252) );
  DFFR_X1 \REGISTERS_reg[36][10]  ( .D(n7490), .CK(CLK), .RN(n3136), .Q(n9979), 
        .QN(n1253) );
  DFFR_X1 \REGISTERS_reg[36][9]  ( .D(n7491), .CK(CLK), .RN(n3136), .Q(n9980), 
        .QN(n1254) );
  DFFR_X1 \REGISTERS_reg[36][8]  ( .D(n7492), .CK(CLK), .RN(n3136), .Q(n9981), 
        .QN(n1255) );
  DFFR_X1 \REGISTERS_reg[36][7]  ( .D(n7493), .CK(CLK), .RN(n3136), .Q(n9982), 
        .QN(n1256) );
  DFFR_X1 \REGISTERS_reg[36][6]  ( .D(n7494), .CK(CLK), .RN(n3136), .Q(n9983), 
        .QN(n1257) );
  DFFR_X1 \REGISTERS_reg[36][5]  ( .D(n7495), .CK(CLK), .RN(n3136), .Q(n9984), 
        .QN(n1258) );
  DFFR_X1 \REGISTERS_reg[36][4]  ( .D(n7496), .CK(CLK), .RN(n3136), .Q(n9985), 
        .QN(n1259) );
  DFFR_X1 \REGISTERS_reg[36][3]  ( .D(n7497), .CK(CLK), .RN(n3135), .Q(n9986), 
        .QN(n1260) );
  DFFR_X1 \REGISTERS_reg[36][2]  ( .D(n7498), .CK(CLK), .RN(n3135), .Q(n9987), 
        .QN(n1261) );
  DFFR_X1 \REGISTERS_reg[36][1]  ( .D(n7499), .CK(CLK), .RN(n3135), .Q(n9988), 
        .QN(n1262) );
  DFFR_X1 \REGISTERS_reg[36][0]  ( .D(n7500), .CK(CLK), .RN(n3135), .Q(n9989), 
        .QN(n1263) );
  DFFR_X1 \REGISTERS_reg[37][31]  ( .D(n7501), .CK(CLK), .RN(n3135), .Q(n9990), 
        .QN(n1264) );
  DFFR_X1 \REGISTERS_reg[37][30]  ( .D(n7502), .CK(CLK), .RN(n3135), .Q(n9991), 
        .QN(n1265) );
  DFFR_X1 \REGISTERS_reg[37][29]  ( .D(n7503), .CK(CLK), .RN(n3135), .Q(n9992), 
        .QN(n1266) );
  DFFR_X1 \REGISTERS_reg[37][28]  ( .D(n7504), .CK(CLK), .RN(n3135), .Q(n9993), 
        .QN(n1267) );
  DFFR_X1 \REGISTERS_reg[37][27]  ( .D(n7505), .CK(CLK), .RN(n3135), .Q(n9994), 
        .QN(n1268) );
  DFFR_X1 \REGISTERS_reg[37][26]  ( .D(n7506), .CK(CLK), .RN(n3135), .Q(n9995), 
        .QN(n1269) );
  DFFR_X1 \REGISTERS_reg[37][25]  ( .D(n7507), .CK(CLK), .RN(n3135), .Q(n9996), 
        .QN(n1270) );
  DFFR_X1 \REGISTERS_reg[37][24]  ( .D(n7508), .CK(CLK), .RN(n3135), .Q(n9997), 
        .QN(n1271) );
  DFFR_X1 \REGISTERS_reg[37][23]  ( .D(n7509), .CK(CLK), .RN(n3134), .Q(n9998), 
        .QN(n1272) );
  DFFR_X1 \REGISTERS_reg[37][22]  ( .D(n7510), .CK(CLK), .RN(n3134), .Q(n9999), 
        .QN(n1273) );
  DFFR_X1 \REGISTERS_reg[37][21]  ( .D(n7511), .CK(CLK), .RN(n3134), .Q(n10000), .QN(n1274) );
  DFFR_X1 \REGISTERS_reg[37][20]  ( .D(n7512), .CK(CLK), .RN(n3134), .Q(n10001), .QN(n1275) );
  DFFR_X1 \REGISTERS_reg[37][19]  ( .D(n7513), .CK(CLK), .RN(n3134), .Q(n10002), .QN(n1276) );
  DFFR_X1 \REGISTERS_reg[37][18]  ( .D(n7514), .CK(CLK), .RN(n3134), .Q(n10003), .QN(n1277) );
  DFFR_X1 \REGISTERS_reg[37][17]  ( .D(n7515), .CK(CLK), .RN(n3134), .Q(n10004), .QN(n1278) );
  DFFR_X1 \REGISTERS_reg[37][16]  ( .D(n7516), .CK(CLK), .RN(n3134), .Q(n10005), .QN(n1279) );
  DFFR_X1 \REGISTERS_reg[37][15]  ( .D(n7517), .CK(CLK), .RN(n3134), .Q(n10006), .QN(n1280) );
  DFFR_X1 \REGISTERS_reg[37][14]  ( .D(n7518), .CK(CLK), .RN(n3134), .Q(n10007), .QN(n1281) );
  DFFR_X1 \REGISTERS_reg[37][13]  ( .D(n7519), .CK(CLK), .RN(n3134), .Q(n10008), .QN(n1282) );
  DFFR_X1 \REGISTERS_reg[37][12]  ( .D(n7520), .CK(CLK), .RN(n3134), .Q(n10009), .QN(n1283) );
  DFFR_X1 \REGISTERS_reg[37][11]  ( .D(n7521), .CK(CLK), .RN(n3132), .Q(n10010), .QN(n1284) );
  DFFR_X1 \REGISTERS_reg[37][10]  ( .D(n7522), .CK(CLK), .RN(n3132), .Q(n10011), .QN(n1285) );
  DFFR_X1 \REGISTERS_reg[37][9]  ( .D(n7523), .CK(CLK), .RN(n3132), .Q(n10012), 
        .QN(n1286) );
  DFFR_X1 \REGISTERS_reg[37][8]  ( .D(n7524), .CK(CLK), .RN(n3132), .Q(n10013), 
        .QN(n1287) );
  DFFR_X1 \REGISTERS_reg[37][7]  ( .D(n7525), .CK(CLK), .RN(n3132), .Q(n10014), 
        .QN(n1288) );
  DFFR_X1 \REGISTERS_reg[37][6]  ( .D(n7526), .CK(CLK), .RN(n3132), .Q(n10015), 
        .QN(n1289) );
  DFFR_X1 \REGISTERS_reg[37][5]  ( .D(n7527), .CK(CLK), .RN(n3132), .Q(n10016), 
        .QN(n1290) );
  DFFR_X1 \REGISTERS_reg[37][4]  ( .D(n7528), .CK(CLK), .RN(n3132), .Q(n10017), 
        .QN(n1291) );
  DFFR_X1 \REGISTERS_reg[37][3]  ( .D(n7529), .CK(CLK), .RN(n3132), .Q(n10018), 
        .QN(n1292) );
  DFFR_X1 \REGISTERS_reg[37][2]  ( .D(n7530), .CK(CLK), .RN(n3132), .Q(n10019), 
        .QN(n1293) );
  DFFR_X1 \REGISTERS_reg[37][1]  ( .D(n7531), .CK(CLK), .RN(n3132), .Q(n10020), 
        .QN(n1294) );
  DFFR_X1 \REGISTERS_reg[37][0]  ( .D(n7532), .CK(CLK), .RN(n3132), .Q(n10021), 
        .QN(n1295) );
  DFFR_X1 \REGISTERS_reg[46][31]  ( .D(n7789), .CK(CLK), .RN(n3096), .Q(n10022), .QN(n1552) );
  DFFR_X1 \REGISTERS_reg[46][30]  ( .D(n7790), .CK(CLK), .RN(n3096), .Q(n10023), .QN(n1553) );
  DFFR_X1 \REGISTERS_reg[46][29]  ( .D(n7791), .CK(CLK), .RN(n3096), .Q(n10024), .QN(n1554) );
  DFFR_X1 \REGISTERS_reg[46][28]  ( .D(n7792), .CK(CLK), .RN(n3096), .Q(n10025), .QN(n1555) );
  DFFR_X1 \REGISTERS_reg[46][27]  ( .D(n7793), .CK(CLK), .RN(n3096), .Q(n10026), .QN(n1556) );
  DFFR_X1 \REGISTERS_reg[46][26]  ( .D(n7794), .CK(CLK), .RN(n3096), .Q(n10027), .QN(n1557) );
  DFFR_X1 \REGISTERS_reg[46][25]  ( .D(n7795), .CK(CLK), .RN(n3096), .Q(n10028), .QN(n1558) );
  DFFR_X1 \REGISTERS_reg[46][24]  ( .D(n7796), .CK(CLK), .RN(n3096), .Q(n10029), .QN(n1559) );
  DFFR_X1 \REGISTERS_reg[46][23]  ( .D(n7797), .CK(CLK), .RN(n3094), .Q(n10030), .QN(n1560) );
  DFFR_X1 \REGISTERS_reg[46][22]  ( .D(n7798), .CK(CLK), .RN(n3094), .Q(n10031), .QN(n1561) );
  DFFR_X1 \REGISTERS_reg[46][21]  ( .D(n7799), .CK(CLK), .RN(n3094), .Q(n10032), .QN(n1562) );
  DFFR_X1 \REGISTERS_reg[46][20]  ( .D(n7800), .CK(CLK), .RN(n3094), .Q(n10033), .QN(n1563) );
  DFFR_X1 \REGISTERS_reg[46][19]  ( .D(n7801), .CK(CLK), .RN(n3094), .Q(n10034), .QN(n1564) );
  DFFR_X1 \REGISTERS_reg[46][18]  ( .D(n7802), .CK(CLK), .RN(n3094), .Q(n10035), .QN(n1565) );
  DFFR_X1 \REGISTERS_reg[46][17]  ( .D(n7803), .CK(CLK), .RN(n3094), .Q(n10036), .QN(n1566) );
  DFFR_X1 \REGISTERS_reg[46][16]  ( .D(n7804), .CK(CLK), .RN(n3094), .Q(n10037), .QN(n1567) );
  DFFR_X1 \REGISTERS_reg[46][15]  ( .D(n7805), .CK(CLK), .RN(n3094), .Q(n10038), .QN(n1568) );
  DFFR_X1 \REGISTERS_reg[46][14]  ( .D(n7806), .CK(CLK), .RN(n3094), .Q(n10039), .QN(n1569) );
  DFFR_X1 \REGISTERS_reg[46][13]  ( .D(n7807), .CK(CLK), .RN(n3094), .Q(n10040), .QN(n1570) );
  DFFR_X1 \REGISTERS_reg[46][12]  ( .D(n7808), .CK(CLK), .RN(n3094), .Q(n10041), .QN(n1571) );
  DFFR_X1 \REGISTERS_reg[46][11]  ( .D(n7809), .CK(CLK), .RN(n3092), .Q(n10042), .QN(n1572) );
  DFFR_X1 \REGISTERS_reg[46][10]  ( .D(n7810), .CK(CLK), .RN(n3092), .Q(n10043), .QN(n1573) );
  DFFR_X1 \REGISTERS_reg[46][9]  ( .D(n7811), .CK(CLK), .RN(n3092), .Q(n10044), 
        .QN(n1574) );
  DFFR_X1 \REGISTERS_reg[46][8]  ( .D(n7812), .CK(CLK), .RN(n3092), .Q(n10045), 
        .QN(n1575) );
  DFFR_X1 \REGISTERS_reg[46][7]  ( .D(n7813), .CK(CLK), .RN(n3092), .Q(n10046), 
        .QN(n1576) );
  DFFR_X1 \REGISTERS_reg[46][6]  ( .D(n7814), .CK(CLK), .RN(n3092), .Q(n10047), 
        .QN(n1577) );
  DFFR_X1 \REGISTERS_reg[46][5]  ( .D(n7815), .CK(CLK), .RN(n3092), .Q(n10048), 
        .QN(n1578) );
  DFFR_X1 \REGISTERS_reg[46][4]  ( .D(n7816), .CK(CLK), .RN(n3092), .Q(n10049), 
        .QN(n1579) );
  DFFR_X1 \REGISTERS_reg[46][3]  ( .D(n7817), .CK(CLK), .RN(n3092), .Q(n10050), 
        .QN(n1580) );
  DFFR_X1 \REGISTERS_reg[46][2]  ( .D(n7818), .CK(CLK), .RN(n3092), .Q(n10051), 
        .QN(n1581) );
  DFFR_X1 \REGISTERS_reg[46][1]  ( .D(n7819), .CK(CLK), .RN(n3092), .Q(n10052), 
        .QN(n1582) );
  DFFR_X1 \REGISTERS_reg[46][0]  ( .D(n7820), .CK(CLK), .RN(n3092), .Q(n10053), 
        .QN(n1583) );
  DFFR_X1 \REGISTERS_reg[47][31]  ( .D(n7821), .CK(CLK), .RN(n3091), .Q(n10054), .QN(n1584) );
  DFFR_X1 \REGISTERS_reg[47][30]  ( .D(n7822), .CK(CLK), .RN(n3091), .Q(n10055), .QN(n1585) );
  DFFR_X1 \REGISTERS_reg[47][29]  ( .D(n7823), .CK(CLK), .RN(n3091), .Q(n10056), .QN(n1586) );
  DFFR_X1 \REGISTERS_reg[47][28]  ( .D(n7824), .CK(CLK), .RN(n3091), .Q(n10057), .QN(n1587) );
  DFFR_X1 \REGISTERS_reg[47][27]  ( .D(n7825), .CK(CLK), .RN(n3091), .Q(n10058), .QN(n1588) );
  DFFR_X1 \REGISTERS_reg[47][26]  ( .D(n7826), .CK(CLK), .RN(n3091), .Q(n10059), .QN(n1589) );
  DFFR_X1 \REGISTERS_reg[47][25]  ( .D(n7827), .CK(CLK), .RN(n3091), .Q(n10060), .QN(n1590) );
  DFFR_X1 \REGISTERS_reg[47][24]  ( .D(n7828), .CK(CLK), .RN(n3091), .Q(n10061), .QN(n1591) );
  DFFR_X1 \REGISTERS_reg[47][23]  ( .D(n7829), .CK(CLK), .RN(n3091), .Q(n10062), .QN(n1592) );
  DFFR_X1 \REGISTERS_reg[47][22]  ( .D(n7830), .CK(CLK), .RN(n3091), .Q(n10063), .QN(n1593) );
  DFFR_X1 \REGISTERS_reg[47][21]  ( .D(n7831), .CK(CLK), .RN(n3091), .Q(n10064), .QN(n1594) );
  DFFR_X1 \REGISTERS_reg[47][20]  ( .D(n7832), .CK(CLK), .RN(n3091), .Q(n10065), .QN(n1595) );
  DFFR_X1 \REGISTERS_reg[47][19]  ( .D(n7833), .CK(CLK), .RN(n3089), .Q(n10066), .QN(n1596) );
  DFFR_X1 \REGISTERS_reg[47][18]  ( .D(n7834), .CK(CLK), .RN(n3089), .Q(n10067), .QN(n1597) );
  DFFR_X1 \REGISTERS_reg[47][17]  ( .D(n7835), .CK(CLK), .RN(n3089), .Q(n10068), .QN(n1598) );
  DFFR_X1 \REGISTERS_reg[47][16]  ( .D(n7836), .CK(CLK), .RN(n3089), .Q(n10069), .QN(n1599) );
  DFFR_X1 \REGISTERS_reg[47][15]  ( .D(n7837), .CK(CLK), .RN(n3089), .Q(n10070), .QN(n1600) );
  DFFR_X1 \REGISTERS_reg[47][14]  ( .D(n7838), .CK(CLK), .RN(n3089), .Q(n10071), .QN(n1601) );
  DFFR_X1 \REGISTERS_reg[47][13]  ( .D(n7839), .CK(CLK), .RN(n3089), .Q(n10072), .QN(n1602) );
  DFFR_X1 \REGISTERS_reg[47][12]  ( .D(n7840), .CK(CLK), .RN(n3089), .Q(n10073), .QN(n1603) );
  DFFR_X1 \REGISTERS_reg[47][11]  ( .D(n7841), .CK(CLK), .RN(n3089), .Q(n10074), .QN(n1604) );
  DFFR_X1 \REGISTERS_reg[47][10]  ( .D(n7842), .CK(CLK), .RN(n3089), .Q(n10075), .QN(n1605) );
  DFFR_X1 \REGISTERS_reg[47][9]  ( .D(n7843), .CK(CLK), .RN(n3089), .Q(n10076), 
        .QN(n1606) );
  DFFR_X1 \REGISTERS_reg[47][8]  ( .D(n7844), .CK(CLK), .RN(n3089), .Q(n10077), 
        .QN(n1607) );
  DFFR_X1 \REGISTERS_reg[47][7]  ( .D(n7845), .CK(CLK), .RN(n3087), .Q(n10078), 
        .QN(n1608) );
  DFFR_X1 \REGISTERS_reg[47][6]  ( .D(n7846), .CK(CLK), .RN(n3087), .Q(n10079), 
        .QN(n1609) );
  DFFR_X1 \REGISTERS_reg[47][5]  ( .D(n7847), .CK(CLK), .RN(n3087), .Q(n10080), 
        .QN(n1610) );
  DFFR_X1 \REGISTERS_reg[47][4]  ( .D(n7848), .CK(CLK), .RN(n3087), .Q(n10081), 
        .QN(n1611) );
  DFFR_X1 \REGISTERS_reg[47][3]  ( .D(n7849), .CK(CLK), .RN(n3087), .Q(n10082), 
        .QN(n1612) );
  DFFR_X1 \REGISTERS_reg[47][2]  ( .D(n7850), .CK(CLK), .RN(n3087), .Q(n10083), 
        .QN(n1613) );
  DFFR_X1 \REGISTERS_reg[47][1]  ( .D(n7851), .CK(CLK), .RN(n3087), .Q(n10084), 
        .QN(n1614) );
  DFFR_X1 \REGISTERS_reg[47][0]  ( .D(n7852), .CK(CLK), .RN(n3087), .Q(n10085), 
        .QN(n1615) );
  DFFR_X1 \REGISTERS_reg[48][31]  ( .D(n7853), .CK(CLK), .RN(n3087), .Q(n10086), .QN(n1616) );
  DFFR_X1 \REGISTERS_reg[48][30]  ( .D(n7854), .CK(CLK), .RN(n3087), .Q(n10087), .QN(n1617) );
  DFFR_X1 \REGISTERS_reg[48][29]  ( .D(n7855), .CK(CLK), .RN(n3087), .Q(n10088), .QN(n1618) );
  DFFR_X1 \REGISTERS_reg[48][28]  ( .D(n7856), .CK(CLK), .RN(n3087), .Q(n10089), .QN(n1619) );
  DFFR_X1 \REGISTERS_reg[48][27]  ( .D(n7857), .CK(CLK), .RN(n3086), .Q(n10090), .QN(n1620) );
  DFFR_X1 \REGISTERS_reg[48][26]  ( .D(n7858), .CK(CLK), .RN(n3086), .Q(n10091), .QN(n1621) );
  DFFR_X1 \REGISTERS_reg[48][25]  ( .D(n7859), .CK(CLK), .RN(n3086), .Q(n10092), .QN(n1622) );
  DFFR_X1 \REGISTERS_reg[48][24]  ( .D(n7860), .CK(CLK), .RN(n3086), .Q(n10093), .QN(n1623) );
  DFFR_X1 \REGISTERS_reg[48][23]  ( .D(n7861), .CK(CLK), .RN(n3086), .Q(n10094), .QN(n1624) );
  DFFR_X1 \REGISTERS_reg[48][22]  ( .D(n7862), .CK(CLK), .RN(n3086), .Q(n10095), .QN(n1625) );
  DFFR_X1 \REGISTERS_reg[48][21]  ( .D(n7863), .CK(CLK), .RN(n3086), .Q(n10096), .QN(n1626) );
  DFFR_X1 \REGISTERS_reg[48][20]  ( .D(n7864), .CK(CLK), .RN(n3086), .Q(n10097), .QN(n1627) );
  DFFR_X1 \REGISTERS_reg[48][19]  ( .D(n7865), .CK(CLK), .RN(n3086), .Q(n10098), .QN(n1628) );
  DFFR_X1 \REGISTERS_reg[48][18]  ( .D(n7866), .CK(CLK), .RN(n3086), .Q(n10099), .QN(n1629) );
  DFFR_X1 \REGISTERS_reg[48][17]  ( .D(n7867), .CK(CLK), .RN(n3086), .Q(n10100), .QN(n1630) );
  DFFR_X1 \REGISTERS_reg[48][16]  ( .D(n7868), .CK(CLK), .RN(n3086), .Q(n10101), .QN(n1631) );
  DFFR_X1 \REGISTERS_reg[48][15]  ( .D(n7869), .CK(CLK), .RN(n3084), .Q(n10102), .QN(n1632) );
  DFFR_X1 \REGISTERS_reg[48][14]  ( .D(n7870), .CK(CLK), .RN(n3084), .Q(n10103), .QN(n1633) );
  DFFR_X1 \REGISTERS_reg[48][13]  ( .D(n7871), .CK(CLK), .RN(n3084), .Q(n10104), .QN(n1634) );
  DFFR_X1 \REGISTERS_reg[48][12]  ( .D(n7872), .CK(CLK), .RN(n3084), .Q(n10105), .QN(n1635) );
  DFFR_X1 \REGISTERS_reg[48][11]  ( .D(n7873), .CK(CLK), .RN(n3084), .Q(n10106), .QN(n1636) );
  DFFR_X1 \REGISTERS_reg[48][10]  ( .D(n7874), .CK(CLK), .RN(n3084), .Q(n10107), .QN(n1637) );
  DFFR_X1 \REGISTERS_reg[48][9]  ( .D(n7875), .CK(CLK), .RN(n3084), .Q(n10108), 
        .QN(n1638) );
  DFFR_X1 \REGISTERS_reg[48][8]  ( .D(n7876), .CK(CLK), .RN(n3084), .Q(n10109), 
        .QN(n1639) );
  DFFR_X1 \REGISTERS_reg[48][7]  ( .D(n7877), .CK(CLK), .RN(n3084), .Q(n10110), 
        .QN(n1640) );
  DFFR_X1 \REGISTERS_reg[48][6]  ( .D(n7878), .CK(CLK), .RN(n3084), .Q(n10111), 
        .QN(n1641) );
  DFFR_X1 \REGISTERS_reg[48][5]  ( .D(n7879), .CK(CLK), .RN(n3084), .Q(n10112), 
        .QN(n1642) );
  DFFR_X1 \REGISTERS_reg[48][4]  ( .D(n7880), .CK(CLK), .RN(n3084), .Q(n10113), 
        .QN(n1643) );
  DFFR_X1 \REGISTERS_reg[48][3]  ( .D(n7881), .CK(CLK), .RN(n3082), .Q(n10114), 
        .QN(n1644) );
  DFFR_X1 \REGISTERS_reg[48][2]  ( .D(n7882), .CK(CLK), .RN(n3082), .Q(n10115), 
        .QN(n1645) );
  DFFR_X1 \REGISTERS_reg[48][1]  ( .D(n7883), .CK(CLK), .RN(n3082), .Q(n10116), 
        .QN(n1646) );
  DFFR_X1 \REGISTERS_reg[48][0]  ( .D(n7884), .CK(CLK), .RN(n3082), .Q(n10117), 
        .QN(n1647) );
  DFFR_X1 \REGISTERS_reg[55][31]  ( .D(n8077), .CK(CLK), .RN(n3056), .Q(n10118), .QN(n1840) );
  DFFR_X1 \REGISTERS_reg[55][30]  ( .D(n8078), .CK(CLK), .RN(n3056), .Q(n10119), .QN(n1841) );
  DFFR_X1 \REGISTERS_reg[55][29]  ( .D(n8079), .CK(CLK), .RN(n3056), .Q(n10120), .QN(n1842) );
  DFFR_X1 \REGISTERS_reg[55][28]  ( .D(n8080), .CK(CLK), .RN(n3056), .Q(n10121), .QN(n1843) );
  DFFR_X1 \REGISTERS_reg[55][27]  ( .D(n8081), .CK(CLK), .RN(n3056), .Q(n10122), .QN(n1844) );
  DFFR_X1 \REGISTERS_reg[55][26]  ( .D(n8082), .CK(CLK), .RN(n3056), .Q(n10123), .QN(n1845) );
  DFFR_X1 \REGISTERS_reg[55][25]  ( .D(n8083), .CK(CLK), .RN(n3056), .Q(n10124), .QN(n1846) );
  DFFR_X1 \REGISTERS_reg[55][24]  ( .D(n8084), .CK(CLK), .RN(n3056), .Q(n10125), .QN(n1847) );
  DFFR_X1 \REGISTERS_reg[55][23]  ( .D(n8085), .CK(CLK), .RN(n3054), .Q(n10126), .QN(n1848) );
  DFFR_X1 \REGISTERS_reg[55][22]  ( .D(n8086), .CK(CLK), .RN(n3054), .Q(n10127), .QN(n1849) );
  DFFR_X1 \REGISTERS_reg[55][21]  ( .D(n8087), .CK(CLK), .RN(n3054), .Q(n10128), .QN(n1850) );
  DFFR_X1 \REGISTERS_reg[55][20]  ( .D(n8088), .CK(CLK), .RN(n3054), .Q(n10129), .QN(n1851) );
  DFFR_X1 \REGISTERS_reg[55][19]  ( .D(n8089), .CK(CLK), .RN(n3054), .Q(n10130), .QN(n1852) );
  DFFR_X1 \REGISTERS_reg[55][18]  ( .D(n8090), .CK(CLK), .RN(n3054), .Q(n10131), .QN(n1853) );
  DFFR_X1 \REGISTERS_reg[55][17]  ( .D(n8091), .CK(CLK), .RN(n3054), .Q(n10132), .QN(n1854) );
  DFFR_X1 \REGISTERS_reg[55][16]  ( .D(n8092), .CK(CLK), .RN(n3054), .Q(n10133), .QN(n1855) );
  DFFR_X1 \REGISTERS_reg[55][15]  ( .D(n8093), .CK(CLK), .RN(n3054), .Q(n10134), .QN(n1856) );
  DFFR_X1 \REGISTERS_reg[55][14]  ( .D(n8094), .CK(CLK), .RN(n3054), .Q(n10135), .QN(n1857) );
  DFFR_X1 \REGISTERS_reg[55][13]  ( .D(n8095), .CK(CLK), .RN(n3054), .Q(n10136), .QN(n1858) );
  DFFR_X1 \REGISTERS_reg[55][12]  ( .D(n8096), .CK(CLK), .RN(n3054), .Q(n10137), .QN(n1859) );
  DFFR_X1 \REGISTERS_reg[55][11]  ( .D(n8097), .CK(CLK), .RN(n3052), .Q(n10138), .QN(n1860) );
  DFFR_X1 \REGISTERS_reg[55][10]  ( .D(n8098), .CK(CLK), .RN(n3052), .Q(n10139), .QN(n1861) );
  DFFR_X1 \REGISTERS_reg[55][9]  ( .D(n8099), .CK(CLK), .RN(n3052), .Q(n10140), 
        .QN(n1862) );
  DFFR_X1 \REGISTERS_reg[55][8]  ( .D(n8100), .CK(CLK), .RN(n3052), .Q(n10141), 
        .QN(n1863) );
  DFFR_X1 \REGISTERS_reg[55][7]  ( .D(n8101), .CK(CLK), .RN(n3052), .Q(n10142), 
        .QN(n1864) );
  DFFR_X1 \REGISTERS_reg[55][6]  ( .D(n8102), .CK(CLK), .RN(n3052), .Q(n10143), 
        .QN(n1865) );
  DFFR_X1 \REGISTERS_reg[55][5]  ( .D(n8103), .CK(CLK), .RN(n3052), .Q(n10144), 
        .QN(n1866) );
  DFFR_X1 \REGISTERS_reg[55][4]  ( .D(n8104), .CK(CLK), .RN(n3052), .Q(n10145), 
        .QN(n1867) );
  DFFR_X1 \REGISTERS_reg[55][3]  ( .D(n8105), .CK(CLK), .RN(n3052), .Q(n10146), 
        .QN(n1868) );
  DFFR_X1 \REGISTERS_reg[55][2]  ( .D(n8106), .CK(CLK), .RN(n3052), .Q(n10147), 
        .QN(n1869) );
  DFFR_X1 \REGISTERS_reg[55][1]  ( .D(n8107), .CK(CLK), .RN(n3052), .Q(n10148), 
        .QN(n1870) );
  DFFR_X1 \REGISTERS_reg[55][0]  ( .D(n8108), .CK(CLK), .RN(n3052), .Q(n10149), 
        .QN(n1871) );
  DFFR_X1 \REGISTERS_reg[56][31]  ( .D(n8109), .CK(CLK), .RN(n3051), .Q(n10150), .QN(n1872) );
  DFFR_X1 \REGISTERS_reg[56][30]  ( .D(n8110), .CK(CLK), .RN(n3051), .Q(n10151), .QN(n1873) );
  DFFR_X1 \REGISTERS_reg[56][29]  ( .D(n8111), .CK(CLK), .RN(n3051), .Q(n10152), .QN(n1874) );
  DFFR_X1 \REGISTERS_reg[56][28]  ( .D(n8112), .CK(CLK), .RN(n3051), .Q(n10153), .QN(n1875) );
  DFFR_X1 \REGISTERS_reg[56][27]  ( .D(n8113), .CK(CLK), .RN(n3051), .Q(n10154), .QN(n1876) );
  DFFR_X1 \REGISTERS_reg[56][26]  ( .D(n8114), .CK(CLK), .RN(n3051), .Q(n10155), .QN(n1877) );
  DFFR_X1 \REGISTERS_reg[56][25]  ( .D(n8115), .CK(CLK), .RN(n3051), .Q(n10156), .QN(n1878) );
  DFFR_X1 \REGISTERS_reg[56][24]  ( .D(n8116), .CK(CLK), .RN(n3051), .Q(n10157), .QN(n1879) );
  DFFR_X1 \REGISTERS_reg[56][23]  ( .D(n8117), .CK(CLK), .RN(n3051), .Q(n10158), .QN(n1880) );
  DFFR_X1 \REGISTERS_reg[56][22]  ( .D(n8118), .CK(CLK), .RN(n3051), .Q(n10159), .QN(n1881) );
  DFFR_X1 \REGISTERS_reg[56][21]  ( .D(n8119), .CK(CLK), .RN(n3051), .Q(n10160), .QN(n1882) );
  DFFR_X1 \REGISTERS_reg[56][20]  ( .D(n8120), .CK(CLK), .RN(n3051), .Q(n10161), .QN(n1883) );
  DFFR_X1 \REGISTERS_reg[56][19]  ( .D(n8121), .CK(CLK), .RN(n3049), .Q(n10162), .QN(n1884) );
  DFFR_X1 \REGISTERS_reg[56][18]  ( .D(n8122), .CK(CLK), .RN(n3049), .Q(n10163), .QN(n1885) );
  DFFR_X1 \REGISTERS_reg[56][17]  ( .D(n8123), .CK(CLK), .RN(n3049), .Q(n10164), .QN(n1886) );
  DFFR_X1 \REGISTERS_reg[56][16]  ( .D(n8124), .CK(CLK), .RN(n3049), .Q(n10165), .QN(n1887) );
  DFFR_X1 \REGISTERS_reg[56][15]  ( .D(n8125), .CK(CLK), .RN(n3049), .Q(n10166), .QN(n1888) );
  DFFR_X1 \REGISTERS_reg[56][14]  ( .D(n8126), .CK(CLK), .RN(n3049), .Q(n10167), .QN(n1889) );
  DFFR_X1 \REGISTERS_reg[56][13]  ( .D(n8127), .CK(CLK), .RN(n3049), .Q(n10168), .QN(n1890) );
  DFFR_X1 \REGISTERS_reg[56][12]  ( .D(n8128), .CK(CLK), .RN(n3049), .Q(n10169), .QN(n1891) );
  DFFR_X1 \REGISTERS_reg[56][11]  ( .D(n8129), .CK(CLK), .RN(n3049), .Q(n10170), .QN(n1892) );
  DFFR_X1 \REGISTERS_reg[56][10]  ( .D(n8130), .CK(CLK), .RN(n3049), .Q(n10171), .QN(n1893) );
  DFFR_X1 \REGISTERS_reg[56][9]  ( .D(n8131), .CK(CLK), .RN(n3049), .Q(n10172), 
        .QN(n1894) );
  DFFR_X1 \REGISTERS_reg[56][8]  ( .D(n8132), .CK(CLK), .RN(n3049), .Q(n10173), 
        .QN(n1895) );
  DFFR_X1 \REGISTERS_reg[56][7]  ( .D(n8133), .CK(CLK), .RN(n3047), .Q(n10174), 
        .QN(n1896) );
  DFFR_X1 \REGISTERS_reg[56][6]  ( .D(n8134), .CK(CLK), .RN(n3047), .Q(n10175), 
        .QN(n1897) );
  DFFR_X1 \REGISTERS_reg[56][5]  ( .D(n8135), .CK(CLK), .RN(n3047), .Q(n10176), 
        .QN(n1898) );
  DFFR_X1 \REGISTERS_reg[56][4]  ( .D(n8136), .CK(CLK), .RN(n3047), .Q(n10177), 
        .QN(n1899) );
  DFFR_X1 \REGISTERS_reg[56][3]  ( .D(n8137), .CK(CLK), .RN(n3047), .Q(n10178), 
        .QN(n1900) );
  DFFR_X1 \REGISTERS_reg[56][2]  ( .D(n8138), .CK(CLK), .RN(n3047), .Q(n10179), 
        .QN(n1901) );
  DFFR_X1 \REGISTERS_reg[56][1]  ( .D(n8139), .CK(CLK), .RN(n3047), .Q(n10180), 
        .QN(n1902) );
  DFFR_X1 \REGISTERS_reg[56][0]  ( .D(n8140), .CK(CLK), .RN(n3047), .Q(n10181), 
        .QN(n1903) );
  DFFR_X1 \REGISTERS_reg[57][31]  ( .D(n8141), .CK(CLK), .RN(n3047), .Q(n10182), .QN(n1904) );
  DFFR_X1 \REGISTERS_reg[57][30]  ( .D(n8142), .CK(CLK), .RN(n3047), .Q(n10183), .QN(n1905) );
  DFFR_X1 \REGISTERS_reg[57][29]  ( .D(n8143), .CK(CLK), .RN(n3047), .Q(n10184), .QN(n1906) );
  DFFR_X1 \REGISTERS_reg[57][28]  ( .D(n8144), .CK(CLK), .RN(n3047), .Q(n10185), .QN(n1907) );
  DFFR_X1 \REGISTERS_reg[57][27]  ( .D(n8145), .CK(CLK), .RN(n3046), .Q(n10186), .QN(n1908) );
  DFFR_X1 \REGISTERS_reg[57][26]  ( .D(n8146), .CK(CLK), .RN(n3046), .Q(n10187), .QN(n1909) );
  DFFR_X1 \REGISTERS_reg[57][25]  ( .D(n8147), .CK(CLK), .RN(n3046), .Q(n10188), .QN(n1910) );
  DFFR_X1 \REGISTERS_reg[57][24]  ( .D(n8148), .CK(CLK), .RN(n3046), .Q(n10189), .QN(n1911) );
  DFFR_X1 \REGISTERS_reg[57][23]  ( .D(n8149), .CK(CLK), .RN(n3046), .Q(n10190), .QN(n1912) );
  DFFR_X1 \REGISTERS_reg[57][22]  ( .D(n8150), .CK(CLK), .RN(n3046), .Q(n10191), .QN(n1913) );
  DFFR_X1 \REGISTERS_reg[57][21]  ( .D(n8151), .CK(CLK), .RN(n3046), .Q(n10192), .QN(n1914) );
  DFFR_X1 \REGISTERS_reg[57][20]  ( .D(n8152), .CK(CLK), .RN(n3046), .Q(n10193), .QN(n1915) );
  DFFR_X1 \REGISTERS_reg[57][19]  ( .D(n8153), .CK(CLK), .RN(n3046), .Q(n10194), .QN(n1916) );
  DFFR_X1 \REGISTERS_reg[57][18]  ( .D(n8154), .CK(CLK), .RN(n3046), .Q(n10195), .QN(n1917) );
  DFFR_X1 \REGISTERS_reg[57][17]  ( .D(n8155), .CK(CLK), .RN(n3046), .Q(n10196), .QN(n1918) );
  DFFR_X1 \REGISTERS_reg[57][16]  ( .D(n8156), .CK(CLK), .RN(n3046), .Q(n10197), .QN(n1919) );
  DFFR_X1 \REGISTERS_reg[57][15]  ( .D(n8157), .CK(CLK), .RN(n3044), .Q(n10198), .QN(n1920) );
  DFFR_X1 \REGISTERS_reg[57][14]  ( .D(n8158), .CK(CLK), .RN(n3044), .Q(n10199), .QN(n1921) );
  DFFR_X1 \REGISTERS_reg[57][13]  ( .D(n8159), .CK(CLK), .RN(n3044), .Q(n10200), .QN(n1922) );
  DFFR_X1 \REGISTERS_reg[57][12]  ( .D(n8160), .CK(CLK), .RN(n3044), .Q(n10201), .QN(n1923) );
  DFFR_X1 \REGISTERS_reg[57][11]  ( .D(n8161), .CK(CLK), .RN(n3044), .Q(n10202), .QN(n1924) );
  DFFR_X1 \REGISTERS_reg[57][10]  ( .D(n8162), .CK(CLK), .RN(n3044), .Q(n10203), .QN(n1925) );
  DFFR_X1 \REGISTERS_reg[57][9]  ( .D(n8163), .CK(CLK), .RN(n3044), .Q(n10204), 
        .QN(n1926) );
  DFFR_X1 \REGISTERS_reg[57][8]  ( .D(n8164), .CK(CLK), .RN(n3044), .Q(n10205), 
        .QN(n1927) );
  DFFR_X1 \REGISTERS_reg[57][7]  ( .D(n8165), .CK(CLK), .RN(n3044), .Q(n10206), 
        .QN(n1928) );
  DFFR_X1 \REGISTERS_reg[57][6]  ( .D(n8166), .CK(CLK), .RN(n3044), .Q(n10207), 
        .QN(n1929) );
  DFFR_X1 \REGISTERS_reg[57][5]  ( .D(n8167), .CK(CLK), .RN(n3044), .Q(n10208), 
        .QN(n1930) );
  DFFR_X1 \REGISTERS_reg[57][4]  ( .D(n8168), .CK(CLK), .RN(n3044), .Q(n10209), 
        .QN(n1931) );
  DFFR_X1 \REGISTERS_reg[57][3]  ( .D(n8169), .CK(CLK), .RN(n3042), .Q(n10210), 
        .QN(n1932) );
  DFFR_X1 \REGISTERS_reg[57][2]  ( .D(n8170), .CK(CLK), .RN(n3042), .Q(n10211), 
        .QN(n1933) );
  DFFR_X1 \REGISTERS_reg[57][1]  ( .D(n8171), .CK(CLK), .RN(n3042), .Q(n10212), 
        .QN(n1934) );
  DFFR_X1 \REGISTERS_reg[57][0]  ( .D(n8172), .CK(CLK), .RN(n3042), .Q(n10213), 
        .QN(n1935) );
  DFFR_X1 \REGISTERS_reg[58][31]  ( .D(n8173), .CK(CLK), .RN(n3042), .Q(n10214), .QN(n1936) );
  DFFR_X1 \REGISTERS_reg[58][30]  ( .D(n8174), .CK(CLK), .RN(n3042), .Q(n10215), .QN(n1937) );
  DFFR_X1 \REGISTERS_reg[58][29]  ( .D(n8175), .CK(CLK), .RN(n3042), .Q(n10216), .QN(n1938) );
  DFFR_X1 \REGISTERS_reg[58][28]  ( .D(n8176), .CK(CLK), .RN(n3042), .Q(n10217), .QN(n1939) );
  DFFR_X1 \REGISTERS_reg[58][27]  ( .D(n8177), .CK(CLK), .RN(n3042), .Q(n10218), .QN(n1940) );
  DFFR_X1 \REGISTERS_reg[58][26]  ( .D(n8178), .CK(CLK), .RN(n3042), .Q(n10219), .QN(n1941) );
  DFFR_X1 \REGISTERS_reg[58][25]  ( .D(n8179), .CK(CLK), .RN(n3042), .Q(n10220), .QN(n1942) );
  DFFR_X1 \REGISTERS_reg[58][24]  ( .D(n8180), .CK(CLK), .RN(n3042), .Q(n10221), .QN(n1943) );
  DFFR_X1 \REGISTERS_reg[58][23]  ( .D(n8181), .CK(CLK), .RN(n3041), .Q(n10222), .QN(n1944) );
  DFFR_X1 \REGISTERS_reg[58][22]  ( .D(n8182), .CK(CLK), .RN(n3041), .Q(n10223), .QN(n1945) );
  DFFR_X1 \REGISTERS_reg[58][21]  ( .D(n8183), .CK(CLK), .RN(n3041), .Q(n10224), .QN(n1946) );
  DFFR_X1 \REGISTERS_reg[58][20]  ( .D(n8184), .CK(CLK), .RN(n3041), .Q(n10225), .QN(n1947) );
  DFFR_X1 \REGISTERS_reg[58][19]  ( .D(n8185), .CK(CLK), .RN(n3041), .Q(n10226), .QN(n1948) );
  DFFR_X1 \REGISTERS_reg[58][18]  ( .D(n8186), .CK(CLK), .RN(n3041), .Q(n10227), .QN(n1949) );
  DFFR_X1 \REGISTERS_reg[58][17]  ( .D(n8187), .CK(CLK), .RN(n3041), .Q(n10228), .QN(n1950) );
  DFFR_X1 \REGISTERS_reg[58][16]  ( .D(n8188), .CK(CLK), .RN(n3041), .Q(n10229), .QN(n1951) );
  DFFR_X1 \REGISTERS_reg[58][15]  ( .D(n8189), .CK(CLK), .RN(n3041), .Q(n10230), .QN(n1952) );
  DFFR_X1 \REGISTERS_reg[58][14]  ( .D(n8190), .CK(CLK), .RN(n3041), .Q(n10231), .QN(n1953) );
  DFFR_X1 \REGISTERS_reg[58][13]  ( .D(n8191), .CK(CLK), .RN(n3041), .Q(n10232), .QN(n1954) );
  DFFR_X1 \REGISTERS_reg[58][12]  ( .D(n8192), .CK(CLK), .RN(n3041), .Q(n10233), .QN(n1955) );
  DFFR_X1 \REGISTERS_reg[58][11]  ( .D(n8193), .CK(CLK), .RN(n3039), .Q(n10234), .QN(n1956) );
  DFFR_X1 \REGISTERS_reg[58][10]  ( .D(n8194), .CK(CLK), .RN(n3039), .Q(n10235), .QN(n1957) );
  DFFR_X1 \REGISTERS_reg[58][9]  ( .D(n8195), .CK(CLK), .RN(n3039), .Q(n10236), 
        .QN(n1958) );
  DFFR_X1 \REGISTERS_reg[58][8]  ( .D(n8196), .CK(CLK), .RN(n3039), .Q(n10237), 
        .QN(n1959) );
  DFFR_X1 \REGISTERS_reg[58][7]  ( .D(n8197), .CK(CLK), .RN(n3039), .Q(n10238), 
        .QN(n1960) );
  DFFR_X1 \REGISTERS_reg[58][6]  ( .D(n8198), .CK(CLK), .RN(n3039), .Q(n10239), 
        .QN(n1961) );
  DFFR_X1 \REGISTERS_reg[58][5]  ( .D(n8199), .CK(CLK), .RN(n3039), .Q(n10240), 
        .QN(n1962) );
  DFFR_X1 \REGISTERS_reg[58][4]  ( .D(n8200), .CK(CLK), .RN(n3039), .Q(n10241), 
        .QN(n1963) );
  DFFR_X1 \REGISTERS_reg[58][3]  ( .D(n8201), .CK(CLK), .RN(n3039), .Q(n10242), 
        .QN(n1964) );
  DFFR_X1 \REGISTERS_reg[58][2]  ( .D(n8202), .CK(CLK), .RN(n3039), .Q(n10243), 
        .QN(n1965) );
  DFFR_X1 \REGISTERS_reg[58][1]  ( .D(n8203), .CK(CLK), .RN(n3039), .Q(n10244), 
        .QN(n1966) );
  DFFR_X1 \REGISTERS_reg[58][0]  ( .D(n8204), .CK(CLK), .RN(n3039), .Q(n10245), 
        .QN(n1967) );
  DFFR_X1 \REGISTERS_reg[59][31]  ( .D(n8205), .CK(CLK), .RN(n3037), .Q(n10246), .QN(n1968) );
  DFFR_X1 \REGISTERS_reg[59][30]  ( .D(n8206), .CK(CLK), .RN(n3037), .Q(n10247), .QN(n1969) );
  DFFR_X1 \REGISTERS_reg[59][29]  ( .D(n8207), .CK(CLK), .RN(n3037), .Q(n10248), .QN(n1970) );
  DFFR_X1 \REGISTERS_reg[59][28]  ( .D(n8208), .CK(CLK), .RN(n3037), .Q(n10249), .QN(n1971) );
  DFFR_X1 \REGISTERS_reg[59][27]  ( .D(n8209), .CK(CLK), .RN(n3037), .Q(n10250), .QN(n1972) );
  DFFR_X1 \REGISTERS_reg[59][26]  ( .D(n8210), .CK(CLK), .RN(n3037), .Q(n10251), .QN(n1973) );
  DFFR_X1 \REGISTERS_reg[59][25]  ( .D(n8211), .CK(CLK), .RN(n3037), .Q(n10252), .QN(n1974) );
  DFFR_X1 \REGISTERS_reg[59][24]  ( .D(n8212), .CK(CLK), .RN(n3037), .Q(n10253), .QN(n1975) );
  DFFR_X1 \REGISTERS_reg[59][23]  ( .D(n8213), .CK(CLK), .RN(n3037), .Q(n10254), .QN(n1976) );
  DFFR_X1 \REGISTERS_reg[59][22]  ( .D(n8214), .CK(CLK), .RN(n3037), .Q(n10255), .QN(n1977) );
  DFFR_X1 \REGISTERS_reg[59][21]  ( .D(n8215), .CK(CLK), .RN(n3037), .Q(n10256), .QN(n1978) );
  DFFR_X1 \REGISTERS_reg[59][20]  ( .D(n8216), .CK(CLK), .RN(n3037), .Q(n10257), .QN(n1979) );
  DFFR_X1 \REGISTERS_reg[59][19]  ( .D(n8217), .CK(CLK), .RN(n3036), .Q(n10258), .QN(n1980) );
  DFFR_X1 \REGISTERS_reg[59][18]  ( .D(n8218), .CK(CLK), .RN(n3036), .Q(n10259), .QN(n1981) );
  DFFR_X1 \REGISTERS_reg[59][17]  ( .D(n8219), .CK(CLK), .RN(n3036), .Q(n10260), .QN(n1982) );
  DFFR_X1 \REGISTERS_reg[59][16]  ( .D(n8220), .CK(CLK), .RN(n3036), .Q(n10261), .QN(n1983) );
  DFFR_X1 \REGISTERS_reg[59][15]  ( .D(n8221), .CK(CLK), .RN(n3036), .Q(n10262), .QN(n1984) );
  DFFR_X1 \REGISTERS_reg[59][14]  ( .D(n8222), .CK(CLK), .RN(n3036), .Q(n10263), .QN(n1985) );
  DFFR_X1 \REGISTERS_reg[59][13]  ( .D(n8223), .CK(CLK), .RN(n3036), .Q(n10264), .QN(n1986) );
  DFFR_X1 \REGISTERS_reg[59][12]  ( .D(n8224), .CK(CLK), .RN(n3036), .Q(n10265), .QN(n1987) );
  DFFR_X1 \REGISTERS_reg[59][11]  ( .D(n8225), .CK(CLK), .RN(n3036), .Q(n10266), .QN(n1988) );
  DFFR_X1 \REGISTERS_reg[59][10]  ( .D(n8226), .CK(CLK), .RN(n3036), .Q(n10267), .QN(n1989) );
  DFFR_X1 \REGISTERS_reg[59][9]  ( .D(n8227), .CK(CLK), .RN(n3036), .Q(n10268), 
        .QN(n1990) );
  DFFR_X1 \REGISTERS_reg[59][8]  ( .D(n8228), .CK(CLK), .RN(n3036), .Q(n10269), 
        .QN(n1991) );
  DFFR_X1 \REGISTERS_reg[59][7]  ( .D(n8229), .CK(CLK), .RN(n3034), .Q(n10270), 
        .QN(n1992) );
  DFFR_X1 \REGISTERS_reg[59][6]  ( .D(n8230), .CK(CLK), .RN(n3034), .Q(n10271), 
        .QN(n1993) );
  DFFR_X1 \REGISTERS_reg[59][5]  ( .D(n8231), .CK(CLK), .RN(n3034), .Q(n10272), 
        .QN(n1994) );
  DFFR_X1 \REGISTERS_reg[59][4]  ( .D(n8232), .CK(CLK), .RN(n3034), .Q(n10273), 
        .QN(n1995) );
  DFFR_X1 \REGISTERS_reg[59][3]  ( .D(n8233), .CK(CLK), .RN(n3034), .Q(n10274), 
        .QN(n1996) );
  DFFR_X1 \REGISTERS_reg[59][2]  ( .D(n8234), .CK(CLK), .RN(n3034), .Q(n10275), 
        .QN(n1997) );
  DFFR_X1 \REGISTERS_reg[59][1]  ( .D(n8235), .CK(CLK), .RN(n3034), .Q(n10276), 
        .QN(n1998) );
  DFFR_X1 \REGISTERS_reg[59][0]  ( .D(n8236), .CK(CLK), .RN(n3034), .Q(n10277), 
        .QN(n1999) );
  DFFR_X1 \REGISTERS_reg[60][31]  ( .D(n8237), .CK(CLK), .RN(n3034), .Q(n10278), .QN(n2000) );
  DFFR_X1 \REGISTERS_reg[60][30]  ( .D(n8238), .CK(CLK), .RN(n3034), .Q(n10279), .QN(n2001) );
  DFFR_X1 \REGISTERS_reg[60][29]  ( .D(n8239), .CK(CLK), .RN(n3034), .Q(n10280), .QN(n2002) );
  DFFR_X1 \REGISTERS_reg[60][28]  ( .D(n8240), .CK(CLK), .RN(n3034), .Q(n10281), .QN(n2003) );
  DFFR_X1 \REGISTERS_reg[60][27]  ( .D(n8241), .CK(CLK), .RN(n3032), .Q(n10282), .QN(n2004) );
  DFFR_X1 \REGISTERS_reg[60][26]  ( .D(n8242), .CK(CLK), .RN(n3032), .Q(n10283), .QN(n2005) );
  DFFR_X1 \REGISTERS_reg[60][25]  ( .D(n8243), .CK(CLK), .RN(n3032), .Q(n10284), .QN(n2006) );
  DFFR_X1 \REGISTERS_reg[60][24]  ( .D(n8244), .CK(CLK), .RN(n3032), .Q(n10285), .QN(n2007) );
  DFFR_X1 \REGISTERS_reg[60][23]  ( .D(n8245), .CK(CLK), .RN(n3032), .Q(n10286), .QN(n2008) );
  DFFR_X1 \REGISTERS_reg[60][22]  ( .D(n8246), .CK(CLK), .RN(n3032), .Q(n10287), .QN(n2009) );
  DFFR_X1 \REGISTERS_reg[60][21]  ( .D(n8247), .CK(CLK), .RN(n3032), .Q(n10288), .QN(n2010) );
  DFFR_X1 \REGISTERS_reg[60][20]  ( .D(n8248), .CK(CLK), .RN(n3032), .Q(n10289), .QN(n2011) );
  DFFR_X1 \REGISTERS_reg[60][19]  ( .D(n8249), .CK(CLK), .RN(n3032), .Q(n10290), .QN(n2012) );
  DFFR_X1 \REGISTERS_reg[60][18]  ( .D(n8250), .CK(CLK), .RN(n3032), .Q(n10291), .QN(n2013) );
  DFFR_X1 \REGISTERS_reg[60][17]  ( .D(n8251), .CK(CLK), .RN(n3032), .Q(n10292), .QN(n2014) );
  DFFR_X1 \REGISTERS_reg[60][16]  ( .D(n8252), .CK(CLK), .RN(n3032), .Q(n10293), .QN(n2015) );
  DFFR_X1 \REGISTERS_reg[60][15]  ( .D(n8253), .CK(CLK), .RN(n3031), .Q(n10294), .QN(n2016) );
  DFFR_X1 \REGISTERS_reg[60][14]  ( .D(n8254), .CK(CLK), .RN(n3031), .Q(n10295), .QN(n2017) );
  DFFR_X1 \REGISTERS_reg[60][13]  ( .D(n8255), .CK(CLK), .RN(n3031), .Q(n10296), .QN(n2018) );
  DFFR_X1 \REGISTERS_reg[60][12]  ( .D(n8256), .CK(CLK), .RN(n3031), .Q(n10297), .QN(n2019) );
  DFFR_X1 \REGISTERS_reg[60][11]  ( .D(n8257), .CK(CLK), .RN(n3031), .Q(n10298), .QN(n2020) );
  DFFR_X1 \REGISTERS_reg[60][10]  ( .D(n8258), .CK(CLK), .RN(n3031), .Q(n10299), .QN(n2021) );
  DFFR_X1 \REGISTERS_reg[60][9]  ( .D(n8259), .CK(CLK), .RN(n3031), .Q(n10300), 
        .QN(n2022) );
  DFFR_X1 \REGISTERS_reg[60][8]  ( .D(n8260), .CK(CLK), .RN(n3031), .Q(n10301), 
        .QN(n2023) );
  DFFR_X1 \REGISTERS_reg[60][7]  ( .D(n8261), .CK(CLK), .RN(n3031), .Q(n10302), 
        .QN(n2024) );
  DFFR_X1 \REGISTERS_reg[60][6]  ( .D(n8262), .CK(CLK), .RN(n3031), .Q(n10303), 
        .QN(n2025) );
  DFFR_X1 \REGISTERS_reg[60][5]  ( .D(n8263), .CK(CLK), .RN(n3031), .Q(n10304), 
        .QN(n2026) );
  DFFR_X1 \REGISTERS_reg[60][4]  ( .D(n8264), .CK(CLK), .RN(n3031), .Q(n10305), 
        .QN(n2027) );
  DFFR_X1 \REGISTERS_reg[60][3]  ( .D(n8265), .CK(CLK), .RN(n3028), .Q(n10306), 
        .QN(n2028) );
  DFFR_X1 \REGISTERS_reg[60][2]  ( .D(n8266), .CK(CLK), .RN(n3028), .Q(n10307), 
        .QN(n2029) );
  DFFR_X1 \REGISTERS_reg[60][1]  ( .D(n8267), .CK(CLK), .RN(n3028), .Q(n10308), 
        .QN(n2030) );
  DFFR_X1 \REGISTERS_reg[60][0]  ( .D(n8268), .CK(CLK), .RN(n3028), .Q(n10309), 
        .QN(n2031) );
  DFFR_X1 \REGISTERS_reg[61][31]  ( .D(n8269), .CK(CLK), .RN(n3028), .Q(n10310), .QN(n2032) );
  DFFR_X1 \REGISTERS_reg[61][30]  ( .D(n8270), .CK(CLK), .RN(n3028), .Q(n10311), .QN(n2033) );
  DFFR_X1 \REGISTERS_reg[61][29]  ( .D(n8271), .CK(CLK), .RN(n3028), .Q(n10312), .QN(n2034) );
  DFFR_X1 \REGISTERS_reg[61][28]  ( .D(n8272), .CK(CLK), .RN(n3028), .Q(n10313), .QN(n2035) );
  DFFR_X1 \REGISTERS_reg[61][27]  ( .D(n8273), .CK(CLK), .RN(n3028), .Q(n10314), .QN(n2036) );
  DFFR_X1 \REGISTERS_reg[61][26]  ( .D(n8274), .CK(CLK), .RN(n3028), .Q(n10315), .QN(n2037) );
  DFFR_X1 \REGISTERS_reg[61][25]  ( .D(n8275), .CK(CLK), .RN(n3028), .Q(n10316), .QN(n2038) );
  DFFR_X1 \REGISTERS_reg[61][24]  ( .D(n8276), .CK(CLK), .RN(n3028), .Q(n10317), .QN(n2039) );
  DFFR_X1 \REGISTERS_reg[61][23]  ( .D(n8277), .CK(CLK), .RN(n3027), .Q(n10318), .QN(n2040) );
  DFFR_X1 \REGISTERS_reg[61][22]  ( .D(n8278), .CK(CLK), .RN(n3027), .Q(n10319), .QN(n2041) );
  DFFR_X1 \REGISTERS_reg[61][21]  ( .D(n8279), .CK(CLK), .RN(n3027), .Q(n10320), .QN(n2042) );
  DFFR_X1 \REGISTERS_reg[61][20]  ( .D(n8280), .CK(CLK), .RN(n3027), .Q(n10321), .QN(n2043) );
  DFFR_X1 \REGISTERS_reg[61][19]  ( .D(n8281), .CK(CLK), .RN(n3027), .Q(n10322), .QN(n2044) );
  DFFR_X1 \REGISTERS_reg[61][18]  ( .D(n8282), .CK(CLK), .RN(n3027), .Q(n10323), .QN(n2045) );
  DFFR_X1 \REGISTERS_reg[61][17]  ( .D(n8283), .CK(CLK), .RN(n3027), .Q(n10324), .QN(n2046) );
  DFFR_X1 \REGISTERS_reg[61][16]  ( .D(n8284), .CK(CLK), .RN(n3027), .Q(n10325), .QN(n2047) );
  DFFR_X1 \REGISTERS_reg[61][15]  ( .D(n8285), .CK(CLK), .RN(n3027), .Q(n10326), .QN(n2048) );
  DFFR_X1 \REGISTERS_reg[61][14]  ( .D(n8286), .CK(CLK), .RN(n3027), .Q(n10327), .QN(n2049) );
  DFFR_X1 \REGISTERS_reg[61][13]  ( .D(n8287), .CK(CLK), .RN(n3027), .Q(n10328), .QN(n2050) );
  DFFR_X1 \REGISTERS_reg[61][12]  ( .D(n8288), .CK(CLK), .RN(n3027), .Q(n10329), .QN(n2051) );
  DFFR_X1 \REGISTERS_reg[61][11]  ( .D(n8289), .CK(CLK), .RN(n3026), .Q(n10330), .QN(n2052) );
  DFFR_X1 \REGISTERS_reg[61][10]  ( .D(n8290), .CK(CLK), .RN(n3026), .Q(n10331), .QN(n2053) );
  DFFR_X1 \REGISTERS_reg[61][9]  ( .D(n8291), .CK(CLK), .RN(n3026), .Q(n10332), 
        .QN(n2054) );
  DFFR_X1 \REGISTERS_reg[61][8]  ( .D(n8292), .CK(CLK), .RN(n3026), .Q(n10333), 
        .QN(n2055) );
  DFFR_X1 \REGISTERS_reg[61][7]  ( .D(n8293), .CK(CLK), .RN(n3026), .Q(n10334), 
        .QN(n2056) );
  DFFR_X1 \REGISTERS_reg[61][6]  ( .D(n8294), .CK(CLK), .RN(n3026), .Q(n10335), 
        .QN(n2057) );
  DFFR_X1 \REGISTERS_reg[61][5]  ( .D(n8295), .CK(CLK), .RN(n3026), .Q(n10336), 
        .QN(n2058) );
  DFFR_X1 \REGISTERS_reg[61][4]  ( .D(n8296), .CK(CLK), .RN(n3026), .Q(n10337), 
        .QN(n2059) );
  DFFR_X1 \REGISTERS_reg[61][3]  ( .D(n8297), .CK(CLK), .RN(n3026), .Q(n10338), 
        .QN(n2060) );
  DFFR_X1 \REGISTERS_reg[61][2]  ( .D(n8298), .CK(CLK), .RN(n3026), .Q(n10339), 
        .QN(n2061) );
  DFFR_X1 \REGISTERS_reg[61][1]  ( .D(n8299), .CK(CLK), .RN(n3026), .Q(n10340), 
        .QN(n2062) );
  DFFR_X1 \REGISTERS_reg[61][0]  ( .D(n8300), .CK(CLK), .RN(n3026), .Q(n10341), 
        .QN(n2063) );
  DFFR_X1 \REGISTERS_reg[62][31]  ( .D(n8301), .CK(CLK), .RN(n2994), .Q(n10342), .QN(n2064) );
  DFFR_X1 \REGISTERS_reg[62][30]  ( .D(n8302), .CK(CLK), .RN(n2992), .Q(n10343), .QN(n2065) );
  DFFR_X1 \REGISTERS_reg[62][29]  ( .D(n8303), .CK(CLK), .RN(n3004), .Q(n10344), .QN(n2066) );
  DFFR_X1 \REGISTERS_reg[62][28]  ( .D(n8304), .CK(CLK), .RN(n3005), .Q(n10345), .QN(n2067) );
  DFFR_X1 \REGISTERS_reg[62][27]  ( .D(n8305), .CK(CLK), .RN(n2993), .Q(n10346), .QN(n2068) );
  DFFR_X1 \REGISTERS_reg[62][26]  ( .D(n8306), .CK(CLK), .RN(n3001), .Q(n10347), .QN(n2069) );
  DFFR_X1 \REGISTERS_reg[62][25]  ( .D(n8307), .CK(CLK), .RN(n3002), .Q(n10348), .QN(n2070) );
  DFFR_X1 \REGISTERS_reg[62][24]  ( .D(n8308), .CK(CLK), .RN(n2999), .Q(n10349), .QN(n2071) );
  DFFR_X1 \REGISTERS_reg[62][23]  ( .D(n8309), .CK(CLK), .RN(n2995), .Q(n10350), .QN(n2072) );
  DFFR_X1 \REGISTERS_reg[62][22]  ( .D(n8310), .CK(CLK), .RN(n3003), .Q(n10351), .QN(n2073) );
  DFFR_X1 \REGISTERS_reg[62][21]  ( .D(n8311), .CK(CLK), .RN(n3000), .Q(n10352), .QN(n2074) );
  DFFR_X1 \REGISTERS_reg[62][20]  ( .D(n8312), .CK(CLK), .RN(n2991), .Q(n10353), .QN(n2075) );
  DFFR_X1 \REGISTERS_reg[62][19]  ( .D(n8313), .CK(CLK), .RN(n3025), .Q(n10354), .QN(n2076) );
  DFFR_X1 \REGISTERS_reg[62][18]  ( .D(n8314), .CK(CLK), .RN(n3025), .Q(n10355), .QN(n2077) );
  DFFR_X1 \REGISTERS_reg[62][17]  ( .D(n8315), .CK(CLK), .RN(n3025), .Q(n10356), .QN(n2078) );
  DFFR_X1 \REGISTERS_reg[62][16]  ( .D(n8316), .CK(CLK), .RN(n3025), .Q(n10357), .QN(n2079) );
  DFFR_X1 \REGISTERS_reg[62][15]  ( .D(n8317), .CK(CLK), .RN(n3025), .Q(n10358), .QN(n2080) );
  DFFR_X1 \REGISTERS_reg[62][14]  ( .D(n8318), .CK(CLK), .RN(n3025), .Q(n10359), .QN(n2081) );
  DFFR_X1 \REGISTERS_reg[62][13]  ( .D(n8319), .CK(CLK), .RN(n3025), .Q(n10360), .QN(n2082) );
  DFFR_X1 \REGISTERS_reg[62][12]  ( .D(n8320), .CK(CLK), .RN(n3025), .Q(n10361), .QN(n2083) );
  DFFR_X1 \REGISTERS_reg[62][11]  ( .D(n8321), .CK(CLK), .RN(n3025), .Q(n10362), .QN(n2084) );
  DFFR_X1 \REGISTERS_reg[62][10]  ( .D(n8322), .CK(CLK), .RN(n3025), .Q(n10363), .QN(n2085) );
  DFFR_X1 \REGISTERS_reg[62][9]  ( .D(n8323), .CK(CLK), .RN(n3025), .Q(n10364), 
        .QN(n2086) );
  DFFR_X1 \REGISTERS_reg[62][8]  ( .D(n8324), .CK(CLK), .RN(n3025), .Q(n10365), 
        .QN(n2087) );
  DFFR_X1 \REGISTERS_reg[62][7]  ( .D(n8325), .CK(CLK), .RN(n3024), .Q(n10366), 
        .QN(n2088) );
  DFFR_X1 \REGISTERS_reg[62][6]  ( .D(n8326), .CK(CLK), .RN(n3024), .Q(n10367), 
        .QN(n2089) );
  DFFR_X1 \REGISTERS_reg[62][5]  ( .D(n8327), .CK(CLK), .RN(n3024), .Q(n10368), 
        .QN(n2090) );
  DFFR_X1 \REGISTERS_reg[62][4]  ( .D(n8328), .CK(CLK), .RN(n3024), .Q(n10369), 
        .QN(n2091) );
  DFFR_X1 \REGISTERS_reg[62][3]  ( .D(n8329), .CK(CLK), .RN(n3024), .Q(n10370), 
        .QN(n2092) );
  DFFR_X1 \REGISTERS_reg[62][2]  ( .D(n8330), .CK(CLK), .RN(n3024), .Q(n10371), 
        .QN(n2093) );
  DFFR_X1 \REGISTERS_reg[62][1]  ( .D(n8331), .CK(CLK), .RN(n3024), .Q(n10372), 
        .QN(n2094) );
  DFFR_X1 \REGISTERS_reg[62][0]  ( .D(n8332), .CK(CLK), .RN(n3024), .Q(n10373), 
        .QN(n2095) );
  DFFR_X1 \REGISTERS_reg[63][31]  ( .D(n8333), .CK(CLK), .RN(n3024), .Q(n10374), .QN(n2096) );
  DFFR_X1 \REGISTERS_reg[63][30]  ( .D(n8334), .CK(CLK), .RN(n3024), .Q(n10375), .QN(n2097) );
  DFFR_X1 \REGISTERS_reg[63][29]  ( .D(n8335), .CK(CLK), .RN(n3024), .Q(n10376), .QN(n2098) );
  DFFR_X1 \REGISTERS_reg[63][28]  ( .D(n8336), .CK(CLK), .RN(n3024), .Q(n10377), .QN(n2099) );
  DFFR_X1 \REGISTERS_reg[63][27]  ( .D(n8337), .CK(CLK), .RN(n3023), .Q(n10378), .QN(n2100) );
  DFFR_X1 \REGISTERS_reg[63][26]  ( .D(n8338), .CK(CLK), .RN(n3023), .Q(n10379), .QN(n2101) );
  DFFR_X1 \REGISTERS_reg[63][25]  ( .D(n8339), .CK(CLK), .RN(n3023), .Q(n10380), .QN(n2102) );
  DFFR_X1 \REGISTERS_reg[63][24]  ( .D(n8340), .CK(CLK), .RN(n3023), .Q(n10381), .QN(n2103) );
  DFFR_X1 \REGISTERS_reg[63][23]  ( .D(n8341), .CK(CLK), .RN(n3023), .Q(n10382), .QN(n2104) );
  DFFR_X1 \REGISTERS_reg[63][22]  ( .D(n8342), .CK(CLK), .RN(n3023), .Q(n10383), .QN(n2105) );
  DFFR_X1 \REGISTERS_reg[63][21]  ( .D(n8343), .CK(CLK), .RN(n3023), .Q(n10384), .QN(n2106) );
  DFFR_X1 \REGISTERS_reg[63][20]  ( .D(n8344), .CK(CLK), .RN(n3023), .Q(n10385), .QN(n2107) );
  DFFR_X1 \REGISTERS_reg[63][19]  ( .D(n8345), .CK(CLK), .RN(n3023), .Q(n10386), .QN(n2108) );
  DFFR_X1 \REGISTERS_reg[63][18]  ( .D(n8346), .CK(CLK), .RN(n3023), .Q(n10387), .QN(n2109) );
  DFFR_X1 \REGISTERS_reg[63][17]  ( .D(n8347), .CK(CLK), .RN(n3023), .Q(n10388), .QN(n2110) );
  DFFR_X1 \REGISTERS_reg[63][16]  ( .D(n8348), .CK(CLK), .RN(n3023), .Q(n10389), .QN(n2111) );
  DFFR_X1 \REGISTERS_reg[63][15]  ( .D(n8349), .CK(CLK), .RN(n3022), .Q(n10390), .QN(n2112) );
  DFFR_X1 \REGISTERS_reg[63][14]  ( .D(n8350), .CK(CLK), .RN(n3022), .Q(n10391), .QN(n2113) );
  DFFR_X1 \REGISTERS_reg[63][13]  ( .D(n8351), .CK(CLK), .RN(n3022), .Q(n10392), .QN(n2114) );
  DFFR_X1 \REGISTERS_reg[63][12]  ( .D(n8352), .CK(CLK), .RN(n3022), .Q(n10393), .QN(n2115) );
  DFFR_X1 \REGISTERS_reg[63][11]  ( .D(n8353), .CK(CLK), .RN(n3022), .Q(n10394), .QN(n2116) );
  DFFR_X1 \REGISTERS_reg[63][10]  ( .D(n8354), .CK(CLK), .RN(n3022), .Q(n10395), .QN(n2117) );
  DFFR_X1 \REGISTERS_reg[63][9]  ( .D(n8355), .CK(CLK), .RN(n3022), .Q(n10396), 
        .QN(n2118) );
  DFFR_X1 \REGISTERS_reg[63][8]  ( .D(n8356), .CK(CLK), .RN(n3022), .Q(n10397), 
        .QN(n2119) );
  DFFR_X1 \REGISTERS_reg[63][7]  ( .D(n8357), .CK(CLK), .RN(n3022), .Q(n10398), 
        .QN(n2120) );
  DFFR_X1 \REGISTERS_reg[63][6]  ( .D(n8358), .CK(CLK), .RN(n3022), .Q(n10399), 
        .QN(n2121) );
  DFFR_X1 \REGISTERS_reg[63][5]  ( .D(n8359), .CK(CLK), .RN(n3022), .Q(n10400), 
        .QN(n2122) );
  DFFR_X1 \REGISTERS_reg[63][4]  ( .D(n8360), .CK(CLK), .RN(n3022), .Q(n10401), 
        .QN(n2123) );
  DFFR_X1 \REGISTERS_reg[63][3]  ( .D(n8361), .CK(CLK), .RN(n3021), .Q(n10402), 
        .QN(n2124) );
  DFFR_X1 \REGISTERS_reg[63][2]  ( .D(n8362), .CK(CLK), .RN(n3021), .Q(n10403), 
        .QN(n2125) );
  DFFR_X1 \REGISTERS_reg[63][1]  ( .D(n8363), .CK(CLK), .RN(n3021), .Q(n10404), 
        .QN(n2126) );
  DFFR_X1 \REGISTERS_reg[63][0]  ( .D(n8364), .CK(CLK), .RN(n3021), .Q(n10405), 
        .QN(n2127) );
  DFFR_X1 \REGISTERS_reg[64][31]  ( .D(n8365), .CK(CLK), .RN(n3021), .Q(n10406), .QN(n2128) );
  DFFR_X1 \REGISTERS_reg[64][30]  ( .D(n8366), .CK(CLK), .RN(n3021), .Q(n10407), .QN(n2129) );
  DFFR_X1 \REGISTERS_reg[64][29]  ( .D(n8367), .CK(CLK), .RN(n3021), .Q(n10408), .QN(n2130) );
  DFFR_X1 \REGISTERS_reg[64][28]  ( .D(n8368), .CK(CLK), .RN(n3021), .Q(n10409), .QN(n2131) );
  DFFR_X1 \REGISTERS_reg[64][27]  ( .D(n8369), .CK(CLK), .RN(n3021), .Q(n10410), .QN(n2132) );
  DFFR_X1 \REGISTERS_reg[64][26]  ( .D(n8370), .CK(CLK), .RN(n3021), .Q(n10411), .QN(n2133) );
  DFFR_X1 \REGISTERS_reg[64][25]  ( .D(n8371), .CK(CLK), .RN(n3021), .Q(n10412), .QN(n2134) );
  DFFR_X1 \REGISTERS_reg[64][24]  ( .D(n8372), .CK(CLK), .RN(n3021), .Q(n10413), .QN(n2135) );
  DFFR_X1 \REGISTERS_reg[64][23]  ( .D(n8373), .CK(CLK), .RN(n3020), .Q(n10414), .QN(n2136) );
  DFFR_X1 \REGISTERS_reg[64][22]  ( .D(n8374), .CK(CLK), .RN(n3020), .Q(n10415), .QN(n2137) );
  DFFR_X1 \REGISTERS_reg[64][21]  ( .D(n8375), .CK(CLK), .RN(n3020), .Q(n10416), .QN(n2138) );
  DFFR_X1 \REGISTERS_reg[64][20]  ( .D(n8376), .CK(CLK), .RN(n3020), .Q(n10417), .QN(n2139) );
  DFFR_X1 \REGISTERS_reg[64][19]  ( .D(n8377), .CK(CLK), .RN(n3020), .Q(n10418), .QN(n2140) );
  DFFR_X1 \REGISTERS_reg[64][18]  ( .D(n8378), .CK(CLK), .RN(n3020), .Q(n10419), .QN(n2141) );
  DFFR_X1 \REGISTERS_reg[64][17]  ( .D(n8379), .CK(CLK), .RN(n3020), .Q(n10420), .QN(n2142) );
  DFFR_X1 \REGISTERS_reg[64][16]  ( .D(n8380), .CK(CLK), .RN(n3020), .Q(n10421), .QN(n2143) );
  DFFR_X1 \REGISTERS_reg[64][15]  ( .D(n8381), .CK(CLK), .RN(n3020), .Q(n10422), .QN(n2144) );
  DFFR_X1 \REGISTERS_reg[64][14]  ( .D(n8382), .CK(CLK), .RN(n3020), .Q(n10423), .QN(n2145) );
  DFFR_X1 \REGISTERS_reg[64][13]  ( .D(n8383), .CK(CLK), .RN(n3020), .Q(n10424), .QN(n2146) );
  DFFR_X1 \REGISTERS_reg[64][12]  ( .D(n8384), .CK(CLK), .RN(n3020), .Q(n10425), .QN(n2147) );
  DFFR_X1 \REGISTERS_reg[64][11]  ( .D(n8385), .CK(CLK), .RN(n3019), .Q(n10426), .QN(n2148) );
  DFFR_X1 \REGISTERS_reg[64][10]  ( .D(n8386), .CK(CLK), .RN(n3019), .Q(n10427), .QN(n2149) );
  DFFR_X1 \REGISTERS_reg[64][9]  ( .D(n8387), .CK(CLK), .RN(n3019), .Q(n10428), 
        .QN(n2150) );
  DFFR_X1 \REGISTERS_reg[64][8]  ( .D(n8388), .CK(CLK), .RN(n3019), .Q(n10429), 
        .QN(n2151) );
  DFFR_X1 \REGISTERS_reg[64][7]  ( .D(n8389), .CK(CLK), .RN(n3019), .Q(n10430), 
        .QN(n2152) );
  DFFR_X1 \REGISTERS_reg[64][6]  ( .D(n8390), .CK(CLK), .RN(n3019), .Q(n10431), 
        .QN(n2153) );
  DFFR_X1 \REGISTERS_reg[64][5]  ( .D(n8391), .CK(CLK), .RN(n3019), .Q(n10432), 
        .QN(n2154) );
  DFFR_X1 \REGISTERS_reg[64][4]  ( .D(n8392), .CK(CLK), .RN(n3019), .Q(n10433), 
        .QN(n2155) );
  DFFR_X1 \REGISTERS_reg[64][3]  ( .D(n8393), .CK(CLK), .RN(n3019), .Q(n10434), 
        .QN(n2156) );
  DFFR_X1 \REGISTERS_reg[64][2]  ( .D(n8394), .CK(CLK), .RN(n3019), .Q(n10435), 
        .QN(n2157) );
  DFFR_X1 \REGISTERS_reg[64][1]  ( .D(n8395), .CK(CLK), .RN(n3019), .Q(n10436), 
        .QN(n2158) );
  DFFR_X1 \REGISTERS_reg[64][0]  ( .D(n8396), .CK(CLK), .RN(n3019), .Q(n10437), 
        .QN(n2159) );
  DFFR_X1 \REGISTERS_reg[65][31]  ( .D(n8397), .CK(CLK), .RN(n3018), .Q(n10438), .QN(n2160) );
  DFFR_X1 \REGISTERS_reg[65][30]  ( .D(n8398), .CK(CLK), .RN(n3018), .Q(n10439), .QN(n2161) );
  DFFR_X1 \REGISTERS_reg[65][29]  ( .D(n8399), .CK(CLK), .RN(n3018), .Q(n10440), .QN(n2162) );
  DFFR_X1 \REGISTERS_reg[65][28]  ( .D(n8400), .CK(CLK), .RN(n3018), .Q(n10441), .QN(n2163) );
  DFFR_X1 \REGISTERS_reg[65][27]  ( .D(n8401), .CK(CLK), .RN(n3018), .Q(n10442), .QN(n2164) );
  DFFR_X1 \REGISTERS_reg[65][26]  ( .D(n8402), .CK(CLK), .RN(n3018), .Q(n10443), .QN(n2165) );
  DFFR_X1 \REGISTERS_reg[65][25]  ( .D(n8403), .CK(CLK), .RN(n3018), .Q(n10444), .QN(n2166) );
  DFFR_X1 \REGISTERS_reg[65][24]  ( .D(n8404), .CK(CLK), .RN(n3018), .Q(n10445), .QN(n2167) );
  DFFR_X1 \REGISTERS_reg[65][23]  ( .D(n8405), .CK(CLK), .RN(n3018), .Q(n10446), .QN(n2168) );
  DFFR_X1 \REGISTERS_reg[65][22]  ( .D(n8406), .CK(CLK), .RN(n3018), .Q(n10447), .QN(n2169) );
  DFFR_X1 \REGISTERS_reg[65][21]  ( .D(n8407), .CK(CLK), .RN(n3018), .Q(n10448), .QN(n2170) );
  DFFR_X1 \REGISTERS_reg[65][20]  ( .D(n8408), .CK(CLK), .RN(n3018), .Q(n10449), .QN(n2171) );
  DFFR_X1 \REGISTERS_reg[65][19]  ( .D(n8409), .CK(CLK), .RN(n3017), .Q(n10450), .QN(n2172) );
  DFFR_X1 \REGISTERS_reg[65][18]  ( .D(n8410), .CK(CLK), .RN(n3017), .Q(n10451), .QN(n2173) );
  DFFR_X1 \REGISTERS_reg[65][17]  ( .D(n8411), .CK(CLK), .RN(n3017), .Q(n10452), .QN(n2174) );
  DFFR_X1 \REGISTERS_reg[65][16]  ( .D(n8412), .CK(CLK), .RN(n3017), .Q(n10453), .QN(n2175) );
  DFFR_X1 \REGISTERS_reg[65][15]  ( .D(n8413), .CK(CLK), .RN(n3017), .Q(n10454), .QN(n2176) );
  DFFR_X1 \REGISTERS_reg[65][14]  ( .D(n8414), .CK(CLK), .RN(n3017), .Q(n10455), .QN(n2177) );
  DFFR_X1 \REGISTERS_reg[65][13]  ( .D(n8415), .CK(CLK), .RN(n3017), .Q(n10456), .QN(n2178) );
  DFFR_X1 \REGISTERS_reg[65][12]  ( .D(n8416), .CK(CLK), .RN(n3017), .Q(n10457), .QN(n2179) );
  DFFR_X1 \REGISTERS_reg[65][11]  ( .D(n8417), .CK(CLK), .RN(n3017), .Q(n10458), .QN(n2180) );
  DFFR_X1 \REGISTERS_reg[65][10]  ( .D(n8418), .CK(CLK), .RN(n3017), .Q(n10459), .QN(n2181) );
  DFFR_X1 \REGISTERS_reg[65][9]  ( .D(n8419), .CK(CLK), .RN(n3017), .Q(n10460), 
        .QN(n2182) );
  DFFR_X1 \REGISTERS_reg[65][8]  ( .D(n8420), .CK(CLK), .RN(n3017), .Q(n10461), 
        .QN(n2183) );
  DFFR_X1 \REGISTERS_reg[65][7]  ( .D(n8421), .CK(CLK), .RN(n3016), .Q(n10462), 
        .QN(n2184) );
  DFFR_X1 \REGISTERS_reg[65][6]  ( .D(n8422), .CK(CLK), .RN(n3016), .Q(n10463), 
        .QN(n2185) );
  DFFR_X1 \REGISTERS_reg[65][5]  ( .D(n8423), .CK(CLK), .RN(n3016), .Q(n10464), 
        .QN(n2186) );
  DFFR_X1 \REGISTERS_reg[65][4]  ( .D(n8424), .CK(CLK), .RN(n3016), .Q(n10465), 
        .QN(n2187) );
  DFFR_X1 \REGISTERS_reg[65][3]  ( .D(n8425), .CK(CLK), .RN(n3016), .Q(n10466), 
        .QN(n2188) );
  DFFR_X1 \REGISTERS_reg[65][2]  ( .D(n8426), .CK(CLK), .RN(n3016), .Q(n10467), 
        .QN(n2189) );
  DFFR_X1 \REGISTERS_reg[65][1]  ( .D(n8427), .CK(CLK), .RN(n3016), .Q(n10468), 
        .QN(n2190) );
  DFFR_X1 \REGISTERS_reg[65][0]  ( .D(n8428), .CK(CLK), .RN(n3016), .Q(n10469), 
        .QN(n2191) );
  DFFR_X1 \REGISTERS_reg[66][31]  ( .D(n8429), .CK(CLK), .RN(n3016), .Q(n10470), .QN(n2192) );
  DFFR_X1 \REGISTERS_reg[66][30]  ( .D(n8430), .CK(CLK), .RN(n3016), .Q(n10471), .QN(n2193) );
  DFFR_X1 \REGISTERS_reg[66][29]  ( .D(n8431), .CK(CLK), .RN(n3016), .Q(n10472), .QN(n2194) );
  DFFR_X1 \REGISTERS_reg[66][28]  ( .D(n8432), .CK(CLK), .RN(n3016), .Q(n10473), .QN(n2195) );
  DFFR_X1 \REGISTERS_reg[66][27]  ( .D(n8433), .CK(CLK), .RN(n3015), .Q(n10474), .QN(n2196) );
  DFFR_X1 \REGISTERS_reg[66][26]  ( .D(n8434), .CK(CLK), .RN(n3015), .Q(n10475), .QN(n2197) );
  DFFR_X1 \REGISTERS_reg[66][25]  ( .D(n8435), .CK(CLK), .RN(n3015), .Q(n10476), .QN(n2198) );
  DFFR_X1 \REGISTERS_reg[66][24]  ( .D(n8436), .CK(CLK), .RN(n3015), .Q(n10477), .QN(n2199) );
  DFFR_X1 \REGISTERS_reg[66][23]  ( .D(n8437), .CK(CLK), .RN(n3015), .Q(n10478), .QN(n2200) );
  DFFR_X1 \REGISTERS_reg[66][22]  ( .D(n8438), .CK(CLK), .RN(n3015), .Q(n10479), .QN(n2201) );
  DFFR_X1 \REGISTERS_reg[66][21]  ( .D(n8439), .CK(CLK), .RN(n3015), .Q(n10480), .QN(n2202) );
  DFFR_X1 \REGISTERS_reg[66][20]  ( .D(n8440), .CK(CLK), .RN(n3015), .Q(n10481), .QN(n2203) );
  DFFR_X1 \REGISTERS_reg[66][19]  ( .D(n8441), .CK(CLK), .RN(n3015), .Q(n10482), .QN(n2204) );
  DFFR_X1 \REGISTERS_reg[66][18]  ( .D(n8442), .CK(CLK), .RN(n3015), .Q(n10483), .QN(n2205) );
  DFFR_X1 \REGISTERS_reg[66][17]  ( .D(n8443), .CK(CLK), .RN(n3015), .Q(n10484), .QN(n2206) );
  DFFR_X1 \REGISTERS_reg[66][16]  ( .D(n8444), .CK(CLK), .RN(n3015), .Q(n10485), .QN(n2207) );
  DFFR_X1 \REGISTERS_reg[66][15]  ( .D(n8445), .CK(CLK), .RN(n3014), .Q(n10486), .QN(n2208) );
  DFFR_X1 \REGISTERS_reg[66][14]  ( .D(n8446), .CK(CLK), .RN(n3014), .Q(n10487), .QN(n2209) );
  DFFR_X1 \REGISTERS_reg[66][13]  ( .D(n8447), .CK(CLK), .RN(n3014), .Q(n10488), .QN(n2210) );
  DFFR_X1 \REGISTERS_reg[66][12]  ( .D(n8448), .CK(CLK), .RN(n3014), .Q(n10489), .QN(n2211) );
  DFFR_X1 \REGISTERS_reg[66][11]  ( .D(n8449), .CK(CLK), .RN(n3014), .Q(n10490), .QN(n2212) );
  DFFR_X1 \REGISTERS_reg[66][10]  ( .D(n8450), .CK(CLK), .RN(n3014), .Q(n10491), .QN(n2213) );
  DFFR_X1 \REGISTERS_reg[66][9]  ( .D(n8451), .CK(CLK), .RN(n3014), .Q(n10492), 
        .QN(n2214) );
  DFFR_X1 \REGISTERS_reg[66][8]  ( .D(n8452), .CK(CLK), .RN(n3014), .Q(n10493), 
        .QN(n2215) );
  DFFR_X1 \REGISTERS_reg[66][7]  ( .D(n8453), .CK(CLK), .RN(n3014), .Q(n10494), 
        .QN(n2216) );
  DFFR_X1 \REGISTERS_reg[66][6]  ( .D(n8454), .CK(CLK), .RN(n3014), .Q(n10495), 
        .QN(n2217) );
  DFFR_X1 \REGISTERS_reg[66][5]  ( .D(n8455), .CK(CLK), .RN(n3014), .Q(n10496), 
        .QN(n2218) );
  DFFR_X1 \REGISTERS_reg[66][4]  ( .D(n8456), .CK(CLK), .RN(n3014), .Q(n10497), 
        .QN(n2219) );
  DFFR_X1 \REGISTERS_reg[66][3]  ( .D(n8457), .CK(CLK), .RN(n3013), .Q(n10498), 
        .QN(n2220) );
  DFFR_X1 \REGISTERS_reg[66][2]  ( .D(n8458), .CK(CLK), .RN(n3013), .Q(n10499), 
        .QN(n2221) );
  DFFR_X1 \REGISTERS_reg[66][1]  ( .D(n8459), .CK(CLK), .RN(n3013), .Q(n10500), 
        .QN(n2222) );
  DFFR_X1 \REGISTERS_reg[66][0]  ( .D(n8460), .CK(CLK), .RN(n3013), .Q(n10501), 
        .QN(n2223) );
  DFFR_X1 \REGISTERS_reg[67][31]  ( .D(n8461), .CK(CLK), .RN(n3013), .Q(n10502), .QN(n2224) );
  DFFR_X1 \REGISTERS_reg[67][30]  ( .D(n8462), .CK(CLK), .RN(n3013), .Q(n10503), .QN(n2225) );
  DFFR_X1 \REGISTERS_reg[67][29]  ( .D(n8463), .CK(CLK), .RN(n3013), .Q(n10504), .QN(n2226) );
  DFFR_X1 \REGISTERS_reg[67][28]  ( .D(n8464), .CK(CLK), .RN(n3013), .Q(n10505), .QN(n2227) );
  DFFR_X1 \REGISTERS_reg[67][27]  ( .D(n8465), .CK(CLK), .RN(n3013), .Q(n10506), .QN(n2228) );
  DFFR_X1 \REGISTERS_reg[67][26]  ( .D(n8466), .CK(CLK), .RN(n3013), .Q(n10507), .QN(n2229) );
  DFFR_X1 \REGISTERS_reg[67][25]  ( .D(n8467), .CK(CLK), .RN(n3013), .Q(n10508), .QN(n2230) );
  DFFR_X1 \REGISTERS_reg[67][24]  ( .D(n8468), .CK(CLK), .RN(n3013), .Q(n10509), .QN(n2231) );
  DFFR_X1 \REGISTERS_reg[67][23]  ( .D(n8469), .CK(CLK), .RN(n3012), .Q(n10510), .QN(n2232) );
  DFFR_X1 \REGISTERS_reg[67][22]  ( .D(n8470), .CK(CLK), .RN(n3012), .Q(n10511), .QN(n2233) );
  DFFR_X1 \REGISTERS_reg[67][21]  ( .D(n8471), .CK(CLK), .RN(n3012), .Q(n10512), .QN(n2234) );
  DFFR_X1 \REGISTERS_reg[67][20]  ( .D(n8472), .CK(CLK), .RN(n3012), .Q(n10513), .QN(n2235) );
  DFFR_X1 \REGISTERS_reg[67][19]  ( .D(n8473), .CK(CLK), .RN(n3012), .Q(n10514), .QN(n2236) );
  DFFR_X1 \REGISTERS_reg[67][18]  ( .D(n8474), .CK(CLK), .RN(n3012), .Q(n10515), .QN(n2237) );
  DFFR_X1 \REGISTERS_reg[67][17]  ( .D(n8475), .CK(CLK), .RN(n3012), .Q(n10516), .QN(n2238) );
  DFFR_X1 \REGISTERS_reg[67][16]  ( .D(n8476), .CK(CLK), .RN(n3012), .Q(n10517), .QN(n2239) );
  DFFR_X1 \REGISTERS_reg[67][15]  ( .D(n8477), .CK(CLK), .RN(n3012), .Q(n10518), .QN(n2240) );
  DFFR_X1 \REGISTERS_reg[67][14]  ( .D(n8478), .CK(CLK), .RN(n3012), .Q(n10519), .QN(n2241) );
  DFFR_X1 \REGISTERS_reg[67][13]  ( .D(n8479), .CK(CLK), .RN(n3012), .Q(n10520), .QN(n2242) );
  DFFR_X1 \REGISTERS_reg[67][12]  ( .D(n8480), .CK(CLK), .RN(n3012), .Q(n10521), .QN(n2243) );
  DFFR_X1 \REGISTERS_reg[67][11]  ( .D(n8481), .CK(CLK), .RN(n3011), .Q(n10522), .QN(n2244) );
  DFFR_X1 \REGISTERS_reg[67][10]  ( .D(n8482), .CK(CLK), .RN(n3011), .Q(n10523), .QN(n2245) );
  DFFR_X1 \REGISTERS_reg[67][9]  ( .D(n8483), .CK(CLK), .RN(n3011), .Q(n10524), 
        .QN(n2246) );
  DFFR_X1 \REGISTERS_reg[67][8]  ( .D(n8484), .CK(CLK), .RN(n3011), .Q(n10525), 
        .QN(n2247) );
  DFFR_X1 \REGISTERS_reg[67][7]  ( .D(n8485), .CK(CLK), .RN(n3011), .Q(n10526), 
        .QN(n2248) );
  DFFR_X1 \REGISTERS_reg[67][6]  ( .D(n8486), .CK(CLK), .RN(n3011), .Q(n10527), 
        .QN(n2249) );
  DFFR_X1 \REGISTERS_reg[67][5]  ( .D(n8487), .CK(CLK), .RN(n3011), .Q(n10528), 
        .QN(n2250) );
  DFFR_X1 \REGISTERS_reg[67][4]  ( .D(n8488), .CK(CLK), .RN(n3011), .Q(n10529), 
        .QN(n2251) );
  DFFR_X1 \REGISTERS_reg[67][3]  ( .D(n8489), .CK(CLK), .RN(n3011), .Q(n10530), 
        .QN(n2252) );
  DFFR_X1 \REGISTERS_reg[67][2]  ( .D(n8490), .CK(CLK), .RN(n3011), .Q(n10531), 
        .QN(n2253) );
  DFFR_X1 \REGISTERS_reg[67][1]  ( .D(n8491), .CK(CLK), .RN(n3011), .Q(n10532), 
        .QN(n2254) );
  DFFR_X1 \REGISTERS_reg[67][0]  ( .D(n8492), .CK(CLK), .RN(n3011), .Q(n10533), 
        .QN(n2255) );
  DFFR_X1 \REGISTERS_reg[68][31]  ( .D(n8493), .CK(CLK), .RN(n3010), .Q(n10534), .QN(n2256) );
  DFFR_X1 \REGISTERS_reg[68][30]  ( .D(n8494), .CK(CLK), .RN(n3010), .Q(n10535), .QN(n2257) );
  DFFR_X1 \REGISTERS_reg[68][29]  ( .D(n8495), .CK(CLK), .RN(n3010), .Q(n10536), .QN(n2258) );
  DFFR_X1 \REGISTERS_reg[68][28]  ( .D(n8496), .CK(CLK), .RN(n3010), .Q(n10537), .QN(n2259) );
  DFFR_X1 \REGISTERS_reg[68][27]  ( .D(n8497), .CK(CLK), .RN(n3010), .Q(n10538), .QN(n2260) );
  DFFR_X1 \REGISTERS_reg[68][26]  ( .D(n8498), .CK(CLK), .RN(n3010), .Q(n10539), .QN(n2261) );
  DFFR_X1 \REGISTERS_reg[68][25]  ( .D(n8499), .CK(CLK), .RN(n3010), .Q(n10540), .QN(n2262) );
  DFFR_X1 \REGISTERS_reg[68][24]  ( .D(n8500), .CK(CLK), .RN(n3010), .Q(n10541), .QN(n2263) );
  DFFR_X1 \REGISTERS_reg[68][23]  ( .D(n8501), .CK(CLK), .RN(n3010), .Q(n10542), .QN(n2264) );
  DFFR_X1 \REGISTERS_reg[68][22]  ( .D(n8502), .CK(CLK), .RN(n3010), .Q(n10543), .QN(n2265) );
  DFFR_X1 \REGISTERS_reg[68][21]  ( .D(n8503), .CK(CLK), .RN(n3010), .Q(n10544), .QN(n2266) );
  DFFR_X1 \REGISTERS_reg[68][20]  ( .D(n8504), .CK(CLK), .RN(n3010), .Q(n10545), .QN(n2267) );
  DFFR_X1 \REGISTERS_reg[68][19]  ( .D(n8505), .CK(CLK), .RN(n3009), .Q(n10546), .QN(n2268) );
  DFFR_X1 \REGISTERS_reg[68][18]  ( .D(n8506), .CK(CLK), .RN(n3009), .Q(n10547), .QN(n2269) );
  DFFR_X1 \REGISTERS_reg[68][17]  ( .D(n8507), .CK(CLK), .RN(n3009), .Q(n10548), .QN(n2270) );
  DFFR_X1 \REGISTERS_reg[68][16]  ( .D(n8508), .CK(CLK), .RN(n3009), .Q(n10549), .QN(n2271) );
  DFFR_X1 \REGISTERS_reg[68][15]  ( .D(n8509), .CK(CLK), .RN(n3009), .Q(n10550), .QN(n2272) );
  DFFR_X1 \REGISTERS_reg[68][14]  ( .D(n8510), .CK(CLK), .RN(n3009), .Q(n10551), .QN(n2273) );
  DFFR_X1 \REGISTERS_reg[68][13]  ( .D(n8511), .CK(CLK), .RN(n3009), .Q(n10552), .QN(n2274) );
  DFFR_X1 \REGISTERS_reg[68][12]  ( .D(n8512), .CK(CLK), .RN(n3009), .Q(n10553), .QN(n2275) );
  DFFR_X1 \REGISTERS_reg[68][11]  ( .D(n8513), .CK(CLK), .RN(n3009), .Q(n10554), .QN(n2276) );
  DFFR_X1 \REGISTERS_reg[68][10]  ( .D(n8514), .CK(CLK), .RN(n3009), .Q(n10555), .QN(n2277) );
  DFFR_X1 \REGISTERS_reg[68][9]  ( .D(n8515), .CK(CLK), .RN(n3009), .Q(n10556), 
        .QN(n2278) );
  DFFR_X1 \REGISTERS_reg[68][8]  ( .D(n8516), .CK(CLK), .RN(n3009), .Q(n10557), 
        .QN(n2279) );
  DFFR_X1 \REGISTERS_reg[68][7]  ( .D(n8517), .CK(CLK), .RN(n3008), .Q(n10558), 
        .QN(n2280) );
  DFFR_X1 \REGISTERS_reg[68][6]  ( .D(n8518), .CK(CLK), .RN(n3008), .Q(n10559), 
        .QN(n2281) );
  DFFR_X1 \REGISTERS_reg[68][5]  ( .D(n8519), .CK(CLK), .RN(n3008), .Q(n10560), 
        .QN(n2282) );
  DFFR_X1 \REGISTERS_reg[68][4]  ( .D(n8520), .CK(CLK), .RN(n3008), .Q(n10561), 
        .QN(n2283) );
  DFFR_X1 \REGISTERS_reg[68][3]  ( .D(n8521), .CK(CLK), .RN(n3008), .Q(n10562), 
        .QN(n2284) );
  DFFR_X1 \REGISTERS_reg[68][2]  ( .D(n8522), .CK(CLK), .RN(n3008), .Q(n10563), 
        .QN(n2285) );
  DFFR_X1 \REGISTERS_reg[68][1]  ( .D(n8523), .CK(CLK), .RN(n3008), .Q(n10564), 
        .QN(n2286) );
  DFFR_X1 \REGISTERS_reg[68][0]  ( .D(n8524), .CK(CLK), .RN(n3008), .Q(n10565), 
        .QN(n2287) );
  DFFR_X1 \REGISTERS_reg[69][31]  ( .D(n8525), .CK(CLK), .RN(n3008), .Q(n10566), .QN(n2288) );
  DFFR_X1 \REGISTERS_reg[69][30]  ( .D(n8526), .CK(CLK), .RN(n3008), .Q(n10567), .QN(n2289) );
  DFFR_X1 \REGISTERS_reg[69][29]  ( .D(n8527), .CK(CLK), .RN(n3008), .Q(n10568), .QN(n2290) );
  DFFR_X1 \REGISTERS_reg[69][28]  ( .D(n8528), .CK(CLK), .RN(n3008), .Q(n10569), .QN(n2291) );
  DFFR_X1 \REGISTERS_reg[69][27]  ( .D(n8529), .CK(CLK), .RN(n3007), .Q(n10570), .QN(n2292) );
  DFFR_X1 \REGISTERS_reg[69][26]  ( .D(n8530), .CK(CLK), .RN(n3007), .Q(n10571), .QN(n2293) );
  DFFR_X1 \REGISTERS_reg[69][25]  ( .D(n8531), .CK(CLK), .RN(n3007), .Q(n10572), .QN(n2294) );
  DFFR_X1 \REGISTERS_reg[69][24]  ( .D(n8532), .CK(CLK), .RN(n3007), .Q(n10573), .QN(n2295) );
  DFFR_X1 \REGISTERS_reg[69][23]  ( .D(n8533), .CK(CLK), .RN(n3007), .Q(n10574), .QN(n2296) );
  DFFR_X1 \REGISTERS_reg[69][22]  ( .D(n8534), .CK(CLK), .RN(n3007), .Q(n10575), .QN(n2297) );
  DFFR_X1 \REGISTERS_reg[69][21]  ( .D(n8535), .CK(CLK), .RN(n3007), .Q(n10576), .QN(n2298) );
  DFFR_X1 \REGISTERS_reg[69][20]  ( .D(n8536), .CK(CLK), .RN(n3007), .Q(n10577), .QN(n2299) );
  DFFR_X1 \REGISTERS_reg[69][19]  ( .D(n8537), .CK(CLK), .RN(n3007), .Q(n10578), .QN(n2300) );
  DFFR_X1 \REGISTERS_reg[69][18]  ( .D(n8538), .CK(CLK), .RN(n3007), .Q(n10579), .QN(n2301) );
  DFFR_X1 \REGISTERS_reg[69][17]  ( .D(n8539), .CK(CLK), .RN(n3007), .Q(n10580), .QN(n2302) );
  DFFR_X1 \REGISTERS_reg[69][16]  ( .D(n8540), .CK(CLK), .RN(n3007), .Q(n10581), .QN(n2303) );
  DFFR_X1 \REGISTERS_reg[69][15]  ( .D(n8541), .CK(CLK), .RN(n3006), .Q(n10582), .QN(n2304) );
  DFFR_X1 \REGISTERS_reg[69][14]  ( .D(n8542), .CK(CLK), .RN(n3006), .Q(n10583), .QN(n2305) );
  DFFR_X1 \REGISTERS_reg[69][13]  ( .D(n8543), .CK(CLK), .RN(n3006), .Q(n10584), .QN(n2306) );
  DFFR_X1 \REGISTERS_reg[69][12]  ( .D(n8544), .CK(CLK), .RN(n3006), .Q(n10585), .QN(n2307) );
  DFFR_X1 \REGISTERS_reg[69][11]  ( .D(n8545), .CK(CLK), .RN(n3006), .Q(n10586), .QN(n2308) );
  DFFR_X1 \REGISTERS_reg[69][10]  ( .D(n8546), .CK(CLK), .RN(n3006), .Q(n10587), .QN(n2309) );
  DFFR_X1 \REGISTERS_reg[69][9]  ( .D(n8547), .CK(CLK), .RN(n3006), .Q(n10588), 
        .QN(n2310) );
  DFFR_X1 \REGISTERS_reg[69][8]  ( .D(n8548), .CK(CLK), .RN(n3006), .Q(n10589), 
        .QN(n2311) );
  DFFR_X1 \REGISTERS_reg[69][7]  ( .D(n8549), .CK(CLK), .RN(n3006), .Q(n10590), 
        .QN(n2312) );
  DFFR_X1 \REGISTERS_reg[69][6]  ( .D(n8550), .CK(CLK), .RN(n3006), .Q(n10591), 
        .QN(n2313) );
  DFFR_X1 \REGISTERS_reg[69][5]  ( .D(n8551), .CK(CLK), .RN(n3006), .Q(n10592), 
        .QN(n2314) );
  DFFR_X1 \REGISTERS_reg[69][4]  ( .D(n8552), .CK(CLK), .RN(n3006), .Q(n10593), 
        .QN(n2315) );
  DFFR_X1 \REGISTERS_reg[69][3]  ( .D(n8553), .CK(CLK), .RN(n3005), .Q(n10594), 
        .QN(n2316) );
  DFFR_X1 \REGISTERS_reg[69][2]  ( .D(n8554), .CK(CLK), .RN(n3005), .Q(n10595), 
        .QN(n2317) );
  DFFR_X1 \REGISTERS_reg[69][1]  ( .D(n8555), .CK(CLK), .RN(n3005), .Q(n10596), 
        .QN(n2318) );
  DFFR_X1 \REGISTERS_reg[69][0]  ( .D(n8556), .CK(CLK), .RN(n3005), .Q(n10597), 
        .QN(n2319) );
  DFFR_X1 \REGISTERS_reg[70][31]  ( .D(n8557), .CK(CLK), .RN(n3005), .Q(n10598), .QN(n2320) );
  DFFR_X1 \REGISTERS_reg[70][30]  ( .D(n8558), .CK(CLK), .RN(n3005), .Q(n10599), .QN(n2321) );
  DFFR_X1 \REGISTERS_reg[70][29]  ( .D(n8559), .CK(CLK), .RN(n3005), .Q(n10600), .QN(n2322) );
  DFFR_X1 \REGISTERS_reg[70][28]  ( .D(n8560), .CK(CLK), .RN(n3005), .Q(n10601), .QN(n2323) );
  DFFR_X1 \REGISTERS_reg[70][27]  ( .D(n8561), .CK(CLK), .RN(n3005), .Q(n10602), .QN(n2324) );
  DFFR_X1 \REGISTERS_reg[70][26]  ( .D(n8562), .CK(CLK), .RN(n3005), .Q(n10603), .QN(n2325) );
  DFFR_X1 \REGISTERS_reg[70][25]  ( .D(n8563), .CK(CLK), .RN(n3005), .Q(n10604), .QN(n2326) );
  DFFR_X1 \REGISTERS_reg[70][24]  ( .D(n8564), .CK(CLK), .RN(n3005), .Q(n10605), .QN(n2327) );
  DFFR_X1 \REGISTERS_reg[70][23]  ( .D(n8565), .CK(CLK), .RN(n3004), .Q(n10606), .QN(n2328) );
  DFFR_X1 \REGISTERS_reg[70][22]  ( .D(n8566), .CK(CLK), .RN(n3004), .Q(n10607), .QN(n2329) );
  DFFR_X1 \REGISTERS_reg[70][21]  ( .D(n8567), .CK(CLK), .RN(n3004), .Q(n10608), .QN(n2330) );
  DFFR_X1 \REGISTERS_reg[70][20]  ( .D(n8568), .CK(CLK), .RN(n3004), .Q(n10609), .QN(n2331) );
  DFFR_X1 \REGISTERS_reg[70][19]  ( .D(n8569), .CK(CLK), .RN(n3004), .Q(n10610), .QN(n2332) );
  DFFR_X1 \REGISTERS_reg[70][18]  ( .D(n8570), .CK(CLK), .RN(n3004), .Q(n10611), .QN(n2333) );
  DFFR_X1 \REGISTERS_reg[70][17]  ( .D(n8571), .CK(CLK), .RN(n3004), .Q(n10612), .QN(n2334) );
  DFFR_X1 \REGISTERS_reg[70][16]  ( .D(n8572), .CK(CLK), .RN(n3004), .Q(n10613), .QN(n2335) );
  DFFR_X1 \REGISTERS_reg[70][15]  ( .D(n8573), .CK(CLK), .RN(n3004), .Q(n10614), .QN(n2336) );
  DFFR_X1 \REGISTERS_reg[70][14]  ( .D(n8574), .CK(CLK), .RN(n3004), .Q(n10615), .QN(n2337) );
  DFFR_X1 \REGISTERS_reg[70][13]  ( .D(n8575), .CK(CLK), .RN(n3004), .Q(n10616), .QN(n2338) );
  DFFR_X1 \REGISTERS_reg[70][12]  ( .D(n8576), .CK(CLK), .RN(n3004), .Q(n10617), .QN(n2339) );
  DFFR_X1 \REGISTERS_reg[70][11]  ( .D(n8577), .CK(CLK), .RN(n3003), .Q(n10618), .QN(n2340) );
  DFFR_X1 \REGISTERS_reg[70][10]  ( .D(n8578), .CK(CLK), .RN(n3003), .Q(n10619), .QN(n2341) );
  DFFR_X1 \REGISTERS_reg[70][9]  ( .D(n8579), .CK(CLK), .RN(n3003), .Q(n10620), 
        .QN(n2342) );
  DFFR_X1 \REGISTERS_reg[70][8]  ( .D(n8580), .CK(CLK), .RN(n3003), .Q(n10621), 
        .QN(n2343) );
  DFFR_X1 \REGISTERS_reg[70][7]  ( .D(n8581), .CK(CLK), .RN(n3003), .Q(n10622), 
        .QN(n2344) );
  DFFR_X1 \REGISTERS_reg[70][6]  ( .D(n8582), .CK(CLK), .RN(n3003), .Q(n10623), 
        .QN(n2345) );
  DFFR_X1 \REGISTERS_reg[70][5]  ( .D(n8583), .CK(CLK), .RN(n3003), .Q(n10624), 
        .QN(n2346) );
  DFFR_X1 \REGISTERS_reg[70][4]  ( .D(n8584), .CK(CLK), .RN(n3003), .Q(n10625), 
        .QN(n2347) );
  DFFR_X1 \REGISTERS_reg[70][3]  ( .D(n8585), .CK(CLK), .RN(n3003), .Q(n10626), 
        .QN(n2348) );
  DFFR_X1 \REGISTERS_reg[70][2]  ( .D(n8586), .CK(CLK), .RN(n3003), .Q(n10627), 
        .QN(n2349) );
  DFFR_X1 \REGISTERS_reg[70][1]  ( .D(n8587), .CK(CLK), .RN(n3003), .Q(n10628), 
        .QN(n2350) );
  DFFR_X1 \REGISTERS_reg[70][0]  ( .D(n8588), .CK(CLK), .RN(n3003), .Q(n10629), 
        .QN(n2351) );
  DFFR_X1 \REGISTERS_reg[71][31]  ( .D(n8589), .CK(CLK), .RN(n3002), .Q(n10630), .QN(n2352) );
  DFFR_X1 \REGISTERS_reg[71][30]  ( .D(n8590), .CK(CLK), .RN(n3002), .Q(n10631), .QN(n2353) );
  DFFR_X1 \REGISTERS_reg[71][29]  ( .D(n8591), .CK(CLK), .RN(n3002), .Q(n10632), .QN(n2354) );
  DFFR_X1 \REGISTERS_reg[71][28]  ( .D(n8592), .CK(CLK), .RN(n3002), .Q(n10633), .QN(n2355) );
  DFFR_X1 \REGISTERS_reg[71][27]  ( .D(n8593), .CK(CLK), .RN(n3002), .Q(n10634), .QN(n2356) );
  DFFR_X1 \REGISTERS_reg[71][26]  ( .D(n8594), .CK(CLK), .RN(n3002), .Q(n10635), .QN(n2357) );
  DFFR_X1 \REGISTERS_reg[71][25]  ( .D(n8595), .CK(CLK), .RN(n3002), .Q(n10636), .QN(n2358) );
  DFFR_X1 \REGISTERS_reg[71][24]  ( .D(n8596), .CK(CLK), .RN(n3002), .Q(n10637), .QN(n2359) );
  DFFR_X1 \REGISTERS_reg[71][23]  ( .D(n8597), .CK(CLK), .RN(n3002), .Q(n10638), .QN(n2360) );
  DFFR_X1 \REGISTERS_reg[71][22]  ( .D(n8598), .CK(CLK), .RN(n3002), .Q(n10639), .QN(n2361) );
  DFFR_X1 \REGISTERS_reg[71][21]  ( .D(n8599), .CK(CLK), .RN(n3002), .Q(n10640), .QN(n2362) );
  DFFR_X1 \REGISTERS_reg[71][20]  ( .D(n8600), .CK(CLK), .RN(n3002), .Q(n10641), .QN(n2363) );
  DFFR_X1 \REGISTERS_reg[71][19]  ( .D(n8601), .CK(CLK), .RN(n3001), .Q(n10642), .QN(n2364) );
  DFFR_X1 \REGISTERS_reg[71][18]  ( .D(n8602), .CK(CLK), .RN(n3001), .Q(n10643), .QN(n2365) );
  DFFR_X1 \REGISTERS_reg[71][17]  ( .D(n8603), .CK(CLK), .RN(n3001), .Q(n10644), .QN(n2366) );
  DFFR_X1 \REGISTERS_reg[71][16]  ( .D(n8604), .CK(CLK), .RN(n3001), .Q(n10645), .QN(n2367) );
  DFFR_X1 \REGISTERS_reg[71][15]  ( .D(n8605), .CK(CLK), .RN(n3001), .Q(n10646), .QN(n2368) );
  DFFR_X1 \REGISTERS_reg[71][14]  ( .D(n8606), .CK(CLK), .RN(n3001), .Q(n10647), .QN(n2369) );
  DFFR_X1 \REGISTERS_reg[71][13]  ( .D(n8607), .CK(CLK), .RN(n3001), .Q(n10648), .QN(n2370) );
  DFFR_X1 \REGISTERS_reg[71][12]  ( .D(n8608), .CK(CLK), .RN(n3001), .Q(n10649), .QN(n2371) );
  DFFR_X1 \REGISTERS_reg[71][11]  ( .D(n8609), .CK(CLK), .RN(n3001), .Q(n10650), .QN(n2372) );
  DFFR_X1 \REGISTERS_reg[71][10]  ( .D(n8610), .CK(CLK), .RN(n3001), .Q(n10651), .QN(n2373) );
  DFFR_X1 \REGISTERS_reg[71][9]  ( .D(n8611), .CK(CLK), .RN(n3001), .Q(n10652), 
        .QN(n2374) );
  DFFR_X1 \REGISTERS_reg[71][8]  ( .D(n8612), .CK(CLK), .RN(n3001), .Q(n10653), 
        .QN(n2375) );
  DFFR_X1 \REGISTERS_reg[71][7]  ( .D(n8613), .CK(CLK), .RN(n3000), .Q(n10654), 
        .QN(n2376) );
  DFFR_X1 \REGISTERS_reg[71][6]  ( .D(n8614), .CK(CLK), .RN(n3000), .Q(n10655), 
        .QN(n2377) );
  DFFR_X1 \REGISTERS_reg[71][5]  ( .D(n8615), .CK(CLK), .RN(n3000), .Q(n10656), 
        .QN(n2378) );
  DFFR_X1 \REGISTERS_reg[71][4]  ( .D(n8616), .CK(CLK), .RN(n3000), .Q(n10657), 
        .QN(n2379) );
  DFFR_X1 \REGISTERS_reg[71][3]  ( .D(n8617), .CK(CLK), .RN(n3000), .Q(n10658), 
        .QN(n2380) );
  DFFR_X1 \REGISTERS_reg[71][2]  ( .D(n8618), .CK(CLK), .RN(n3000), .Q(n10659), 
        .QN(n2381) );
  DFFR_X1 \REGISTERS_reg[71][1]  ( .D(n8619), .CK(CLK), .RN(n3000), .Q(n10660), 
        .QN(n2382) );
  DFFR_X1 \REGISTERS_reg[71][0]  ( .D(n8620), .CK(CLK), .RN(n3000), .Q(n10661), 
        .QN(n2383) );
  DFFR_X1 \REGISTERS_reg[72][31]  ( .D(n8621), .CK(CLK), .RN(n3000), .Q(n10662), .QN(n2384) );
  DFFR_X1 \REGISTERS_reg[72][30]  ( .D(n8622), .CK(CLK), .RN(n3000), .Q(n10663), .QN(n2385) );
  DFFR_X1 \REGISTERS_reg[72][29]  ( .D(n8623), .CK(CLK), .RN(n3000), .Q(n10664), .QN(n2386) );
  DFFR_X1 \REGISTERS_reg[72][28]  ( .D(n8624), .CK(CLK), .RN(n3000), .Q(n10665), .QN(n2387) );
  DFFR_X1 \REGISTERS_reg[72][27]  ( .D(n8625), .CK(CLK), .RN(n2999), .Q(n10666), .QN(n2388) );
  DFFR_X1 \REGISTERS_reg[72][26]  ( .D(n8626), .CK(CLK), .RN(n2999), .Q(n10667), .QN(n2389) );
  DFFR_X1 \REGISTERS_reg[72][25]  ( .D(n8627), .CK(CLK), .RN(n2999), .Q(n10668), .QN(n2390) );
  DFFR_X1 \REGISTERS_reg[72][24]  ( .D(n8628), .CK(CLK), .RN(n2999), .Q(n10669), .QN(n2391) );
  DFFR_X1 \REGISTERS_reg[72][23]  ( .D(n8629), .CK(CLK), .RN(n2999), .Q(n10670), .QN(n2392) );
  DFFR_X1 \REGISTERS_reg[72][22]  ( .D(n8630), .CK(CLK), .RN(n2999), .Q(n10671), .QN(n2393) );
  DFFR_X1 \REGISTERS_reg[72][21]  ( .D(n8631), .CK(CLK), .RN(n2999), .Q(n10672), .QN(n2394) );
  DFFR_X1 \REGISTERS_reg[72][20]  ( .D(n8632), .CK(CLK), .RN(n2999), .Q(n10673), .QN(n2395) );
  DFFR_X1 \REGISTERS_reg[72][19]  ( .D(n8633), .CK(CLK), .RN(n2999), .Q(n10674), .QN(n2396) );
  DFFR_X1 \REGISTERS_reg[72][18]  ( .D(n8634), .CK(CLK), .RN(n2999), .Q(n10675), .QN(n2397) );
  DFFR_X1 \REGISTERS_reg[72][17]  ( .D(n8635), .CK(CLK), .RN(n2999), .Q(n10676), .QN(n2398) );
  DFFR_X1 \REGISTERS_reg[72][16]  ( .D(n8636), .CK(CLK), .RN(n2999), .Q(n10677), .QN(n2399) );
  DFFR_X1 \REGISTERS_reg[72][15]  ( .D(n8637), .CK(CLK), .RN(n2998), .Q(n10678), .QN(n2400) );
  DFFR_X1 \REGISTERS_reg[72][14]  ( .D(n8638), .CK(CLK), .RN(n2998), .Q(n10679), .QN(n2401) );
  DFFR_X1 \REGISTERS_reg[72][13]  ( .D(n8639), .CK(CLK), .RN(n2998), .Q(n10680), .QN(n2402) );
  DFFR_X1 \REGISTERS_reg[72][12]  ( .D(n8640), .CK(CLK), .RN(n2998), .Q(n10681), .QN(n2403) );
  DFFR_X1 \REGISTERS_reg[72][11]  ( .D(n8641), .CK(CLK), .RN(n2998), .Q(n10682), .QN(n2404) );
  DFFR_X1 \REGISTERS_reg[72][10]  ( .D(n8642), .CK(CLK), .RN(n2998), .Q(n10683), .QN(n2405) );
  DFFR_X1 \REGISTERS_reg[72][9]  ( .D(n8643), .CK(CLK), .RN(n2998), .Q(n10684), 
        .QN(n2406) );
  DFFR_X1 \REGISTERS_reg[72][8]  ( .D(n8644), .CK(CLK), .RN(n2998), .Q(n10685), 
        .QN(n2407) );
  DFFR_X1 \REGISTERS_reg[72][7]  ( .D(n8645), .CK(CLK), .RN(n2998), .Q(n10686), 
        .QN(n2408) );
  DFFR_X1 \REGISTERS_reg[72][6]  ( .D(n8646), .CK(CLK), .RN(n2998), .Q(n10687), 
        .QN(n2409) );
  DFFR_X1 \REGISTERS_reg[72][5]  ( .D(n8647), .CK(CLK), .RN(n2998), .Q(n10688), 
        .QN(n2410) );
  DFFR_X1 \REGISTERS_reg[72][4]  ( .D(n8648), .CK(CLK), .RN(n2998), .Q(n10689), 
        .QN(n2411) );
  DFFR_X1 \REGISTERS_reg[72][3]  ( .D(n8649), .CK(CLK), .RN(n2997), .Q(n10690), 
        .QN(n2412) );
  DFFR_X1 \REGISTERS_reg[72][2]  ( .D(n8650), .CK(CLK), .RN(n2997), .Q(n10691), 
        .QN(n2413) );
  DFFR_X1 \REGISTERS_reg[72][1]  ( .D(n8651), .CK(CLK), .RN(n2997), .Q(n10692), 
        .QN(n2414) );
  DFFR_X1 \REGISTERS_reg[72][0]  ( .D(n8652), .CK(CLK), .RN(n2997), .Q(n10693), 
        .QN(n2415) );
  DFFR_X1 \REGISTERS_reg[73][31]  ( .D(n8653), .CK(CLK), .RN(n2997), .Q(n10694), .QN(n2416) );
  DFFR_X1 \REGISTERS_reg[73][30]  ( .D(n8654), .CK(CLK), .RN(n2997), .Q(n10695), .QN(n2417) );
  DFFR_X1 \REGISTERS_reg[73][29]  ( .D(n8655), .CK(CLK), .RN(n2997), .Q(n10696), .QN(n2418) );
  DFFR_X1 \REGISTERS_reg[73][28]  ( .D(n8656), .CK(CLK), .RN(n2997), .Q(n10697), .QN(n2419) );
  DFFR_X1 \REGISTERS_reg[73][27]  ( .D(n8657), .CK(CLK), .RN(n2997), .Q(n10698), .QN(n2420) );
  DFFR_X1 \REGISTERS_reg[73][26]  ( .D(n8658), .CK(CLK), .RN(n2997), .Q(n10699), .QN(n2421) );
  DFFR_X1 \REGISTERS_reg[73][25]  ( .D(n8659), .CK(CLK), .RN(n2997), .Q(n10700), .QN(n2422) );
  DFFR_X1 \REGISTERS_reg[73][24]  ( .D(n8660), .CK(CLK), .RN(n2997), .Q(n10701), .QN(n2423) );
  DFFR_X1 \REGISTERS_reg[73][23]  ( .D(n8661), .CK(CLK), .RN(n2995), .Q(n10702), .QN(n2424) );
  DFFR_X1 \REGISTERS_reg[73][22]  ( .D(n8662), .CK(CLK), .RN(n2995), .Q(n10703), .QN(n2425) );
  DFFR_X1 \REGISTERS_reg[73][21]  ( .D(n8663), .CK(CLK), .RN(n2995), .Q(n10704), .QN(n2426) );
  DFFR_X1 \REGISTERS_reg[73][20]  ( .D(n8664), .CK(CLK), .RN(n2995), .Q(n10705), .QN(n2427) );
  DFFR_X1 \REGISTERS_reg[73][19]  ( .D(n8665), .CK(CLK), .RN(n2995), .Q(n10706), .QN(n2428) );
  DFFR_X1 \REGISTERS_reg[73][18]  ( .D(n8666), .CK(CLK), .RN(n2995), .Q(n10707), .QN(n2429) );
  DFFR_X1 \REGISTERS_reg[73][17]  ( .D(n8667), .CK(CLK), .RN(n2995), .Q(n10708), .QN(n2430) );
  DFFR_X1 \REGISTERS_reg[73][16]  ( .D(n8668), .CK(CLK), .RN(n2995), .Q(n10709), .QN(n2431) );
  DFFR_X1 \REGISTERS_reg[73][15]  ( .D(n8669), .CK(CLK), .RN(n2995), .Q(n10710), .QN(n2432) );
  DFFR_X1 \REGISTERS_reg[73][14]  ( .D(n8670), .CK(CLK), .RN(n2995), .Q(n10711), .QN(n2433) );
  DFFR_X1 \REGISTERS_reg[73][13]  ( .D(n8671), .CK(CLK), .RN(n2995), .Q(n10712), .QN(n2434) );
  DFFR_X1 \REGISTERS_reg[73][12]  ( .D(n8672), .CK(CLK), .RN(n2995), .Q(n10713), .QN(n2435) );
  DFFR_X1 \REGISTERS_reg[73][11]  ( .D(n8673), .CK(CLK), .RN(n2994), .Q(n10714), .QN(n2436) );
  DFFR_X1 \REGISTERS_reg[73][10]  ( .D(n8674), .CK(CLK), .RN(n2994), .Q(n10715), .QN(n2437) );
  DFFR_X1 \REGISTERS_reg[73][9]  ( .D(n8675), .CK(CLK), .RN(n2994), .Q(n10716), 
        .QN(n2438) );
  DFFR_X1 \REGISTERS_reg[73][8]  ( .D(n8676), .CK(CLK), .RN(n2994), .Q(n10717), 
        .QN(n2439) );
  DFFR_X1 \REGISTERS_reg[73][7]  ( .D(n8677), .CK(CLK), .RN(n2994), .Q(n10718), 
        .QN(n2440) );
  DFFR_X1 \REGISTERS_reg[73][6]  ( .D(n8678), .CK(CLK), .RN(n2994), .Q(n10719), 
        .QN(n2441) );
  DFFR_X1 \REGISTERS_reg[73][5]  ( .D(n8679), .CK(CLK), .RN(n2994), .Q(n10720), 
        .QN(n2442) );
  DFFR_X1 \REGISTERS_reg[73][4]  ( .D(n8680), .CK(CLK), .RN(n2994), .Q(n10721), 
        .QN(n2443) );
  DFFR_X1 \REGISTERS_reg[73][3]  ( .D(n8681), .CK(CLK), .RN(n2994), .Q(n10722), 
        .QN(n2444) );
  DFFR_X1 \REGISTERS_reg[73][2]  ( .D(n8682), .CK(CLK), .RN(n2994), .Q(n10723), 
        .QN(n2445) );
  DFFR_X1 \REGISTERS_reg[73][1]  ( .D(n8683), .CK(CLK), .RN(n2994), .Q(n10724), 
        .QN(n2446) );
  DFFR_X1 \REGISTERS_reg[73][0]  ( .D(n8684), .CK(CLK), .RN(n2994), .Q(n10725), 
        .QN(n2447) );
  DFFR_X1 \REGISTERS_reg[74][31]  ( .D(n8685), .CK(CLK), .RN(n2993), .Q(n10726), .QN(n2448) );
  DFFR_X1 \REGISTERS_reg[74][30]  ( .D(n8686), .CK(CLK), .RN(n2993), .Q(n10727), .QN(n2449) );
  DFFR_X1 \REGISTERS_reg[74][29]  ( .D(n8687), .CK(CLK), .RN(n2993), .Q(n10728), .QN(n2450) );
  DFFR_X1 \REGISTERS_reg[74][28]  ( .D(n8688), .CK(CLK), .RN(n2993), .Q(n10729), .QN(n2451) );
  DFFR_X1 \REGISTERS_reg[74][27]  ( .D(n8689), .CK(CLK), .RN(n2993), .Q(n10730), .QN(n2452) );
  DFFR_X1 \REGISTERS_reg[74][26]  ( .D(n8690), .CK(CLK), .RN(n2993), .Q(n10731), .QN(n2453) );
  DFFR_X1 \REGISTERS_reg[74][25]  ( .D(n8691), .CK(CLK), .RN(n2993), .Q(n10732), .QN(n2454) );
  DFFR_X1 \REGISTERS_reg[74][24]  ( .D(n8692), .CK(CLK), .RN(n2993), .Q(n10733), .QN(n2455) );
  DFFR_X1 \REGISTERS_reg[74][23]  ( .D(n8693), .CK(CLK), .RN(n2993), .Q(n10734), .QN(n2456) );
  DFFR_X1 \REGISTERS_reg[74][22]  ( .D(n8694), .CK(CLK), .RN(n2993), .Q(n10735), .QN(n2457) );
  DFFR_X1 \REGISTERS_reg[74][21]  ( .D(n8695), .CK(CLK), .RN(n2993), .Q(n10736), .QN(n2458) );
  DFFR_X1 \REGISTERS_reg[74][20]  ( .D(n8696), .CK(CLK), .RN(n2993), .Q(n10737), .QN(n2459) );
  DFFR_X1 \REGISTERS_reg[74][19]  ( .D(n8697), .CK(CLK), .RN(n2992), .Q(n10738), .QN(n2460) );
  DFFR_X1 \REGISTERS_reg[74][18]  ( .D(n8698), .CK(CLK), .RN(n2992), .Q(n10739), .QN(n2461) );
  DFFR_X1 \REGISTERS_reg[74][17]  ( .D(n8699), .CK(CLK), .RN(n2992), .Q(n10740), .QN(n2462) );
  DFFR_X1 \REGISTERS_reg[74][16]  ( .D(n8700), .CK(CLK), .RN(n2992), .Q(n10741), .QN(n2463) );
  DFFR_X1 \REGISTERS_reg[74][15]  ( .D(n8701), .CK(CLK), .RN(n2992), .Q(n10742), .QN(n2464) );
  DFFR_X1 \REGISTERS_reg[74][14]  ( .D(n8702), .CK(CLK), .RN(n2992), .Q(n10743), .QN(n2465) );
  DFFR_X1 \REGISTERS_reg[74][13]  ( .D(n8703), .CK(CLK), .RN(n2992), .Q(n10744), .QN(n2466) );
  DFFR_X1 \REGISTERS_reg[74][12]  ( .D(n8704), .CK(CLK), .RN(n2992), .Q(n10745), .QN(n2467) );
  DFFR_X1 \REGISTERS_reg[74][11]  ( .D(n8705), .CK(CLK), .RN(n2992), .Q(n10746), .QN(n2468) );
  DFFR_X1 \REGISTERS_reg[74][10]  ( .D(n8706), .CK(CLK), .RN(n2992), .Q(n10747), .QN(n2469) );
  DFFR_X1 \REGISTERS_reg[74][9]  ( .D(n8707), .CK(CLK), .RN(n2992), .Q(n10748), 
        .QN(n2470) );
  DFFR_X1 \REGISTERS_reg[74][8]  ( .D(n8708), .CK(CLK), .RN(n2992), .Q(n10749), 
        .QN(n2471) );
  DFFR_X1 \REGISTERS_reg[74][7]  ( .D(n8709), .CK(CLK), .RN(n2991), .Q(n10750), 
        .QN(n2472) );
  DFFR_X1 \REGISTERS_reg[74][6]  ( .D(n8710), .CK(CLK), .RN(n2991), .Q(n10751), 
        .QN(n2473) );
  DFFR_X1 \REGISTERS_reg[74][5]  ( .D(n8711), .CK(CLK), .RN(n2991), .Q(n10752), 
        .QN(n2474) );
  DFFR_X1 \REGISTERS_reg[74][4]  ( .D(n8712), .CK(CLK), .RN(n2991), .Q(n10753), 
        .QN(n2475) );
  DFFR_X1 \REGISTERS_reg[74][3]  ( .D(n8713), .CK(CLK), .RN(n2991), .Q(n10754), 
        .QN(n2476) );
  DFFR_X1 \REGISTERS_reg[74][2]  ( .D(n8714), .CK(CLK), .RN(n2991), .Q(n10755), 
        .QN(n2477) );
  DFFR_X1 \REGISTERS_reg[74][1]  ( .D(n8715), .CK(CLK), .RN(n2991), .Q(n10756), 
        .QN(n2478) );
  DFFR_X1 \REGISTERS_reg[74][0]  ( .D(n8716), .CK(CLK), .RN(n2991), .Q(n10757), 
        .QN(n2479) );
  DFFR_X1 \REGISTERS_reg[75][31]  ( .D(n8717), .CK(CLK), .RN(n2991), .Q(n10758), .QN(n2480) );
  DFFR_X1 \REGISTERS_reg[75][30]  ( .D(n8718), .CK(CLK), .RN(n2991), .Q(n10759), .QN(n2481) );
  DFFR_X1 \REGISTERS_reg[75][29]  ( .D(n8719), .CK(CLK), .RN(n2991), .Q(n10760), .QN(n2482) );
  DFFR_X1 \REGISTERS_reg[75][28]  ( .D(n8720), .CK(CLK), .RN(n2991), .Q(n10761), .QN(n2483) );
  DFFR_X1 \REGISTERS_reg[75][27]  ( .D(n8721), .CK(CLK), .RN(n2990), .Q(n10762), .QN(n2484) );
  DFFR_X1 \REGISTERS_reg[75][26]  ( .D(n8722), .CK(CLK), .RN(n2990), .Q(n10763), .QN(n2485) );
  DFFR_X1 \REGISTERS_reg[75][25]  ( .D(n8723), .CK(CLK), .RN(n2990), .Q(n10764), .QN(n2486) );
  DFFR_X1 \REGISTERS_reg[75][24]  ( .D(n8724), .CK(CLK), .RN(n2990), .Q(n10765), .QN(n2487) );
  DFFR_X1 \REGISTERS_reg[75][23]  ( .D(n8725), .CK(CLK), .RN(n2990), .Q(n10766), .QN(n2488) );
  DFFR_X1 \REGISTERS_reg[75][22]  ( .D(n8726), .CK(CLK), .RN(n2990), .Q(n10767), .QN(n2489) );
  DFFR_X1 \REGISTERS_reg[75][21]  ( .D(n8727), .CK(CLK), .RN(n2990), .Q(n10768), .QN(n2490) );
  DFFR_X1 \REGISTERS_reg[75][20]  ( .D(n8728), .CK(CLK), .RN(n2990), .Q(n10769), .QN(n2491) );
  DFFR_X1 \REGISTERS_reg[75][19]  ( .D(n8729), .CK(CLK), .RN(n2990), .Q(n10770), .QN(n2492) );
  DFFR_X1 \REGISTERS_reg[75][18]  ( .D(n8730), .CK(CLK), .RN(n2990), .Q(n10771), .QN(n2493) );
  DFFR_X1 \REGISTERS_reg[75][17]  ( .D(n8731), .CK(CLK), .RN(n2990), .Q(n10772), .QN(n2494) );
  DFFR_X1 \REGISTERS_reg[75][16]  ( .D(n8732), .CK(CLK), .RN(n2990), .Q(n10773), .QN(n2495) );
  DFFR_X1 \REGISTERS_reg[75][15]  ( .D(n8733), .CK(CLK), .RN(n2989), .Q(n10774), .QN(n2496) );
  DFFR_X1 \REGISTERS_reg[75][14]  ( .D(n8734), .CK(CLK), .RN(n2989), .Q(n10775), .QN(n2497) );
  DFFR_X1 \REGISTERS_reg[75][13]  ( .D(n8735), .CK(CLK), .RN(n2989), .Q(n10776), .QN(n2498) );
  DFFR_X1 \REGISTERS_reg[75][12]  ( .D(n8736), .CK(CLK), .RN(n2989), .Q(n10777), .QN(n2499) );
  DFFR_X1 \REGISTERS_reg[75][11]  ( .D(n8737), .CK(CLK), .RN(n2989), .Q(n10778), .QN(n2500) );
  DFFR_X1 \REGISTERS_reg[75][10]  ( .D(n8738), .CK(CLK), .RN(n2989), .Q(n10779), .QN(n2501) );
  DFFR_X1 \REGISTERS_reg[75][9]  ( .D(n8739), .CK(CLK), .RN(n2989), .Q(n10780), 
        .QN(n2502) );
  DFFR_X1 \REGISTERS_reg[75][8]  ( .D(n8740), .CK(CLK), .RN(n2989), .Q(n10781), 
        .QN(n2503) );
  DFFR_X1 \REGISTERS_reg[75][7]  ( .D(n8741), .CK(CLK), .RN(n2989), .Q(n10782), 
        .QN(n2504) );
  DFFR_X1 \REGISTERS_reg[75][6]  ( .D(n8742), .CK(CLK), .RN(n2989), .Q(n10783), 
        .QN(n2505) );
  DFFR_X1 \REGISTERS_reg[75][5]  ( .D(n8743), .CK(CLK), .RN(n2989), .Q(n10784), 
        .QN(n2506) );
  DFFR_X1 \REGISTERS_reg[75][4]  ( .D(n8744), .CK(CLK), .RN(n2989), .Q(n10785), 
        .QN(n2507) );
  DFFR_X1 \REGISTERS_reg[75][3]  ( .D(n8745), .CK(CLK), .RN(n2988), .Q(n10786), 
        .QN(n2508) );
  DFFR_X1 \REGISTERS_reg[75][2]  ( .D(n8746), .CK(CLK), .RN(n2988), .Q(n10787), 
        .QN(n2509) );
  DFFR_X1 \REGISTERS_reg[75][1]  ( .D(n8747), .CK(CLK), .RN(n2988), .Q(n10788), 
        .QN(n2510) );
  DFFR_X1 \REGISTERS_reg[75][0]  ( .D(n8748), .CK(CLK), .RN(n2988), .Q(n10789), 
        .QN(n2511) );
  DFFR_X1 \REGISTERS_reg[76][31]  ( .D(n8749), .CK(CLK), .RN(n2988), .Q(n10790), .QN(n2512) );
  DFFR_X1 \REGISTERS_reg[76][30]  ( .D(n8750), .CK(CLK), .RN(n2988), .Q(n10791), .QN(n2513) );
  DFFR_X1 \REGISTERS_reg[76][29]  ( .D(n8751), .CK(CLK), .RN(n2988), .Q(n10792), .QN(n2514) );
  DFFR_X1 \REGISTERS_reg[76][28]  ( .D(n8752), .CK(CLK), .RN(n2988), .Q(n10793), .QN(n2515) );
  DFFR_X1 \REGISTERS_reg[76][27]  ( .D(n8753), .CK(CLK), .RN(n2988), .Q(n10794), .QN(n2516) );
  DFFR_X1 \REGISTERS_reg[76][26]  ( .D(n8754), .CK(CLK), .RN(n2988), .Q(n10795), .QN(n2517) );
  DFFR_X1 \REGISTERS_reg[76][25]  ( .D(n8755), .CK(CLK), .RN(n2988), .Q(n10796), .QN(n2518) );
  DFFR_X1 \REGISTERS_reg[76][24]  ( .D(n8756), .CK(CLK), .RN(n2988), .Q(n10797), .QN(n2519) );
  DFFR_X1 \REGISTERS_reg[76][23]  ( .D(n8757), .CK(CLK), .RN(n2987), .Q(n10798), .QN(n2520) );
  DFFR_X1 \REGISTERS_reg[76][22]  ( .D(n8758), .CK(CLK), .RN(n2987), .Q(n10799), .QN(n2521) );
  DFFR_X1 \REGISTERS_reg[76][21]  ( .D(n8759), .CK(CLK), .RN(n2987), .Q(n10800), .QN(n2522) );
  DFFR_X1 \REGISTERS_reg[76][20]  ( .D(n8760), .CK(CLK), .RN(n2987), .Q(n10801), .QN(n2523) );
  DFFR_X1 \REGISTERS_reg[76][19]  ( .D(n8761), .CK(CLK), .RN(n2987), .Q(n10802), .QN(n2524) );
  DFFR_X1 \REGISTERS_reg[76][18]  ( .D(n8762), .CK(CLK), .RN(n2987), .Q(n10803), .QN(n2525) );
  DFFR_X1 \REGISTERS_reg[76][17]  ( .D(n8763), .CK(CLK), .RN(n2987), .Q(n10804), .QN(n2526) );
  DFFR_X1 \REGISTERS_reg[76][16]  ( .D(n8764), .CK(CLK), .RN(n2987), .Q(n10805), .QN(n2527) );
  DFFR_X1 \REGISTERS_reg[76][15]  ( .D(n8765), .CK(CLK), .RN(n2987), .Q(n10806), .QN(n2528) );
  DFFR_X1 \REGISTERS_reg[76][14]  ( .D(n8766), .CK(CLK), .RN(n2987), .Q(n10807), .QN(n2529) );
  DFFR_X1 \REGISTERS_reg[76][13]  ( .D(n8767), .CK(CLK), .RN(n2987), .Q(n10808), .QN(n2530) );
  DFFR_X1 \REGISTERS_reg[76][12]  ( .D(n8768), .CK(CLK), .RN(n2987), .Q(n10809), .QN(n2531) );
  DFFR_X1 \REGISTERS_reg[76][11]  ( .D(n8769), .CK(CLK), .RN(n2986), .Q(n10810), .QN(n2532) );
  DFFR_X1 \REGISTERS_reg[76][10]  ( .D(n8770), .CK(CLK), .RN(n2986), .Q(n10811), .QN(n2533) );
  DFFR_X1 \REGISTERS_reg[76][9]  ( .D(n8771), .CK(CLK), .RN(n2986), .Q(n10812), 
        .QN(n2534) );
  DFFR_X1 \REGISTERS_reg[76][8]  ( .D(n8772), .CK(CLK), .RN(n2986), .Q(n10813), 
        .QN(n2535) );
  DFFR_X1 \REGISTERS_reg[76][7]  ( .D(n8773), .CK(CLK), .RN(n2986), .Q(n10814), 
        .QN(n2536) );
  DFFR_X1 \REGISTERS_reg[76][6]  ( .D(n8774), .CK(CLK), .RN(n2986), .Q(n10815), 
        .QN(n2537) );
  DFFR_X1 \REGISTERS_reg[76][5]  ( .D(n8775), .CK(CLK), .RN(n2986), .Q(n10816), 
        .QN(n2538) );
  DFFR_X1 \REGISTERS_reg[76][4]  ( .D(n8776), .CK(CLK), .RN(n2986), .Q(n10817), 
        .QN(n2539) );
  DFFR_X1 \REGISTERS_reg[76][3]  ( .D(n8777), .CK(CLK), .RN(n2986), .Q(n10818), 
        .QN(n2540) );
  DFFR_X1 \REGISTERS_reg[76][2]  ( .D(n8778), .CK(CLK), .RN(n2986), .Q(n10819), 
        .QN(n2541) );
  DFFR_X1 \REGISTERS_reg[76][1]  ( .D(n8779), .CK(CLK), .RN(n2986), .Q(n10820), 
        .QN(n2542) );
  DFFR_X1 \REGISTERS_reg[76][0]  ( .D(n8780), .CK(CLK), .RN(n2986), .Q(n10821), 
        .QN(n2543) );
  DFFR_X1 \REGISTERS_reg[79][31]  ( .D(n8845), .CK(CLK), .RN(n2980), .Q(n10822), .QN(n2608) );
  DFFR_X1 \REGISTERS_reg[79][30]  ( .D(n8846), .CK(CLK), .RN(n2980), .Q(n10823), .QN(n2609) );
  DFFR_X1 \REGISTERS_reg[79][29]  ( .D(n8847), .CK(CLK), .RN(n2980), .Q(n10824), .QN(n2610) );
  DFFR_X1 \REGISTERS_reg[79][28]  ( .D(n8848), .CK(CLK), .RN(n2980), .Q(n10825), .QN(n2611) );
  DFFR_X1 \REGISTERS_reg[79][27]  ( .D(n8849), .CK(CLK), .RN(n2980), .Q(n10826), .QN(n2612) );
  DFFR_X1 \REGISTERS_reg[79][26]  ( .D(n8850), .CK(CLK), .RN(n2980), .Q(n10827), .QN(n2613) );
  DFFR_X1 \REGISTERS_reg[79][25]  ( .D(n8851), .CK(CLK), .RN(n2980), .Q(n10828), .QN(n2614) );
  DFFR_X1 \REGISTERS_reg[79][24]  ( .D(n8852), .CK(CLK), .RN(n2980), .Q(n10829), .QN(n2615) );
  DFFR_X1 \REGISTERS_reg[79][23]  ( .D(n8853), .CK(CLK), .RN(n2979), .Q(n10830), .QN(n2616) );
  DFFR_X1 \REGISTERS_reg[79][22]  ( .D(n8854), .CK(CLK), .RN(n2979), .Q(n10831), .QN(n2617) );
  DFFR_X1 \REGISTERS_reg[79][21]  ( .D(n8855), .CK(CLK), .RN(n2979), .Q(n10832), .QN(n2618) );
  DFFR_X1 \REGISTERS_reg[79][20]  ( .D(n8856), .CK(CLK), .RN(n2979), .Q(n10833), .QN(n2619) );
  DFFR_X1 \REGISTERS_reg[79][19]  ( .D(n8857), .CK(CLK), .RN(n2979), .Q(n10834), .QN(n2620) );
  DFFR_X1 \REGISTERS_reg[79][18]  ( .D(n8858), .CK(CLK), .RN(n2979), .Q(n10835), .QN(n2621) );
  DFFR_X1 \REGISTERS_reg[79][17]  ( .D(n8859), .CK(CLK), .RN(n2979), .Q(n10836), .QN(n2622) );
  DFFR_X1 \REGISTERS_reg[79][16]  ( .D(n8860), .CK(CLK), .RN(n2979), .Q(n10837), .QN(n2623) );
  DFFR_X1 \REGISTERS_reg[79][15]  ( .D(n8861), .CK(CLK), .RN(n2979), .Q(n10838), .QN(n2624) );
  DFFR_X1 \REGISTERS_reg[79][14]  ( .D(n8862), .CK(CLK), .RN(n2979), .Q(n10839), .QN(n2625) );
  DFFR_X1 \REGISTERS_reg[79][13]  ( .D(n8863), .CK(CLK), .RN(n2979), .Q(n10840), .QN(n2626) );
  DFFR_X1 \REGISTERS_reg[79][12]  ( .D(n8864), .CK(CLK), .RN(n2979), .Q(n10841), .QN(n2627) );
  DFFR_X1 \REGISTERS_reg[79][11]  ( .D(n8865), .CK(CLK), .RN(n2978), .Q(n10842), .QN(n2628) );
  DFFR_X1 \REGISTERS_reg[79][10]  ( .D(n8866), .CK(CLK), .RN(n2978), .Q(n10843), .QN(n2629) );
  DFFR_X1 \REGISTERS_reg[79][9]  ( .D(n8867), .CK(CLK), .RN(n2978), .Q(n10844), 
        .QN(n2630) );
  DFFR_X1 \REGISTERS_reg[79][8]  ( .D(n8868), .CK(CLK), .RN(n2978), .Q(n10845), 
        .QN(n2631) );
  DFFR_X1 \REGISTERS_reg[79][7]  ( .D(n8869), .CK(CLK), .RN(n2978), .Q(n10846), 
        .QN(n2632) );
  DFFR_X1 \REGISTERS_reg[79][6]  ( .D(n8870), .CK(CLK), .RN(n2978), .Q(n10847), 
        .QN(n2633) );
  DFFR_X1 \REGISTERS_reg[79][5]  ( .D(n8871), .CK(CLK), .RN(n2978), .Q(n10848), 
        .QN(n2634) );
  DFFR_X1 \REGISTERS_reg[79][4]  ( .D(n8872), .CK(CLK), .RN(n2978), .Q(n10849), 
        .QN(n2635) );
  DFFR_X1 \REGISTERS_reg[79][3]  ( .D(n8873), .CK(CLK), .RN(n2978), .Q(n10850), 
        .QN(n2636) );
  DFFR_X1 \REGISTERS_reg[79][2]  ( .D(n8874), .CK(CLK), .RN(n2978), .Q(n10851), 
        .QN(n2637) );
  DFFR_X1 \REGISTERS_reg[79][1]  ( .D(n8875), .CK(CLK), .RN(n2978), .Q(n10852), 
        .QN(n2638) );
  DFFR_X1 \REGISTERS_reg[79][0]  ( .D(n8876), .CK(CLK), .RN(n2978), .Q(n10853), 
        .QN(n2639) );
  DFFR_X1 \REGISTERS_reg[80][31]  ( .D(n8877), .CK(CLK), .RN(n2977), .Q(n10854), .QN(n2640) );
  DFFR_X1 \REGISTERS_reg[80][30]  ( .D(n8878), .CK(CLK), .RN(n2977), .Q(n10855), .QN(n2641) );
  DFFR_X1 \REGISTERS_reg[80][29]  ( .D(n8879), .CK(CLK), .RN(n2977), .Q(n10856), .QN(n2642) );
  DFFR_X1 \REGISTERS_reg[80][28]  ( .D(n8880), .CK(CLK), .RN(n2977), .Q(n10857), .QN(n2643) );
  DFFR_X1 \REGISTERS_reg[80][27]  ( .D(n8881), .CK(CLK), .RN(n2977), .Q(n10858), .QN(n2644) );
  DFFR_X1 \REGISTERS_reg[80][26]  ( .D(n8882), .CK(CLK), .RN(n2977), .Q(n10859), .QN(n2645) );
  DFFR_X1 \REGISTERS_reg[80][25]  ( .D(n8883), .CK(CLK), .RN(n2977), .Q(n10860), .QN(n2646) );
  DFFR_X1 \REGISTERS_reg[80][24]  ( .D(n8884), .CK(CLK), .RN(n2977), .Q(n10861), .QN(n2647) );
  DFFR_X1 \REGISTERS_reg[80][23]  ( .D(n8885), .CK(CLK), .RN(n2977), .Q(n10862), .QN(n2648) );
  DFFR_X1 \REGISTERS_reg[80][22]  ( .D(n8886), .CK(CLK), .RN(n2977), .Q(n10863), .QN(n2649) );
  DFFR_X1 \REGISTERS_reg[80][21]  ( .D(n8887), .CK(CLK), .RN(n2977), .Q(n10864), .QN(n2650) );
  DFFR_X1 \REGISTERS_reg[80][20]  ( .D(n8888), .CK(CLK), .RN(n2977), .Q(n10865), .QN(n2651) );
  DFFR_X1 \REGISTERS_reg[80][19]  ( .D(n8889), .CK(CLK), .RN(n2976), .Q(n10866), .QN(n2652) );
  DFFR_X1 \REGISTERS_reg[80][18]  ( .D(n8890), .CK(CLK), .RN(n2976), .Q(n10867), .QN(n2653) );
  DFFR_X1 \REGISTERS_reg[80][17]  ( .D(n8891), .CK(CLK), .RN(n2976), .Q(n10868), .QN(n2654) );
  DFFR_X1 \REGISTERS_reg[80][16]  ( .D(n8892), .CK(CLK), .RN(n2976), .Q(n10869), .QN(n2655) );
  DFFR_X1 \REGISTERS_reg[80][15]  ( .D(n8893), .CK(CLK), .RN(n2976), .Q(n10870), .QN(n2656) );
  DFFR_X1 \REGISTERS_reg[80][14]  ( .D(n8894), .CK(CLK), .RN(n2976), .Q(n10871), .QN(n2657) );
  DFFR_X1 \REGISTERS_reg[80][13]  ( .D(n8895), .CK(CLK), .RN(n2976), .Q(n10872), .QN(n2658) );
  DFFR_X1 \REGISTERS_reg[80][12]  ( .D(n8896), .CK(CLK), .RN(n2976), .Q(n10873), .QN(n2659) );
  DFFR_X1 \REGISTERS_reg[80][11]  ( .D(n8897), .CK(CLK), .RN(n2976), .Q(n10874), .QN(n2660) );
  DFFR_X1 \REGISTERS_reg[80][10]  ( .D(n8898), .CK(CLK), .RN(n2976), .Q(n10875), .QN(n2661) );
  DFFR_X1 \REGISTERS_reg[80][9]  ( .D(n8899), .CK(CLK), .RN(n2976), .Q(n10876), 
        .QN(n2662) );
  DFFR_X1 \REGISTERS_reg[80][8]  ( .D(n8900), .CK(CLK), .RN(n2976), .Q(n10877), 
        .QN(n2663) );
  DFFR_X1 \REGISTERS_reg[80][7]  ( .D(n8901), .CK(CLK), .RN(n2975), .Q(n10878), 
        .QN(n2664) );
  DFFR_X1 \REGISTERS_reg[80][6]  ( .D(n8902), .CK(CLK), .RN(n2975), .Q(n10879), 
        .QN(n2665) );
  DFFR_X1 \REGISTERS_reg[80][5]  ( .D(n8903), .CK(CLK), .RN(n2975), .Q(n10880), 
        .QN(n2666) );
  DFFR_X1 \REGISTERS_reg[80][4]  ( .D(n8904), .CK(CLK), .RN(n2975), .Q(n10881), 
        .QN(n2667) );
  DFFR_X1 \REGISTERS_reg[80][3]  ( .D(n8905), .CK(CLK), .RN(n2975), .Q(n10882), 
        .QN(n2668) );
  DFFR_X1 \REGISTERS_reg[80][2]  ( .D(n8906), .CK(CLK), .RN(n2975), .Q(n10883), 
        .QN(n2669) );
  DFFR_X1 \REGISTERS_reg[80][1]  ( .D(n8907), .CK(CLK), .RN(n2975), .Q(n10884), 
        .QN(n2670) );
  DFFR_X1 \REGISTERS_reg[80][0]  ( .D(n8908), .CK(CLK), .RN(n2975), .Q(n10885), 
        .QN(n2671) );
  DFFR_X1 \REGISTERS_reg[81][31]  ( .D(n8909), .CK(CLK), .RN(n2975), .Q(n10886), .QN(n2672) );
  DFFR_X1 \REGISTERS_reg[81][30]  ( .D(n8910), .CK(CLK), .RN(n2975), .Q(n10887), .QN(n2673) );
  DFFR_X1 \REGISTERS_reg[81][29]  ( .D(n8911), .CK(CLK), .RN(n2975), .Q(n10888), .QN(n2674) );
  DFFR_X1 \REGISTERS_reg[81][28]  ( .D(n8912), .CK(CLK), .RN(n2975), .Q(n10889), .QN(n2675) );
  DFFR_X1 \REGISTERS_reg[81][27]  ( .D(n8913), .CK(CLK), .RN(n2974), .Q(n10890), .QN(n2676) );
  DFFR_X1 \REGISTERS_reg[81][26]  ( .D(n8914), .CK(CLK), .RN(n2974), .Q(n10891), .QN(n2677) );
  DFFR_X1 \REGISTERS_reg[81][25]  ( .D(n8915), .CK(CLK), .RN(n2974), .Q(n10892), .QN(n2678) );
  DFFR_X1 \REGISTERS_reg[81][24]  ( .D(n8916), .CK(CLK), .RN(n2974), .Q(n10893), .QN(n2679) );
  DFFR_X1 \REGISTERS_reg[81][23]  ( .D(n8917), .CK(CLK), .RN(n2974), .Q(n10894), .QN(n2680) );
  DFFR_X1 \REGISTERS_reg[81][22]  ( .D(n8918), .CK(CLK), .RN(n2974), .Q(n10895), .QN(n2681) );
  DFFR_X1 \REGISTERS_reg[81][21]  ( .D(n8919), .CK(CLK), .RN(n2974), .Q(n10896), .QN(n2682) );
  DFFR_X1 \REGISTERS_reg[81][20]  ( .D(n8920), .CK(CLK), .RN(n2974), .Q(n10897), .QN(n2683) );
  DFFR_X1 \REGISTERS_reg[81][19]  ( .D(n8921), .CK(CLK), .RN(n2974), .Q(n10898), .QN(n2684) );
  DFFR_X1 \REGISTERS_reg[81][18]  ( .D(n8922), .CK(CLK), .RN(n2974), .Q(n10899), .QN(n2685) );
  DFFR_X1 \REGISTERS_reg[81][17]  ( .D(n8923), .CK(CLK), .RN(n2974), .Q(n10900), .QN(n2686) );
  DFFR_X1 \REGISTERS_reg[81][16]  ( .D(n8924), .CK(CLK), .RN(n2974), .Q(n10901), .QN(n2687) );
  DFFR_X1 \REGISTERS_reg[81][15]  ( .D(n8925), .CK(CLK), .RN(n2973), .Q(n10902), .QN(n2688) );
  DFFR_X1 \REGISTERS_reg[81][14]  ( .D(n8926), .CK(CLK), .RN(n2973), .Q(n10903), .QN(n2689) );
  DFFR_X1 \REGISTERS_reg[81][13]  ( .D(n8927), .CK(CLK), .RN(n2973), .Q(n10904), .QN(n2690) );
  DFFR_X1 \REGISTERS_reg[81][12]  ( .D(n8928), .CK(CLK), .RN(n2973), .Q(n10905), .QN(n2691) );
  DFFR_X1 \REGISTERS_reg[81][11]  ( .D(n8929), .CK(CLK), .RN(n2973), .Q(n10906), .QN(n2692) );
  DFFR_X1 \REGISTERS_reg[81][10]  ( .D(n8930), .CK(CLK), .RN(n2973), .Q(n10907), .QN(n2693) );
  DFFR_X1 \REGISTERS_reg[81][9]  ( .D(n8931), .CK(CLK), .RN(n2973), .Q(n10908), 
        .QN(n2694) );
  DFFR_X1 \REGISTERS_reg[81][8]  ( .D(n8932), .CK(CLK), .RN(n2973), .Q(n10909), 
        .QN(n2695) );
  DFFR_X1 \REGISTERS_reg[81][7]  ( .D(n8933), .CK(CLK), .RN(n2973), .Q(n10910), 
        .QN(n2696) );
  DFFR_X1 \REGISTERS_reg[81][6]  ( .D(n8934), .CK(CLK), .RN(n2973), .Q(n10911), 
        .QN(n2697) );
  DFFR_X1 \REGISTERS_reg[81][5]  ( .D(n8935), .CK(CLK), .RN(n2973), .Q(n10912), 
        .QN(n2698) );
  DFFR_X1 \REGISTERS_reg[81][4]  ( .D(n8936), .CK(CLK), .RN(n2973), .Q(n10913), 
        .QN(n2699) );
  DFFR_X1 \REGISTERS_reg[81][3]  ( .D(n8937), .CK(CLK), .RN(n2972), .Q(n10914), 
        .QN(n2700) );
  DFFR_X1 \REGISTERS_reg[81][2]  ( .D(n8938), .CK(CLK), .RN(n2972), .Q(n10915), 
        .QN(n2701) );
  DFFR_X1 \REGISTERS_reg[81][1]  ( .D(n8939), .CK(CLK), .RN(n2972), .Q(n10916), 
        .QN(n2702) );
  DFFR_X1 \REGISTERS_reg[81][0]  ( .D(n8940), .CK(CLK), .RN(n2972), .Q(n10917), 
        .QN(n2703) );
  DLH_X1 \OUT2_reg[31]  ( .G(n1791), .D(N8767), .Q(OUT2[31]) );
  DLH_X1 \OUT1_reg[31]  ( .G(n1794), .D(N8734), .Q(OUT1[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(n1791), .D(N8766), .Q(OUT2[30]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n1794), .D(N8733), .Q(OUT1[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(n1791), .D(N8765), .Q(OUT2[29]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n1794), .D(N8732), .Q(OUT1[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(n1791), .D(N8764), .Q(OUT2[28]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n1794), .D(N8731), .Q(OUT1[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(n1791), .D(N8763), .Q(OUT2[27]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n1794), .D(N8730), .Q(OUT1[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(n1791), .D(N8762), .Q(OUT2[26]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n1794), .D(N8729), .Q(OUT1[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(n1791), .D(N8761), .Q(OUT2[25]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n1794), .D(N8728), .Q(OUT1[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(n1791), .D(N8760), .Q(OUT2[24]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n1794), .D(N8727), .Q(OUT1[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(n1791), .D(N8759), .Q(OUT2[23]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n1794), .D(N8726), .Q(OUT1[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(n1791), .D(N8758), .Q(OUT2[22]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n1794), .D(N8725), .Q(OUT1[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(n1791), .D(N8757), .Q(OUT2[21]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n1794), .D(N8724), .Q(OUT1[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(n1792), .D(N8756), .Q(OUT2[20]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n1795), .D(N8723), .Q(OUT1[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(n1792), .D(N8755), .Q(OUT2[19]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n1795), .D(N8722), .Q(OUT1[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(n1792), .D(N8754), .Q(OUT2[18]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n1795), .D(N8721), .Q(OUT1[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(n1792), .D(N8753), .Q(OUT2[17]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n1795), .D(N8720), .Q(OUT1[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(n1792), .D(N8752), .Q(OUT2[16]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n1795), .D(N8719), .Q(OUT1[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(n1792), .D(N8751), .Q(OUT2[15]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n1795), .D(N8718), .Q(OUT1[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(n1792), .D(N8750), .Q(OUT2[14]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n1795), .D(N8717), .Q(OUT1[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(n1792), .D(N8749), .Q(OUT2[13]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n1795), .D(N8716), .Q(OUT1[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(n1792), .D(N8748), .Q(OUT2[12]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n1795), .D(N8715), .Q(OUT1[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(n1792), .D(N8747), .Q(OUT2[11]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n1795), .D(N8714), .Q(OUT1[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(n1792), .D(N8746), .Q(OUT2[10]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n1795), .D(N8713), .Q(OUT1[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(n1793), .D(N8745), .Q(OUT2[9]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n1796), .D(N8712), .Q(OUT1[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(n1793), .D(N8744), .Q(OUT2[8]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n1796), .D(N8711), .Q(OUT1[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(n1793), .D(N8743), .Q(OUT2[7]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n1796), .D(N8710), .Q(OUT1[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(n1793), .D(N8742), .Q(OUT2[6]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n1796), .D(N8709), .Q(OUT1[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(n1793), .D(N8741), .Q(OUT2[5]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n1796), .D(N8708), .Q(OUT1[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(n1793), .D(N8740), .Q(OUT2[4]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n1796), .D(N8707), .Q(OUT1[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(n1793), .D(N8739), .Q(OUT2[3]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n1796), .D(N8706), .Q(OUT1[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(n1793), .D(N8738), .Q(OUT2[2]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n1796), .D(N8705), .Q(OUT1[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(n1793), .D(N8737), .Q(OUT2[1]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n1796), .D(N8704), .Q(OUT1[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(n1793), .D(N8736), .Q(OUT2[0]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n1796), .D(N8703), .Q(OUT1[0]) );
  windRF_M8_N8_F5_NBIT32_DW01_add_1 add_66_C130 ( .A({CWP[6:4], N8790, N8789, 
        N8788, N8787}), .B({1'b0, 1'b0, ADD_RD2[4:3], N8570, N8569, N8568}), 
        .CI(1'b0), .SUM({N8567, N8566, N8565, N8564, N8563, N8562, N8561}) );
  windRF_M8_N8_F5_NBIT32_DW01_add_3 add_66_C126 ( .A({CWP[6:4], N8790, N8789, 
        N8788, N8787}), .B({1'b0, 1'b0, ADD_RD1[4:3], N8426, N8425, N8424}), 
        .CI(1'b0), .SUM({N8423, N8422, N8421, N8420, N8419, N8418, N8417}) );
  windRF_M8_N8_F5_NBIT32_DW01_add_5 add_66_C91 ( .A({CWP[6:4], N8790, N8789, 
        N8788, N8787}), .B({1'b0, 1'b0, ADD_WR[4:3], N2162, N2161, N2160}), 
        .CI(1'b0), .SUM({N2159, N2158, N2157, N2156, N2155, N2154, N2153}) );
  DFFR_X1 \REGISTERS_reg[87][31]  ( .D(n9101), .CK(CLK), .RN(RESET), .Q(
        \REGISTERS[87][31] ) );
  DFFR_X1 \REGISTERS_reg[87][30]  ( .D(n9102), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[87][30] ) );
  DFFR_X1 \REGISTERS_reg[87][29]  ( .D(n9103), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[87][29] ) );
  DFFR_X1 \REGISTERS_reg[87][28]  ( .D(n9104), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[87][28] ) );
  DFFR_X1 \REGISTERS_reg[87][27]  ( .D(n9105), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][27] ) );
  DFFR_X1 \REGISTERS_reg[87][26]  ( .D(n9106), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][26] ) );
  DFFR_X1 \REGISTERS_reg[87][25]  ( .D(n9107), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][25] ) );
  DFFR_X1 \REGISTERS_reg[87][24]  ( .D(n9108), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][24] ) );
  DFFR_X1 \REGISTERS_reg[87][23]  ( .D(n9109), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][23] ) );
  DFFR_X1 \REGISTERS_reg[87][22]  ( .D(n9110), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][22] ) );
  DFFR_X1 \REGISTERS_reg[87][21]  ( .D(n9111), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][21] ) );
  DFFR_X1 \REGISTERS_reg[87][20]  ( .D(n9112), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][20] ) );
  DFFR_X1 \REGISTERS_reg[87][19]  ( .D(n9113), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][19] ) );
  DFFR_X1 \REGISTERS_reg[87][18]  ( .D(n9114), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][18] ) );
  DFFR_X1 \REGISTERS_reg[87][17]  ( .D(n9115), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][17] ) );
  DFFR_X1 \REGISTERS_reg[87][16]  ( .D(n9116), .CK(CLK), .RN(n2958), .Q(
        \REGISTERS[87][16] ) );
  DFFR_X1 \REGISTERS_reg[87][15]  ( .D(n9117), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][15] ) );
  DFFR_X1 \REGISTERS_reg[87][14]  ( .D(n9118), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][14] ) );
  DFFR_X1 \REGISTERS_reg[87][13]  ( .D(n9119), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][13] ) );
  DFFR_X1 \REGISTERS_reg[87][12]  ( .D(n9120), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][12] ) );
  DFFR_X1 \REGISTERS_reg[87][11]  ( .D(n9121), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][11] ) );
  DFFR_X1 \REGISTERS_reg[87][10]  ( .D(n9122), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][10] ) );
  DFFR_X1 \REGISTERS_reg[87][9]  ( .D(n9123), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][9] ) );
  DFFR_X1 \REGISTERS_reg[87][8]  ( .D(n9124), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][8] ) );
  DFFR_X1 \REGISTERS_reg[87][7]  ( .D(n9125), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][7] ) );
  DFFR_X1 \REGISTERS_reg[87][6]  ( .D(n9126), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][6] ) );
  DFFR_X1 \REGISTERS_reg[87][5]  ( .D(n9127), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][5] ) );
  DFFR_X1 \REGISTERS_reg[87][4]  ( .D(n9128), .CK(CLK), .RN(n2957), .Q(
        \REGISTERS[87][4] ) );
  DFFR_X1 \REGISTERS_reg[87][3]  ( .D(n9129), .CK(CLK), .RN(n2956), .Q(
        \REGISTERS[87][3] ) );
  DFFR_X1 \REGISTERS_reg[87][2]  ( .D(n9130), .CK(CLK), .RN(n2956), .Q(
        \REGISTERS[87][2] ) );
  DFFR_X1 \REGISTERS_reg[87][1]  ( .D(n9131), .CK(CLK), .RN(n2956), .Q(
        \REGISTERS[87][1] ) );
  DFFR_X1 \REGISTERS_reg[87][0]  ( .D(n9132), .CK(CLK), .RN(n2956), .Q(
        \REGISTERS[87][0] ) );
  DFFR_X1 \REGISTERS_reg[86][31]  ( .D(n9069), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][31] ) );
  DFFR_X1 \REGISTERS_reg[86][30]  ( .D(n9070), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][30] ) );
  DFFR_X1 \REGISTERS_reg[86][29]  ( .D(n9071), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][29] ) );
  DFFR_X1 \REGISTERS_reg[86][28]  ( .D(n9072), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][28] ) );
  DFFR_X1 \REGISTERS_reg[86][27]  ( .D(n9073), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][27] ) );
  DFFR_X1 \REGISTERS_reg[86][26]  ( .D(n9074), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][26] ) );
  DFFR_X1 \REGISTERS_reg[86][25]  ( .D(n9075), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][25] ) );
  DFFR_X1 \REGISTERS_reg[86][24]  ( .D(n9076), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][24] ) );
  DFFR_X1 \REGISTERS_reg[86][23]  ( .D(n9077), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][23] ) );
  DFFR_X1 \REGISTERS_reg[86][22]  ( .D(n9078), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][22] ) );
  DFFR_X1 \REGISTERS_reg[86][21]  ( .D(n9079), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][21] ) );
  DFFR_X1 \REGISTERS_reg[86][20]  ( .D(n9080), .CK(CLK), .RN(n2961), .Q(
        \REGISTERS[86][20] ) );
  DFFR_X1 \REGISTERS_reg[86][19]  ( .D(n9081), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][19] ) );
  DFFR_X1 \REGISTERS_reg[86][18]  ( .D(n9082), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][18] ) );
  DFFR_X1 \REGISTERS_reg[86][17]  ( .D(n9083), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][17] ) );
  DFFR_X1 \REGISTERS_reg[86][16]  ( .D(n9084), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][16] ) );
  DFFR_X1 \REGISTERS_reg[86][15]  ( .D(n9085), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][15] ) );
  DFFR_X1 \REGISTERS_reg[86][14]  ( .D(n9086), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][14] ) );
  DFFR_X1 \REGISTERS_reg[86][13]  ( .D(n9087), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][13] ) );
  DFFR_X1 \REGISTERS_reg[86][12]  ( .D(n9088), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][12] ) );
  DFFR_X1 \REGISTERS_reg[86][11]  ( .D(n9089), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][11] ) );
  DFFR_X1 \REGISTERS_reg[86][10]  ( .D(n9090), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][10] ) );
  DFFR_X1 \REGISTERS_reg[86][9]  ( .D(n9091), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][9] ) );
  DFFR_X1 \REGISTERS_reg[86][8]  ( .D(n9092), .CK(CLK), .RN(n2960), .Q(
        \REGISTERS[86][8] ) );
  DFFR_X1 \REGISTERS_reg[86][7]  ( .D(n9093), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[86][7] ) );
  DFFR_X1 \REGISTERS_reg[86][6]  ( .D(n9094), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[86][6] ) );
  DFFR_X1 \REGISTERS_reg[86][5]  ( .D(n9095), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[86][5] ) );
  DFFR_X1 \REGISTERS_reg[86][4]  ( .D(n9096), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[86][4] ) );
  DFFR_X1 \REGISTERS_reg[86][3]  ( .D(n9097), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[86][3] ) );
  DFFR_X1 \REGISTERS_reg[86][2]  ( .D(n9098), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[86][2] ) );
  DFFR_X1 \REGISTERS_reg[86][1]  ( .D(n9099), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[86][1] ) );
  DFFR_X1 \REGISTERS_reg[86][0]  ( .D(n9100), .CK(CLK), .RN(n2959), .Q(
        \REGISTERS[86][0] ) );
  DFFR_X1 \REGISTERS_reg[85][31]  ( .D(n9037), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[85][31] ) );
  DFFR_X1 \REGISTERS_reg[85][30]  ( .D(n9038), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[85][30] ) );
  DFFR_X1 \REGISTERS_reg[85][29]  ( .D(n9039), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[85][29] ) );
  DFFR_X1 \REGISTERS_reg[85][28]  ( .D(n9040), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[85][28] ) );
  DFFR_X1 \REGISTERS_reg[85][27]  ( .D(n9041), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[85][27] ) );
  DFFR_X1 \REGISTERS_reg[85][26]  ( .D(n9042), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[85][26] ) );
  DFFR_X1 \REGISTERS_reg[85][25]  ( .D(n9043), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[85][25] ) );
  DFFR_X1 \REGISTERS_reg[85][24]  ( .D(n9044), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[85][24] ) );
  DFFR_X1 \REGISTERS_reg[85][23]  ( .D(n9045), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][23] ) );
  DFFR_X1 \REGISTERS_reg[85][22]  ( .D(n9046), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][22] ) );
  DFFR_X1 \REGISTERS_reg[85][21]  ( .D(n9047), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][21] ) );
  DFFR_X1 \REGISTERS_reg[85][20]  ( .D(n9048), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][20] ) );
  DFFR_X1 \REGISTERS_reg[85][19]  ( .D(n9049), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][19] ) );
  DFFR_X1 \REGISTERS_reg[85][18]  ( .D(n9050), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][18] ) );
  DFFR_X1 \REGISTERS_reg[85][17]  ( .D(n9051), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][17] ) );
  DFFR_X1 \REGISTERS_reg[85][16]  ( .D(n9052), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][16] ) );
  DFFR_X1 \REGISTERS_reg[85][15]  ( .D(n9053), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][15] ) );
  DFFR_X1 \REGISTERS_reg[85][14]  ( .D(n9054), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][14] ) );
  DFFR_X1 \REGISTERS_reg[85][13]  ( .D(n9055), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][13] ) );
  DFFR_X1 \REGISTERS_reg[85][12]  ( .D(n9056), .CK(CLK), .RN(n2963), .Q(
        \REGISTERS[85][12] ) );
  DFFR_X1 \REGISTERS_reg[85][11]  ( .D(n9057), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][11] ) );
  DFFR_X1 \REGISTERS_reg[85][10]  ( .D(n9058), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][10] ) );
  DFFR_X1 \REGISTERS_reg[85][9]  ( .D(n9059), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][9] ) );
  DFFR_X1 \REGISTERS_reg[85][8]  ( .D(n9060), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][8] ) );
  DFFR_X1 \REGISTERS_reg[85][7]  ( .D(n9061), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][7] ) );
  DFFR_X1 \REGISTERS_reg[85][6]  ( .D(n9062), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][6] ) );
  DFFR_X1 \REGISTERS_reg[85][5]  ( .D(n9063), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][5] ) );
  DFFR_X1 \REGISTERS_reg[85][4]  ( .D(n9064), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][4] ) );
  DFFR_X1 \REGISTERS_reg[85][3]  ( .D(n9065), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][3] ) );
  DFFR_X1 \REGISTERS_reg[85][2]  ( .D(n9066), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][2] ) );
  DFFR_X1 \REGISTERS_reg[85][1]  ( .D(n9067), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][1] ) );
  DFFR_X1 \REGISTERS_reg[85][0]  ( .D(n9068), .CK(CLK), .RN(n2962), .Q(
        \REGISTERS[85][0] ) );
  DFFR_X1 \REGISTERS_reg[84][31]  ( .D(n9005), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[84][31] ) );
  DFFR_X1 \REGISTERS_reg[84][30]  ( .D(n9006), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[84][30] ) );
  DFFR_X1 \REGISTERS_reg[84][29]  ( .D(n9007), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[84][29] ) );
  DFFR_X1 \REGISTERS_reg[84][28]  ( .D(n9008), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[84][28] ) );
  DFFR_X1 \REGISTERS_reg[84][27]  ( .D(n9009), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][27] ) );
  DFFR_X1 \REGISTERS_reg[84][26]  ( .D(n9010), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][26] ) );
  DFFR_X1 \REGISTERS_reg[84][25]  ( .D(n9011), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][25] ) );
  DFFR_X1 \REGISTERS_reg[84][24]  ( .D(n9012), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][24] ) );
  DFFR_X1 \REGISTERS_reg[84][23]  ( .D(n9013), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][23] ) );
  DFFR_X1 \REGISTERS_reg[84][22]  ( .D(n9014), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][22] ) );
  DFFR_X1 \REGISTERS_reg[84][21]  ( .D(n9015), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][21] ) );
  DFFR_X1 \REGISTERS_reg[84][20]  ( .D(n9016), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][20] ) );
  DFFR_X1 \REGISTERS_reg[84][19]  ( .D(n9017), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][19] ) );
  DFFR_X1 \REGISTERS_reg[84][18]  ( .D(n9018), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][18] ) );
  DFFR_X1 \REGISTERS_reg[84][17]  ( .D(n9019), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][17] ) );
  DFFR_X1 \REGISTERS_reg[84][16]  ( .D(n9020), .CK(CLK), .RN(n2966), .Q(
        \REGISTERS[84][16] ) );
  DFFR_X1 \REGISTERS_reg[84][15]  ( .D(n9021), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][15] ) );
  DFFR_X1 \REGISTERS_reg[84][14]  ( .D(n9022), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][14] ) );
  DFFR_X1 \REGISTERS_reg[84][13]  ( .D(n9023), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][13] ) );
  DFFR_X1 \REGISTERS_reg[84][12]  ( .D(n9024), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][12] ) );
  DFFR_X1 \REGISTERS_reg[84][11]  ( .D(n9025), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][11] ) );
  DFFR_X1 \REGISTERS_reg[84][10]  ( .D(n9026), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][10] ) );
  DFFR_X1 \REGISTERS_reg[84][9]  ( .D(n9027), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][9] ) );
  DFFR_X1 \REGISTERS_reg[84][8]  ( .D(n9028), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][8] ) );
  DFFR_X1 \REGISTERS_reg[84][7]  ( .D(n9029), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][7] ) );
  DFFR_X1 \REGISTERS_reg[84][6]  ( .D(n9030), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][6] ) );
  DFFR_X1 \REGISTERS_reg[84][5]  ( .D(n9031), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][5] ) );
  DFFR_X1 \REGISTERS_reg[84][4]  ( .D(n9032), .CK(CLK), .RN(n2965), .Q(
        \REGISTERS[84][4] ) );
  DFFR_X1 \REGISTERS_reg[84][3]  ( .D(n9033), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[84][3] ) );
  DFFR_X1 \REGISTERS_reg[84][2]  ( .D(n9034), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[84][2] ) );
  DFFR_X1 \REGISTERS_reg[84][1]  ( .D(n9035), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[84][1] ) );
  DFFR_X1 \REGISTERS_reg[84][0]  ( .D(n9036), .CK(CLK), .RN(n2964), .Q(
        \REGISTERS[84][0] ) );
  DFFR_X1 \REGISTERS_reg[83][31]  ( .D(n8973), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][31] ) );
  DFFR_X1 \REGISTERS_reg[83][30]  ( .D(n8974), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][30] ) );
  DFFR_X1 \REGISTERS_reg[83][29]  ( .D(n8975), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][29] ) );
  DFFR_X1 \REGISTERS_reg[83][28]  ( .D(n8976), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][28] ) );
  DFFR_X1 \REGISTERS_reg[83][27]  ( .D(n8977), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][27] ) );
  DFFR_X1 \REGISTERS_reg[83][26]  ( .D(n8978), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][26] ) );
  DFFR_X1 \REGISTERS_reg[83][25]  ( .D(n8979), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][25] ) );
  DFFR_X1 \REGISTERS_reg[83][24]  ( .D(n8980), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][24] ) );
  DFFR_X1 \REGISTERS_reg[83][23]  ( .D(n8981), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][23] ) );
  DFFR_X1 \REGISTERS_reg[83][22]  ( .D(n8982), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][22] ) );
  DFFR_X1 \REGISTERS_reg[83][21]  ( .D(n8983), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][21] ) );
  DFFR_X1 \REGISTERS_reg[83][20]  ( .D(n8984), .CK(CLK), .RN(n2969), .Q(
        \REGISTERS[83][20] ) );
  DFFR_X1 \REGISTERS_reg[83][19]  ( .D(n8985), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][19] ) );
  DFFR_X1 \REGISTERS_reg[83][18]  ( .D(n8986), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][18] ) );
  DFFR_X1 \REGISTERS_reg[83][17]  ( .D(n8987), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][17] ) );
  DFFR_X1 \REGISTERS_reg[83][16]  ( .D(n8988), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][16] ) );
  DFFR_X1 \REGISTERS_reg[83][15]  ( .D(n8989), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][15] ) );
  DFFR_X1 \REGISTERS_reg[83][14]  ( .D(n8990), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][14] ) );
  DFFR_X1 \REGISTERS_reg[83][13]  ( .D(n8991), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][13] ) );
  DFFR_X1 \REGISTERS_reg[83][12]  ( .D(n8992), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][12] ) );
  DFFR_X1 \REGISTERS_reg[83][11]  ( .D(n8993), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][11] ) );
  DFFR_X1 \REGISTERS_reg[83][10]  ( .D(n8994), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][10] ) );
  DFFR_X1 \REGISTERS_reg[83][9]  ( .D(n8995), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][9] ) );
  DFFR_X1 \REGISTERS_reg[83][8]  ( .D(n8996), .CK(CLK), .RN(n2968), .Q(
        \REGISTERS[83][8] ) );
  DFFR_X1 \REGISTERS_reg[83][7]  ( .D(n8997), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[83][7] ) );
  DFFR_X1 \REGISTERS_reg[83][6]  ( .D(n8998), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[83][6] ) );
  DFFR_X1 \REGISTERS_reg[83][5]  ( .D(n8999), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[83][5] ) );
  DFFR_X1 \REGISTERS_reg[83][4]  ( .D(n9000), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[83][4] ) );
  DFFR_X1 \REGISTERS_reg[83][3]  ( .D(n9001), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[83][3] ) );
  DFFR_X1 \REGISTERS_reg[83][2]  ( .D(n9002), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[83][2] ) );
  DFFR_X1 \REGISTERS_reg[83][1]  ( .D(n9003), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[83][1] ) );
  DFFR_X1 \REGISTERS_reg[83][0]  ( .D(n9004), .CK(CLK), .RN(n2967), .Q(
        \REGISTERS[83][0] ) );
  DFFR_X1 \REGISTERS_reg[82][31]  ( .D(n8941), .CK(CLK), .RN(n2972), .Q(
        \REGISTERS[82][31] ) );
  DFFR_X1 \REGISTERS_reg[82][30]  ( .D(n8942), .CK(CLK), .RN(n2972), .Q(
        \REGISTERS[82][30] ) );
  DFFR_X1 \REGISTERS_reg[82][29]  ( .D(n8943), .CK(CLK), .RN(n2972), .Q(
        \REGISTERS[82][29] ) );
  DFFR_X1 \REGISTERS_reg[82][28]  ( .D(n8944), .CK(CLK), .RN(n2972), .Q(
        \REGISTERS[82][28] ) );
  DFFR_X1 \REGISTERS_reg[82][27]  ( .D(n8945), .CK(CLK), .RN(n2972), .Q(
        \REGISTERS[82][27] ) );
  DFFR_X1 \REGISTERS_reg[82][26]  ( .D(n8946), .CK(CLK), .RN(n2972), .Q(
        \REGISTERS[82][26] ) );
  DFFR_X1 \REGISTERS_reg[82][25]  ( .D(n8947), .CK(CLK), .RN(n2972), .Q(
        \REGISTERS[82][25] ) );
  DFFR_X1 \REGISTERS_reg[82][24]  ( .D(n8948), .CK(CLK), .RN(n2972), .Q(
        \REGISTERS[82][24] ) );
  DFFR_X1 \REGISTERS_reg[82][23]  ( .D(n8949), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][23] ) );
  DFFR_X1 \REGISTERS_reg[82][22]  ( .D(n8950), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][22] ) );
  DFFR_X1 \REGISTERS_reg[82][21]  ( .D(n8951), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][21] ) );
  DFFR_X1 \REGISTERS_reg[82][20]  ( .D(n8952), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][20] ) );
  DFFR_X1 \REGISTERS_reg[82][19]  ( .D(n8953), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][19] ) );
  DFFR_X1 \REGISTERS_reg[82][18]  ( .D(n8954), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][18] ) );
  DFFR_X1 \REGISTERS_reg[82][17]  ( .D(n8955), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][17] ) );
  DFFR_X1 \REGISTERS_reg[82][16]  ( .D(n8956), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][16] ) );
  DFFR_X1 \REGISTERS_reg[82][15]  ( .D(n8957), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][15] ) );
  DFFR_X1 \REGISTERS_reg[82][14]  ( .D(n8958), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][14] ) );
  DFFR_X1 \REGISTERS_reg[82][13]  ( .D(n8959), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][13] ) );
  DFFR_X1 \REGISTERS_reg[82][12]  ( .D(n8960), .CK(CLK), .RN(n2971), .Q(
        \REGISTERS[82][12] ) );
  DFFR_X1 \REGISTERS_reg[82][11]  ( .D(n8961), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][11] ) );
  DFFR_X1 \REGISTERS_reg[82][10]  ( .D(n8962), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][10] ) );
  DFFR_X1 \REGISTERS_reg[82][9]  ( .D(n8963), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][9] ) );
  DFFR_X1 \REGISTERS_reg[82][8]  ( .D(n8964), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][8] ) );
  DFFR_X1 \REGISTERS_reg[82][7]  ( .D(n8965), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][7] ) );
  DFFR_X1 \REGISTERS_reg[82][6]  ( .D(n8966), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][6] ) );
  DFFR_X1 \REGISTERS_reg[82][5]  ( .D(n8967), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][5] ) );
  DFFR_X1 \REGISTERS_reg[82][4]  ( .D(n8968), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][4] ) );
  DFFR_X1 \REGISTERS_reg[82][3]  ( .D(n8969), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][3] ) );
  DFFR_X1 \REGISTERS_reg[82][2]  ( .D(n8970), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][2] ) );
  DFFR_X1 \REGISTERS_reg[82][1]  ( .D(n8971), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][1] ) );
  DFFR_X1 \REGISTERS_reg[82][0]  ( .D(n8972), .CK(CLK), .RN(n2970), .Q(
        \REGISTERS[82][0] ) );
  DFFR_X1 \REGISTERS_reg[78][31]  ( .D(n8813), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[78][31] ) );
  DFFR_X1 \REGISTERS_reg[78][30]  ( .D(n8814), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[78][30] ) );
  DFFR_X1 \REGISTERS_reg[78][29]  ( .D(n8815), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[78][29] ) );
  DFFR_X1 \REGISTERS_reg[78][28]  ( .D(n8816), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[78][28] ) );
  DFFR_X1 \REGISTERS_reg[78][27]  ( .D(n8817), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][27] ) );
  DFFR_X1 \REGISTERS_reg[78][26]  ( .D(n8818), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][26] ) );
  DFFR_X1 \REGISTERS_reg[78][25]  ( .D(n8819), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][25] ) );
  DFFR_X1 \REGISTERS_reg[78][24]  ( .D(n8820), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][24] ) );
  DFFR_X1 \REGISTERS_reg[78][23]  ( .D(n8821), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][23] ) );
  DFFR_X1 \REGISTERS_reg[78][22]  ( .D(n8822), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][22] ) );
  DFFR_X1 \REGISTERS_reg[78][21]  ( .D(n8823), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][21] ) );
  DFFR_X1 \REGISTERS_reg[78][20]  ( .D(n8824), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][20] ) );
  DFFR_X1 \REGISTERS_reg[78][19]  ( .D(n8825), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][19] ) );
  DFFR_X1 \REGISTERS_reg[78][18]  ( .D(n8826), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][18] ) );
  DFFR_X1 \REGISTERS_reg[78][17]  ( .D(n8827), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][17] ) );
  DFFR_X1 \REGISTERS_reg[78][16]  ( .D(n8828), .CK(CLK), .RN(n2982), .Q(
        \REGISTERS[78][16] ) );
  DFFR_X1 \REGISTERS_reg[78][15]  ( .D(n8829), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][15] ) );
  DFFR_X1 \REGISTERS_reg[78][14]  ( .D(n8830), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][14] ) );
  DFFR_X1 \REGISTERS_reg[78][13]  ( .D(n8831), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][13] ) );
  DFFR_X1 \REGISTERS_reg[78][12]  ( .D(n8832), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][12] ) );
  DFFR_X1 \REGISTERS_reg[78][11]  ( .D(n8833), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][11] ) );
  DFFR_X1 \REGISTERS_reg[78][10]  ( .D(n8834), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][10] ) );
  DFFR_X1 \REGISTERS_reg[78][9]  ( .D(n8835), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][9] ) );
  DFFR_X1 \REGISTERS_reg[78][8]  ( .D(n8836), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][8] ) );
  DFFR_X1 \REGISTERS_reg[78][7]  ( .D(n8837), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][7] ) );
  DFFR_X1 \REGISTERS_reg[78][6]  ( .D(n8838), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][6] ) );
  DFFR_X1 \REGISTERS_reg[78][5]  ( .D(n8839), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][5] ) );
  DFFR_X1 \REGISTERS_reg[78][4]  ( .D(n8840), .CK(CLK), .RN(n2981), .Q(
        \REGISTERS[78][4] ) );
  DFFR_X1 \REGISTERS_reg[78][3]  ( .D(n8841), .CK(CLK), .RN(n2980), .Q(
        \REGISTERS[78][3] ) );
  DFFR_X1 \REGISTERS_reg[78][2]  ( .D(n8842), .CK(CLK), .RN(n2980), .Q(
        \REGISTERS[78][2] ) );
  DFFR_X1 \REGISTERS_reg[78][1]  ( .D(n8843), .CK(CLK), .RN(n2980), .Q(
        \REGISTERS[78][1] ) );
  DFFR_X1 \REGISTERS_reg[78][0]  ( .D(n8844), .CK(CLK), .RN(n2980), .Q(
        \REGISTERS[78][0] ) );
  DFFR_X1 \REGISTERS_reg[77][31]  ( .D(n8781), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][31] ) );
  DFFR_X1 \REGISTERS_reg[77][30]  ( .D(n8782), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][30] ) );
  DFFR_X1 \REGISTERS_reg[77][29]  ( .D(n8783), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][29] ) );
  DFFR_X1 \REGISTERS_reg[77][28]  ( .D(n8784), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][28] ) );
  DFFR_X1 \REGISTERS_reg[77][27]  ( .D(n8785), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][27] ) );
  DFFR_X1 \REGISTERS_reg[77][26]  ( .D(n8786), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][26] ) );
  DFFR_X1 \REGISTERS_reg[77][25]  ( .D(n8787), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][25] ) );
  DFFR_X1 \REGISTERS_reg[77][24]  ( .D(n8788), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][24] ) );
  DFFR_X1 \REGISTERS_reg[77][23]  ( .D(n8789), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][23] ) );
  DFFR_X1 \REGISTERS_reg[77][22]  ( .D(n8790), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][22] ) );
  DFFR_X1 \REGISTERS_reg[77][21]  ( .D(n8791), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][21] ) );
  DFFR_X1 \REGISTERS_reg[77][20]  ( .D(n8792), .CK(CLK), .RN(n2985), .Q(
        \REGISTERS[77][20] ) );
  DFFR_X1 \REGISTERS_reg[77][19]  ( .D(n8793), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][19] ) );
  DFFR_X1 \REGISTERS_reg[77][18]  ( .D(n8794), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][18] ) );
  DFFR_X1 \REGISTERS_reg[77][17]  ( .D(n8795), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][17] ) );
  DFFR_X1 \REGISTERS_reg[77][16]  ( .D(n8796), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][16] ) );
  DFFR_X1 \REGISTERS_reg[77][15]  ( .D(n8797), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][15] ) );
  DFFR_X1 \REGISTERS_reg[77][14]  ( .D(n8798), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][14] ) );
  DFFR_X1 \REGISTERS_reg[77][13]  ( .D(n8799), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][13] ) );
  DFFR_X1 \REGISTERS_reg[77][12]  ( .D(n8800), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][12] ) );
  DFFR_X1 \REGISTERS_reg[77][11]  ( .D(n8801), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][11] ) );
  DFFR_X1 \REGISTERS_reg[77][10]  ( .D(n8802), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][10] ) );
  DFFR_X1 \REGISTERS_reg[77][9]  ( .D(n8803), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][9] ) );
  DFFR_X1 \REGISTERS_reg[77][8]  ( .D(n8804), .CK(CLK), .RN(n2984), .Q(
        \REGISTERS[77][8] ) );
  DFFR_X1 \REGISTERS_reg[77][7]  ( .D(n8805), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[77][7] ) );
  DFFR_X1 \REGISTERS_reg[77][6]  ( .D(n8806), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[77][6] ) );
  DFFR_X1 \REGISTERS_reg[77][5]  ( .D(n8807), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[77][5] ) );
  DFFR_X1 \REGISTERS_reg[77][4]  ( .D(n8808), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[77][4] ) );
  DFFR_X1 \REGISTERS_reg[77][3]  ( .D(n8809), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[77][3] ) );
  DFFR_X1 \REGISTERS_reg[77][2]  ( .D(n8810), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[77][2] ) );
  DFFR_X1 \REGISTERS_reg[77][1]  ( .D(n8811), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[77][1] ) );
  DFFR_X1 \REGISTERS_reg[77][0]  ( .D(n8812), .CK(CLK), .RN(n2983), .Q(
        \REGISTERS[77][0] ) );
  DFFR_X1 \REGISTERS_reg[54][31]  ( .D(n8045), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[54][31] ) );
  DFFR_X1 \REGISTERS_reg[54][30]  ( .D(n8046), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[54][30] ) );
  DFFR_X1 \REGISTERS_reg[54][29]  ( .D(n8047), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[54][29] ) );
  DFFR_X1 \REGISTERS_reg[54][28]  ( .D(n8048), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[54][28] ) );
  DFFR_X1 \REGISTERS_reg[54][27]  ( .D(n8049), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][27] ) );
  DFFR_X1 \REGISTERS_reg[54][26]  ( .D(n8050), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][26] ) );
  DFFR_X1 \REGISTERS_reg[54][25]  ( .D(n8051), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][25] ) );
  DFFR_X1 \REGISTERS_reg[54][24]  ( .D(n8052), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][24] ) );
  DFFR_X1 \REGISTERS_reg[54][23]  ( .D(n8053), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][23] ) );
  DFFR_X1 \REGISTERS_reg[54][22]  ( .D(n8054), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][22] ) );
  DFFR_X1 \REGISTERS_reg[54][21]  ( .D(n8055), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][21] ) );
  DFFR_X1 \REGISTERS_reg[54][20]  ( .D(n8056), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][20] ) );
  DFFR_X1 \REGISTERS_reg[54][19]  ( .D(n8057), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][19] ) );
  DFFR_X1 \REGISTERS_reg[54][18]  ( .D(n8058), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][18] ) );
  DFFR_X1 \REGISTERS_reg[54][17]  ( .D(n8059), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][17] ) );
  DFFR_X1 \REGISTERS_reg[54][16]  ( .D(n8060), .CK(CLK), .RN(n3059), .Q(
        \REGISTERS[54][16] ) );
  DFFR_X1 \REGISTERS_reg[54][15]  ( .D(n8061), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][15] ) );
  DFFR_X1 \REGISTERS_reg[54][14]  ( .D(n8062), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][14] ) );
  DFFR_X1 \REGISTERS_reg[54][13]  ( .D(n8063), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][13] ) );
  DFFR_X1 \REGISTERS_reg[54][12]  ( .D(n8064), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][12] ) );
  DFFR_X1 \REGISTERS_reg[54][11]  ( .D(n8065), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][11] ) );
  DFFR_X1 \REGISTERS_reg[54][10]  ( .D(n8066), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][10] ) );
  DFFR_X1 \REGISTERS_reg[54][9]  ( .D(n8067), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][9] ) );
  DFFR_X1 \REGISTERS_reg[54][8]  ( .D(n8068), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][8] ) );
  DFFR_X1 \REGISTERS_reg[54][7]  ( .D(n8069), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][7] ) );
  DFFR_X1 \REGISTERS_reg[54][6]  ( .D(n8070), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][6] ) );
  DFFR_X1 \REGISTERS_reg[54][5]  ( .D(n8071), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][5] ) );
  DFFR_X1 \REGISTERS_reg[54][4]  ( .D(n8072), .CK(CLK), .RN(n3057), .Q(
        \REGISTERS[54][4] ) );
  DFFR_X1 \REGISTERS_reg[54][3]  ( .D(n8073), .CK(CLK), .RN(n3056), .Q(
        \REGISTERS[54][3] ) );
  DFFR_X1 \REGISTERS_reg[54][2]  ( .D(n8074), .CK(CLK), .RN(n3056), .Q(
        \REGISTERS[54][2] ) );
  DFFR_X1 \REGISTERS_reg[54][1]  ( .D(n8075), .CK(CLK), .RN(n3056), .Q(
        \REGISTERS[54][1] ) );
  DFFR_X1 \REGISTERS_reg[54][0]  ( .D(n8076), .CK(CLK), .RN(n3056), .Q(
        \REGISTERS[54][0] ) );
  DFFR_X1 \REGISTERS_reg[53][31]  ( .D(n8013), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][31] ) );
  DFFR_X1 \REGISTERS_reg[53][30]  ( .D(n8014), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][30] ) );
  DFFR_X1 \REGISTERS_reg[53][29]  ( .D(n8015), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][29] ) );
  DFFR_X1 \REGISTERS_reg[53][28]  ( .D(n8016), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][28] ) );
  DFFR_X1 \REGISTERS_reg[53][27]  ( .D(n8017), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][27] ) );
  DFFR_X1 \REGISTERS_reg[53][26]  ( .D(n8018), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][26] ) );
  DFFR_X1 \REGISTERS_reg[53][25]  ( .D(n8019), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][25] ) );
  DFFR_X1 \REGISTERS_reg[53][24]  ( .D(n8020), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][24] ) );
  DFFR_X1 \REGISTERS_reg[53][23]  ( .D(n8021), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][23] ) );
  DFFR_X1 \REGISTERS_reg[53][22]  ( .D(n8022), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][22] ) );
  DFFR_X1 \REGISTERS_reg[53][21]  ( .D(n8023), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][21] ) );
  DFFR_X1 \REGISTERS_reg[53][20]  ( .D(n8024), .CK(CLK), .RN(n3064), .Q(
        \REGISTERS[53][20] ) );
  DFFR_X1 \REGISTERS_reg[53][19]  ( .D(n8025), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][19] ) );
  DFFR_X1 \REGISTERS_reg[53][18]  ( .D(n8026), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][18] ) );
  DFFR_X1 \REGISTERS_reg[53][17]  ( .D(n8027), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][17] ) );
  DFFR_X1 \REGISTERS_reg[53][16]  ( .D(n8028), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][16] ) );
  DFFR_X1 \REGISTERS_reg[53][15]  ( .D(n8029), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][15] ) );
  DFFR_X1 \REGISTERS_reg[53][14]  ( .D(n8030), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][14] ) );
  DFFR_X1 \REGISTERS_reg[53][13]  ( .D(n8031), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][13] ) );
  DFFR_X1 \REGISTERS_reg[53][12]  ( .D(n8032), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][12] ) );
  DFFR_X1 \REGISTERS_reg[53][11]  ( .D(n8033), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][11] ) );
  DFFR_X1 \REGISTERS_reg[53][10]  ( .D(n8034), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][10] ) );
  DFFR_X1 \REGISTERS_reg[53][9]  ( .D(n8035), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][9] ) );
  DFFR_X1 \REGISTERS_reg[53][8]  ( .D(n8036), .CK(CLK), .RN(n3062), .Q(
        \REGISTERS[53][8] ) );
  DFFR_X1 \REGISTERS_reg[53][7]  ( .D(n8037), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[53][7] ) );
  DFFR_X1 \REGISTERS_reg[53][6]  ( .D(n8038), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[53][6] ) );
  DFFR_X1 \REGISTERS_reg[53][5]  ( .D(n8039), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[53][5] ) );
  DFFR_X1 \REGISTERS_reg[53][4]  ( .D(n8040), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[53][4] ) );
  DFFR_X1 \REGISTERS_reg[53][3]  ( .D(n8041), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[53][3] ) );
  DFFR_X1 \REGISTERS_reg[53][2]  ( .D(n8042), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[53][2] ) );
  DFFR_X1 \REGISTERS_reg[53][1]  ( .D(n8043), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[53][1] ) );
  DFFR_X1 \REGISTERS_reg[53][0]  ( .D(n8044), .CK(CLK), .RN(n3061), .Q(
        \REGISTERS[53][0] ) );
  DFFR_X1 \REGISTERS_reg[52][31]  ( .D(n7981), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[52][31] ) );
  DFFR_X1 \REGISTERS_reg[52][30]  ( .D(n7982), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[52][30] ) );
  DFFR_X1 \REGISTERS_reg[52][29]  ( .D(n7983), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[52][29] ) );
  DFFR_X1 \REGISTERS_reg[52][28]  ( .D(n7984), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[52][28] ) );
  DFFR_X1 \REGISTERS_reg[52][27]  ( .D(n7985), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[52][27] ) );
  DFFR_X1 \REGISTERS_reg[52][26]  ( .D(n7986), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[52][26] ) );
  DFFR_X1 \REGISTERS_reg[52][25]  ( .D(n7987), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[52][25] ) );
  DFFR_X1 \REGISTERS_reg[52][24]  ( .D(n7988), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[52][24] ) );
  DFFR_X1 \REGISTERS_reg[52][23]  ( .D(n7989), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][23] ) );
  DFFR_X1 \REGISTERS_reg[52][22]  ( .D(n7990), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][22] ) );
  DFFR_X1 \REGISTERS_reg[52][21]  ( .D(n7991), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][21] ) );
  DFFR_X1 \REGISTERS_reg[52][20]  ( .D(n7992), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][20] ) );
  DFFR_X1 \REGISTERS_reg[52][19]  ( .D(n7993), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][19] ) );
  DFFR_X1 \REGISTERS_reg[52][18]  ( .D(n7994), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][18] ) );
  DFFR_X1 \REGISTERS_reg[52][17]  ( .D(n7995), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][17] ) );
  DFFR_X1 \REGISTERS_reg[52][16]  ( .D(n7996), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][16] ) );
  DFFR_X1 \REGISTERS_reg[52][15]  ( .D(n7997), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][15] ) );
  DFFR_X1 \REGISTERS_reg[52][14]  ( .D(n7998), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][14] ) );
  DFFR_X1 \REGISTERS_reg[52][13]  ( .D(n7999), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][13] ) );
  DFFR_X1 \REGISTERS_reg[52][12]  ( .D(n8000), .CK(CLK), .RN(n3067), .Q(
        \REGISTERS[52][12] ) );
  DFFR_X1 \REGISTERS_reg[52][11]  ( .D(n8001), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][11] ) );
  DFFR_X1 \REGISTERS_reg[52][10]  ( .D(n8002), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][10] ) );
  DFFR_X1 \REGISTERS_reg[52][9]  ( .D(n8003), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][9] ) );
  DFFR_X1 \REGISTERS_reg[52][8]  ( .D(n8004), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][8] ) );
  DFFR_X1 \REGISTERS_reg[52][7]  ( .D(n8005), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][7] ) );
  DFFR_X1 \REGISTERS_reg[52][6]  ( .D(n8006), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][6] ) );
  DFFR_X1 \REGISTERS_reg[52][5]  ( .D(n8007), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][5] ) );
  DFFR_X1 \REGISTERS_reg[52][4]  ( .D(n8008), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][4] ) );
  DFFR_X1 \REGISTERS_reg[52][3]  ( .D(n8009), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][3] ) );
  DFFR_X1 \REGISTERS_reg[52][2]  ( .D(n8010), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][2] ) );
  DFFR_X1 \REGISTERS_reg[52][1]  ( .D(n8011), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][1] ) );
  DFFR_X1 \REGISTERS_reg[52][0]  ( .D(n8012), .CK(CLK), .RN(n3066), .Q(
        \REGISTERS[52][0] ) );
  DFFR_X1 \REGISTERS_reg[51][31]  ( .D(n7949), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[51][31] ) );
  DFFR_X1 \REGISTERS_reg[51][30]  ( .D(n7950), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[51][30] ) );
  DFFR_X1 \REGISTERS_reg[51][29]  ( .D(n7951), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[51][29] ) );
  DFFR_X1 \REGISTERS_reg[51][28]  ( .D(n7952), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[51][28] ) );
  DFFR_X1 \REGISTERS_reg[51][27]  ( .D(n7953), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][27] ) );
  DFFR_X1 \REGISTERS_reg[51][26]  ( .D(n7954), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][26] ) );
  DFFR_X1 \REGISTERS_reg[51][25]  ( .D(n7955), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][25] ) );
  DFFR_X1 \REGISTERS_reg[51][24]  ( .D(n7956), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][24] ) );
  DFFR_X1 \REGISTERS_reg[51][23]  ( .D(n7957), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][23] ) );
  DFFR_X1 \REGISTERS_reg[51][22]  ( .D(n7958), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][22] ) );
  DFFR_X1 \REGISTERS_reg[51][21]  ( .D(n7959), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][21] ) );
  DFFR_X1 \REGISTERS_reg[51][20]  ( .D(n7960), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][20] ) );
  DFFR_X1 \REGISTERS_reg[51][19]  ( .D(n7961), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][19] ) );
  DFFR_X1 \REGISTERS_reg[51][18]  ( .D(n7962), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][18] ) );
  DFFR_X1 \REGISTERS_reg[51][17]  ( .D(n7963), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][17] ) );
  DFFR_X1 \REGISTERS_reg[51][16]  ( .D(n7964), .CK(CLK), .RN(n3072), .Q(
        \REGISTERS[51][16] ) );
  DFFR_X1 \REGISTERS_reg[51][15]  ( .D(n7965), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][15] ) );
  DFFR_X1 \REGISTERS_reg[51][14]  ( .D(n7966), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][14] ) );
  DFFR_X1 \REGISTERS_reg[51][13]  ( .D(n7967), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][13] ) );
  DFFR_X1 \REGISTERS_reg[51][12]  ( .D(n7968), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][12] ) );
  DFFR_X1 \REGISTERS_reg[51][11]  ( .D(n7969), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][11] ) );
  DFFR_X1 \REGISTERS_reg[51][10]  ( .D(n7970), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][10] ) );
  DFFR_X1 \REGISTERS_reg[51][9]  ( .D(n7971), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][9] ) );
  DFFR_X1 \REGISTERS_reg[51][8]  ( .D(n7972), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][8] ) );
  DFFR_X1 \REGISTERS_reg[51][7]  ( .D(n7973), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][7] ) );
  DFFR_X1 \REGISTERS_reg[51][6]  ( .D(n7974), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][6] ) );
  DFFR_X1 \REGISTERS_reg[51][5]  ( .D(n7975), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][5] ) );
  DFFR_X1 \REGISTERS_reg[51][4]  ( .D(n7976), .CK(CLK), .RN(n3071), .Q(
        \REGISTERS[51][4] ) );
  DFFR_X1 \REGISTERS_reg[51][3]  ( .D(n7977), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[51][3] ) );
  DFFR_X1 \REGISTERS_reg[51][2]  ( .D(n7978), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[51][2] ) );
  DFFR_X1 \REGISTERS_reg[51][1]  ( .D(n7979), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[51][1] ) );
  DFFR_X1 \REGISTERS_reg[51][0]  ( .D(n7980), .CK(CLK), .RN(n3069), .Q(
        \REGISTERS[51][0] ) );
  DFFR_X1 \REGISTERS_reg[50][31]  ( .D(n7917), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][31] ) );
  DFFR_X1 \REGISTERS_reg[50][30]  ( .D(n7918), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][30] ) );
  DFFR_X1 \REGISTERS_reg[50][29]  ( .D(n7919), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][29] ) );
  DFFR_X1 \REGISTERS_reg[50][28]  ( .D(n7920), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][28] ) );
  DFFR_X1 \REGISTERS_reg[50][27]  ( .D(n7921), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][27] ) );
  DFFR_X1 \REGISTERS_reg[50][26]  ( .D(n7922), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][26] ) );
  DFFR_X1 \REGISTERS_reg[50][25]  ( .D(n7923), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][25] ) );
  DFFR_X1 \REGISTERS_reg[50][24]  ( .D(n7924), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][24] ) );
  DFFR_X1 \REGISTERS_reg[50][23]  ( .D(n7925), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][23] ) );
  DFFR_X1 \REGISTERS_reg[50][22]  ( .D(n7926), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][22] ) );
  DFFR_X1 \REGISTERS_reg[50][21]  ( .D(n7927), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][21] ) );
  DFFR_X1 \REGISTERS_reg[50][20]  ( .D(n7928), .CK(CLK), .RN(n3077), .Q(
        \REGISTERS[50][20] ) );
  DFFR_X1 \REGISTERS_reg[50][19]  ( .D(n7929), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][19] ) );
  DFFR_X1 \REGISTERS_reg[50][18]  ( .D(n7930), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][18] ) );
  DFFR_X1 \REGISTERS_reg[50][17]  ( .D(n7931), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][17] ) );
  DFFR_X1 \REGISTERS_reg[50][16]  ( .D(n7932), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][16] ) );
  DFFR_X1 \REGISTERS_reg[50][15]  ( .D(n7933), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][15] ) );
  DFFR_X1 \REGISTERS_reg[50][14]  ( .D(n7934), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][14] ) );
  DFFR_X1 \REGISTERS_reg[50][13]  ( .D(n7935), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][13] ) );
  DFFR_X1 \REGISTERS_reg[50][12]  ( .D(n7936), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][12] ) );
  DFFR_X1 \REGISTERS_reg[50][11]  ( .D(n7937), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][11] ) );
  DFFR_X1 \REGISTERS_reg[50][10]  ( .D(n7938), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][10] ) );
  DFFR_X1 \REGISTERS_reg[50][9]  ( .D(n7939), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][9] ) );
  DFFR_X1 \REGISTERS_reg[50][8]  ( .D(n7940), .CK(CLK), .RN(n3076), .Q(
        \REGISTERS[50][8] ) );
  DFFR_X1 \REGISTERS_reg[50][7]  ( .D(n7941), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[50][7] ) );
  DFFR_X1 \REGISTERS_reg[50][6]  ( .D(n7942), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[50][6] ) );
  DFFR_X1 \REGISTERS_reg[50][5]  ( .D(n7943), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[50][5] ) );
  DFFR_X1 \REGISTERS_reg[50][4]  ( .D(n7944), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[50][4] ) );
  DFFR_X1 \REGISTERS_reg[50][3]  ( .D(n7945), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[50][3] ) );
  DFFR_X1 \REGISTERS_reg[50][2]  ( .D(n7946), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[50][2] ) );
  DFFR_X1 \REGISTERS_reg[50][1]  ( .D(n7947), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[50][1] ) );
  DFFR_X1 \REGISTERS_reg[50][0]  ( .D(n7948), .CK(CLK), .RN(n3074), .Q(
        \REGISTERS[50][0] ) );
  DFFR_X1 \REGISTERS_reg[49][31]  ( .D(n7885), .CK(CLK), .RN(n3082), .Q(
        \REGISTERS[49][31] ) );
  DFFR_X1 \REGISTERS_reg[49][30]  ( .D(n7886), .CK(CLK), .RN(n3082), .Q(
        \REGISTERS[49][30] ) );
  DFFR_X1 \REGISTERS_reg[49][29]  ( .D(n7887), .CK(CLK), .RN(n3082), .Q(
        \REGISTERS[49][29] ) );
  DFFR_X1 \REGISTERS_reg[49][28]  ( .D(n7888), .CK(CLK), .RN(n3082), .Q(
        \REGISTERS[49][28] ) );
  DFFR_X1 \REGISTERS_reg[49][27]  ( .D(n7889), .CK(CLK), .RN(n3082), .Q(
        \REGISTERS[49][27] ) );
  DFFR_X1 \REGISTERS_reg[49][26]  ( .D(n7890), .CK(CLK), .RN(n3082), .Q(
        \REGISTERS[49][26] ) );
  DFFR_X1 \REGISTERS_reg[49][25]  ( .D(n7891), .CK(CLK), .RN(n3082), .Q(
        \REGISTERS[49][25] ) );
  DFFR_X1 \REGISTERS_reg[49][24]  ( .D(n7892), .CK(CLK), .RN(n3082), .Q(
        \REGISTERS[49][24] ) );
  DFFR_X1 \REGISTERS_reg[49][23]  ( .D(n7893), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][23] ) );
  DFFR_X1 \REGISTERS_reg[49][22]  ( .D(n7894), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][22] ) );
  DFFR_X1 \REGISTERS_reg[49][21]  ( .D(n7895), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][21] ) );
  DFFR_X1 \REGISTERS_reg[49][20]  ( .D(n7896), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][20] ) );
  DFFR_X1 \REGISTERS_reg[49][19]  ( .D(n7897), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][19] ) );
  DFFR_X1 \REGISTERS_reg[49][18]  ( .D(n7898), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][18] ) );
  DFFR_X1 \REGISTERS_reg[49][17]  ( .D(n7899), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][17] ) );
  DFFR_X1 \REGISTERS_reg[49][16]  ( .D(n7900), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][16] ) );
  DFFR_X1 \REGISTERS_reg[49][15]  ( .D(n7901), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][15] ) );
  DFFR_X1 \REGISTERS_reg[49][14]  ( .D(n7902), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][14] ) );
  DFFR_X1 \REGISTERS_reg[49][13]  ( .D(n7903), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][13] ) );
  DFFR_X1 \REGISTERS_reg[49][12]  ( .D(n7904), .CK(CLK), .RN(n3081), .Q(
        \REGISTERS[49][12] ) );
  DFFR_X1 \REGISTERS_reg[49][11]  ( .D(n7905), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][11] ) );
  DFFR_X1 \REGISTERS_reg[49][10]  ( .D(n7906), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][10] ) );
  DFFR_X1 \REGISTERS_reg[49][9]  ( .D(n7907), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][9] ) );
  DFFR_X1 \REGISTERS_reg[49][8]  ( .D(n7908), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][8] ) );
  DFFR_X1 \REGISTERS_reg[49][7]  ( .D(n7909), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][7] ) );
  DFFR_X1 \REGISTERS_reg[49][6]  ( .D(n7910), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][6] ) );
  DFFR_X1 \REGISTERS_reg[49][5]  ( .D(n7911), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][5] ) );
  DFFR_X1 \REGISTERS_reg[49][4]  ( .D(n7912), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][4] ) );
  DFFR_X1 \REGISTERS_reg[49][3]  ( .D(n7913), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][3] ) );
  DFFR_X1 \REGISTERS_reg[49][2]  ( .D(n7914), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][2] ) );
  DFFR_X1 \REGISTERS_reg[49][1]  ( .D(n7915), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][1] ) );
  DFFR_X1 \REGISTERS_reg[49][0]  ( .D(n7916), .CK(CLK), .RN(n3079), .Q(
        \REGISTERS[49][0] ) );
  DFFR_X1 \REGISTERS_reg[45][31]  ( .D(n7757), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[45][31] ) );
  DFFR_X1 \REGISTERS_reg[45][30]  ( .D(n7758), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[45][30] ) );
  DFFR_X1 \REGISTERS_reg[45][29]  ( .D(n7759), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[45][29] ) );
  DFFR_X1 \REGISTERS_reg[45][28]  ( .D(n7760), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[45][28] ) );
  DFFR_X1 \REGISTERS_reg[45][27]  ( .D(n7761), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][27] ) );
  DFFR_X1 \REGISTERS_reg[45][26]  ( .D(n7762), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][26] ) );
  DFFR_X1 \REGISTERS_reg[45][25]  ( .D(n7763), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][25] ) );
  DFFR_X1 \REGISTERS_reg[45][24]  ( .D(n7764), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][24] ) );
  DFFR_X1 \REGISTERS_reg[45][23]  ( .D(n7765), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][23] ) );
  DFFR_X1 \REGISTERS_reg[45][22]  ( .D(n7766), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][22] ) );
  DFFR_X1 \REGISTERS_reg[45][21]  ( .D(n7767), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][21] ) );
  DFFR_X1 \REGISTERS_reg[45][20]  ( .D(n7768), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][20] ) );
  DFFR_X1 \REGISTERS_reg[45][19]  ( .D(n7769), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][19] ) );
  DFFR_X1 \REGISTERS_reg[45][18]  ( .D(n7770), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][18] ) );
  DFFR_X1 \REGISTERS_reg[45][17]  ( .D(n7771), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][17] ) );
  DFFR_X1 \REGISTERS_reg[45][16]  ( .D(n7772), .CK(CLK), .RN(n3099), .Q(
        \REGISTERS[45][16] ) );
  DFFR_X1 \REGISTERS_reg[45][15]  ( .D(n7773), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][15] ) );
  DFFR_X1 \REGISTERS_reg[45][14]  ( .D(n7774), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][14] ) );
  DFFR_X1 \REGISTERS_reg[45][13]  ( .D(n7775), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][13] ) );
  DFFR_X1 \REGISTERS_reg[45][12]  ( .D(n7776), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][12] ) );
  DFFR_X1 \REGISTERS_reg[45][11]  ( .D(n7777), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][11] ) );
  DFFR_X1 \REGISTERS_reg[45][10]  ( .D(n7778), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][10] ) );
  DFFR_X1 \REGISTERS_reg[45][9]  ( .D(n7779), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][9] ) );
  DFFR_X1 \REGISTERS_reg[45][8]  ( .D(n7780), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][8] ) );
  DFFR_X1 \REGISTERS_reg[45][7]  ( .D(n7781), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][7] ) );
  DFFR_X1 \REGISTERS_reg[45][6]  ( .D(n7782), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][6] ) );
  DFFR_X1 \REGISTERS_reg[45][5]  ( .D(n7783), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][5] ) );
  DFFR_X1 \REGISTERS_reg[45][4]  ( .D(n7784), .CK(CLK), .RN(n3097), .Q(
        \REGISTERS[45][4] ) );
  DFFR_X1 \REGISTERS_reg[45][3]  ( .D(n7785), .CK(CLK), .RN(n3096), .Q(
        \REGISTERS[45][3] ) );
  DFFR_X1 \REGISTERS_reg[45][2]  ( .D(n7786), .CK(CLK), .RN(n3096), .Q(
        \REGISTERS[45][2] ) );
  DFFR_X1 \REGISTERS_reg[45][1]  ( .D(n7787), .CK(CLK), .RN(n3096), .Q(
        \REGISTERS[45][1] ) );
  DFFR_X1 \REGISTERS_reg[45][0]  ( .D(n7788), .CK(CLK), .RN(n3096), .Q(
        \REGISTERS[45][0] ) );
  DFFR_X1 \REGISTERS_reg[44][31]  ( .D(n7725), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][31] ) );
  DFFR_X1 \REGISTERS_reg[44][30]  ( .D(n7726), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][30] ) );
  DFFR_X1 \REGISTERS_reg[44][29]  ( .D(n7727), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][29] ) );
  DFFR_X1 \REGISTERS_reg[44][28]  ( .D(n7728), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][28] ) );
  DFFR_X1 \REGISTERS_reg[44][27]  ( .D(n7729), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][27] ) );
  DFFR_X1 \REGISTERS_reg[44][26]  ( .D(n7730), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][26] ) );
  DFFR_X1 \REGISTERS_reg[44][25]  ( .D(n7731), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][25] ) );
  DFFR_X1 \REGISTERS_reg[44][24]  ( .D(n7732), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][24] ) );
  DFFR_X1 \REGISTERS_reg[44][23]  ( .D(n7733), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][23] ) );
  DFFR_X1 \REGISTERS_reg[44][22]  ( .D(n7734), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][22] ) );
  DFFR_X1 \REGISTERS_reg[44][21]  ( .D(n7735), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][21] ) );
  DFFR_X1 \REGISTERS_reg[44][20]  ( .D(n7736), .CK(CLK), .RN(n3104), .Q(
        \REGISTERS[44][20] ) );
  DFFR_X1 \REGISTERS_reg[44][19]  ( .D(n7737), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][19] ) );
  DFFR_X1 \REGISTERS_reg[44][18]  ( .D(n7738), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][18] ) );
  DFFR_X1 \REGISTERS_reg[44][17]  ( .D(n7739), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][17] ) );
  DFFR_X1 \REGISTERS_reg[44][16]  ( .D(n7740), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][16] ) );
  DFFR_X1 \REGISTERS_reg[44][15]  ( .D(n7741), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][15] ) );
  DFFR_X1 \REGISTERS_reg[44][14]  ( .D(n7742), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][14] ) );
  DFFR_X1 \REGISTERS_reg[44][13]  ( .D(n7743), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][13] ) );
  DFFR_X1 \REGISTERS_reg[44][12]  ( .D(n7744), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][12] ) );
  DFFR_X1 \REGISTERS_reg[44][11]  ( .D(n7745), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][11] ) );
  DFFR_X1 \REGISTERS_reg[44][10]  ( .D(n7746), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][10] ) );
  DFFR_X1 \REGISTERS_reg[44][9]  ( .D(n7747), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][9] ) );
  DFFR_X1 \REGISTERS_reg[44][8]  ( .D(n7748), .CK(CLK), .RN(n3102), .Q(
        \REGISTERS[44][8] ) );
  DFFR_X1 \REGISTERS_reg[44][7]  ( .D(n7749), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[44][7] ) );
  DFFR_X1 \REGISTERS_reg[44][6]  ( .D(n7750), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[44][6] ) );
  DFFR_X1 \REGISTERS_reg[44][5]  ( .D(n7751), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[44][5] ) );
  DFFR_X1 \REGISTERS_reg[44][4]  ( .D(n7752), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[44][4] ) );
  DFFR_X1 \REGISTERS_reg[44][3]  ( .D(n7753), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[44][3] ) );
  DFFR_X1 \REGISTERS_reg[44][2]  ( .D(n7754), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[44][2] ) );
  DFFR_X1 \REGISTERS_reg[44][1]  ( .D(n7755), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[44][1] ) );
  DFFR_X1 \REGISTERS_reg[44][0]  ( .D(n7756), .CK(CLK), .RN(n3101), .Q(
        \REGISTERS[44][0] ) );
  DFFR_X1 \REGISTERS_reg[43][31]  ( .D(n7693), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[43][31] ) );
  DFFR_X1 \REGISTERS_reg[43][30]  ( .D(n7694), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[43][30] ) );
  DFFR_X1 \REGISTERS_reg[43][29]  ( .D(n7695), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[43][29] ) );
  DFFR_X1 \REGISTERS_reg[43][28]  ( .D(n7696), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[43][28] ) );
  DFFR_X1 \REGISTERS_reg[43][27]  ( .D(n7697), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[43][27] ) );
  DFFR_X1 \REGISTERS_reg[43][26]  ( .D(n7698), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[43][26] ) );
  DFFR_X1 \REGISTERS_reg[43][25]  ( .D(n7699), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[43][25] ) );
  DFFR_X1 \REGISTERS_reg[43][24]  ( .D(n7700), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[43][24] ) );
  DFFR_X1 \REGISTERS_reg[43][23]  ( .D(n7701), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][23] ) );
  DFFR_X1 \REGISTERS_reg[43][22]  ( .D(n7702), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][22] ) );
  DFFR_X1 \REGISTERS_reg[43][21]  ( .D(n7703), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][21] ) );
  DFFR_X1 \REGISTERS_reg[43][20]  ( .D(n7704), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][20] ) );
  DFFR_X1 \REGISTERS_reg[43][19]  ( .D(n7705), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][19] ) );
  DFFR_X1 \REGISTERS_reg[43][18]  ( .D(n7706), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][18] ) );
  DFFR_X1 \REGISTERS_reg[43][17]  ( .D(n7707), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][17] ) );
  DFFR_X1 \REGISTERS_reg[43][16]  ( .D(n7708), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][16] ) );
  DFFR_X1 \REGISTERS_reg[43][15]  ( .D(n7709), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][15] ) );
  DFFR_X1 \REGISTERS_reg[43][14]  ( .D(n7710), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][14] ) );
  DFFR_X1 \REGISTERS_reg[43][13]  ( .D(n7711), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][13] ) );
  DFFR_X1 \REGISTERS_reg[43][12]  ( .D(n7712), .CK(CLK), .RN(n3111), .Q(
        \REGISTERS[43][12] ) );
  DFFR_X1 \REGISTERS_reg[43][11]  ( .D(n7713), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][11] ) );
  DFFR_X1 \REGISTERS_reg[43][10]  ( .D(n7714), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][10] ) );
  DFFR_X1 \REGISTERS_reg[43][9]  ( .D(n7715), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][9] ) );
  DFFR_X1 \REGISTERS_reg[43][8]  ( .D(n7716), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][8] ) );
  DFFR_X1 \REGISTERS_reg[43][7]  ( .D(n7717), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][7] ) );
  DFFR_X1 \REGISTERS_reg[43][6]  ( .D(n7718), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][6] ) );
  DFFR_X1 \REGISTERS_reg[43][5]  ( .D(n7719), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][5] ) );
  DFFR_X1 \REGISTERS_reg[43][4]  ( .D(n7720), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][4] ) );
  DFFR_X1 \REGISTERS_reg[43][3]  ( .D(n7721), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][3] ) );
  DFFR_X1 \REGISTERS_reg[43][2]  ( .D(n7722), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][2] ) );
  DFFR_X1 \REGISTERS_reg[43][1]  ( .D(n7723), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][1] ) );
  DFFR_X1 \REGISTERS_reg[43][0]  ( .D(n7724), .CK(CLK), .RN(n3110), .Q(
        \REGISTERS[43][0] ) );
  DFFR_X1 \REGISTERS_reg[42][31]  ( .D(n7661), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[42][31] ) );
  DFFR_X1 \REGISTERS_reg[42][30]  ( .D(n7662), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[42][30] ) );
  DFFR_X1 \REGISTERS_reg[42][29]  ( .D(n7663), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[42][29] ) );
  DFFR_X1 \REGISTERS_reg[42][28]  ( .D(n7664), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[42][28] ) );
  DFFR_X1 \REGISTERS_reg[42][27]  ( .D(n7665), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][27] ) );
  DFFR_X1 \REGISTERS_reg[42][26]  ( .D(n7666), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][26] ) );
  DFFR_X1 \REGISTERS_reg[42][25]  ( .D(n7667), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][25] ) );
  DFFR_X1 \REGISTERS_reg[42][24]  ( .D(n7668), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][24] ) );
  DFFR_X1 \REGISTERS_reg[42][23]  ( .D(n7669), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][23] ) );
  DFFR_X1 \REGISTERS_reg[42][22]  ( .D(n7670), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][22] ) );
  DFFR_X1 \REGISTERS_reg[42][21]  ( .D(n7671), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][21] ) );
  DFFR_X1 \REGISTERS_reg[42][20]  ( .D(n7672), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][20] ) );
  DFFR_X1 \REGISTERS_reg[42][19]  ( .D(n7673), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][19] ) );
  DFFR_X1 \REGISTERS_reg[42][18]  ( .D(n7674), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][18] ) );
  DFFR_X1 \REGISTERS_reg[42][17]  ( .D(n7675), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][17] ) );
  DFFR_X1 \REGISTERS_reg[42][16]  ( .D(n7676), .CK(CLK), .RN(n3116), .Q(
        \REGISTERS[42][16] ) );
  DFFR_X1 \REGISTERS_reg[42][15]  ( .D(n7677), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][15] ) );
  DFFR_X1 \REGISTERS_reg[42][14]  ( .D(n7678), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][14] ) );
  DFFR_X1 \REGISTERS_reg[42][13]  ( .D(n7679), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][13] ) );
  DFFR_X1 \REGISTERS_reg[42][12]  ( .D(n7680), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][12] ) );
  DFFR_X1 \REGISTERS_reg[42][11]  ( .D(n7681), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][11] ) );
  DFFR_X1 \REGISTERS_reg[42][10]  ( .D(n7682), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][10] ) );
  DFFR_X1 \REGISTERS_reg[42][9]  ( .D(n7683), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][9] ) );
  DFFR_X1 \REGISTERS_reg[42][8]  ( .D(n7684), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][8] ) );
  DFFR_X1 \REGISTERS_reg[42][7]  ( .D(n7685), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][7] ) );
  DFFR_X1 \REGISTERS_reg[42][6]  ( .D(n7686), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][6] ) );
  DFFR_X1 \REGISTERS_reg[42][5]  ( .D(n7687), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][5] ) );
  DFFR_X1 \REGISTERS_reg[42][4]  ( .D(n7688), .CK(CLK), .RN(n3115), .Q(
        \REGISTERS[42][4] ) );
  DFFR_X1 \REGISTERS_reg[42][3]  ( .D(n7689), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[42][3] ) );
  DFFR_X1 \REGISTERS_reg[42][2]  ( .D(n7690), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[42][2] ) );
  DFFR_X1 \REGISTERS_reg[42][1]  ( .D(n7691), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[42][1] ) );
  DFFR_X1 \REGISTERS_reg[42][0]  ( .D(n7692), .CK(CLK), .RN(n3113), .Q(
        \REGISTERS[42][0] ) );
  DFFR_X1 \REGISTERS_reg[41][31]  ( .D(n7629), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][31] ) );
  DFFR_X1 \REGISTERS_reg[41][30]  ( .D(n7630), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][30] ) );
  DFFR_X1 \REGISTERS_reg[41][29]  ( .D(n7631), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][29] ) );
  DFFR_X1 \REGISTERS_reg[41][28]  ( .D(n7632), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][28] ) );
  DFFR_X1 \REGISTERS_reg[41][27]  ( .D(n7633), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][27] ) );
  DFFR_X1 \REGISTERS_reg[41][26]  ( .D(n7634), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][26] ) );
  DFFR_X1 \REGISTERS_reg[41][25]  ( .D(n7635), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][25] ) );
  DFFR_X1 \REGISTERS_reg[41][24]  ( .D(n7636), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][24] ) );
  DFFR_X1 \REGISTERS_reg[41][23]  ( .D(n7637), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][23] ) );
  DFFR_X1 \REGISTERS_reg[41][22]  ( .D(n7638), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][22] ) );
  DFFR_X1 \REGISTERS_reg[41][21]  ( .D(n7639), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][21] ) );
  DFFR_X1 \REGISTERS_reg[41][20]  ( .D(n7640), .CK(CLK), .RN(n3120), .Q(
        \REGISTERS[41][20] ) );
  DFFR_X1 \REGISTERS_reg[41][19]  ( .D(n7641), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][19] ) );
  DFFR_X1 \REGISTERS_reg[41][18]  ( .D(n7642), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][18] ) );
  DFFR_X1 \REGISTERS_reg[41][17]  ( .D(n7643), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][17] ) );
  DFFR_X1 \REGISTERS_reg[41][16]  ( .D(n7644), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][16] ) );
  DFFR_X1 \REGISTERS_reg[41][15]  ( .D(n7645), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][15] ) );
  DFFR_X1 \REGISTERS_reg[41][14]  ( .D(n7646), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][14] ) );
  DFFR_X1 \REGISTERS_reg[41][13]  ( .D(n7647), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][13] ) );
  DFFR_X1 \REGISTERS_reg[41][12]  ( .D(n7648), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][12] ) );
  DFFR_X1 \REGISTERS_reg[41][11]  ( .D(n7649), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][11] ) );
  DFFR_X1 \REGISTERS_reg[41][10]  ( .D(n7650), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][10] ) );
  DFFR_X1 \REGISTERS_reg[41][9]  ( .D(n7651), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][9] ) );
  DFFR_X1 \REGISTERS_reg[41][8]  ( .D(n7652), .CK(CLK), .RN(n3119), .Q(
        \REGISTERS[41][8] ) );
  DFFR_X1 \REGISTERS_reg[41][7]  ( .D(n7653), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[41][7] ) );
  DFFR_X1 \REGISTERS_reg[41][6]  ( .D(n7654), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[41][6] ) );
  DFFR_X1 \REGISTERS_reg[41][5]  ( .D(n7655), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[41][5] ) );
  DFFR_X1 \REGISTERS_reg[41][4]  ( .D(n7656), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[41][4] ) );
  DFFR_X1 \REGISTERS_reg[41][3]  ( .D(n7657), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[41][3] ) );
  DFFR_X1 \REGISTERS_reg[41][2]  ( .D(n7658), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[41][2] ) );
  DFFR_X1 \REGISTERS_reg[41][1]  ( .D(n7659), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[41][1] ) );
  DFFR_X1 \REGISTERS_reg[41][0]  ( .D(n7660), .CK(CLK), .RN(n3118), .Q(
        \REGISTERS[41][0] ) );
  DFFR_X1 \REGISTERS_reg[40][31]  ( .D(n7597), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[40][31] ) );
  DFFR_X1 \REGISTERS_reg[40][30]  ( .D(n7598), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[40][30] ) );
  DFFR_X1 \REGISTERS_reg[40][29]  ( .D(n7599), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[40][29] ) );
  DFFR_X1 \REGISTERS_reg[40][28]  ( .D(n7600), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[40][28] ) );
  DFFR_X1 \REGISTERS_reg[40][27]  ( .D(n7601), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[40][27] ) );
  DFFR_X1 \REGISTERS_reg[40][26]  ( .D(n7602), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[40][26] ) );
  DFFR_X1 \REGISTERS_reg[40][25]  ( .D(n7603), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[40][25] ) );
  DFFR_X1 \REGISTERS_reg[40][24]  ( .D(n7604), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[40][24] ) );
  DFFR_X1 \REGISTERS_reg[40][23]  ( .D(n7605), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][23] ) );
  DFFR_X1 \REGISTERS_reg[40][22]  ( .D(n7606), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][22] ) );
  DFFR_X1 \REGISTERS_reg[40][21]  ( .D(n7607), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][21] ) );
  DFFR_X1 \REGISTERS_reg[40][20]  ( .D(n7608), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][20] ) );
  DFFR_X1 \REGISTERS_reg[40][19]  ( .D(n7609), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][19] ) );
  DFFR_X1 \REGISTERS_reg[40][18]  ( .D(n7610), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][18] ) );
  DFFR_X1 \REGISTERS_reg[40][17]  ( .D(n7611), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][17] ) );
  DFFR_X1 \REGISTERS_reg[40][16]  ( .D(n7612), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][16] ) );
  DFFR_X1 \REGISTERS_reg[40][15]  ( .D(n7613), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][15] ) );
  DFFR_X1 \REGISTERS_reg[40][14]  ( .D(n7614), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][14] ) );
  DFFR_X1 \REGISTERS_reg[40][13]  ( .D(n7615), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][13] ) );
  DFFR_X1 \REGISTERS_reg[40][12]  ( .D(n7616), .CK(CLK), .RN(n3123), .Q(
        \REGISTERS[40][12] ) );
  DFFR_X1 \REGISTERS_reg[40][11]  ( .D(n7617), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][11] ) );
  DFFR_X1 \REGISTERS_reg[40][10]  ( .D(n7618), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][10] ) );
  DFFR_X1 \REGISTERS_reg[40][9]  ( .D(n7619), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][9] ) );
  DFFR_X1 \REGISTERS_reg[40][8]  ( .D(n7620), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][8] ) );
  DFFR_X1 \REGISTERS_reg[40][7]  ( .D(n7621), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][7] ) );
  DFFR_X1 \REGISTERS_reg[40][6]  ( .D(n7622), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][6] ) );
  DFFR_X1 \REGISTERS_reg[40][5]  ( .D(n7623), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][5] ) );
  DFFR_X1 \REGISTERS_reg[40][4]  ( .D(n7624), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][4] ) );
  DFFR_X1 \REGISTERS_reg[40][3]  ( .D(n7625), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][3] ) );
  DFFR_X1 \REGISTERS_reg[40][2]  ( .D(n7626), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][2] ) );
  DFFR_X1 \REGISTERS_reg[40][1]  ( .D(n7627), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][1] ) );
  DFFR_X1 \REGISTERS_reg[40][0]  ( .D(n7628), .CK(CLK), .RN(n3122), .Q(
        \REGISTERS[40][0] ) );
  DFFR_X1 \REGISTERS_reg[39][31]  ( .D(n7565), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[39][31] ) );
  DFFR_X1 \REGISTERS_reg[39][30]  ( .D(n7566), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[39][30] ) );
  DFFR_X1 \REGISTERS_reg[39][29]  ( .D(n7567), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[39][29] ) );
  DFFR_X1 \REGISTERS_reg[39][28]  ( .D(n7568), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[39][28] ) );
  DFFR_X1 \REGISTERS_reg[39][27]  ( .D(n7569), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][27] ) );
  DFFR_X1 \REGISTERS_reg[39][26]  ( .D(n7570), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][26] ) );
  DFFR_X1 \REGISTERS_reg[39][25]  ( .D(n7571), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][25] ) );
  DFFR_X1 \REGISTERS_reg[39][24]  ( .D(n7572), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][24] ) );
  DFFR_X1 \REGISTERS_reg[39][23]  ( .D(n7573), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][23] ) );
  DFFR_X1 \REGISTERS_reg[39][22]  ( .D(n7574), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][22] ) );
  DFFR_X1 \REGISTERS_reg[39][21]  ( .D(n7575), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][21] ) );
  DFFR_X1 \REGISTERS_reg[39][20]  ( .D(n7576), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][20] ) );
  DFFR_X1 \REGISTERS_reg[39][19]  ( .D(n7577), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][19] ) );
  DFFR_X1 \REGISTERS_reg[39][18]  ( .D(n7578), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][18] ) );
  DFFR_X1 \REGISTERS_reg[39][17]  ( .D(n7579), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][17] ) );
  DFFR_X1 \REGISTERS_reg[39][16]  ( .D(n7580), .CK(CLK), .RN(n3127), .Q(
        \REGISTERS[39][16] ) );
  DFFR_X1 \REGISTERS_reg[39][15]  ( .D(n7581), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][15] ) );
  DFFR_X1 \REGISTERS_reg[39][14]  ( .D(n7582), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][14] ) );
  DFFR_X1 \REGISTERS_reg[39][13]  ( .D(n7583), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][13] ) );
  DFFR_X1 \REGISTERS_reg[39][12]  ( .D(n7584), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][12] ) );
  DFFR_X1 \REGISTERS_reg[39][11]  ( .D(n7585), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][11] ) );
  DFFR_X1 \REGISTERS_reg[39][10]  ( .D(n7586), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][10] ) );
  DFFR_X1 \REGISTERS_reg[39][9]  ( .D(n7587), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][9] ) );
  DFFR_X1 \REGISTERS_reg[39][8]  ( .D(n7588), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][8] ) );
  DFFR_X1 \REGISTERS_reg[39][7]  ( .D(n7589), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][7] ) );
  DFFR_X1 \REGISTERS_reg[39][6]  ( .D(n7590), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][6] ) );
  DFFR_X1 \REGISTERS_reg[39][5]  ( .D(n7591), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][5] ) );
  DFFR_X1 \REGISTERS_reg[39][4]  ( .D(n7592), .CK(CLK), .RN(n3126), .Q(
        \REGISTERS[39][4] ) );
  DFFR_X1 \REGISTERS_reg[39][3]  ( .D(n7593), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[39][3] ) );
  DFFR_X1 \REGISTERS_reg[39][2]  ( .D(n7594), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[39][2] ) );
  DFFR_X1 \REGISTERS_reg[39][1]  ( .D(n7595), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[39][1] ) );
  DFFR_X1 \REGISTERS_reg[39][0]  ( .D(n7596), .CK(CLK), .RN(n3124), .Q(
        \REGISTERS[39][0] ) );
  DFFR_X1 \REGISTERS_reg[38][31]  ( .D(n7533), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][31] ) );
  DFFR_X1 \REGISTERS_reg[38][30]  ( .D(n7534), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][30] ) );
  DFFR_X1 \REGISTERS_reg[38][29]  ( .D(n7535), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][29] ) );
  DFFR_X1 \REGISTERS_reg[38][28]  ( .D(n7536), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][28] ) );
  DFFR_X1 \REGISTERS_reg[38][27]  ( .D(n7537), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][27] ) );
  DFFR_X1 \REGISTERS_reg[38][26]  ( .D(n7538), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][26] ) );
  DFFR_X1 \REGISTERS_reg[38][25]  ( .D(n7539), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][25] ) );
  DFFR_X1 \REGISTERS_reg[38][24]  ( .D(n7540), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][24] ) );
  DFFR_X1 \REGISTERS_reg[38][23]  ( .D(n7541), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][23] ) );
  DFFR_X1 \REGISTERS_reg[38][22]  ( .D(n7542), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][22] ) );
  DFFR_X1 \REGISTERS_reg[38][21]  ( .D(n7543), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][21] ) );
  DFFR_X1 \REGISTERS_reg[38][20]  ( .D(n7544), .CK(CLK), .RN(n3131), .Q(
        \REGISTERS[38][20] ) );
  DFFR_X1 \REGISTERS_reg[38][19]  ( .D(n7545), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][19] ) );
  DFFR_X1 \REGISTERS_reg[38][18]  ( .D(n7546), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][18] ) );
  DFFR_X1 \REGISTERS_reg[38][17]  ( .D(n7547), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][17] ) );
  DFFR_X1 \REGISTERS_reg[38][16]  ( .D(n7548), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][16] ) );
  DFFR_X1 \REGISTERS_reg[38][15]  ( .D(n7549), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][15] ) );
  DFFR_X1 \REGISTERS_reg[38][14]  ( .D(n7550), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][14] ) );
  DFFR_X1 \REGISTERS_reg[38][13]  ( .D(n7551), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][13] ) );
  DFFR_X1 \REGISTERS_reg[38][12]  ( .D(n7552), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][12] ) );
  DFFR_X1 \REGISTERS_reg[38][11]  ( .D(n7553), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][11] ) );
  DFFR_X1 \REGISTERS_reg[38][10]  ( .D(n7554), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][10] ) );
  DFFR_X1 \REGISTERS_reg[38][9]  ( .D(n7555), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][9] ) );
  DFFR_X1 \REGISTERS_reg[38][8]  ( .D(n7556), .CK(CLK), .RN(n3130), .Q(
        \REGISTERS[38][8] ) );
  DFFR_X1 \REGISTERS_reg[38][7]  ( .D(n7557), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[38][7] ) );
  DFFR_X1 \REGISTERS_reg[38][6]  ( .D(n7558), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[38][6] ) );
  DFFR_X1 \REGISTERS_reg[38][5]  ( .D(n7559), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[38][5] ) );
  DFFR_X1 \REGISTERS_reg[38][4]  ( .D(n7560), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[38][4] ) );
  DFFR_X1 \REGISTERS_reg[38][3]  ( .D(n7561), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[38][3] ) );
  DFFR_X1 \REGISTERS_reg[38][2]  ( .D(n7562), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[38][2] ) );
  DFFR_X1 \REGISTERS_reg[38][1]  ( .D(n7563), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[38][1] ) );
  DFFR_X1 \REGISTERS_reg[38][0]  ( .D(n7564), .CK(CLK), .RN(n3128), .Q(
        \REGISTERS[38][0] ) );
  DFFR_X1 \REGISTERS_reg[34][31]  ( .D(n7405), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[34][31] ) );
  DFFR_X1 \REGISTERS_reg[34][30]  ( .D(n7406), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[34][30] ) );
  DFFR_X1 \REGISTERS_reg[34][29]  ( .D(n7407), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[34][29] ) );
  DFFR_X1 \REGISTERS_reg[34][28]  ( .D(n7408), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[34][28] ) );
  DFFR_X1 \REGISTERS_reg[34][27]  ( .D(n7409), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[34][27] ) );
  DFFR_X1 \REGISTERS_reg[34][26]  ( .D(n7410), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[34][26] ) );
  DFFR_X1 \REGISTERS_reg[34][25]  ( .D(n7411), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[34][25] ) );
  DFFR_X1 \REGISTERS_reg[34][24]  ( .D(n7412), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[34][24] ) );
  DFFR_X1 \REGISTERS_reg[34][23]  ( .D(n7413), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][23] ) );
  DFFR_X1 \REGISTERS_reg[34][22]  ( .D(n7414), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][22] ) );
  DFFR_X1 \REGISTERS_reg[34][21]  ( .D(n7415), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][21] ) );
  DFFR_X1 \REGISTERS_reg[34][20]  ( .D(n7416), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][20] ) );
  DFFR_X1 \REGISTERS_reg[34][19]  ( .D(n7417), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][19] ) );
  DFFR_X1 \REGISTERS_reg[34][18]  ( .D(n7418), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][18] ) );
  DFFR_X1 \REGISTERS_reg[34][17]  ( .D(n7419), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][17] ) );
  DFFR_X1 \REGISTERS_reg[34][16]  ( .D(n7420), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][16] ) );
  DFFR_X1 \REGISTERS_reg[34][15]  ( .D(n7421), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][15] ) );
  DFFR_X1 \REGISTERS_reg[34][14]  ( .D(n7422), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][14] ) );
  DFFR_X1 \REGISTERS_reg[34][13]  ( .D(n7423), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][13] ) );
  DFFR_X1 \REGISTERS_reg[34][12]  ( .D(n7424), .CK(CLK), .RN(n3144), .Q(
        \REGISTERS[34][12] ) );
  DFFR_X1 \REGISTERS_reg[34][11]  ( .D(n7425), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][11] ) );
  DFFR_X1 \REGISTERS_reg[34][10]  ( .D(n7426), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][10] ) );
  DFFR_X1 \REGISTERS_reg[34][9]  ( .D(n7427), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][9] ) );
  DFFR_X1 \REGISTERS_reg[34][8]  ( .D(n7428), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][8] ) );
  DFFR_X1 \REGISTERS_reg[34][7]  ( .D(n7429), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][7] ) );
  DFFR_X1 \REGISTERS_reg[34][6]  ( .D(n7430), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][6] ) );
  DFFR_X1 \REGISTERS_reg[34][5]  ( .D(n7431), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][5] ) );
  DFFR_X1 \REGISTERS_reg[34][4]  ( .D(n7432), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][4] ) );
  DFFR_X1 \REGISTERS_reg[34][3]  ( .D(n7433), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][3] ) );
  DFFR_X1 \REGISTERS_reg[34][2]  ( .D(n7434), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][2] ) );
  DFFR_X1 \REGISTERS_reg[34][1]  ( .D(n7435), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][1] ) );
  DFFR_X1 \REGISTERS_reg[34][0]  ( .D(n7436), .CK(CLK), .RN(n3143), .Q(
        \REGISTERS[34][0] ) );
  DFFR_X1 \REGISTERS_reg[33][31]  ( .D(n7373), .CK(CLK), .RN(n3150), .Q(
        \REGISTERS[33][31] ) );
  DFFR_X1 \REGISTERS_reg[33][30]  ( .D(n7374), .CK(CLK), .RN(n3150), .Q(
        \REGISTERS[33][30] ) );
  DFFR_X1 \REGISTERS_reg[33][29]  ( .D(n7375), .CK(CLK), .RN(n3150), .Q(
        \REGISTERS[33][29] ) );
  DFFR_X1 \REGISTERS_reg[33][28]  ( .D(n7376), .CK(CLK), .RN(n3150), .Q(
        \REGISTERS[33][28] ) );
  DFFR_X1 \REGISTERS_reg[33][27]  ( .D(n7377), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][27] ) );
  DFFR_X1 \REGISTERS_reg[33][26]  ( .D(n7378), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][26] ) );
  DFFR_X1 \REGISTERS_reg[33][25]  ( .D(n7379), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][25] ) );
  DFFR_X1 \REGISTERS_reg[33][24]  ( .D(n7380), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][24] ) );
  DFFR_X1 \REGISTERS_reg[33][23]  ( .D(n7381), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][23] ) );
  DFFR_X1 \REGISTERS_reg[33][22]  ( .D(n7382), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][22] ) );
  DFFR_X1 \REGISTERS_reg[33][21]  ( .D(n7383), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][21] ) );
  DFFR_X1 \REGISTERS_reg[33][20]  ( .D(n7384), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][20] ) );
  DFFR_X1 \REGISTERS_reg[33][19]  ( .D(n7385), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][19] ) );
  DFFR_X1 \REGISTERS_reg[33][18]  ( .D(n7386), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][18] ) );
  DFFR_X1 \REGISTERS_reg[33][17]  ( .D(n7387), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][17] ) );
  DFFR_X1 \REGISTERS_reg[33][16]  ( .D(n7388), .CK(CLK), .RN(n3148), .Q(
        \REGISTERS[33][16] ) );
  DFFR_X1 \REGISTERS_reg[33][15]  ( .D(n7389), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][15] ) );
  DFFR_X1 \REGISTERS_reg[33][14]  ( .D(n7390), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][14] ) );
  DFFR_X1 \REGISTERS_reg[33][13]  ( .D(n7391), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][13] ) );
  DFFR_X1 \REGISTERS_reg[33][12]  ( .D(n7392), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][12] ) );
  DFFR_X1 \REGISTERS_reg[33][11]  ( .D(n7393), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][11] ) );
  DFFR_X1 \REGISTERS_reg[33][10]  ( .D(n7394), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][10] ) );
  DFFR_X1 \REGISTERS_reg[33][9]  ( .D(n7395), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][9] ) );
  DFFR_X1 \REGISTERS_reg[33][8]  ( .D(n7396), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][8] ) );
  DFFR_X1 \REGISTERS_reg[33][7]  ( .D(n7397), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][7] ) );
  DFFR_X1 \REGISTERS_reg[33][6]  ( .D(n7398), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][6] ) );
  DFFR_X1 \REGISTERS_reg[33][5]  ( .D(n7399), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][5] ) );
  DFFR_X1 \REGISTERS_reg[33][4]  ( .D(n7400), .CK(CLK), .RN(n3147), .Q(
        \REGISTERS[33][4] ) );
  DFFR_X1 \REGISTERS_reg[33][3]  ( .D(n7401), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[33][3] ) );
  DFFR_X1 \REGISTERS_reg[33][2]  ( .D(n7402), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[33][2] ) );
  DFFR_X1 \REGISTERS_reg[33][1]  ( .D(n7403), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[33][1] ) );
  DFFR_X1 \REGISTERS_reg[33][0]  ( .D(n7404), .CK(CLK), .RN(n3146), .Q(
        \REGISTERS[33][0] ) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n6989), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[21][31] ) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n6990), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[21][30] ) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n6991), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[21][29] ) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n6992), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[21][28] ) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n6993), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][27] ) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n6994), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][26] ) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n6995), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][25] ) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n6996), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][24] ) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n6997), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][23] ) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n6998), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][22] ) );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n6999), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][21] ) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n7000), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][20] ) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n7001), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][19] ) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n7002), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][18] ) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n7003), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][17] ) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n7004), .CK(CLK), .RN(n3192), .Q(
        \REGISTERS[21][16] ) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n7005), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][15] ) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n7006), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][14] ) );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n7007), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][13] ) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n7008), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][12] ) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n7009), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][11] ) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n7010), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][10] ) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n7011), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][9] ) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n7012), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][8] ) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n7013), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][7] ) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n7014), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][6] ) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n7015), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][5] ) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n7016), .CK(CLK), .RN(n3191), .Q(
        \REGISTERS[21][4] ) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n7017), .CK(CLK), .RN(n3189), .Q(
        \REGISTERS[21][3] ) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n7018), .CK(CLK), .RN(n3189), .Q(
        \REGISTERS[21][2] ) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n7019), .CK(CLK), .RN(n3189), .Q(
        \REGISTERS[21][1] ) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n7020), .CK(CLK), .RN(n3189), .Q(
        \REGISTERS[21][0] ) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n6957), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][31] ) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n6958), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][30] ) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n6959), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][29] ) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n6960), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][28] ) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n6961), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][27] ) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n6962), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][26] ) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n6963), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][25] ) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n6964), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][24] ) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n6965), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][23] ) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n6966), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][22] ) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n6967), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][21] ) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n6968), .CK(CLK), .RN(n3196), .Q(
        \REGISTERS[20][20] ) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n6969), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][19] ) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n6970), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][18] ) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n6971), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][17] ) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n6972), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][16] ) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n6973), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][15] ) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n6974), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][14] ) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n6975), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][13] ) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n6976), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][12] ) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n6977), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][11] ) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n6978), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][10] ) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n6979), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][9] ) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n6980), .CK(CLK), .RN(n3195), .Q(
        \REGISTERS[20][8] ) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n6981), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[20][7] ) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n6982), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[20][6] ) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n6983), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[20][5] ) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n6984), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[20][4] ) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n6985), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[20][3] ) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n6986), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[20][2] ) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n6987), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[20][1] ) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n6988), .CK(CLK), .RN(n3193), .Q(
        \REGISTERS[20][0] ) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n6925), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[19][31] ) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n6926), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[19][30] ) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n6927), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[19][29] ) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n6928), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[19][28] ) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n6929), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[19][27] ) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n6930), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[19][26] ) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n6931), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[19][25] ) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n6932), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[19][24] ) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n6933), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][23] ) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n6934), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][22] ) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n6935), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][21] ) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n6936), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][20] ) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n6937), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][19] ) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n6938), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][18] ) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n6939), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][17] ) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n6940), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][16] ) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n6941), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][15] ) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n6942), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][14] ) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n6943), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][13] ) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n6944), .CK(CLK), .RN(n3199), .Q(
        \REGISTERS[19][12] ) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n6945), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][11] ) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n6946), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][10] ) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n6947), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][9] ) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n6948), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][8] ) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n6949), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][7] ) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n6950), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][6] ) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n6951), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][5] ) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n6952), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][4] ) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n6953), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][3] ) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n6954), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][2] ) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n6955), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][1] ) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n6956), .CK(CLK), .RN(n3197), .Q(
        \REGISTERS[19][0] ) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n6893), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[18][31] ) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n6894), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[18][30] ) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n6895), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[18][29] ) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n6896), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[18][28] ) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n6897), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][27] ) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n6898), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][26] ) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n6899), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][25] ) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n6900), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][24] ) );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n6901), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][23] ) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n6902), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][22] ) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n6903), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][21] ) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n6904), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][20] ) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n6905), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][19] ) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n6906), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][18] ) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n6907), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][17] ) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n6908), .CK(CLK), .RN(n3203), .Q(
        \REGISTERS[18][16] ) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n6909), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][15] ) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n6910), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][14] ) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n6911), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][13] ) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n6912), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][12] ) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n6913), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][11] ) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n6914), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][10] ) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n6915), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][9] ) );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n6916), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][8] ) );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n6917), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][7] ) );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n6918), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][6] ) );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n6919), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][5] ) );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n6920), .CK(CLK), .RN(n3201), .Q(
        \REGISTERS[18][4] ) );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n6921), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[18][3] ) );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n6922), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[18][2] ) );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n6923), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[18][1] ) );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n6924), .CK(CLK), .RN(n3200), .Q(
        \REGISTERS[18][0] ) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n6861), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][31] ) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n6862), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][30] ) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n6863), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][29] ) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n6864), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][28] ) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n6865), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][27] ) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n6866), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][26] ) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n6867), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][25] ) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n6868), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][24] ) );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n6869), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][23] ) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n6870), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][22] ) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n6871), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][21] ) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n6872), .CK(CLK), .RN(n3207), .Q(
        \REGISTERS[17][20] ) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n6873), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][19] ) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n6874), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][18] ) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n6875), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][17] ) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n6876), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][16] ) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n6877), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][15] ) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n6878), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][14] ) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n6879), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][13] ) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n6880), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][12] ) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n6881), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][11] ) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n6882), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][10] ) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n6883), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][9] ) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n6884), .CK(CLK), .RN(n3205), .Q(
        \REGISTERS[17][8] ) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n6885), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[17][7] ) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n6886), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[17][6] ) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n6887), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[17][5] ) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n6888), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[17][4] ) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n6889), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[17][3] ) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n6890), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[17][2] ) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n6891), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[17][1] ) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n6892), .CK(CLK), .RN(n3204), .Q(
        \REGISTERS[17][0] ) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n6829), .CK(CLK), .RN(n3211), .Q(
        \REGISTERS[16][31] ) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n6830), .CK(CLK), .RN(n3211), .Q(
        \REGISTERS[16][30] ) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n6831), .CK(CLK), .RN(n3211), .Q(
        \REGISTERS[16][29] ) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n6832), .CK(CLK), .RN(n3211), .Q(
        \REGISTERS[16][28] ) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n6833), .CK(CLK), .RN(n3211), .Q(
        \REGISTERS[16][27] ) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n6834), .CK(CLK), .RN(n3211), .Q(
        \REGISTERS[16][26] ) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n6835), .CK(CLK), .RN(n3211), .Q(
        \REGISTERS[16][25] ) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n6836), .CK(CLK), .RN(n3211), .Q(
        \REGISTERS[16][24] ) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n6837), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][23] ) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n6838), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][22] ) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n6839), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][21] ) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n6840), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][20] ) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n6841), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][19] ) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n6842), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][18] ) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n6843), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][17] ) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n6844), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][16] ) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n6845), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][15] ) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n6846), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][14] ) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n6847), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][13] ) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n6848), .CK(CLK), .RN(n3209), .Q(
        \REGISTERS[16][12] ) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n6849), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][11] ) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n6850), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][10] ) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n6851), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][9] ) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n6852), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][8] ) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n6853), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][7] ) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n6854), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][6] ) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n6855), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][5] ) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n6856), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][4] ) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n6857), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][3] ) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n6858), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][2] ) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n6859), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][1] ) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n6860), .CK(CLK), .RN(n3208), .Q(
        \REGISTERS[16][0] ) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n6701), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[12][31] ) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n6702), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[12][30] ) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n6703), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[12][29] ) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n6704), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[12][28] ) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n6705), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][27] ) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n6706), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][26] ) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n6707), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][25] ) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n6708), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][24] ) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n6709), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][23] ) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n6710), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][22] ) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n6711), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][21] ) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n6712), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][20] ) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n6713), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][19] ) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n6714), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][18] ) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n6715), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][17] ) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n6716), .CK(CLK), .RN(n3224), .Q(
        \REGISTERS[12][16] ) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n6717), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][15] ) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n6718), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][14] ) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n6719), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][13] ) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n6720), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][12] ) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n6721), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][11] ) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n6722), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][10] ) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n6723), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][9] ) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n6724), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][8] ) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n6725), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][7] ) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n6726), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][6] ) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n6727), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][5] ) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n6728), .CK(CLK), .RN(n3223), .Q(
        \REGISTERS[12][4] ) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n6729), .CK(CLK), .RN(n3221), .Q(
        \REGISTERS[12][3] ) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n6730), .CK(CLK), .RN(n3221), .Q(
        \REGISTERS[12][2] ) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n6731), .CK(CLK), .RN(n3221), .Q(
        \REGISTERS[12][1] ) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n6732), .CK(CLK), .RN(n3221), .Q(
        \REGISTERS[12][0] ) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n6669), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][31] ) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n6670), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][30] ) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n6671), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][29] ) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n6672), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][28] ) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n6673), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][27] ) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n6674), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][26] ) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n6675), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][25] ) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n6676), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][24] ) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n6677), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][23] ) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n6678), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][22] ) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n6679), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][21] ) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n6680), .CK(CLK), .RN(n3228), .Q(
        \REGISTERS[11][20] ) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n6681), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][19] ) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n6682), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][18] ) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n6683), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][17] ) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n6684), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][16] ) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n6685), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][15] ) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n6686), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][14] ) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n6687), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][13] ) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n6688), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][12] ) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n6689), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][11] ) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n6690), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][10] ) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n6691), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][9] ) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n6692), .CK(CLK), .RN(n3227), .Q(
        \REGISTERS[11][8] ) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n6693), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[11][7] ) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n6694), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[11][6] ) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n6695), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[11][5] ) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n6696), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[11][4] ) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n6697), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[11][3] ) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n6698), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[11][2] ) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n6699), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[11][1] ) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n6700), .CK(CLK), .RN(n3225), .Q(
        \REGISTERS[11][0] ) );
  DFFR_X1 \CWP_reg[6]  ( .D(n9133), .CK(CLK), .RN(n2970), .Q(CWP[6]), .QN(
        n2898) );
  DFFR_X1 \CWP_reg[5]  ( .D(n9134), .CK(CLK), .RN(n2969), .Q(CWP[5]), .QN(
        n2916) );
  DFFR_X1 \CWP_reg[4]  ( .D(n9135), .CK(CLK), .RN(n2968), .Q(CWP[4]), .QN(
        N8791) );
  DFFR_X1 \CWP_reg[3]  ( .D(n9136), .CK(CLK), .RN(n2967), .Q(N8790), .QN(n2918) );
  DFFR_X1 \CWP_reg[2]  ( .D(n9137), .CK(CLK), .RN(n2966), .Q(N8789), .QN(n2919) );
  DFFR_X1 \CWP_reg[1]  ( .D(n9138), .CK(CLK), .RN(n2965), .Q(N8788), .QN(n2920) );
  DFFR_X1 \CWP_reg[0]  ( .D(n9139), .CK(CLK), .RN(n2964), .Q(N8787), .QN(n2921) );
  AOI22_X1 U3 ( .A1(N8430), .A2(n10918), .B1(N8423), .B2(N8415), .ZN(n6266) );
  AOI22_X1 U4 ( .A1(N8574), .A2(n10919), .B1(N8567), .B2(N8559), .ZN(n4823) );
  NOR2_X1 U5 ( .A1(n3378), .A2(n6314), .ZN(n6249) );
  NOR2_X1 U6 ( .A1(n3387), .A2(n4871), .ZN(n4806) );
  AOI22_X1 U7 ( .A1(N2165), .A2(n3391), .B1(N2158), .B2(N2151), .ZN(n3108) );
  AOI22_X1 U8 ( .A1(N2166), .A2(n3391), .B1(N2159), .B2(N2151), .ZN(n3107) );
  XOR2_X1 U9 ( .A(CWP[5]), .B(CWP[4]), .Z(n1) );
  NOR2_X1 U10 ( .A1(n3378), .A2(n3379), .ZN(n6247) );
  NOR2_X1 U11 ( .A1(n3387), .A2(n3388), .ZN(n4804) );
  NAND4_X1 U12 ( .A1(n3106), .A2(n3107), .A3(n3108), .A4(n3109), .ZN(n3029) );
  NAND4_X1 U13 ( .A1(n3106), .A2(n3108), .A3(n3109), .A4(n3365), .ZN(n3309) );
  NAND4_X1 U14 ( .A1(n3106), .A2(n3107), .A3(n3109), .A4(n3366), .ZN(n3179) );
  NAND4_X1 U15 ( .A1(n3106), .A2(n3107), .A3(n3368), .A4(n3366), .ZN(n3244) );
  NAND4_X1 U16 ( .A1(n3106), .A2(n3107), .A3(n3108), .A4(n3368), .ZN(n3114) );
  NOR2_X1 U17 ( .A1(n6265), .A2(n6264), .ZN(n6296) );
  NOR2_X1 U18 ( .A1(n4822), .A2(n4821), .ZN(n4853) );
  NOR2_X1 U20 ( .A1(n3376), .A2(n6264), .ZN(n6283) );
  NOR2_X1 U21 ( .A1(n3385), .A2(n4821), .ZN(n4840) );
  NOR2_X1 U22 ( .A1(n6314), .A2(n6315), .ZN(n6251) );
  NOR2_X1 U24 ( .A1(n4871), .A2(n4872), .ZN(n4808) );
  NOR2_X1 U25 ( .A1(n3379), .A2(n6315), .ZN(n6250) );
  NOR2_X1 U26 ( .A1(n3388), .A2(n4872), .ZN(n4807) );
  INV_X1 U27 ( .A(N2166), .ZN(N2165) );
  BUF_X1 U28 ( .A(n3345), .Z(n3301) );
  BUF_X1 U30 ( .A(n3347), .Z(n3300) );
  BUF_X1 U31 ( .A(n3347), .Z(n3298) );
  BUF_X1 U32 ( .A(n3347), .Z(n3297) );
  BUF_X1 U33 ( .A(n3349), .Z(n3296) );
  BUF_X1 U34 ( .A(n3349), .Z(n3293) );
  BUF_X1 U35 ( .A(n3350), .Z(n3292) );
  BUF_X1 U36 ( .A(n3350), .Z(n3290) );
  BUF_X1 U37 ( .A(n3350), .Z(n3289) );
  BUF_X1 U38 ( .A(n3352), .Z(n3288) );
  BUF_X1 U39 ( .A(n3349), .Z(n3294) );
  BUF_X1 U40 ( .A(n3334), .Z(n3331) );
  BUF_X1 U41 ( .A(n3334), .Z(n3330) );
  BUF_X1 U42 ( .A(n3335), .Z(n3329) );
  BUF_X1 U43 ( .A(n3335), .Z(n3327) );
  BUF_X1 U44 ( .A(n3335), .Z(n3326) );
  BUF_X1 U45 ( .A(n3337), .Z(n3325) );
  BUF_X1 U46 ( .A(n3337), .Z(n3323) );
  BUF_X1 U47 ( .A(n3337), .Z(n3322) );
  BUF_X1 U48 ( .A(n3338), .Z(n3321) );
  BUF_X1 U49 ( .A(n3338), .Z(n3319) );
  BUF_X1 U50 ( .A(n3339), .Z(n3317) );
  BUF_X1 U51 ( .A(n3339), .Z(n3315) );
  BUF_X1 U52 ( .A(n3339), .Z(n3314) );
  BUF_X1 U53 ( .A(n3341), .Z(n3313) );
  BUF_X1 U54 ( .A(n3341), .Z(n3311) );
  BUF_X1 U55 ( .A(n3341), .Z(n3310) );
  BUF_X1 U56 ( .A(n3344), .Z(n3308) );
  BUF_X1 U57 ( .A(n3344), .Z(n3306) );
  BUF_X1 U58 ( .A(n3344), .Z(n3305) );
  BUF_X1 U59 ( .A(n3345), .Z(n3304) );
  BUF_X1 U60 ( .A(n3338), .Z(n3318) );
  BUF_X1 U61 ( .A(n3352), .Z(n3286) );
  BUF_X1 U62 ( .A(n3361), .Z(n3265) );
  BUF_X1 U63 ( .A(n3355), .Z(n3277) );
  BUF_X1 U64 ( .A(n3361), .Z(n3266) );
  BUF_X1 U65 ( .A(n3355), .Z(n3278) );
  BUF_X1 U66 ( .A(n3361), .Z(n3268) );
  BUF_X1 U67 ( .A(n3355), .Z(n3280) );
  BUF_X1 U68 ( .A(n3360), .Z(n3269) );
  BUF_X1 U69 ( .A(n3354), .Z(n3281) );
  BUF_X1 U70 ( .A(n3360), .Z(n3270) );
  BUF_X1 U71 ( .A(n3354), .Z(n3282) );
  BUF_X1 U72 ( .A(n3360), .Z(n3272) );
  BUF_X1 U73 ( .A(n3354), .Z(n3284) );
  BUF_X1 U74 ( .A(n3357), .Z(n3273) );
  BUF_X1 U75 ( .A(n3352), .Z(n3285) );
  BUF_X1 U76 ( .A(n3357), .Z(n3274) );
  BUF_X1 U77 ( .A(n3357), .Z(n3276) );
  BUF_X1 U78 ( .A(n3345), .Z(n3302) );
  BUF_X1 U79 ( .A(n3334), .Z(n3333) );
  BUF_X1 U80 ( .A(n4887), .Z(n716) );
  BUF_X1 U81 ( .A(n3444), .Z(n1428) );
  BUF_X1 U82 ( .A(n4887), .Z(n717) );
  BUF_X1 U83 ( .A(n3444), .Z(n1429) );
  BUF_X1 U84 ( .A(n4888), .Z(n713) );
  BUF_X1 U85 ( .A(n3445), .Z(n1425) );
  BUF_X1 U86 ( .A(n4888), .Z(n714) );
  BUF_X1 U87 ( .A(n3445), .Z(n1426) );
  BUF_X1 U88 ( .A(n4887), .Z(n718) );
  BUF_X1 U89 ( .A(n3444), .Z(n1430) );
  BUF_X1 U90 ( .A(n4957), .Z(n464) );
  BUF_X1 U91 ( .A(n3514), .Z(n1176) );
  BUF_X1 U92 ( .A(n4957), .Z(n465) );
  BUF_X1 U93 ( .A(n3514), .Z(n1177) );
  BUF_X1 U94 ( .A(n4927), .Z(n623) );
  BUF_X1 U95 ( .A(n4964), .Z(n446) );
  BUF_X1 U96 ( .A(n4995), .Z(n28) );
  BUF_X1 U97 ( .A(n3484), .Z(n1335) );
  BUF_X1 U98 ( .A(n3521), .Z(n1158) );
  BUF_X1 U99 ( .A(n3552), .Z(n740) );
  BUF_X1 U100 ( .A(n4927), .Z(n624) );
  BUF_X1 U101 ( .A(n4964), .Z(n447) );
  BUF_X1 U102 ( .A(n4995), .Z(n29) );
  BUF_X1 U103 ( .A(n3484), .Z(n1336) );
  BUF_X1 U104 ( .A(n3521), .Z(n1159) );
  BUF_X1 U105 ( .A(n3552), .Z(n741) );
  BUF_X1 U106 ( .A(n4888), .Z(n715) );
  BUF_X1 U107 ( .A(n3445), .Z(n1427) );
  BUF_X1 U108 ( .A(n4909), .Z(n654) );
  BUF_X1 U109 ( .A(n3466), .Z(n1366) );
  BUF_X1 U110 ( .A(n4909), .Z(n653) );
  BUF_X1 U111 ( .A(n3466), .Z(n1365) );
  BUF_X1 U112 ( .A(n4957), .Z(n466) );
  BUF_X1 U113 ( .A(n3514), .Z(n1178) );
  BUF_X1 U114 ( .A(n4927), .Z(n625) );
  BUF_X1 U115 ( .A(n4964), .Z(n448) );
  BUF_X1 U116 ( .A(n4995), .Z(n30) );
  BUF_X1 U117 ( .A(n3484), .Z(n1337) );
  BUF_X1 U118 ( .A(n3521), .Z(n1160) );
  BUF_X1 U119 ( .A(n3552), .Z(n742) );
  BUF_X1 U120 ( .A(n4909), .Z(n655) );
  BUF_X1 U121 ( .A(n3466), .Z(n1367) );
  BUF_X1 U122 ( .A(n3354), .Z(n3361) );
  BUF_X1 U123 ( .A(n3363), .Z(n3355) );
  BUF_X1 U124 ( .A(n3352), .Z(n3360) );
  BUF_X1 U125 ( .A(n3347), .Z(n3354) );
  BUF_X1 U126 ( .A(n3349), .Z(n3357) );
  BUF_X1 U127 ( .A(n3363), .Z(n3347) );
  BUF_X1 U128 ( .A(n3363), .Z(n3350) );
  BUF_X1 U129 ( .A(n3363), .Z(n3349) );
  BUF_X1 U130 ( .A(n3341), .Z(n3337) );
  BUF_X1 U131 ( .A(n3344), .Z(n3339) );
  BUF_X1 U132 ( .A(n3333), .Z(n3341) );
  BUF_X1 U133 ( .A(n3333), .Z(n3344) );
  BUF_X1 U134 ( .A(n3335), .Z(n3338) );
  BUF_X1 U135 ( .A(n3350), .Z(n3352) );
  BUF_X1 U136 ( .A(n3334), .Z(n3345) );
  BUF_X1 U137 ( .A(n3355), .Z(n3334) );
  BUF_X1 U138 ( .A(n3361), .Z(n3335) );
  NAND2_X1 U139 ( .A1(n3383), .A2(n3343), .ZN(n3030) );
  BUF_X1 U140 ( .A(n4980), .Z(n70) );
  BUF_X1 U141 ( .A(n3537), .Z(n782) );
  BUF_X1 U142 ( .A(n4980), .Z(n71) );
  BUF_X1 U143 ( .A(n3537), .Z(n783) );
  BUF_X1 U144 ( .A(n4918), .Z(n650) );
  BUF_X1 U145 ( .A(n3475), .Z(n1362) );
  BUF_X1 U146 ( .A(n4918), .Z(n651) );
  BUF_X1 U147 ( .A(n3475), .Z(n1363) );
  BUF_X1 U148 ( .A(n4949), .Z(n488) );
  BUF_X1 U149 ( .A(n3506), .Z(n1296) );
  BUF_X1 U150 ( .A(n4949), .Z(n489) );
  BUF_X1 U151 ( .A(n3506), .Z(n1297) );
  BUF_X1 U152 ( .A(n4919), .Z(n647) );
  BUF_X1 U153 ( .A(n3476), .Z(n1359) );
  BUF_X1 U154 ( .A(n4919), .Z(n648) );
  BUF_X1 U155 ( .A(n3476), .Z(n1360) );
  BUF_X1 U156 ( .A(n4950), .Z(n485) );
  BUF_X1 U157 ( .A(n4981), .Z(n67) );
  BUF_X1 U158 ( .A(n3507), .Z(n1197) );
  BUF_X1 U159 ( .A(n3538), .Z(n779) );
  BUF_X1 U160 ( .A(n4950), .Z(n486) );
  BUF_X1 U161 ( .A(n4981), .Z(n68) );
  BUF_X1 U162 ( .A(n3507), .Z(n1198) );
  BUF_X1 U163 ( .A(n3538), .Z(n780) );
  BUF_X1 U164 ( .A(n4898), .Z(n683) );
  BUF_X1 U165 ( .A(n4929), .Z(n617) );
  BUF_X1 U166 ( .A(n4960), .Z(n455) );
  BUF_X1 U167 ( .A(n4991), .Z(n37) );
  BUF_X1 U168 ( .A(n3455), .Z(n1395) );
  BUF_X1 U169 ( .A(n3486), .Z(n1329) );
  BUF_X1 U170 ( .A(n3517), .Z(n1167) );
  BUF_X1 U171 ( .A(n3548), .Z(n749) );
  BUF_X1 U172 ( .A(n4898), .Z(n684) );
  BUF_X1 U173 ( .A(n4929), .Z(n618) );
  BUF_X1 U174 ( .A(n4960), .Z(n456) );
  BUF_X1 U175 ( .A(n4991), .Z(n38) );
  BUF_X1 U176 ( .A(n3455), .Z(n1396) );
  BUF_X1 U177 ( .A(n3486), .Z(n1330) );
  BUF_X1 U178 ( .A(n3517), .Z(n1168) );
  BUF_X1 U179 ( .A(n3548), .Z(n750) );
  BUF_X1 U180 ( .A(n4904), .Z(n668) );
  BUF_X1 U181 ( .A(n4907), .Z(n659) );
  BUF_X1 U182 ( .A(n4935), .Z(n602) );
  BUF_X1 U183 ( .A(n4938), .Z(n593) );
  BUF_X1 U184 ( .A(n4966), .Z(n440) );
  BUF_X1 U185 ( .A(n4969), .Z(n79) );
  BUF_X1 U186 ( .A(n4997), .Z(n22) );
  BUF_X1 U187 ( .A(n5000), .Z(n12) );
  BUF_X1 U188 ( .A(n3461), .Z(n1380) );
  BUF_X1 U189 ( .A(n3464), .Z(n1371) );
  BUF_X1 U190 ( .A(n3492), .Z(n1314) );
  BUF_X1 U191 ( .A(n3495), .Z(n1305) );
  BUF_X1 U192 ( .A(n3523), .Z(n1152) );
  BUF_X1 U194 ( .A(n3526), .Z(n1143) );
  BUF_X1 U195 ( .A(n3554), .Z(n734) );
  BUF_X1 U196 ( .A(n3557), .Z(n725) );
  BUF_X1 U197 ( .A(n4904), .Z(n669) );
  BUF_X1 U198 ( .A(n4907), .Z(n660) );
  BUF_X1 U199 ( .A(n4935), .Z(n603) );
  BUF_X1 U200 ( .A(n4938), .Z(n594) );
  BUF_X1 U201 ( .A(n4966), .Z(n441) );
  BUF_X1 U202 ( .A(n4969), .Z(n432) );
  BUF_X1 U203 ( .A(n4997), .Z(n23) );
  BUF_X1 U204 ( .A(n5000), .Z(n13) );
  BUF_X1 U205 ( .A(n3461), .Z(n1381) );
  BUF_X1 U206 ( .A(n3464), .Z(n1372) );
  BUF_X1 U207 ( .A(n3492), .Z(n1315) );
  BUF_X1 U208 ( .A(n3495), .Z(n1306) );
  BUF_X1 U209 ( .A(n3523), .Z(n1153) );
  BUF_X1 U210 ( .A(n3526), .Z(n1144) );
  BUF_X1 U211 ( .A(n3554), .Z(n735) );
  BUF_X1 U212 ( .A(n3557), .Z(n726) );
  BUF_X1 U213 ( .A(n4899), .Z(n680) );
  BUF_X1 U214 ( .A(n4930), .Z(n614) );
  BUF_X1 U215 ( .A(n4961), .Z(n452) );
  BUF_X1 U216 ( .A(n4992), .Z(n34) );
  BUF_X1 U217 ( .A(n3456), .Z(n1392) );
  BUF_X1 U218 ( .A(n3487), .Z(n1326) );
  BUF_X1 U219 ( .A(n3518), .Z(n1164) );
  BUF_X1 U220 ( .A(n3549), .Z(n746) );
  BUF_X1 U221 ( .A(n4899), .Z(n681) );
  BUF_X1 U222 ( .A(n4930), .Z(n615) );
  BUF_X1 U223 ( .A(n4961), .Z(n453) );
  BUF_X1 U224 ( .A(n4992), .Z(n35) );
  BUF_X1 U225 ( .A(n3456), .Z(n1393) );
  BUF_X1 U226 ( .A(n3487), .Z(n1327) );
  BUF_X1 U228 ( .A(n3518), .Z(n1165) );
  BUF_X1 U229 ( .A(n3549), .Z(n747) );
  BUF_X1 U230 ( .A(n4891), .Z(n704) );
  BUF_X1 U231 ( .A(n3448), .Z(n1416) );
  BUF_X1 U232 ( .A(n4891), .Z(n705) );
  BUF_X1 U233 ( .A(n3448), .Z(n1417) );
  BUF_X1 U234 ( .A(n4990), .Z(n40) );
  BUF_X1 U235 ( .A(n4996), .Z(n25) );
  BUF_X1 U236 ( .A(n3547), .Z(n752) );
  BUF_X1 U237 ( .A(n3553), .Z(n737) );
  BUF_X1 U238 ( .A(n4990), .Z(n41) );
  BUF_X1 U239 ( .A(n4996), .Z(n26) );
  BUF_X1 U240 ( .A(n3547), .Z(n753) );
  BUF_X1 U241 ( .A(n3553), .Z(n738) );
  BUF_X1 U242 ( .A(n4894), .Z(n695) );
  BUF_X1 U243 ( .A(n4897), .Z(n686) );
  BUF_X1 U244 ( .A(n4903), .Z(n671) );
  BUF_X1 U245 ( .A(n4922), .Z(n638) );
  BUF_X1 U246 ( .A(n4925), .Z(n629) );
  BUF_X1 U247 ( .A(n4928), .Z(n620) );
  BUF_X1 U248 ( .A(n4934), .Z(n605) );
  BUF_X1 U249 ( .A(n4953), .Z(n476) );
  BUF_X1 U250 ( .A(n4956), .Z(n467) );
  BUF_X1 U251 ( .A(n4959), .Z(n458) );
  BUF_X1 U252 ( .A(n4965), .Z(n443) );
  BUF_X1 U253 ( .A(n4984), .Z(n58) );
  BUF_X1 U254 ( .A(n4987), .Z(n49) );
  BUF_X1 U255 ( .A(n3451), .Z(n1407) );
  BUF_X1 U256 ( .A(n3454), .Z(n1398) );
  BUF_X1 U257 ( .A(n3460), .Z(n1383) );
  BUF_X1 U258 ( .A(n3479), .Z(n1350) );
  BUF_X1 U259 ( .A(n3482), .Z(n1341) );
  BUF_X1 U260 ( .A(n3485), .Z(n1332) );
  BUF_X1 U261 ( .A(n3491), .Z(n1317) );
  BUF_X1 U262 ( .A(n3510), .Z(n1188) );
  BUF_X1 U263 ( .A(n3513), .Z(n1179) );
  BUF_X1 U264 ( .A(n3516), .Z(n1170) );
  BUF_X1 U265 ( .A(n3522), .Z(n1155) );
  BUF_X1 U266 ( .A(n3541), .Z(n770) );
  BUF_X1 U267 ( .A(n3544), .Z(n761) );
  BUF_X1 U268 ( .A(n4894), .Z(n696) );
  BUF_X1 U269 ( .A(n4897), .Z(n687) );
  BUF_X1 U270 ( .A(n4903), .Z(n672) );
  BUF_X1 U271 ( .A(n4922), .Z(n639) );
  BUF_X1 U272 ( .A(n4925), .Z(n630) );
  BUF_X1 U273 ( .A(n4928), .Z(n621) );
  BUF_X1 U274 ( .A(n4934), .Z(n606) );
  BUF_X1 U275 ( .A(n4953), .Z(n477) );
  BUF_X1 U276 ( .A(n4956), .Z(n468) );
  BUF_X1 U277 ( .A(n4959), .Z(n459) );
  BUF_X1 U278 ( .A(n4965), .Z(n444) );
  BUF_X1 U279 ( .A(n4984), .Z(n59) );
  BUF_X1 U280 ( .A(n4987), .Z(n50) );
  BUF_X1 U281 ( .A(n3451), .Z(n1408) );
  BUF_X1 U282 ( .A(n3454), .Z(n1399) );
  BUF_X1 U283 ( .A(n3460), .Z(n1384) );
  BUF_X1 U284 ( .A(n3479), .Z(n1351) );
  BUF_X1 U285 ( .A(n3482), .Z(n1342) );
  BUF_X1 U286 ( .A(n3485), .Z(n1333) );
  BUF_X1 U287 ( .A(n3491), .Z(n1318) );
  BUF_X1 U288 ( .A(n3510), .Z(n1189) );
  BUF_X1 U289 ( .A(n3513), .Z(n1180) );
  BUF_X1 U290 ( .A(n3516), .Z(n1171) );
  BUF_X1 U291 ( .A(n3522), .Z(n1156) );
  BUF_X1 U292 ( .A(n3541), .Z(n771) );
  BUF_X1 U293 ( .A(n3544), .Z(n762) );
  BUF_X1 U294 ( .A(n4980), .Z(n72) );
  BUF_X1 U295 ( .A(n3537), .Z(n1136) );
  BUF_X1 U296 ( .A(n4918), .Z(n652) );
  BUF_X1 U297 ( .A(n3475), .Z(n1364) );
  BUF_X1 U298 ( .A(n4949), .Z(n490) );
  BUF_X1 U299 ( .A(n3506), .Z(n1298) );
  BUF_X1 U300 ( .A(n4905), .Z(n666) );
  BUF_X1 U301 ( .A(n4908), .Z(n657) );
  BUF_X1 U302 ( .A(n4936), .Z(n600) );
  BUF_X1 U303 ( .A(n4939), .Z(n495) );
  BUF_X1 U304 ( .A(n4967), .Z(n438) );
  BUF_X1 U305 ( .A(n4970), .Z(n77) );
  BUF_X1 U306 ( .A(n4998), .Z(n20) );
  BUF_X1 U307 ( .A(n5001), .Z(n9) );
  BUF_X1 U308 ( .A(n3462), .Z(n1378) );
  BUF_X1 U309 ( .A(n3465), .Z(n1369) );
  BUF_X1 U310 ( .A(n3493), .Z(n1312) );
  BUF_X1 U311 ( .A(n3496), .Z(n1303) );
  BUF_X1 U312 ( .A(n3524), .Z(n1150) );
  BUF_X1 U313 ( .A(n3527), .Z(n1141) );
  BUF_X1 U314 ( .A(n3555), .Z(n732) );
  BUF_X1 U315 ( .A(n3558), .Z(n723) );
  BUF_X1 U316 ( .A(n4905), .Z(n665) );
  BUF_X1 U317 ( .A(n4908), .Z(n656) );
  BUF_X1 U318 ( .A(n4936), .Z(n599) );
  BUF_X1 U319 ( .A(n4939), .Z(n494) );
  BUF_X1 U320 ( .A(n4967), .Z(n437) );
  BUF_X1 U321 ( .A(n4970), .Z(n76) );
  BUF_X1 U322 ( .A(n4998), .Z(n19) );
  BUF_X1 U323 ( .A(n5001), .Z(n8) );
  BUF_X1 U324 ( .A(n3462), .Z(n1377) );
  BUF_X1 U325 ( .A(n3465), .Z(n1368) );
  BUF_X1 U326 ( .A(n3493), .Z(n1311) );
  BUF_X1 U327 ( .A(n3496), .Z(n1302) );
  BUF_X1 U328 ( .A(n3524), .Z(n1149) );
  BUF_X1 U329 ( .A(n3527), .Z(n1140) );
  BUF_X1 U330 ( .A(n3555), .Z(n731) );
  BUF_X1 U331 ( .A(n3558), .Z(n722) );
  BUF_X1 U332 ( .A(n4889), .Z(n710) );
  BUF_X1 U333 ( .A(n3446), .Z(n1422) );
  BUF_X1 U334 ( .A(n4889), .Z(n711) );
  BUF_X1 U335 ( .A(n3446), .Z(n1423) );
  BUF_X1 U336 ( .A(n4985), .Z(n55) );
  BUF_X1 U337 ( .A(n4988), .Z(n46) );
  BUF_X1 U338 ( .A(n3542), .Z(n767) );
  BUF_X1 U339 ( .A(n3545), .Z(n758) );
  BUF_X1 U340 ( .A(n4985), .Z(n56) );
  BUF_X1 U341 ( .A(n4988), .Z(n47) );
  BUF_X1 U342 ( .A(n3542), .Z(n768) );
  BUF_X1 U343 ( .A(n3545), .Z(n759) );
  BUF_X1 U344 ( .A(n4892), .Z(n701) );
  BUF_X1 U345 ( .A(n3449), .Z(n1413) );
  BUF_X1 U346 ( .A(n4892), .Z(n702) );
  BUF_X1 U347 ( .A(n3449), .Z(n1414) );
  BUF_X1 U348 ( .A(n4895), .Z(n692) );
  BUF_X1 U349 ( .A(n4901), .Z(n677) );
  BUF_X1 U350 ( .A(n4920), .Z(n644) );
  BUF_X1 U351 ( .A(n4923), .Z(n635) );
  BUF_X1 U352 ( .A(n4926), .Z(n626) );
  BUF_X1 U353 ( .A(n4932), .Z(n611) );
  BUF_X1 U354 ( .A(n4951), .Z(n482) );
  BUF_X1 U355 ( .A(n4954), .Z(n473) );
  BUF_X1 U356 ( .A(n4963), .Z(n449) );
  BUF_X1 U357 ( .A(n4982), .Z(n64) );
  BUF_X1 U358 ( .A(n4994), .Z(n31) );
  BUF_X1 U359 ( .A(n3452), .Z(n1404) );
  BUF_X1 U360 ( .A(n3458), .Z(n1389) );
  BUF_X1 U361 ( .A(n3477), .Z(n1356) );
  BUF_X1 U362 ( .A(n3480), .Z(n1347) );
  BUF_X1 U363 ( .A(n3483), .Z(n1338) );
  BUF_X1 U364 ( .A(n3489), .Z(n1323) );
  BUF_X1 U365 ( .A(n3508), .Z(n1194) );
  BUF_X1 U366 ( .A(n3511), .Z(n1185) );
  BUF_X1 U367 ( .A(n3520), .Z(n1161) );
  BUF_X1 U368 ( .A(n3539), .Z(n776) );
  BUF_X1 U369 ( .A(n3551), .Z(n743) );
  BUF_X1 U370 ( .A(n4895), .Z(n693) );
  BUF_X1 U371 ( .A(n4901), .Z(n678) );
  BUF_X1 U372 ( .A(n4920), .Z(n645) );
  BUF_X1 U373 ( .A(n4923), .Z(n636) );
  BUF_X1 U374 ( .A(n4926), .Z(n627) );
  BUF_X1 U375 ( .A(n4932), .Z(n612) );
  BUF_X1 U376 ( .A(n4951), .Z(n483) );
  BUF_X1 U377 ( .A(n4954), .Z(n474) );
  BUF_X1 U378 ( .A(n4963), .Z(n450) );
  BUF_X1 U379 ( .A(n4982), .Z(n65) );
  BUF_X1 U380 ( .A(n4994), .Z(n32) );
  BUF_X1 U381 ( .A(n3452), .Z(n1405) );
  BUF_X1 U382 ( .A(n3458), .Z(n1390) );
  BUF_X1 U383 ( .A(n3477), .Z(n1357) );
  BUF_X1 U384 ( .A(n3480), .Z(n1348) );
  BUF_X1 U385 ( .A(n3483), .Z(n1339) );
  BUF_X1 U386 ( .A(n3489), .Z(n1324) );
  BUF_X1 U387 ( .A(n3508), .Z(n1195) );
  BUF_X1 U388 ( .A(n3511), .Z(n1186) );
  BUF_X1 U389 ( .A(n3520), .Z(n1162) );
  BUF_X1 U390 ( .A(n3539), .Z(n777) );
  BUF_X1 U391 ( .A(n3551), .Z(n744) );
  BUF_X1 U392 ( .A(n4986), .Z(n52) );
  BUF_X1 U393 ( .A(n4989), .Z(n43) );
  BUF_X1 U394 ( .A(n3543), .Z(n764) );
  BUF_X1 U395 ( .A(n3546), .Z(n755) );
  BUF_X1 U396 ( .A(n4986), .Z(n53) );
  BUF_X1 U397 ( .A(n4989), .Z(n44) );
  BUF_X1 U398 ( .A(n3543), .Z(n765) );
  BUF_X1 U399 ( .A(n3546), .Z(n756) );
  BUF_X1 U400 ( .A(n4890), .Z(n707) );
  BUF_X1 U401 ( .A(n4893), .Z(n698) );
  BUF_X1 U402 ( .A(n4983), .Z(n61) );
  BUF_X1 U403 ( .A(n3540), .Z(n773) );
  BUF_X1 U404 ( .A(n4893), .Z(n699) );
  BUF_X1 U405 ( .A(n4983), .Z(n62) );
  BUF_X1 U406 ( .A(n3540), .Z(n774) );
  BUF_X1 U407 ( .A(n4896), .Z(n689) );
  BUF_X1 U408 ( .A(n4902), .Z(n674) );
  BUF_X1 U409 ( .A(n4921), .Z(n641) );
  BUF_X1 U410 ( .A(n4924), .Z(n632) );
  BUF_X1 U411 ( .A(n4933), .Z(n608) );
  BUF_X1 U412 ( .A(n4952), .Z(n479) );
  BUF_X1 U413 ( .A(n4955), .Z(n470) );
  BUF_X1 U414 ( .A(n4958), .Z(n461) );
  BUF_X1 U415 ( .A(n3447), .Z(n1419) );
  BUF_X1 U416 ( .A(n3450), .Z(n1410) );
  BUF_X1 U417 ( .A(n3453), .Z(n1401) );
  BUF_X1 U418 ( .A(n3459), .Z(n1386) );
  BUF_X1 U419 ( .A(n3478), .Z(n1353) );
  BUF_X1 U420 ( .A(n3481), .Z(n1344) );
  BUF_X1 U421 ( .A(n3490), .Z(n1320) );
  BUF_X1 U422 ( .A(n3509), .Z(n1191) );
  BUF_X1 U423 ( .A(n3512), .Z(n1182) );
  BUF_X1 U424 ( .A(n3515), .Z(n1173) );
  BUF_X1 U425 ( .A(n4890), .Z(n708) );
  BUF_X1 U426 ( .A(n4896), .Z(n690) );
  BUF_X1 U427 ( .A(n4902), .Z(n675) );
  BUF_X1 U428 ( .A(n4921), .Z(n642) );
  BUF_X1 U429 ( .A(n4924), .Z(n633) );
  BUF_X1 U430 ( .A(n4933), .Z(n609) );
  BUF_X1 U431 ( .A(n4952), .Z(n480) );
  BUF_X1 U432 ( .A(n4955), .Z(n471) );
  BUF_X1 U433 ( .A(n4958), .Z(n462) );
  BUF_X1 U434 ( .A(n3447), .Z(n1420) );
  BUF_X1 U435 ( .A(n3450), .Z(n1411) );
  BUF_X1 U436 ( .A(n3453), .Z(n1402) );
  BUF_X1 U437 ( .A(n3459), .Z(n1387) );
  BUF_X1 U438 ( .A(n3478), .Z(n1354) );
  BUF_X1 U439 ( .A(n3481), .Z(n1345) );
  BUF_X1 U440 ( .A(n3490), .Z(n1321) );
  BUF_X1 U441 ( .A(n3509), .Z(n1192) );
  BUF_X1 U442 ( .A(n3512), .Z(n1183) );
  BUF_X1 U443 ( .A(n3515), .Z(n1174) );
  BUF_X1 U444 ( .A(n4919), .Z(n649) );
  BUF_X1 U445 ( .A(n3476), .Z(n1361) );
  BUF_X1 U446 ( .A(n4950), .Z(n487) );
  BUF_X1 U447 ( .A(n4981), .Z(n69) );
  BUF_X1 U448 ( .A(n3538), .Z(n781) );
  BUF_X1 U449 ( .A(n3507), .Z(n1199) );
  BUF_X1 U450 ( .A(n4906), .Z(n663) );
  BUF_X1 U451 ( .A(n4937), .Z(n597) );
  BUF_X1 U452 ( .A(n4940), .Z(n492) );
  BUF_X1 U453 ( .A(n4968), .Z(n435) );
  BUF_X1 U454 ( .A(n4971), .Z(n74) );
  BUF_X1 U455 ( .A(n4999), .Z(n16) );
  BUF_X1 U456 ( .A(n5002), .Z(n5) );
  BUF_X1 U457 ( .A(n3463), .Z(n1375) );
  BUF_X1 U458 ( .A(n3494), .Z(n1309) );
  BUF_X1 U459 ( .A(n3497), .Z(n1300) );
  BUF_X1 U460 ( .A(n3525), .Z(n1147) );
  BUF_X1 U461 ( .A(n3528), .Z(n1138) );
  BUF_X1 U462 ( .A(n3556), .Z(n729) );
  BUF_X1 U463 ( .A(n3559), .Z(n720) );
  BUF_X1 U464 ( .A(n4906), .Z(n662) );
  BUF_X1 U465 ( .A(n4937), .Z(n596) );
  BUF_X1 U466 ( .A(n4940), .Z(n491) );
  BUF_X1 U467 ( .A(n4968), .Z(n434) );
  BUF_X1 U468 ( .A(n4971), .Z(n73) );
  BUF_X1 U469 ( .A(n4999), .Z(n15) );
  BUF_X1 U470 ( .A(n5002), .Z(n4) );
  BUF_X1 U471 ( .A(n3463), .Z(n1374) );
  BUF_X1 U472 ( .A(n3494), .Z(n1308) );
  BUF_X1 U473 ( .A(n3497), .Z(n1299) );
  BUF_X1 U474 ( .A(n3525), .Z(n1146) );
  BUF_X1 U475 ( .A(n3528), .Z(n1137) );
  BUF_X1 U476 ( .A(n3556), .Z(n728) );
  BUF_X1 U477 ( .A(n3559), .Z(n719) );
  BUF_X1 U478 ( .A(n4898), .Z(n685) );
  BUF_X1 U479 ( .A(n4929), .Z(n619) );
  BUF_X1 U480 ( .A(n4960), .Z(n457) );
  BUF_X1 U481 ( .A(n4991), .Z(n39) );
  BUF_X1 U482 ( .A(n3455), .Z(n1397) );
  BUF_X1 U483 ( .A(n3486), .Z(n1331) );
  BUF_X1 U484 ( .A(n3517), .Z(n1169) );
  BUF_X1 U485 ( .A(n3548), .Z(n751) );
  BUF_X1 U486 ( .A(n4904), .Z(n670) );
  BUF_X1 U487 ( .A(n4907), .Z(n661) );
  BUF_X1 U488 ( .A(n4935), .Z(n604) );
  BUF_X1 U489 ( .A(n4938), .Z(n595) );
  BUF_X1 U490 ( .A(n4966), .Z(n442) );
  BUF_X1 U491 ( .A(n4969), .Z(n433) );
  BUF_X1 U492 ( .A(n4997), .Z(n24) );
  BUF_X1 U493 ( .A(n5000), .Z(n14) );
  BUF_X1 U494 ( .A(n3461), .Z(n1382) );
  BUF_X1 U495 ( .A(n3464), .Z(n1373) );
  BUF_X1 U496 ( .A(n3492), .Z(n1316) );
  BUF_X1 U497 ( .A(n3495), .Z(n1307) );
  BUF_X1 U498 ( .A(n3523), .Z(n1154) );
  BUF_X1 U499 ( .A(n3526), .Z(n1145) );
  BUF_X1 U500 ( .A(n3554), .Z(n736) );
  BUF_X1 U501 ( .A(n3557), .Z(n727) );
  BUF_X1 U502 ( .A(n4899), .Z(n682) );
  BUF_X1 U503 ( .A(n4930), .Z(n616) );
  BUF_X1 U504 ( .A(n4961), .Z(n454) );
  BUF_X1 U505 ( .A(n4992), .Z(n36) );
  BUF_X1 U506 ( .A(n3456), .Z(n1394) );
  BUF_X1 U507 ( .A(n3487), .Z(n1328) );
  BUF_X1 U508 ( .A(n3518), .Z(n1166) );
  BUF_X1 U509 ( .A(n3549), .Z(n748) );
  BUF_X1 U510 ( .A(n3103), .Z(n1744) );
  BUF_X1 U511 ( .A(n3103), .Z(n1743) );
  BUF_X1 U512 ( .A(n3098), .Z(n1747) );
  BUF_X1 U513 ( .A(n3098), .Z(n1746) );
  BUF_X1 U514 ( .A(n3093), .Z(n1750) );
  BUF_X1 U515 ( .A(n3093), .Z(n1749) );
  BUF_X1 U516 ( .A(n3088), .Z(n1753) );
  BUF_X1 U517 ( .A(n3088), .Z(n1752) );
  BUF_X1 U518 ( .A(n3083), .Z(n1756) );
  BUF_X1 U519 ( .A(n3083), .Z(n1755) );
  BUF_X1 U520 ( .A(n3078), .Z(n1759) );
  BUF_X1 U521 ( .A(n3078), .Z(n1758) );
  BUF_X1 U522 ( .A(n3073), .Z(n1762) );
  BUF_X1 U523 ( .A(n3073), .Z(n1761) );
  BUF_X1 U524 ( .A(n3068), .Z(n1765) );
  BUF_X1 U525 ( .A(n3068), .Z(n1764) );
  BUF_X1 U526 ( .A(n3063), .Z(n1768) );
  BUF_X1 U527 ( .A(n3063), .Z(n1767) );
  BUF_X1 U528 ( .A(n3058), .Z(n1771) );
  BUF_X1 U529 ( .A(n3058), .Z(n1770) );
  BUF_X1 U530 ( .A(n3053), .Z(n1774) );
  BUF_X1 U531 ( .A(n3053), .Z(n1773) );
  BUF_X1 U532 ( .A(n3048), .Z(n1777) );
  BUF_X1 U533 ( .A(n3048), .Z(n1776) );
  BUF_X1 U534 ( .A(n3043), .Z(n1780) );
  BUF_X1 U535 ( .A(n3043), .Z(n1779) );
  BUF_X1 U536 ( .A(n3038), .Z(n1783) );
  BUF_X1 U537 ( .A(n3038), .Z(n1782) );
  BUF_X1 U538 ( .A(n3033), .Z(n1786) );
  BUF_X1 U539 ( .A(n3033), .Z(n1785) );
  BUF_X1 U540 ( .A(n2996), .Z(n1789) );
  BUF_X1 U541 ( .A(n2996), .Z(n1788) );
  BUF_X1 U542 ( .A(n3303), .Z(n1504) );
  BUF_X1 U543 ( .A(n3303), .Z(n1503) );
  BUF_X1 U544 ( .A(n3299), .Z(n1507) );
  BUF_X1 U545 ( .A(n3299), .Z(n1506) );
  BUF_X1 U546 ( .A(n3295), .Z(n1510) );
  BUF_X1 U547 ( .A(n3295), .Z(n1509) );
  BUF_X1 U548 ( .A(n3291), .Z(n1513) );
  BUF_X1 U549 ( .A(n3291), .Z(n1512) );
  BUF_X1 U550 ( .A(n3287), .Z(n1516) );
  BUF_X1 U551 ( .A(n3287), .Z(n1515) );
  BUF_X1 U552 ( .A(n3283), .Z(n1519) );
  BUF_X1 U553 ( .A(n3283), .Z(n1518) );
  BUF_X1 U554 ( .A(n3279), .Z(n1522) );
  BUF_X1 U555 ( .A(n3279), .Z(n1521) );
  BUF_X1 U556 ( .A(n3275), .Z(n1525) );
  BUF_X1 U557 ( .A(n3275), .Z(n1524) );
  BUF_X1 U558 ( .A(n3271), .Z(n1528) );
  BUF_X1 U559 ( .A(n3271), .Z(n1527) );
  BUF_X1 U560 ( .A(n3267), .Z(n1531) );
  BUF_X1 U561 ( .A(n3267), .Z(n1530) );
  BUF_X1 U562 ( .A(n3263), .Z(n1534) );
  BUF_X1 U563 ( .A(n3263), .Z(n1533) );
  BUF_X1 U564 ( .A(n3259), .Z(n1537) );
  BUF_X1 U565 ( .A(n3259), .Z(n1536) );
  BUF_X1 U566 ( .A(n3255), .Z(n1540) );
  BUF_X1 U567 ( .A(n3255), .Z(n1539) );
  BUF_X1 U568 ( .A(n3251), .Z(n1543) );
  BUF_X1 U569 ( .A(n3251), .Z(n1542) );
  BUF_X1 U570 ( .A(n3247), .Z(n1546) );
  BUF_X1 U571 ( .A(n3247), .Z(n1545) );
  BUF_X1 U572 ( .A(n3242), .Z(n1549) );
  BUF_X1 U573 ( .A(n3242), .Z(n1548) );
  BUF_X1 U574 ( .A(n3238), .Z(n1648) );
  BUF_X1 U575 ( .A(n3238), .Z(n1551) );
  BUF_X1 U576 ( .A(n3234), .Z(n1651) );
  BUF_X1 U577 ( .A(n3234), .Z(n1650) );
  BUF_X1 U578 ( .A(n3230), .Z(n1654) );
  BUF_X1 U579 ( .A(n3230), .Z(n1653) );
  BUF_X1 U580 ( .A(n3226), .Z(n1657) );
  BUF_X1 U581 ( .A(n3226), .Z(n1656) );
  BUF_X1 U582 ( .A(n3222), .Z(n1660) );
  BUF_X1 U583 ( .A(n3222), .Z(n1659) );
  BUF_X1 U584 ( .A(n3218), .Z(n1663) );
  BUF_X1 U585 ( .A(n3218), .Z(n1662) );
  BUF_X1 U586 ( .A(n3214), .Z(n1666) );
  BUF_X1 U587 ( .A(n3214), .Z(n1665) );
  BUF_X1 U588 ( .A(n3210), .Z(n1669) );
  BUF_X1 U589 ( .A(n3210), .Z(n1668) );
  BUF_X1 U590 ( .A(n3206), .Z(n1672) );
  BUF_X1 U591 ( .A(n3206), .Z(n1671) );
  BUF_X1 U592 ( .A(n3202), .Z(n1675) );
  BUF_X1 U593 ( .A(n3202), .Z(n1674) );
  BUF_X1 U594 ( .A(n3198), .Z(n1678) );
  BUF_X1 U595 ( .A(n3198), .Z(n1677) );
  BUF_X1 U596 ( .A(n3194), .Z(n1681) );
  BUF_X1 U597 ( .A(n3194), .Z(n1680) );
  BUF_X1 U598 ( .A(n3190), .Z(n1684) );
  BUF_X1 U599 ( .A(n3190), .Z(n1683) );
  BUF_X1 U600 ( .A(n3186), .Z(n1687) );
  BUF_X1 U601 ( .A(n3186), .Z(n1686) );
  BUF_X1 U602 ( .A(n3182), .Z(n1690) );
  BUF_X1 U603 ( .A(n3182), .Z(n1689) );
  BUF_X1 U604 ( .A(n3177), .Z(n1693) );
  BUF_X1 U605 ( .A(n3177), .Z(n1692) );
  BUF_X1 U606 ( .A(n3173), .Z(n1696) );
  BUF_X1 U607 ( .A(n3173), .Z(n1695) );
  BUF_X1 U608 ( .A(n3169), .Z(n1699) );
  BUF_X1 U609 ( .A(n3169), .Z(n1698) );
  BUF_X1 U610 ( .A(n3165), .Z(n1702) );
  BUF_X1 U611 ( .A(n3165), .Z(n1701) );
  BUF_X1 U612 ( .A(n3161), .Z(n1705) );
  BUF_X1 U613 ( .A(n3161), .Z(n1704) );
  BUF_X1 U614 ( .A(n3157), .Z(n1708) );
  BUF_X1 U615 ( .A(n3157), .Z(n1707) );
  BUF_X1 U616 ( .A(n3153), .Z(n1711) );
  BUF_X1 U617 ( .A(n3153), .Z(n1710) );
  BUF_X1 U618 ( .A(n3149), .Z(n1714) );
  BUF_X1 U619 ( .A(n3149), .Z(n1713) );
  BUF_X1 U620 ( .A(n3145), .Z(n1717) );
  BUF_X1 U621 ( .A(n3145), .Z(n1716) );
  BUF_X1 U622 ( .A(n3141), .Z(n1720) );
  BUF_X1 U623 ( .A(n3141), .Z(n1719) );
  BUF_X1 U624 ( .A(n3137), .Z(n1723) );
  BUF_X1 U625 ( .A(n3137), .Z(n1722) );
  BUF_X1 U626 ( .A(n3133), .Z(n1726) );
  BUF_X1 U627 ( .A(n3133), .Z(n1725) );
  BUF_X1 U628 ( .A(n3129), .Z(n1729) );
  BUF_X1 U629 ( .A(n3129), .Z(n1728) );
  BUF_X1 U630 ( .A(n3125), .Z(n1732) );
  BUF_X1 U631 ( .A(n3125), .Z(n1731) );
  BUF_X1 U632 ( .A(n3121), .Z(n1735) );
  BUF_X1 U633 ( .A(n3121), .Z(n1734) );
  BUF_X1 U634 ( .A(n3117), .Z(n1738) );
  BUF_X1 U635 ( .A(n3117), .Z(n1737) );
  BUF_X1 U636 ( .A(n3112), .Z(n1741) );
  BUF_X1 U637 ( .A(n3112), .Z(n1740) );
  BUF_X1 U638 ( .A(n3375), .Z(n1456) );
  BUF_X1 U639 ( .A(n3375), .Z(n1455) );
  BUF_X1 U640 ( .A(n3371), .Z(n1459) );
  BUF_X1 U641 ( .A(n3371), .Z(n1458) );
  BUF_X1 U642 ( .A(n3367), .Z(n1462) );
  BUF_X1 U643 ( .A(n3367), .Z(n1461) );
  BUF_X1 U644 ( .A(n3362), .Z(n1465) );
  BUF_X1 U645 ( .A(n3362), .Z(n1464) );
  BUF_X1 U646 ( .A(n3356), .Z(n1468) );
  BUF_X1 U647 ( .A(n3356), .Z(n1467) );
  BUF_X1 U648 ( .A(n3351), .Z(n1471) );
  BUF_X1 U649 ( .A(n3351), .Z(n1470) );
  BUF_X1 U650 ( .A(n3346), .Z(n1474) );
  BUF_X1 U651 ( .A(n3346), .Z(n1473) );
  BUF_X1 U652 ( .A(n3340), .Z(n1477) );
  BUF_X1 U653 ( .A(n3340), .Z(n1476) );
  BUF_X1 U654 ( .A(n3336), .Z(n1480) );
  BUF_X1 U655 ( .A(n3336), .Z(n1479) );
  BUF_X1 U656 ( .A(n3332), .Z(n1483) );
  BUF_X1 U657 ( .A(n3332), .Z(n1482) );
  BUF_X1 U658 ( .A(n3328), .Z(n1486) );
  BUF_X1 U659 ( .A(n3328), .Z(n1485) );
  BUF_X1 U660 ( .A(n3324), .Z(n1489) );
  BUF_X1 U661 ( .A(n3324), .Z(n1488) );
  BUF_X1 U662 ( .A(n3320), .Z(n1492) );
  BUF_X1 U663 ( .A(n3320), .Z(n1491) );
  BUF_X1 U664 ( .A(n3316), .Z(n1495) );
  BUF_X1 U665 ( .A(n3316), .Z(n1494) );
  BUF_X1 U666 ( .A(n3312), .Z(n1498) );
  BUF_X1 U667 ( .A(n3312), .Z(n1497) );
  BUF_X1 U668 ( .A(n3307), .Z(n1501) );
  BUF_X1 U669 ( .A(n3307), .Z(n1500) );
  BUF_X1 U670 ( .A(n3413), .Z(n1432) );
  BUF_X1 U671 ( .A(n3413), .Z(n1431) );
  BUF_X1 U672 ( .A(n3409), .Z(n1435) );
  BUF_X1 U673 ( .A(n3409), .Z(n1434) );
  BUF_X1 U674 ( .A(n3403), .Z(n1438) );
  BUF_X1 U675 ( .A(n3403), .Z(n1437) );
  BUF_X1 U676 ( .A(n3398), .Z(n1441) );
  BUF_X1 U677 ( .A(n3398), .Z(n1440) );
  BUF_X1 U678 ( .A(n3394), .Z(n1444) );
  BUF_X1 U679 ( .A(n3394), .Z(n1443) );
  BUF_X1 U680 ( .A(n3390), .Z(n1447) );
  BUF_X1 U681 ( .A(n3390), .Z(n1446) );
  BUF_X1 U682 ( .A(n3386), .Z(n1450) );
  BUF_X1 U683 ( .A(n3386), .Z(n1449) );
  BUF_X1 U684 ( .A(n3380), .Z(n1453) );
  BUF_X1 U685 ( .A(n3380), .Z(n1452) );
  BUF_X1 U686 ( .A(n4891), .Z(n706) );
  BUF_X1 U687 ( .A(n3448), .Z(n1418) );
  BUF_X1 U688 ( .A(n4990), .Z(n42) );
  BUF_X1 U689 ( .A(n4996), .Z(n27) );
  BUF_X1 U690 ( .A(n3547), .Z(n754) );
  BUF_X1 U691 ( .A(n3553), .Z(n739) );
  BUF_X1 U692 ( .A(n4894), .Z(n697) );
  BUF_X1 U693 ( .A(n4984), .Z(n60) );
  BUF_X1 U694 ( .A(n3451), .Z(n1409) );
  BUF_X1 U695 ( .A(n3541), .Z(n772) );
  BUF_X1 U696 ( .A(n4897), .Z(n688) );
  BUF_X1 U697 ( .A(n4903), .Z(n673) );
  BUF_X1 U698 ( .A(n4922), .Z(n640) );
  BUF_X1 U699 ( .A(n4925), .Z(n631) );
  BUF_X1 U700 ( .A(n4928), .Z(n622) );
  BUF_X1 U701 ( .A(n4934), .Z(n607) );
  BUF_X1 U702 ( .A(n4953), .Z(n478) );
  BUF_X1 U703 ( .A(n4956), .Z(n469) );
  BUF_X1 U704 ( .A(n4959), .Z(n460) );
  BUF_X1 U705 ( .A(n4965), .Z(n445) );
  BUF_X1 U706 ( .A(n4987), .Z(n51) );
  BUF_X1 U707 ( .A(n3454), .Z(n1400) );
  BUF_X1 U708 ( .A(n3460), .Z(n1385) );
  BUF_X1 U709 ( .A(n3479), .Z(n1352) );
  BUF_X1 U710 ( .A(n3482), .Z(n1343) );
  BUF_X1 U711 ( .A(n3485), .Z(n1334) );
  BUF_X1 U712 ( .A(n3491), .Z(n1319) );
  BUF_X1 U713 ( .A(n3510), .Z(n1190) );
  BUF_X1 U714 ( .A(n3513), .Z(n1181) );
  BUF_X1 U715 ( .A(n3516), .Z(n1172) );
  BUF_X1 U716 ( .A(n3522), .Z(n1157) );
  BUF_X1 U717 ( .A(n3544), .Z(n763) );
  BUF_X1 U718 ( .A(n4905), .Z(n667) );
  BUF_X1 U719 ( .A(n4908), .Z(n658) );
  BUF_X1 U720 ( .A(n4936), .Z(n601) );
  BUF_X1 U721 ( .A(n4939), .Z(n592) );
  BUF_X1 U722 ( .A(n4967), .Z(n439) );
  BUF_X1 U723 ( .A(n4970), .Z(n78) );
  BUF_X1 U724 ( .A(n4998), .Z(n21) );
  BUF_X1 U725 ( .A(n5001), .Z(n10) );
  BUF_X1 U726 ( .A(n3462), .Z(n1379) );
  BUF_X1 U727 ( .A(n3465), .Z(n1370) );
  BUF_X1 U728 ( .A(n3493), .Z(n1313) );
  BUF_X1 U729 ( .A(n3496), .Z(n1304) );
  BUF_X1 U730 ( .A(n3524), .Z(n1151) );
  BUF_X1 U731 ( .A(n3527), .Z(n1142) );
  BUF_X1 U732 ( .A(n3555), .Z(n733) );
  BUF_X1 U733 ( .A(n3558), .Z(n724) );
  BUF_X1 U734 ( .A(n4889), .Z(n712) );
  BUF_X1 U735 ( .A(n3446), .Z(n1424) );
  BUF_X1 U736 ( .A(n4985), .Z(n57) );
  BUF_X1 U737 ( .A(n4988), .Z(n48) );
  BUF_X1 U738 ( .A(n3542), .Z(n769) );
  BUF_X1 U739 ( .A(n3545), .Z(n760) );
  BUF_X1 U740 ( .A(n4892), .Z(n703) );
  BUF_X1 U741 ( .A(n3449), .Z(n1415) );
  BUF_X1 U742 ( .A(n4932), .Z(n613) );
  BUF_X1 U743 ( .A(n3489), .Z(n1325) );
  BUF_X1 U744 ( .A(n4895), .Z(n694) );
  BUF_X1 U745 ( .A(n4901), .Z(n679) );
  BUF_X1 U746 ( .A(n4920), .Z(n646) );
  BUF_X1 U747 ( .A(n4923), .Z(n637) );
  BUF_X1 U748 ( .A(n4926), .Z(n628) );
  BUF_X1 U749 ( .A(n4951), .Z(n484) );
  BUF_X1 U750 ( .A(n4954), .Z(n475) );
  BUF_X1 U751 ( .A(n4963), .Z(n451) );
  BUF_X1 U752 ( .A(n4982), .Z(n66) );
  BUF_X1 U753 ( .A(n3539), .Z(n778) );
  BUF_X1 U754 ( .A(n4994), .Z(n33) );
  BUF_X1 U755 ( .A(n3452), .Z(n1406) );
  BUF_X1 U756 ( .A(n3458), .Z(n1391) );
  BUF_X1 U757 ( .A(n3477), .Z(n1358) );
  BUF_X1 U758 ( .A(n3480), .Z(n1349) );
  BUF_X1 U759 ( .A(n3483), .Z(n1340) );
  BUF_X1 U760 ( .A(n3508), .Z(n1196) );
  BUF_X1 U761 ( .A(n3511), .Z(n1187) );
  BUF_X1 U762 ( .A(n3520), .Z(n1163) );
  BUF_X1 U763 ( .A(n3551), .Z(n745) );
  BUF_X1 U764 ( .A(n4986), .Z(n54) );
  BUF_X1 U765 ( .A(n4989), .Z(n45) );
  BUF_X1 U766 ( .A(n3543), .Z(n766) );
  BUF_X1 U767 ( .A(n3546), .Z(n757) );
  BUF_X1 U768 ( .A(n4893), .Z(n700) );
  BUF_X1 U769 ( .A(n4983), .Z(n63) );
  BUF_X1 U770 ( .A(n3450), .Z(n1412) );
  BUF_X1 U771 ( .A(n3540), .Z(n775) );
  BUF_X1 U772 ( .A(n4890), .Z(n709) );
  BUF_X1 U773 ( .A(n3447), .Z(n1421) );
  BUF_X1 U774 ( .A(n4896), .Z(n691) );
  BUF_X1 U775 ( .A(n4902), .Z(n676) );
  BUF_X1 U776 ( .A(n4921), .Z(n643) );
  BUF_X1 U777 ( .A(n4924), .Z(n634) );
  BUF_X1 U778 ( .A(n4933), .Z(n610) );
  BUF_X1 U779 ( .A(n4952), .Z(n481) );
  BUF_X1 U780 ( .A(n4955), .Z(n472) );
  BUF_X1 U781 ( .A(n4958), .Z(n463) );
  BUF_X1 U782 ( .A(n3453), .Z(n1403) );
  BUF_X1 U783 ( .A(n3459), .Z(n1388) );
  BUF_X1 U784 ( .A(n3478), .Z(n1355) );
  BUF_X1 U785 ( .A(n3481), .Z(n1346) );
  BUF_X1 U786 ( .A(n3490), .Z(n1322) );
  BUF_X1 U787 ( .A(n3509), .Z(n1193) );
  BUF_X1 U788 ( .A(n3512), .Z(n1184) );
  BUF_X1 U789 ( .A(n3515), .Z(n1175) );
  BUF_X1 U790 ( .A(n5002), .Z(n6) );
  BUF_X1 U791 ( .A(n3559), .Z(n721) );
  BUF_X1 U792 ( .A(n4906), .Z(n664) );
  BUF_X1 U793 ( .A(n4937), .Z(n598) );
  BUF_X1 U794 ( .A(n4940), .Z(n493) );
  BUF_X1 U795 ( .A(n4968), .Z(n436) );
  BUF_X1 U796 ( .A(n4971), .Z(n75) );
  BUF_X1 U797 ( .A(n4999), .Z(n18) );
  BUF_X1 U798 ( .A(n3463), .Z(n1376) );
  BUF_X1 U799 ( .A(n3494), .Z(n1310) );
  BUF_X1 U800 ( .A(n3497), .Z(n1301) );
  BUF_X1 U801 ( .A(n3525), .Z(n1148) );
  BUF_X1 U802 ( .A(n3528), .Z(n1139) );
  BUF_X1 U803 ( .A(n3556), .Z(n730) );
  NAND2_X1 U804 ( .A1(n6247), .A2(n6312), .ZN(n4995) );
  NAND2_X1 U805 ( .A1(n4804), .A2(n4869), .ZN(n3552) );
  BUF_X1 U806 ( .A(n3103), .Z(n1745) );
  BUF_X1 U807 ( .A(n3098), .Z(n1748) );
  BUF_X1 U808 ( .A(n3093), .Z(n1751) );
  BUF_X1 U809 ( .A(n3088), .Z(n1754) );
  BUF_X1 U810 ( .A(n3083), .Z(n1757) );
  BUF_X1 U811 ( .A(n3078), .Z(n1760) );
  BUF_X1 U812 ( .A(n3073), .Z(n1763) );
  BUF_X1 U813 ( .A(n3068), .Z(n1766) );
  BUF_X1 U814 ( .A(n3063), .Z(n1769) );
  BUF_X1 U815 ( .A(n3058), .Z(n1772) );
  BUF_X1 U816 ( .A(n3053), .Z(n1775) );
  BUF_X1 U817 ( .A(n3048), .Z(n1778) );
  BUF_X1 U818 ( .A(n3043), .Z(n1781) );
  BUF_X1 U819 ( .A(n3038), .Z(n1784) );
  BUF_X1 U820 ( .A(n3033), .Z(n1787) );
  BUF_X1 U821 ( .A(n2996), .Z(n1790) );
  BUF_X1 U822 ( .A(n3303), .Z(n1505) );
  BUF_X1 U823 ( .A(n3299), .Z(n1508) );
  BUF_X1 U824 ( .A(n3295), .Z(n1511) );
  BUF_X1 U825 ( .A(n3291), .Z(n1514) );
  BUF_X1 U826 ( .A(n3287), .Z(n1517) );
  BUF_X1 U827 ( .A(n3283), .Z(n1520) );
  BUF_X1 U828 ( .A(n3279), .Z(n1523) );
  BUF_X1 U829 ( .A(n3275), .Z(n1526) );
  BUF_X1 U830 ( .A(n3271), .Z(n1529) );
  BUF_X1 U831 ( .A(n3267), .Z(n1532) );
  BUF_X1 U832 ( .A(n3263), .Z(n1535) );
  BUF_X1 U833 ( .A(n3259), .Z(n1538) );
  BUF_X1 U834 ( .A(n3255), .Z(n1541) );
  BUF_X1 U835 ( .A(n3251), .Z(n1544) );
  BUF_X1 U836 ( .A(n3247), .Z(n1547) );
  BUF_X1 U837 ( .A(n3242), .Z(n1550) );
  BUF_X1 U838 ( .A(n3238), .Z(n1649) );
  BUF_X1 U839 ( .A(n3234), .Z(n1652) );
  BUF_X1 U840 ( .A(n3230), .Z(n1655) );
  BUF_X1 U841 ( .A(n3226), .Z(n1658) );
  BUF_X1 U842 ( .A(n3222), .Z(n1661) );
  BUF_X1 U843 ( .A(n3218), .Z(n1664) );
  BUF_X1 U844 ( .A(n3214), .Z(n1667) );
  BUF_X1 U845 ( .A(n3210), .Z(n1670) );
  BUF_X1 U846 ( .A(n3206), .Z(n1673) );
  BUF_X1 U847 ( .A(n3202), .Z(n1676) );
  BUF_X1 U848 ( .A(n3198), .Z(n1679) );
  BUF_X1 U849 ( .A(n3194), .Z(n1682) );
  BUF_X1 U850 ( .A(n3190), .Z(n1685) );
  BUF_X1 U851 ( .A(n3186), .Z(n1688) );
  BUF_X1 U852 ( .A(n3182), .Z(n1691) );
  BUF_X1 U853 ( .A(n3177), .Z(n1694) );
  BUF_X1 U854 ( .A(n3173), .Z(n1697) );
  BUF_X1 U855 ( .A(n3169), .Z(n1700) );
  BUF_X1 U856 ( .A(n3165), .Z(n1703) );
  BUF_X1 U857 ( .A(n3161), .Z(n1706) );
  BUF_X1 U858 ( .A(n3157), .Z(n1709) );
  BUF_X1 U859 ( .A(n3153), .Z(n1712) );
  BUF_X1 U860 ( .A(n3149), .Z(n1715) );
  BUF_X1 U861 ( .A(n3145), .Z(n1718) );
  BUF_X1 U862 ( .A(n3141), .Z(n1721) );
  BUF_X1 U863 ( .A(n3137), .Z(n1724) );
  BUF_X1 U864 ( .A(n3133), .Z(n1727) );
  BUF_X1 U865 ( .A(n3129), .Z(n1730) );
  BUF_X1 U866 ( .A(n3125), .Z(n1733) );
  BUF_X1 U867 ( .A(n3121), .Z(n1736) );
  BUF_X1 U868 ( .A(n3117), .Z(n1739) );
  BUF_X1 U869 ( .A(n3112), .Z(n1742) );
  BUF_X1 U870 ( .A(n3375), .Z(n1457) );
  BUF_X1 U871 ( .A(n3371), .Z(n1460) );
  BUF_X1 U872 ( .A(n3367), .Z(n1463) );
  BUF_X1 U873 ( .A(n3362), .Z(n1466) );
  BUF_X1 U874 ( .A(n3356), .Z(n1469) );
  BUF_X1 U875 ( .A(n3351), .Z(n1472) );
  BUF_X1 U876 ( .A(n3346), .Z(n1475) );
  BUF_X1 U877 ( .A(n3340), .Z(n1478) );
  BUF_X1 U878 ( .A(n3336), .Z(n1481) );
  BUF_X1 U879 ( .A(n3332), .Z(n1484) );
  BUF_X1 U880 ( .A(n3328), .Z(n1487) );
  BUF_X1 U881 ( .A(n3324), .Z(n1490) );
  BUF_X1 U882 ( .A(n3320), .Z(n1493) );
  BUF_X1 U883 ( .A(n3316), .Z(n1496) );
  BUF_X1 U884 ( .A(n3312), .Z(n1499) );
  BUF_X1 U885 ( .A(n3307), .Z(n1502) );
  BUF_X1 U886 ( .A(n3413), .Z(n1433) );
  BUF_X1 U887 ( .A(n3409), .Z(n1436) );
  BUF_X1 U888 ( .A(n3403), .Z(n1439) );
  BUF_X1 U889 ( .A(n3398), .Z(n1442) );
  BUF_X1 U890 ( .A(n3394), .Z(n1445) );
  BUF_X1 U891 ( .A(n3390), .Z(n1448) );
  BUF_X1 U892 ( .A(n3386), .Z(n1451) );
  BUF_X1 U893 ( .A(n3380), .Z(n1454) );
  NAND2_X1 U894 ( .A1(n6248), .A2(n6247), .ZN(n4887) );
  NAND2_X1 U895 ( .A1(n6246), .A2(n6247), .ZN(n4888) );
  NAND2_X1 U896 ( .A1(n6281), .A2(n6247), .ZN(n4927) );
  NAND2_X1 U897 ( .A1(n6298), .A2(n6247), .ZN(n4957) );
  NAND2_X1 U898 ( .A1(n6300), .A2(n6247), .ZN(n4964) );
  NAND2_X1 U899 ( .A1(n4805), .A2(n4804), .ZN(n3444) );
  NAND2_X1 U900 ( .A1(n4803), .A2(n4804), .ZN(n3445) );
  NAND2_X1 U901 ( .A1(n4838), .A2(n4804), .ZN(n3484) );
  NAND2_X1 U902 ( .A1(n4855), .A2(n4804), .ZN(n3514) );
  NAND2_X1 U903 ( .A1(n4857), .A2(n4804), .ZN(n3521) );
  AND2_X1 U904 ( .A1(n6268), .A2(n6247), .ZN(n4909) );
  AND2_X1 U905 ( .A1(n4825), .A2(n4804), .ZN(n3466) );
  INV_X1 U906 ( .A(n2955), .ZN(n3363) );
  NOR2_X1 U907 ( .A1(n3372), .A2(n3373), .ZN(n3343) );
  NOR2_X1 U908 ( .A1(n3369), .A2(n3370), .ZN(n3383) );
  NAND2_X1 U909 ( .A1(n3400), .A2(n3358), .ZN(n3065) );
  NAND2_X1 U910 ( .A1(n3400), .A2(n3353), .ZN(n3060) );
  NAND2_X1 U911 ( .A1(n3400), .A2(n3348), .ZN(n3055) );
  NAND2_X1 U912 ( .A1(n3400), .A2(n3343), .ZN(n3050) );
  NAND2_X1 U913 ( .A1(n3358), .A2(n3383), .ZN(n3045) );
  NAND2_X1 U914 ( .A1(n3353), .A2(n3383), .ZN(n3040) );
  NAND2_X1 U915 ( .A1(n3348), .A2(n3383), .ZN(n3035) );
  NOR2_X1 U916 ( .A1(n3029), .A2(n3105), .ZN(n3103) );
  NOR2_X1 U917 ( .A1(n3029), .A2(n3100), .ZN(n3098) );
  NOR2_X1 U918 ( .A1(n3029), .A2(n3095), .ZN(n3093) );
  NOR2_X1 U919 ( .A1(n3029), .A2(n3090), .ZN(n3088) );
  NOR2_X1 U920 ( .A1(n3029), .A2(n3085), .ZN(n3083) );
  NOR2_X1 U921 ( .A1(n3029), .A2(n3080), .ZN(n3078) );
  NOR2_X1 U922 ( .A1(n3029), .A2(n3075), .ZN(n3073) );
  NOR2_X1 U923 ( .A1(n3029), .A2(n3070), .ZN(n3068) );
  NOR2_X1 U924 ( .A1(n3029), .A2(n3065), .ZN(n3063) );
  NOR2_X1 U925 ( .A1(n3029), .A2(n3060), .ZN(n3058) );
  NOR2_X1 U926 ( .A1(n3029), .A2(n3055), .ZN(n3053) );
  NOR2_X1 U927 ( .A1(n3029), .A2(n3050), .ZN(n3048) );
  NOR2_X1 U928 ( .A1(n3029), .A2(n3045), .ZN(n3043) );
  NOR2_X1 U929 ( .A1(n3029), .A2(n3040), .ZN(n3038) );
  NOR2_X1 U930 ( .A1(n3029), .A2(n3035), .ZN(n3033) );
  NOR2_X1 U931 ( .A1(n3029), .A2(n3030), .ZN(n2996) );
  NAND2_X1 U932 ( .A1(n3364), .A2(n3358), .ZN(n3105) );
  NAND2_X1 U933 ( .A1(n3364), .A2(n3353), .ZN(n3100) );
  NAND2_X1 U934 ( .A1(n3342), .A2(n3358), .ZN(n3085) );
  NAND2_X1 U935 ( .A1(n3342), .A2(n3353), .ZN(n3080) );
  NAND2_X1 U936 ( .A1(n3364), .A2(n3348), .ZN(n3095) );
  NAND2_X1 U937 ( .A1(n3342), .A2(n3348), .ZN(n3075) );
  NAND2_X1 U938 ( .A1(n3364), .A2(n3343), .ZN(n3090) );
  NAND2_X1 U939 ( .A1(n3342), .A2(n3343), .ZN(n3070) );
  NOR2_X1 U940 ( .A1(n3105), .A2(n3244), .ZN(n3303) );
  NOR2_X1 U941 ( .A1(n3100), .A2(n3244), .ZN(n3299) );
  NOR2_X1 U942 ( .A1(n3095), .A2(n3244), .ZN(n3295) );
  NOR2_X1 U943 ( .A1(n3090), .A2(n3244), .ZN(n3291) );
  NOR2_X1 U944 ( .A1(n3085), .A2(n3244), .ZN(n3287) );
  NOR2_X1 U945 ( .A1(n3080), .A2(n3244), .ZN(n3283) );
  NOR2_X1 U946 ( .A1(n3075), .A2(n3244), .ZN(n3279) );
  NOR2_X1 U947 ( .A1(n3070), .A2(n3244), .ZN(n3275) );
  NOR2_X1 U948 ( .A1(n3065), .A2(n3244), .ZN(n3271) );
  NOR2_X1 U949 ( .A1(n3060), .A2(n3244), .ZN(n3267) );
  NOR2_X1 U950 ( .A1(n3055), .A2(n3244), .ZN(n3263) );
  NOR2_X1 U951 ( .A1(n3050), .A2(n3244), .ZN(n3259) );
  NOR2_X1 U952 ( .A1(n3045), .A2(n3244), .ZN(n3255) );
  NOR2_X1 U953 ( .A1(n3040), .A2(n3244), .ZN(n3251) );
  NOR2_X1 U954 ( .A1(n3035), .A2(n3244), .ZN(n3247) );
  NOR2_X1 U955 ( .A1(n3030), .A2(n3244), .ZN(n3242) );
  NOR2_X1 U956 ( .A1(n3105), .A2(n3179), .ZN(n3238) );
  NOR2_X1 U957 ( .A1(n3100), .A2(n3179), .ZN(n3234) );
  NOR2_X1 U958 ( .A1(n3095), .A2(n3179), .ZN(n3230) );
  NOR2_X1 U959 ( .A1(n3090), .A2(n3179), .ZN(n3226) );
  NOR2_X1 U960 ( .A1(n3085), .A2(n3179), .ZN(n3222) );
  NOR2_X1 U961 ( .A1(n3080), .A2(n3179), .ZN(n3218) );
  NOR2_X1 U962 ( .A1(n3075), .A2(n3179), .ZN(n3214) );
  NOR2_X1 U963 ( .A1(n3070), .A2(n3179), .ZN(n3210) );
  NOR2_X1 U964 ( .A1(n3065), .A2(n3179), .ZN(n3206) );
  NOR2_X1 U965 ( .A1(n3060), .A2(n3179), .ZN(n3202) );
  NOR2_X1 U966 ( .A1(n3055), .A2(n3179), .ZN(n3198) );
  NOR2_X1 U967 ( .A1(n3050), .A2(n3179), .ZN(n3194) );
  NOR2_X1 U968 ( .A1(n3045), .A2(n3179), .ZN(n3190) );
  NOR2_X1 U969 ( .A1(n3040), .A2(n3179), .ZN(n3186) );
  NOR2_X1 U970 ( .A1(n3035), .A2(n3179), .ZN(n3182) );
  NOR2_X1 U971 ( .A1(n3030), .A2(n3179), .ZN(n3177) );
  NOR2_X1 U972 ( .A1(n3105), .A2(n3114), .ZN(n3173) );
  NOR2_X1 U973 ( .A1(n3100), .A2(n3114), .ZN(n3169) );
  NOR2_X1 U974 ( .A1(n3095), .A2(n3114), .ZN(n3165) );
  NOR2_X1 U975 ( .A1(n3090), .A2(n3114), .ZN(n3161) );
  NOR2_X1 U976 ( .A1(n3085), .A2(n3114), .ZN(n3157) );
  NOR2_X1 U977 ( .A1(n3080), .A2(n3114), .ZN(n3153) );
  NOR2_X1 U978 ( .A1(n3075), .A2(n3114), .ZN(n3149) );
  NOR2_X1 U979 ( .A1(n3070), .A2(n3114), .ZN(n3145) );
  NOR2_X1 U980 ( .A1(n3065), .A2(n3114), .ZN(n3141) );
  NOR2_X1 U981 ( .A1(n3060), .A2(n3114), .ZN(n3137) );
  NOR2_X1 U982 ( .A1(n3055), .A2(n3114), .ZN(n3133) );
  NOR2_X1 U983 ( .A1(n3050), .A2(n3114), .ZN(n3129) );
  NOR2_X1 U984 ( .A1(n3045), .A2(n3114), .ZN(n3125) );
  NOR2_X1 U985 ( .A1(n3040), .A2(n3114), .ZN(n3121) );
  NOR2_X1 U986 ( .A1(n3035), .A2(n3114), .ZN(n3117) );
  NOR2_X1 U987 ( .A1(n3030), .A2(n3114), .ZN(n3112) );
  NOR2_X1 U988 ( .A1(n3105), .A2(n3309), .ZN(n3375) );
  NOR2_X1 U989 ( .A1(n3100), .A2(n3309), .ZN(n3371) );
  NOR2_X1 U990 ( .A1(n3095), .A2(n3309), .ZN(n3367) );
  NOR2_X1 U991 ( .A1(n3090), .A2(n3309), .ZN(n3362) );
  NOR2_X1 U992 ( .A1(n3085), .A2(n3309), .ZN(n3356) );
  NOR2_X1 U993 ( .A1(n3080), .A2(n3309), .ZN(n3351) );
  NOR2_X1 U994 ( .A1(n3075), .A2(n3309), .ZN(n3346) );
  NOR2_X1 U995 ( .A1(n3070), .A2(n3309), .ZN(n3340) );
  NOR2_X1 U996 ( .A1(n3065), .A2(n3309), .ZN(n3336) );
  NOR2_X1 U997 ( .A1(n3060), .A2(n3309), .ZN(n3332) );
  NOR2_X1 U998 ( .A1(n3055), .A2(n3309), .ZN(n3328) );
  NOR2_X1 U999 ( .A1(n3050), .A2(n3309), .ZN(n3324) );
  NOR2_X1 U1000 ( .A1(n3045), .A2(n3309), .ZN(n3320) );
  NOR2_X1 U1001 ( .A1(n3040), .A2(n3309), .ZN(n3316) );
  NOR2_X1 U1002 ( .A1(n3035), .A2(n3309), .ZN(n3312) );
  NOR2_X1 U1003 ( .A1(n3030), .A2(n3309), .ZN(n3307) );
  AND2_X1 U1004 ( .A1(n6309), .A2(n6251), .ZN(n6260) );
  AND2_X1 U1005 ( .A1(n4866), .A2(n4808), .ZN(n4817) );
  NOR2_X1 U1006 ( .A1(n3065), .A2(n3382), .ZN(n3413) );
  NOR2_X1 U1007 ( .A1(n3060), .A2(n3382), .ZN(n3409) );
  NOR2_X1 U1008 ( .A1(n3055), .A2(n3382), .ZN(n3403) );
  NOR2_X1 U1009 ( .A1(n3050), .A2(n3382), .ZN(n3398) );
  NOR2_X1 U1010 ( .A1(n3045), .A2(n3382), .ZN(n3394) );
  NOR2_X1 U1011 ( .A1(n3040), .A2(n3382), .ZN(n3390) );
  NOR2_X1 U1012 ( .A1(n3035), .A2(n3382), .ZN(n3386) );
  NOR2_X1 U1013 ( .A1(n3030), .A2(n3382), .ZN(n3380) );
  AND2_X1 U1014 ( .A1(n6310), .A2(n6251), .ZN(n6261) );
  AND2_X1 U1015 ( .A1(n4867), .A2(n4808), .ZN(n4818) );
  AND2_X1 U1016 ( .A1(n6310), .A2(n6249), .ZN(n6256) );
  AND2_X1 U1017 ( .A1(n4867), .A2(n4806), .ZN(n4813) );
  AND2_X1 U1018 ( .A1(n6310), .A2(n6247), .ZN(n6255) );
  AND2_X1 U1019 ( .A1(n6309), .A2(n6247), .ZN(n6257) );
  AND2_X1 U1020 ( .A1(n4867), .A2(n4804), .ZN(n4812) );
  AND2_X1 U1021 ( .A1(n4866), .A2(n4804), .ZN(n4814) );
  AND2_X1 U1022 ( .A1(n6309), .A2(n6250), .ZN(n6259) );
  AND2_X1 U1023 ( .A1(n4866), .A2(n4807), .ZN(n4816) );
  AND2_X1 U1024 ( .A1(n6309), .A2(n6249), .ZN(n6262) );
  AND2_X1 U1025 ( .A1(n4866), .A2(n4806), .ZN(n4819) );
  AND2_X1 U1026 ( .A1(n6310), .A2(n6250), .ZN(n6263) );
  AND2_X1 U1027 ( .A1(n4867), .A2(n4807), .ZN(n4820) );
  NAND2_X1 U1028 ( .A1(n6296), .A2(n6257), .ZN(n4953) );
  NAND2_X1 U1029 ( .A1(n6296), .A2(n6256), .ZN(n4951) );
  NAND2_X1 U1030 ( .A1(n6296), .A2(n6262), .ZN(n4952) );
  NAND2_X1 U1031 ( .A1(n6296), .A2(n6263), .ZN(n4956) );
  NAND2_X1 U1032 ( .A1(n6296), .A2(n6259), .ZN(n4954) );
  NAND2_X1 U1033 ( .A1(n6296), .A2(n6261), .ZN(n4955) );
  NAND2_X1 U1034 ( .A1(n6296), .A2(n6260), .ZN(n4959) );
  NAND2_X1 U1035 ( .A1(n6296), .A2(n6287), .ZN(n4949) );
  NAND2_X1 U1036 ( .A1(n6296), .A2(n6255), .ZN(n4950) );
  NAND2_X1 U1037 ( .A1(n4853), .A2(n4814), .ZN(n3510) );
  NAND2_X1 U1038 ( .A1(n4853), .A2(n4813), .ZN(n3508) );
  NAND2_X1 U1039 ( .A1(n4853), .A2(n4819), .ZN(n3509) );
  NAND2_X1 U1040 ( .A1(n4853), .A2(n4820), .ZN(n3513) );
  NAND2_X1 U1041 ( .A1(n4853), .A2(n4816), .ZN(n3511) );
  NAND2_X1 U1042 ( .A1(n4853), .A2(n4818), .ZN(n3512) );
  NAND2_X1 U1043 ( .A1(n4853), .A2(n4817), .ZN(n3516) );
  NAND2_X1 U1044 ( .A1(n4853), .A2(n4844), .ZN(n3506) );
  NAND2_X1 U1045 ( .A1(n4853), .A2(n4812), .ZN(n3507) );
  NAND2_X1 U1046 ( .A1(n6248), .A2(n6249), .ZN(n4891) );
  NAND2_X1 U1047 ( .A1(n6246), .A2(n6249), .ZN(n4889) );
  NAND2_X1 U1048 ( .A1(n6298), .A2(n6249), .ZN(n4980) );
  NAND2_X1 U1049 ( .A1(n4805), .A2(n4806), .ZN(n3448) );
  NAND2_X1 U1050 ( .A1(n4803), .A2(n4806), .ZN(n3446) );
  NAND2_X1 U1051 ( .A1(n4855), .A2(n4806), .ZN(n3537) );
  BUF_X1 U1052 ( .A(n1797), .Z(n1800) );
  BUF_X1 U1053 ( .A(n1808), .Z(n1811) );
  BUF_X1 U1054 ( .A(n1819), .Z(n1822) );
  BUF_X1 U1055 ( .A(n1830), .Z(n1833) );
  BUF_X1 U1056 ( .A(n2545), .Z(n2548) );
  BUF_X1 U1057 ( .A(n2556), .Z(n2559) );
  BUF_X1 U1058 ( .A(n2567), .Z(n2570) );
  BUF_X1 U1059 ( .A(n2578), .Z(n2581) );
  BUF_X1 U1060 ( .A(n2589), .Z(n2592) );
  BUF_X1 U1061 ( .A(n2600), .Z(n2603) );
  BUF_X1 U1062 ( .A(n2707), .Z(n2710) );
  BUF_X1 U1063 ( .A(n2718), .Z(n2721) );
  BUF_X1 U1064 ( .A(n2729), .Z(n2732) );
  BUF_X1 U1065 ( .A(n2740), .Z(n2743) );
  BUF_X1 U1066 ( .A(n2751), .Z(n2754) );
  BUF_X1 U1067 ( .A(n2762), .Z(n2765) );
  BUF_X1 U1068 ( .A(n2773), .Z(n2776) );
  BUF_X1 U1069 ( .A(n2784), .Z(n2787) );
  BUF_X1 U1070 ( .A(n2795), .Z(n2798) );
  BUF_X1 U1071 ( .A(n2806), .Z(n2809) );
  BUF_X1 U1072 ( .A(n2817), .Z(n2820) );
  BUF_X1 U1073 ( .A(n2828), .Z(n2831) );
  BUF_X1 U1074 ( .A(n2839), .Z(n2842) );
  BUF_X1 U1075 ( .A(n2850), .Z(n2853) );
  BUF_X1 U1076 ( .A(n2861), .Z(n2864) );
  BUF_X1 U1077 ( .A(n2872), .Z(n2875) );
  BUF_X1 U1078 ( .A(n2883), .Z(n2886) );
  BUF_X1 U1079 ( .A(n2894), .Z(n2897) );
  BUF_X1 U1080 ( .A(n2906), .Z(n2909) );
  BUF_X1 U1081 ( .A(n2922), .Z(n2925) );
  BUF_X1 U1082 ( .A(n2933), .Z(n2936) );
  BUF_X1 U1083 ( .A(n2944), .Z(n2947) );
  BUF_X1 U1084 ( .A(n1797), .Z(n1801) );
  BUF_X1 U1085 ( .A(n1808), .Z(n1812) );
  BUF_X1 U1086 ( .A(n1819), .Z(n1823) );
  BUF_X1 U1087 ( .A(n1830), .Z(n1834) );
  BUF_X1 U1088 ( .A(n2545), .Z(n2549) );
  BUF_X1 U1089 ( .A(n2556), .Z(n2560) );
  BUF_X1 U1090 ( .A(n2567), .Z(n2571) );
  BUF_X1 U1091 ( .A(n2578), .Z(n2582) );
  BUF_X1 U1092 ( .A(n2589), .Z(n2593) );
  BUF_X1 U1093 ( .A(n2600), .Z(n2604) );
  BUF_X1 U1094 ( .A(n2707), .Z(n2711) );
  BUF_X1 U1095 ( .A(n2718), .Z(n2722) );
  BUF_X1 U1096 ( .A(n2729), .Z(n2733) );
  BUF_X1 U1097 ( .A(n2740), .Z(n2744) );
  BUF_X1 U1098 ( .A(n2751), .Z(n2755) );
  BUF_X1 U1099 ( .A(n2762), .Z(n2766) );
  BUF_X1 U1100 ( .A(n2773), .Z(n2777) );
  BUF_X1 U1101 ( .A(n2784), .Z(n2788) );
  BUF_X1 U1102 ( .A(n2795), .Z(n2799) );
  BUF_X1 U1103 ( .A(n2806), .Z(n2810) );
  BUF_X1 U1104 ( .A(n2817), .Z(n2821) );
  BUF_X1 U1105 ( .A(n2828), .Z(n2832) );
  BUF_X1 U1106 ( .A(n2839), .Z(n2843) );
  BUF_X1 U1107 ( .A(n2850), .Z(n2854) );
  BUF_X1 U1108 ( .A(n2861), .Z(n2865) );
  BUF_X1 U1109 ( .A(n2872), .Z(n2876) );
  BUF_X1 U1110 ( .A(n2883), .Z(n2887) );
  BUF_X1 U1111 ( .A(n2894), .Z(n2899) );
  BUF_X1 U1112 ( .A(n2906), .Z(n2910) );
  BUF_X1 U1113 ( .A(n2922), .Z(n2926) );
  BUF_X1 U1114 ( .A(n2933), .Z(n2937) );
  BUF_X1 U1115 ( .A(n2944), .Z(n2948) );
  BUF_X1 U1116 ( .A(n1797), .Z(n1802) );
  BUF_X1 U1117 ( .A(n1808), .Z(n1813) );
  BUF_X1 U1118 ( .A(n1819), .Z(n1824) );
  BUF_X1 U1119 ( .A(n1830), .Z(n1835) );
  BUF_X1 U1120 ( .A(n2545), .Z(n2550) );
  BUF_X1 U1121 ( .A(n2556), .Z(n2561) );
  BUF_X1 U1122 ( .A(n2567), .Z(n2572) );
  BUF_X1 U1123 ( .A(n2578), .Z(n2583) );
  BUF_X1 U1124 ( .A(n2589), .Z(n2594) );
  BUF_X1 U1125 ( .A(n2600), .Z(n2605) );
  BUF_X1 U1126 ( .A(n2707), .Z(n2712) );
  BUF_X1 U1127 ( .A(n2718), .Z(n2723) );
  BUF_X1 U1128 ( .A(n2729), .Z(n2734) );
  BUF_X1 U1129 ( .A(n2740), .Z(n2745) );
  BUF_X1 U1130 ( .A(n2751), .Z(n2756) );
  BUF_X1 U1131 ( .A(n2762), .Z(n2767) );
  BUF_X1 U1132 ( .A(n2773), .Z(n2778) );
  BUF_X1 U1133 ( .A(n2784), .Z(n2789) );
  BUF_X1 U1134 ( .A(n2795), .Z(n2800) );
  BUF_X1 U1135 ( .A(n2806), .Z(n2811) );
  BUF_X1 U1136 ( .A(n2817), .Z(n2822) );
  BUF_X1 U1137 ( .A(n2828), .Z(n2833) );
  BUF_X1 U1138 ( .A(n2839), .Z(n2844) );
  BUF_X1 U1139 ( .A(n2850), .Z(n2855) );
  BUF_X1 U1140 ( .A(n2861), .Z(n2866) );
  BUF_X1 U1141 ( .A(n2872), .Z(n2877) );
  BUF_X1 U1142 ( .A(n2883), .Z(n2888) );
  BUF_X1 U1143 ( .A(n2894), .Z(n2900) );
  BUF_X1 U1144 ( .A(n2906), .Z(n2911) );
  BUF_X1 U1145 ( .A(n2922), .Z(n2927) );
  BUF_X1 U1146 ( .A(n2933), .Z(n2938) );
  BUF_X1 U1147 ( .A(n2944), .Z(n2949) );
  BUF_X1 U1148 ( .A(n1798), .Z(n1803) );
  BUF_X1 U1149 ( .A(n1809), .Z(n1814) );
  BUF_X1 U1150 ( .A(n1820), .Z(n1825) );
  BUF_X1 U1151 ( .A(n1831), .Z(n1836) );
  BUF_X1 U1152 ( .A(n2546), .Z(n2551) );
  BUF_X1 U1153 ( .A(n2557), .Z(n2562) );
  BUF_X1 U1154 ( .A(n2568), .Z(n2573) );
  BUF_X1 U1155 ( .A(n2579), .Z(n2584) );
  BUF_X1 U1156 ( .A(n2590), .Z(n2595) );
  BUF_X1 U1157 ( .A(n2601), .Z(n2606) );
  BUF_X1 U1158 ( .A(n2708), .Z(n2713) );
  BUF_X1 U1159 ( .A(n2719), .Z(n2724) );
  BUF_X1 U1160 ( .A(n2730), .Z(n2735) );
  BUF_X1 U1161 ( .A(n2741), .Z(n2746) );
  BUF_X1 U1162 ( .A(n2752), .Z(n2757) );
  BUF_X1 U1163 ( .A(n2763), .Z(n2768) );
  BUF_X1 U1164 ( .A(n2774), .Z(n2779) );
  BUF_X1 U1165 ( .A(n2785), .Z(n2790) );
  BUF_X1 U1166 ( .A(n2796), .Z(n2801) );
  BUF_X1 U1167 ( .A(n2807), .Z(n2812) );
  BUF_X1 U1168 ( .A(n2818), .Z(n2823) );
  BUF_X1 U1169 ( .A(n2829), .Z(n2834) );
  BUF_X1 U1170 ( .A(n2840), .Z(n2845) );
  BUF_X1 U1171 ( .A(n2851), .Z(n2856) );
  BUF_X1 U1172 ( .A(n2862), .Z(n2867) );
  BUF_X1 U1173 ( .A(n2873), .Z(n2878) );
  BUF_X1 U1174 ( .A(n2884), .Z(n2889) );
  BUF_X1 U1175 ( .A(n2895), .Z(n2901) );
  BUF_X1 U1176 ( .A(n2907), .Z(n2912) );
  BUF_X1 U1177 ( .A(n2923), .Z(n2928) );
  BUF_X1 U1178 ( .A(n2934), .Z(n2939) );
  BUF_X1 U1179 ( .A(n2945), .Z(n2950) );
  BUF_X1 U1180 ( .A(n1798), .Z(n1804) );
  BUF_X1 U1181 ( .A(n1809), .Z(n1815) );
  BUF_X1 U1182 ( .A(n1820), .Z(n1826) );
  BUF_X1 U1183 ( .A(n1831), .Z(n1837) );
  BUF_X1 U1184 ( .A(n2546), .Z(n2552) );
  BUF_X1 U1185 ( .A(n2557), .Z(n2563) );
  BUF_X1 U1186 ( .A(n2568), .Z(n2574) );
  BUF_X1 U1187 ( .A(n2579), .Z(n2585) );
  BUF_X1 U1188 ( .A(n2590), .Z(n2596) );
  BUF_X1 U1189 ( .A(n2601), .Z(n2607) );
  BUF_X1 U1190 ( .A(n2708), .Z(n2714) );
  BUF_X1 U1191 ( .A(n2719), .Z(n2725) );
  BUF_X1 U1192 ( .A(n2730), .Z(n2736) );
  BUF_X1 U1193 ( .A(n2741), .Z(n2747) );
  BUF_X1 U1194 ( .A(n2752), .Z(n2758) );
  BUF_X1 U1195 ( .A(n2763), .Z(n2769) );
  BUF_X1 U1196 ( .A(n2774), .Z(n2780) );
  BUF_X1 U1197 ( .A(n2785), .Z(n2791) );
  BUF_X1 U1198 ( .A(n2796), .Z(n2802) );
  BUF_X1 U1199 ( .A(n2807), .Z(n2813) );
  BUF_X1 U1200 ( .A(n2818), .Z(n2824) );
  BUF_X1 U1201 ( .A(n2829), .Z(n2835) );
  BUF_X1 U1202 ( .A(n2840), .Z(n2846) );
  BUF_X1 U1203 ( .A(n2851), .Z(n2857) );
  BUF_X1 U1204 ( .A(n2862), .Z(n2868) );
  BUF_X1 U1205 ( .A(n2873), .Z(n2879) );
  BUF_X1 U1206 ( .A(n2884), .Z(n2890) );
  BUF_X1 U1207 ( .A(n2895), .Z(n2902) );
  BUF_X1 U1208 ( .A(n2907), .Z(n2913) );
  BUF_X1 U1209 ( .A(n2923), .Z(n2929) );
  BUF_X1 U1210 ( .A(n2934), .Z(n2940) );
  BUF_X1 U1211 ( .A(n2945), .Z(n2951) );
  BUF_X1 U1212 ( .A(n1798), .Z(n1805) );
  BUF_X1 U1213 ( .A(n1809), .Z(n1816) );
  BUF_X1 U1214 ( .A(n1820), .Z(n1827) );
  BUF_X1 U1215 ( .A(n1831), .Z(n1838) );
  BUF_X1 U1216 ( .A(n2546), .Z(n2553) );
  BUF_X1 U1217 ( .A(n2557), .Z(n2564) );
  BUF_X1 U1218 ( .A(n2568), .Z(n2575) );
  BUF_X1 U1219 ( .A(n2579), .Z(n2586) );
  BUF_X1 U1220 ( .A(n2590), .Z(n2597) );
  BUF_X1 U1221 ( .A(n2601), .Z(n2704) );
  BUF_X1 U1222 ( .A(n2708), .Z(n2715) );
  BUF_X1 U1223 ( .A(n2719), .Z(n2726) );
  BUF_X1 U1224 ( .A(n2730), .Z(n2737) );
  BUF_X1 U1225 ( .A(n2741), .Z(n2748) );
  BUF_X1 U1226 ( .A(n2752), .Z(n2759) );
  BUF_X1 U1227 ( .A(n2763), .Z(n2770) );
  BUF_X1 U1228 ( .A(n2774), .Z(n2781) );
  BUF_X1 U1229 ( .A(n2785), .Z(n2792) );
  BUF_X1 U1230 ( .A(n2796), .Z(n2803) );
  BUF_X1 U1231 ( .A(n2807), .Z(n2814) );
  BUF_X1 U1232 ( .A(n2818), .Z(n2825) );
  BUF_X1 U1233 ( .A(n2829), .Z(n2836) );
  BUF_X1 U1234 ( .A(n2840), .Z(n2847) );
  BUF_X1 U1235 ( .A(n2851), .Z(n2858) );
  BUF_X1 U1236 ( .A(n2862), .Z(n2869) );
  BUF_X1 U1237 ( .A(n2873), .Z(n2880) );
  BUF_X1 U1238 ( .A(n2884), .Z(n2891) );
  BUF_X1 U1239 ( .A(n2895), .Z(n2903) );
  BUF_X1 U1240 ( .A(n2907), .Z(n2914) );
  BUF_X1 U1241 ( .A(n2923), .Z(n2930) );
  BUF_X1 U1242 ( .A(n2934), .Z(n2941) );
  BUF_X1 U1243 ( .A(n2945), .Z(n2952) );
  BUF_X1 U1244 ( .A(n1799), .Z(n1806) );
  BUF_X1 U1245 ( .A(n1810), .Z(n1817) );
  BUF_X1 U1246 ( .A(n1821), .Z(n1828) );
  BUF_X1 U1247 ( .A(n1832), .Z(n1839) );
  BUF_X1 U1248 ( .A(n2547), .Z(n2554) );
  BUF_X1 U1249 ( .A(n2558), .Z(n2565) );
  BUF_X1 U1250 ( .A(n2569), .Z(n2576) );
  BUF_X1 U1251 ( .A(n2580), .Z(n2587) );
  BUF_X1 U1252 ( .A(n2591), .Z(n2598) );
  BUF_X1 U1253 ( .A(n2602), .Z(n2705) );
  BUF_X1 U1254 ( .A(n2709), .Z(n2716) );
  BUF_X1 U1255 ( .A(n2720), .Z(n2727) );
  BUF_X1 U1256 ( .A(n2731), .Z(n2738) );
  BUF_X1 U1257 ( .A(n2742), .Z(n2749) );
  BUF_X1 U1258 ( .A(n2753), .Z(n2760) );
  BUF_X1 U1259 ( .A(n2764), .Z(n2771) );
  BUF_X1 U1260 ( .A(n2775), .Z(n2782) );
  BUF_X1 U1261 ( .A(n2786), .Z(n2793) );
  BUF_X1 U1262 ( .A(n2797), .Z(n2804) );
  BUF_X1 U1263 ( .A(n2808), .Z(n2815) );
  BUF_X1 U1264 ( .A(n2819), .Z(n2826) );
  BUF_X1 U1265 ( .A(n2830), .Z(n2837) );
  BUF_X1 U1266 ( .A(n2841), .Z(n2848) );
  BUF_X1 U1267 ( .A(n2852), .Z(n2859) );
  BUF_X1 U1268 ( .A(n2863), .Z(n2870) );
  BUF_X1 U1269 ( .A(n2874), .Z(n2881) );
  BUF_X1 U1270 ( .A(n2885), .Z(n2892) );
  BUF_X1 U1271 ( .A(n2896), .Z(n2904) );
  BUF_X1 U1272 ( .A(n2908), .Z(n2915) );
  BUF_X1 U1273 ( .A(n2924), .Z(n2931) );
  BUF_X1 U1274 ( .A(n2935), .Z(n2942) );
  BUF_X1 U1275 ( .A(n2946), .Z(n2953) );
  BUF_X1 U1276 ( .A(n1799), .Z(n1807) );
  BUF_X1 U1277 ( .A(n1810), .Z(n1818) );
  BUF_X1 U1278 ( .A(n1821), .Z(n1829) );
  BUF_X1 U1279 ( .A(n1832), .Z(n2544) );
  BUF_X1 U1280 ( .A(n2547), .Z(n2555) );
  BUF_X1 U1281 ( .A(n2558), .Z(n2566) );
  BUF_X1 U1282 ( .A(n2569), .Z(n2577) );
  BUF_X1 U1283 ( .A(n2580), .Z(n2588) );
  BUF_X1 U1284 ( .A(n2591), .Z(n2599) );
  BUF_X1 U1285 ( .A(n2602), .Z(n2706) );
  BUF_X1 U1286 ( .A(n2709), .Z(n2717) );
  BUF_X1 U1287 ( .A(n2720), .Z(n2728) );
  BUF_X1 U1288 ( .A(n2731), .Z(n2739) );
  BUF_X1 U1289 ( .A(n2742), .Z(n2750) );
  BUF_X1 U1290 ( .A(n2753), .Z(n2761) );
  BUF_X1 U1291 ( .A(n2764), .Z(n2772) );
  BUF_X1 U1292 ( .A(n2775), .Z(n2783) );
  BUF_X1 U1293 ( .A(n2786), .Z(n2794) );
  BUF_X1 U1294 ( .A(n2797), .Z(n2805) );
  BUF_X1 U1295 ( .A(n2808), .Z(n2816) );
  BUF_X1 U1296 ( .A(n2819), .Z(n2827) );
  BUF_X1 U1297 ( .A(n2830), .Z(n2838) );
  BUF_X1 U1298 ( .A(n2841), .Z(n2849) );
  BUF_X1 U1299 ( .A(n2852), .Z(n2860) );
  BUF_X1 U1300 ( .A(n2863), .Z(n2871) );
  BUF_X1 U1301 ( .A(n2874), .Z(n2882) );
  BUF_X1 U1302 ( .A(n2885), .Z(n2893) );
  BUF_X1 U1303 ( .A(n2896), .Z(n2905) );
  BUF_X1 U1304 ( .A(n2908), .Z(n2917) );
  BUF_X1 U1305 ( .A(n2924), .Z(n2932) );
  BUF_X1 U1306 ( .A(n2935), .Z(n2943) );
  BUF_X1 U1307 ( .A(n2946), .Z(n2954) );
  NAND2_X1 U1308 ( .A1(n6247), .A2(n6313), .ZN(n4994) );
  NAND2_X1 U1309 ( .A1(n4804), .A2(n4870), .ZN(n3551) );
  AND2_X1 U1310 ( .A1(n6252), .A2(n6254), .ZN(n6248) );
  AND2_X1 U1311 ( .A1(n6252), .A2(n6253), .ZN(n6246) );
  AND2_X1 U1312 ( .A1(n4809), .A2(n4811), .ZN(n4805) );
  AND2_X1 U1313 ( .A1(n4809), .A2(n4810), .ZN(n4803) );
  AND2_X1 U1314 ( .A1(n6254), .A2(n6297), .ZN(n6298) );
  AND2_X1 U1315 ( .A1(n4811), .A2(n4854), .ZN(n4855) );
  NAND2_X1 U1316 ( .A1(n6297), .A2(n6287), .ZN(n4987) );
  NAND2_X1 U1317 ( .A1(n4854), .A2(n4844), .ZN(n3544) );
  NAND2_X1 U1318 ( .A1(n6283), .A2(n6284), .ZN(n4934) );
  NAND2_X1 U1319 ( .A1(n6283), .A2(n6285), .ZN(n4933) );
  NAND2_X1 U1320 ( .A1(n6283), .A2(n6261), .ZN(n4965) );
  NAND2_X1 U1321 ( .A1(n6283), .A2(n6260), .ZN(n4963) );
  NAND2_X1 U1322 ( .A1(n4840), .A2(n4841), .ZN(n3491) );
  NAND2_X1 U1323 ( .A1(n4840), .A2(n4842), .ZN(n3490) );
  NAND2_X1 U1324 ( .A1(n4840), .A2(n4818), .ZN(n3522) );
  NAND2_X1 U1325 ( .A1(n4840), .A2(n4817), .ZN(n3520) );
  NAND2_X1 U1326 ( .A1(n6255), .A2(n3374), .ZN(n4985) );
  NAND2_X1 U1327 ( .A1(n6257), .A2(n3374), .ZN(n4986) );
  NAND2_X1 U1328 ( .A1(n6256), .A2(n3374), .ZN(n4990) );
  NAND2_X1 U1329 ( .A1(n6262), .A2(n3374), .ZN(n4988) );
  NAND2_X1 U1330 ( .A1(n6263), .A2(n3374), .ZN(n4989) );
  NAND2_X1 U1331 ( .A1(n6260), .A2(n3374), .ZN(n4996) );
  NAND2_X1 U1332 ( .A1(n4812), .A2(n3384), .ZN(n3542) );
  NAND2_X1 U1333 ( .A1(n4814), .A2(n3384), .ZN(n3543) );
  NAND2_X1 U1334 ( .A1(n4813), .A2(n3384), .ZN(n3547) );
  NAND2_X1 U1335 ( .A1(n4819), .A2(n3384), .ZN(n3545) );
  NAND2_X1 U1336 ( .A1(n4820), .A2(n3384), .ZN(n3546) );
  NAND2_X1 U1337 ( .A1(n4817), .A2(n3384), .ZN(n3553) );
  NAND2_X1 U1338 ( .A1(n6252), .A2(n6255), .ZN(n4897) );
  NAND2_X1 U1339 ( .A1(n6252), .A2(n6257), .ZN(n4895) );
  NAND2_X1 U1340 ( .A1(n6252), .A2(n6256), .ZN(n4896) );
  NAND2_X1 U1341 ( .A1(n6252), .A2(n6259), .ZN(n4903) );
  NAND2_X1 U1342 ( .A1(n6252), .A2(n6261), .ZN(n4901) );
  NAND2_X1 U1343 ( .A1(n6252), .A2(n6260), .ZN(n4902) );
  NAND2_X1 U1344 ( .A1(n4809), .A2(n4812), .ZN(n3454) );
  NAND2_X1 U1345 ( .A1(n4809), .A2(n4814), .ZN(n3452) );
  NAND2_X1 U1346 ( .A1(n4809), .A2(n4813), .ZN(n3453) );
  NAND2_X1 U1347 ( .A1(n4809), .A2(n4816), .ZN(n3460) );
  NAND2_X1 U1348 ( .A1(n4809), .A2(n4818), .ZN(n3458) );
  NAND2_X1 U1349 ( .A1(n4809), .A2(n4817), .ZN(n3459) );
  NAND2_X1 U1350 ( .A1(n6248), .A2(n6251), .ZN(n4892) );
  NAND2_X1 U1351 ( .A1(n6246), .A2(n6251), .ZN(n4893) );
  NAND2_X1 U1352 ( .A1(n6267), .A2(n6251), .ZN(n4918) );
  NAND2_X1 U1353 ( .A1(n6268), .A2(n6251), .ZN(n4919) );
  NAND2_X1 U1354 ( .A1(n6298), .A2(n6251), .ZN(n4983) );
  NAND2_X1 U1355 ( .A1(n4805), .A2(n4808), .ZN(n3449) );
  NAND2_X1 U1356 ( .A1(n4803), .A2(n4808), .ZN(n3450) );
  NAND2_X1 U1357 ( .A1(n4824), .A2(n4808), .ZN(n3475) );
  NAND2_X1 U1358 ( .A1(n4825), .A2(n4808), .ZN(n3476) );
  NAND2_X1 U1359 ( .A1(n4855), .A2(n4808), .ZN(n3540) );
  NAND2_X1 U1360 ( .A1(n6248), .A2(n6250), .ZN(n4890) );
  NAND2_X1 U1361 ( .A1(n6246), .A2(n6250), .ZN(n4894) );
  NAND2_X1 U1362 ( .A1(n6281), .A2(n6250), .ZN(n4932) );
  NAND2_X1 U1363 ( .A1(n6298), .A2(n6250), .ZN(n4984) );
  NAND2_X1 U1364 ( .A1(n4805), .A2(n4807), .ZN(n3447) );
  NAND2_X1 U1365 ( .A1(n4803), .A2(n4807), .ZN(n3451) );
  NAND2_X1 U1366 ( .A1(n4838), .A2(n4807), .ZN(n3489) );
  NAND2_X1 U1367 ( .A1(n4855), .A2(n4807), .ZN(n3541) );
  AND2_X1 U1368 ( .A1(n6283), .A2(n6254), .ZN(n6281) );
  AND2_X1 U1369 ( .A1(n4840), .A2(n4811), .ZN(n4838) );
  NAND2_X1 U1370 ( .A1(n6286), .A2(n6297), .ZN(n4958) );
  NAND2_X1 U1371 ( .A1(n6285), .A2(n6297), .ZN(n4982) );
  NAND2_X1 U1372 ( .A1(n6284), .A2(n6297), .ZN(n4981) );
  NAND2_X1 U1373 ( .A1(n4843), .A2(n4854), .ZN(n3515) );
  NAND2_X1 U1374 ( .A1(n4842), .A2(n4854), .ZN(n3539) );
  NAND2_X1 U1375 ( .A1(n4841), .A2(n4854), .ZN(n3538) );
  BUF_X1 U1376 ( .A(RESET), .Z(n2955) );
  NAND2_X1 U1377 ( .A1(n6279), .A2(n6260), .ZN(n4926) );
  NAND2_X1 U1378 ( .A1(n4836), .A2(n4817), .ZN(n3483) );
  NAND2_X1 U1379 ( .A1(n6279), .A2(n6261), .ZN(n4928) );
  NAND2_X1 U1380 ( .A1(n4836), .A2(n4818), .ZN(n3485) );
  NAND2_X1 U1381 ( .A1(n6279), .A2(n6256), .ZN(n4921) );
  NAND2_X1 U1382 ( .A1(n4836), .A2(n4813), .ZN(n3478) );
  NAND2_X1 U1383 ( .A1(n6279), .A2(n6255), .ZN(n4922) );
  NAND2_X1 U1384 ( .A1(n6279), .A2(n6257), .ZN(n4920) );
  NAND2_X1 U1385 ( .A1(n4836), .A2(n4812), .ZN(n3479) );
  NAND2_X1 U1386 ( .A1(n4836), .A2(n4814), .ZN(n3477) );
  NAND2_X1 U1387 ( .A1(n6279), .A2(n6259), .ZN(n4924) );
  NAND2_X1 U1388 ( .A1(n4836), .A2(n4816), .ZN(n3481) );
  NAND2_X1 U1389 ( .A1(n6279), .A2(n6262), .ZN(n4925) );
  NAND2_X1 U1390 ( .A1(n4836), .A2(n4819), .ZN(n3482) );
  NAND2_X1 U1391 ( .A1(n6279), .A2(n6263), .ZN(n4923) );
  NAND2_X1 U1392 ( .A1(n4836), .A2(n4820), .ZN(n3480) );
  AND2_X1 U1393 ( .A1(n6249), .A2(n6312), .ZN(n5002) );
  AND2_X1 U1394 ( .A1(n6249), .A2(n6313), .ZN(n5000) );
  AND2_X1 U1395 ( .A1(n4806), .A2(n4869), .ZN(n3559) );
  AND2_X1 U1396 ( .A1(n4806), .A2(n4870), .ZN(n3557) );
  AND2_X1 U1397 ( .A1(n6296), .A2(n6254), .ZN(n6300) );
  AND2_X1 U1398 ( .A1(n4853), .A2(n4811), .ZN(n4857) );
  AND2_X1 U1399 ( .A1(n6316), .A2(n3381), .ZN(n6312) );
  AND2_X1 U1400 ( .A1(n4873), .A2(n3389), .ZN(n4869) );
  AND2_X1 U1401 ( .A1(n6253), .A2(n6249), .ZN(n6284) );
  AND2_X1 U1402 ( .A1(n4810), .A2(n4806), .ZN(n4841) );
  AND2_X1 U1403 ( .A1(n6268), .A2(n6249), .ZN(n4904) );
  AND2_X1 U1404 ( .A1(n6267), .A2(n6249), .ZN(n4908) );
  AND2_X1 U1405 ( .A1(n6281), .A2(n6249), .ZN(n4929) );
  AND2_X1 U1406 ( .A1(n6300), .A2(n6249), .ZN(n4971) );
  AND2_X1 U1407 ( .A1(n4825), .A2(n4806), .ZN(n3461) );
  AND2_X1 U1408 ( .A1(n4824), .A2(n4806), .ZN(n3465) );
  AND2_X1 U1409 ( .A1(n4838), .A2(n4806), .ZN(n3486) );
  AND2_X1 U1410 ( .A1(n4857), .A2(n4806), .ZN(n3528) );
  AND2_X1 U1411 ( .A1(n6253), .A2(n6251), .ZN(n6287) );
  AND2_X1 U1412 ( .A1(n4810), .A2(n4808), .ZN(n4844) );
  AND2_X1 U1413 ( .A1(n6296), .A2(n6285), .ZN(n4968) );
  AND2_X1 U1414 ( .A1(n6296), .A2(n6284), .ZN(n4970) );
  AND2_X1 U1415 ( .A1(n6296), .A2(n6286), .ZN(n4969) );
  AND2_X1 U1416 ( .A1(n4853), .A2(n4842), .ZN(n3525) );
  AND2_X1 U1417 ( .A1(n4853), .A2(n4841), .ZN(n3527) );
  AND2_X1 U1418 ( .A1(n4853), .A2(n4843), .ZN(n3526) );
  AND2_X1 U1419 ( .A1(n6251), .A2(n6312), .ZN(n4998) );
  AND2_X1 U1420 ( .A1(n4808), .A2(n4869), .ZN(n3555) );
  AND2_X1 U1421 ( .A1(n6283), .A2(n6262), .ZN(n4936) );
  AND2_X1 U1422 ( .A1(n6283), .A2(n6256), .ZN(n4937) );
  AND2_X1 U1423 ( .A1(n6283), .A2(n6257), .ZN(n4935) );
  AND2_X1 U1424 ( .A1(n6283), .A2(n6255), .ZN(n4939) );
  AND2_X1 U1425 ( .A1(n6283), .A2(n6287), .ZN(n4940) );
  AND2_X1 U1426 ( .A1(n6283), .A2(n6286), .ZN(n4930) );
  AND2_X1 U1427 ( .A1(n6283), .A2(n6259), .ZN(n4960) );
  AND2_X1 U1428 ( .A1(n6283), .A2(n6263), .ZN(n4961) );
  AND2_X1 U1429 ( .A1(n4840), .A2(n4819), .ZN(n3493) );
  AND2_X1 U1430 ( .A1(n4840), .A2(n4813), .ZN(n3494) );
  AND2_X1 U1431 ( .A1(n4840), .A2(n4814), .ZN(n3492) );
  AND2_X1 U1432 ( .A1(n4840), .A2(n4812), .ZN(n3496) );
  AND2_X1 U1433 ( .A1(n4840), .A2(n4844), .ZN(n3497) );
  AND2_X1 U1434 ( .A1(n4840), .A2(n4843), .ZN(n3487) );
  AND2_X1 U1435 ( .A1(n4840), .A2(n4816), .ZN(n3517) );
  AND2_X1 U1436 ( .A1(n4840), .A2(n4820), .ZN(n3518) );
  AND2_X1 U1437 ( .A1(n6250), .A2(n6312), .ZN(n4997) );
  AND2_X1 U1438 ( .A1(n6250), .A2(n6313), .ZN(n5001) );
  AND2_X1 U1439 ( .A1(n4807), .A2(n4869), .ZN(n3554) );
  AND2_X1 U1440 ( .A1(n4807), .A2(n4870), .ZN(n3558) );
  AND2_X1 U1441 ( .A1(n6267), .A2(n6247), .ZN(n4907) );
  AND2_X1 U1442 ( .A1(n4824), .A2(n4804), .ZN(n3464) );
  AND2_X1 U1443 ( .A1(n6252), .A2(n6263), .ZN(n4898) );
  AND2_X1 U1444 ( .A1(n6252), .A2(n6262), .ZN(n4899) );
  AND2_X1 U1445 ( .A1(n4809), .A2(n4820), .ZN(n3455) );
  AND2_X1 U1446 ( .A1(n4809), .A2(n4819), .ZN(n3456) );
  AND2_X1 U1447 ( .A1(n6281), .A2(n6251), .ZN(n4938) );
  AND2_X1 U1448 ( .A1(n6300), .A2(n6251), .ZN(n4967) );
  AND2_X1 U1449 ( .A1(n6313), .A2(n6251), .ZN(n4999) );
  AND2_X1 U1450 ( .A1(n4838), .A2(n4808), .ZN(n3495) );
  AND2_X1 U1451 ( .A1(n4857), .A2(n4808), .ZN(n3524) );
  AND2_X1 U1452 ( .A1(n4870), .A2(n4808), .ZN(n3556) );
  AND2_X1 U1453 ( .A1(n6253), .A2(n6250), .ZN(n6285) );
  AND2_X1 U1454 ( .A1(n4810), .A2(n4807), .ZN(n4842) );
  AND2_X1 U1455 ( .A1(n6268), .A2(n6250), .ZN(n4905) );
  AND2_X1 U1456 ( .A1(n6267), .A2(n6250), .ZN(n4906) );
  AND2_X1 U1457 ( .A1(n6300), .A2(n6250), .ZN(n4966) );
  AND2_X1 U1458 ( .A1(n4825), .A2(n4807), .ZN(n3462) );
  AND2_X1 U1459 ( .A1(n4824), .A2(n4807), .ZN(n3463) );
  AND2_X1 U1460 ( .A1(n4857), .A2(n4807), .ZN(n3523) );
  AND2_X1 U1461 ( .A1(n6277), .A2(n3381), .ZN(n6268) );
  AND2_X1 U1462 ( .A1(n4834), .A2(n3389), .ZN(n4825) );
  AND2_X1 U1463 ( .A1(n6261), .A2(n3374), .ZN(n4991) );
  AND2_X1 U1464 ( .A1(n6259), .A2(n3374), .ZN(n4992) );
  AND2_X1 U1465 ( .A1(n4818), .A2(n3384), .ZN(n3548) );
  AND2_X1 U1466 ( .A1(n4816), .A2(n3384), .ZN(n3549) );
  AND2_X1 U1467 ( .A1(n6253), .A2(n6247), .ZN(n6286) );
  AND2_X1 U1468 ( .A1(n4810), .A2(n4804), .ZN(n4843) );
  INV_X1 U1469 ( .A(n3419), .ZN(n3392) );
  NAND4_X1 U1470 ( .A1(n3106), .A2(n3108), .A3(n3368), .A4(n3365), .ZN(n3382)
         );
  NOR2_X1 U1471 ( .A1(n3376), .A2(n6266), .ZN(n6297) );
  NOR2_X1 U1472 ( .A1(n3385), .A2(n4823), .ZN(n4854) );
  NOR2_X1 U1473 ( .A1(n3405), .A2(n3406), .ZN(n3358) );
  NOR2_X1 U1474 ( .A1(n3373), .A2(n3406), .ZN(n3353) );
  NOR2_X1 U1475 ( .A1(n3372), .A2(n3405), .ZN(n3348) );
  NOR2_X1 U1476 ( .A1(n3377), .A2(n3359), .ZN(n3364) );
  NOR2_X1 U1477 ( .A1(n3370), .A2(n3359), .ZN(n3342) );
  NOR2_X1 U1478 ( .A1(n3369), .A2(n3377), .ZN(n3400) );
  INV_X1 U1479 ( .A(N8415), .ZN(n10918) );
  INV_X1 U1480 ( .A(N8559), .ZN(n10919) );
  INV_X1 U1481 ( .A(N2151), .ZN(n3391) );
  AND3_X1 U1482 ( .A1(n6264), .A2(n6265), .A3(n6266), .ZN(n6252) );
  AND3_X1 U1483 ( .A1(n4821), .A2(n4822), .A3(n4823), .ZN(n4809) );
  INV_X1 U1484 ( .A(n6266), .ZN(n3374) );
  INV_X1 U1485 ( .A(n4823), .ZN(n3384) );
  NOR2_X1 U1486 ( .A1(n6278), .A2(n6280), .ZN(n6309) );
  NOR2_X1 U1487 ( .A1(n4835), .A2(n4837), .ZN(n4866) );
  NOR2_X1 U1488 ( .A1(n3381), .A2(n6280), .ZN(n6310) );
  NOR2_X1 U1489 ( .A1(n3389), .A2(n4837), .ZN(n4867) );
  INV_X1 U1490 ( .A(n3109), .ZN(n3368) );
  INV_X1 U1491 ( .A(n3108), .ZN(n3366) );
  INV_X1 U1492 ( .A(n3107), .ZN(n3365) );
  AND2_X1 U1493 ( .A1(n6264), .A2(n3376), .ZN(n6279) );
  AND2_X1 U1494 ( .A1(n4821), .A2(n3385), .ZN(n4836) );
  INV_X1 U1495 ( .A(n6265), .ZN(n3376) );
  INV_X1 U1496 ( .A(n4822), .ZN(n3385) );
  INV_X1 U1497 ( .A(n6314), .ZN(n3379) );
  INV_X1 U1498 ( .A(n4871), .ZN(n3388) );
  NOR2_X1 U1499 ( .A1(n6265), .A2(n6266), .ZN(n6316) );
  NOR2_X1 U1500 ( .A1(n4822), .A2(n4823), .ZN(n4873) );
  INV_X1 U1501 ( .A(n6315), .ZN(n3378) );
  INV_X1 U1502 ( .A(n4872), .ZN(n3387) );
  INV_X1 U1503 ( .A(n6278), .ZN(n3381) );
  INV_X1 U1504 ( .A(n4835), .ZN(n3389) );
  AND2_X1 U1505 ( .A1(n6280), .A2(n3381), .ZN(n6253) );
  AND2_X1 U1506 ( .A1(n4837), .A2(n3389), .ZN(n4810) );
  AND2_X1 U1507 ( .A1(n6278), .A2(n6316), .ZN(n6313) );
  AND2_X1 U1508 ( .A1(n4835), .A2(n4873), .ZN(n4870) );
  BUF_X1 U1509 ( .A(N8702), .Z(n1795) );
  BUF_X1 U1510 ( .A(N8735), .Z(n1792) );
  BUF_X1 U1511 ( .A(N8702), .Z(n1794) );
  BUF_X1 U1512 ( .A(N8735), .Z(n1791) );
  AND2_X1 U1513 ( .A1(n6277), .A2(n6278), .ZN(n6267) );
  AND2_X1 U1514 ( .A1(n4834), .A2(n4835), .ZN(n4824) );
  BUF_X1 U1515 ( .A(N8702), .Z(n1796) );
  BUF_X1 U1516 ( .A(N8735), .Z(n1793) );
  AND2_X1 U1517 ( .A1(n6280), .A2(n6278), .ZN(n6254) );
  AND2_X1 U1518 ( .A1(n4837), .A2(n4835), .ZN(n4811) );
  INV_X1 U1519 ( .A(n3405), .ZN(n3373) );
  INV_X1 U1520 ( .A(n3377), .ZN(n3370) );
  INV_X1 U1521 ( .A(n3406), .ZN(n3372) );
  INV_X1 U1522 ( .A(n3359), .ZN(n3369) );
  AND3_X1 U1523 ( .A1(n6279), .A2(n6280), .A3(n6266), .ZN(n6277) );
  AND3_X1 U1524 ( .A1(n4836), .A2(n4837), .A3(n4823), .ZN(n4834) );
  NOR2_X1 U1525 ( .A1(n3265), .A2(n6233), .ZN(N8703) );
  NOR4_X1 U1526 ( .A1(n6234), .A2(n6235), .A3(n6236), .A4(n6237), .ZN(n6233)
         );
  NAND4_X1 U1527 ( .A1(n6301), .A2(n6302), .A3(n6303), .A4(n6304), .ZN(n6234)
         );
  NAND4_X1 U1528 ( .A1(n6288), .A2(n6289), .A3(n6290), .A4(n6291), .ZN(n6235)
         );
  NOR2_X1 U1529 ( .A1(n3276), .A2(n4790), .ZN(N8736) );
  NOR4_X1 U1530 ( .A1(n4791), .A2(n4792), .A3(n4793), .A4(n4794), .ZN(n4790)
         );
  NAND4_X1 U1531 ( .A1(n4858), .A2(n4859), .A3(n4860), .A4(n4861), .ZN(n4791)
         );
  NAND4_X1 U1532 ( .A1(n4845), .A2(n4846), .A3(n4847), .A4(n4848), .ZN(n4792)
         );
  NOR2_X1 U1533 ( .A1(n3265), .A2(n6192), .ZN(N8704) );
  NOR4_X1 U1534 ( .A1(n6193), .A2(n6194), .A3(n6195), .A4(n6196), .ZN(n6192)
         );
  NAND4_X1 U1535 ( .A1(n6224), .A2(n6225), .A3(n6226), .A4(n6227), .ZN(n6193)
         );
  NAND4_X1 U1536 ( .A1(n6215), .A2(n6216), .A3(n6217), .A4(n6218), .ZN(n6194)
         );
  NOR2_X1 U1537 ( .A1(n3276), .A2(n4749), .ZN(N8737) );
  NOR4_X1 U1538 ( .A1(n4750), .A2(n4751), .A3(n4752), .A4(n4753), .ZN(n4749)
         );
  NAND4_X1 U1539 ( .A1(n4781), .A2(n4782), .A3(n4783), .A4(n4784), .ZN(n4750)
         );
  NAND4_X1 U1540 ( .A1(n4772), .A2(n4773), .A3(n4774), .A4(n4775), .ZN(n4751)
         );
  NOR2_X1 U1541 ( .A1(n3265), .A2(n6151), .ZN(N8705) );
  NOR4_X1 U1542 ( .A1(n6152), .A2(n6153), .A3(n6154), .A4(n6155), .ZN(n6151)
         );
  NAND4_X1 U1543 ( .A1(n6183), .A2(n6184), .A3(n6185), .A4(n6186), .ZN(n6152)
         );
  NAND4_X1 U1544 ( .A1(n6174), .A2(n6175), .A3(n6176), .A4(n6177), .ZN(n6153)
         );
  NOR2_X1 U1545 ( .A1(n3276), .A2(n4708), .ZN(N8738) );
  NOR4_X1 U1546 ( .A1(n4709), .A2(n4710), .A3(n4711), .A4(n4712), .ZN(n4708)
         );
  NAND4_X1 U1547 ( .A1(n4740), .A2(n4741), .A3(n4742), .A4(n4743), .ZN(n4709)
         );
  NAND4_X1 U1548 ( .A1(n4731), .A2(n4732), .A3(n4733), .A4(n4734), .ZN(n4710)
         );
  NOR2_X1 U1549 ( .A1(n3265), .A2(n6110), .ZN(N8706) );
  NOR4_X1 U1550 ( .A1(n6111), .A2(n6112), .A3(n6113), .A4(n6114), .ZN(n6110)
         );
  NAND4_X1 U1551 ( .A1(n6142), .A2(n6143), .A3(n6144), .A4(n6145), .ZN(n6111)
         );
  NAND4_X1 U1552 ( .A1(n6133), .A2(n6134), .A3(n6135), .A4(n6136), .ZN(n6112)
         );
  NOR2_X1 U1553 ( .A1(n3277), .A2(n4667), .ZN(N8739) );
  NOR4_X1 U1554 ( .A1(n4668), .A2(n4669), .A3(n4670), .A4(n4671), .ZN(n4667)
         );
  NAND4_X1 U1555 ( .A1(n4699), .A2(n4700), .A3(n4701), .A4(n4702), .ZN(n4668)
         );
  NAND4_X1 U1556 ( .A1(n4690), .A2(n4691), .A3(n4692), .A4(n4693), .ZN(n4669)
         );
  NOR2_X1 U1557 ( .A1(n3266), .A2(n6069), .ZN(N8707) );
  NOR4_X1 U1558 ( .A1(n6070), .A2(n6071), .A3(n6072), .A4(n6073), .ZN(n6069)
         );
  NAND4_X1 U1559 ( .A1(n6101), .A2(n6102), .A3(n6103), .A4(n6104), .ZN(n6070)
         );
  NAND4_X1 U1560 ( .A1(n6092), .A2(n6093), .A3(n6094), .A4(n6095), .ZN(n6071)
         );
  NOR2_X1 U1561 ( .A1(n3277), .A2(n4626), .ZN(N8740) );
  NOR4_X1 U1562 ( .A1(n4627), .A2(n4628), .A3(n4629), .A4(n4630), .ZN(n4626)
         );
  NAND4_X1 U1563 ( .A1(n4658), .A2(n4659), .A3(n4660), .A4(n4661), .ZN(n4627)
         );
  NAND4_X1 U1564 ( .A1(n4649), .A2(n4650), .A3(n4651), .A4(n4652), .ZN(n4628)
         );
  NOR2_X1 U1565 ( .A1(n3266), .A2(n6028), .ZN(N8708) );
  NOR4_X1 U1566 ( .A1(n6029), .A2(n6030), .A3(n6031), .A4(n6032), .ZN(n6028)
         );
  NAND4_X1 U1567 ( .A1(n6060), .A2(n6061), .A3(n6062), .A4(n6063), .ZN(n6029)
         );
  NAND4_X1 U1568 ( .A1(n6051), .A2(n6052), .A3(n6053), .A4(n6054), .ZN(n6030)
         );
  NOR2_X1 U1569 ( .A1(n3277), .A2(n4585), .ZN(N8741) );
  NOR4_X1 U1570 ( .A1(n4586), .A2(n4587), .A3(n4588), .A4(n4589), .ZN(n4585)
         );
  NAND4_X1 U1571 ( .A1(n4617), .A2(n4618), .A3(n4619), .A4(n4620), .ZN(n4586)
         );
  NAND4_X1 U1572 ( .A1(n4608), .A2(n4609), .A3(n4610), .A4(n4611), .ZN(n4587)
         );
  NOR2_X1 U1573 ( .A1(n3266), .A2(n5987), .ZN(N8709) );
  NOR4_X1 U1574 ( .A1(n5988), .A2(n5989), .A3(n5990), .A4(n5991), .ZN(n5987)
         );
  NAND4_X1 U1575 ( .A1(n6019), .A2(n6020), .A3(n6021), .A4(n6022), .ZN(n5988)
         );
  NAND4_X1 U1576 ( .A1(n6010), .A2(n6011), .A3(n6012), .A4(n6013), .ZN(n5989)
         );
  NOR2_X1 U1577 ( .A1(n3277), .A2(n4544), .ZN(N8742) );
  NOR4_X1 U1578 ( .A1(n4545), .A2(n4546), .A3(n4547), .A4(n4548), .ZN(n4544)
         );
  NAND4_X1 U1579 ( .A1(n4576), .A2(n4577), .A3(n4578), .A4(n4579), .ZN(n4545)
         );
  NAND4_X1 U1580 ( .A1(n4567), .A2(n4568), .A3(n4569), .A4(n4570), .ZN(n4546)
         );
  NOR2_X1 U1581 ( .A1(n3266), .A2(n5946), .ZN(N8710) );
  NOR4_X1 U1582 ( .A1(n5947), .A2(n5948), .A3(n5949), .A4(n5950), .ZN(n5946)
         );
  NAND4_X1 U1583 ( .A1(n5978), .A2(n5979), .A3(n5980), .A4(n5981), .ZN(n5947)
         );
  NAND4_X1 U1584 ( .A1(n5969), .A2(n5970), .A3(n5971), .A4(n5972), .ZN(n5948)
         );
  NOR2_X1 U1585 ( .A1(n3278), .A2(n4503), .ZN(N8743) );
  NOR4_X1 U1586 ( .A1(n4504), .A2(n4505), .A3(n4506), .A4(n4507), .ZN(n4503)
         );
  NAND4_X1 U1587 ( .A1(n4535), .A2(n4536), .A3(n4537), .A4(n4538), .ZN(n4504)
         );
  NAND4_X1 U1588 ( .A1(n4526), .A2(n4527), .A3(n4528), .A4(n4529), .ZN(n4505)
         );
  NOR2_X1 U1589 ( .A1(n3268), .A2(n5905), .ZN(N8711) );
  NOR4_X1 U1590 ( .A1(n5906), .A2(n5907), .A3(n5908), .A4(n5909), .ZN(n5905)
         );
  NAND4_X1 U1591 ( .A1(n5937), .A2(n5938), .A3(n5939), .A4(n5940), .ZN(n5906)
         );
  NAND4_X1 U1592 ( .A1(n5928), .A2(n5929), .A3(n5930), .A4(n5931), .ZN(n5907)
         );
  NOR2_X1 U1593 ( .A1(n3278), .A2(n4462), .ZN(N8744) );
  NOR4_X1 U1594 ( .A1(n4463), .A2(n4464), .A3(n4465), .A4(n4466), .ZN(n4462)
         );
  NAND4_X1 U1595 ( .A1(n4494), .A2(n4495), .A3(n4496), .A4(n4497), .ZN(n4463)
         );
  NAND4_X1 U1596 ( .A1(n4485), .A2(n4486), .A3(n4487), .A4(n4488), .ZN(n4464)
         );
  NOR2_X1 U1597 ( .A1(n3268), .A2(n5864), .ZN(N8712) );
  NOR4_X1 U1598 ( .A1(n5865), .A2(n5866), .A3(n5867), .A4(n5868), .ZN(n5864)
         );
  NAND4_X1 U1599 ( .A1(n5896), .A2(n5897), .A3(n5898), .A4(n5899), .ZN(n5865)
         );
  NAND4_X1 U1600 ( .A1(n5887), .A2(n5888), .A3(n5889), .A4(n5890), .ZN(n5866)
         );
  NOR2_X1 U1601 ( .A1(n3278), .A2(n4421), .ZN(N8745) );
  NOR4_X1 U1602 ( .A1(n4422), .A2(n4423), .A3(n4424), .A4(n4425), .ZN(n4421)
         );
  NAND4_X1 U1603 ( .A1(n4453), .A2(n4454), .A3(n4455), .A4(n4456), .ZN(n4422)
         );
  NAND4_X1 U1604 ( .A1(n4444), .A2(n4445), .A3(n4446), .A4(n4447), .ZN(n4423)
         );
  NOR2_X1 U1605 ( .A1(n3268), .A2(n5823), .ZN(N8713) );
  NOR4_X1 U1606 ( .A1(n5824), .A2(n5825), .A3(n5826), .A4(n5827), .ZN(n5823)
         );
  NAND4_X1 U1607 ( .A1(n5855), .A2(n5856), .A3(n5857), .A4(n5858), .ZN(n5824)
         );
  NAND4_X1 U1608 ( .A1(n5846), .A2(n5847), .A3(n5848), .A4(n5849), .ZN(n5825)
         );
  NOR2_X1 U1609 ( .A1(n3278), .A2(n4380), .ZN(N8746) );
  NOR4_X1 U1610 ( .A1(n4381), .A2(n4382), .A3(n4383), .A4(n4384), .ZN(n4380)
         );
  NAND4_X1 U1611 ( .A1(n4412), .A2(n4413), .A3(n4414), .A4(n4415), .ZN(n4381)
         );
  NAND4_X1 U1612 ( .A1(n4403), .A2(n4404), .A3(n4405), .A4(n4406), .ZN(n4382)
         );
  NOR2_X1 U1613 ( .A1(n3268), .A2(n5782), .ZN(N8714) );
  NOR4_X1 U1614 ( .A1(n5783), .A2(n5784), .A3(n5785), .A4(n5786), .ZN(n5782)
         );
  NAND4_X1 U1615 ( .A1(n5814), .A2(n5815), .A3(n5816), .A4(n5817), .ZN(n5783)
         );
  NAND4_X1 U1616 ( .A1(n5805), .A2(n5806), .A3(n5807), .A4(n5808), .ZN(n5784)
         );
  NOR2_X1 U1617 ( .A1(n3280), .A2(n4339), .ZN(N8747) );
  NOR4_X1 U1618 ( .A1(n4340), .A2(n4341), .A3(n4342), .A4(n4343), .ZN(n4339)
         );
  NAND4_X1 U1619 ( .A1(n4371), .A2(n4372), .A3(n4373), .A4(n4374), .ZN(n4340)
         );
  NAND4_X1 U1620 ( .A1(n4362), .A2(n4363), .A3(n4364), .A4(n4365), .ZN(n4341)
         );
  NOR2_X1 U1621 ( .A1(n3269), .A2(n5741), .ZN(N8715) );
  NOR4_X1 U1622 ( .A1(n5742), .A2(n5743), .A3(n5744), .A4(n5745), .ZN(n5741)
         );
  NAND4_X1 U1623 ( .A1(n5773), .A2(n5774), .A3(n5775), .A4(n5776), .ZN(n5742)
         );
  NAND4_X1 U1624 ( .A1(n5764), .A2(n5765), .A3(n5766), .A4(n5767), .ZN(n5743)
         );
  NOR2_X1 U1625 ( .A1(n3280), .A2(n4298), .ZN(N8748) );
  NOR4_X1 U1626 ( .A1(n4299), .A2(n4300), .A3(n4301), .A4(n4302), .ZN(n4298)
         );
  NAND4_X1 U1627 ( .A1(n4330), .A2(n4331), .A3(n4332), .A4(n4333), .ZN(n4299)
         );
  NAND4_X1 U1628 ( .A1(n4321), .A2(n4322), .A3(n4323), .A4(n4324), .ZN(n4300)
         );
  NOR2_X1 U1629 ( .A1(n3269), .A2(n5700), .ZN(N8716) );
  NOR4_X1 U1630 ( .A1(n5701), .A2(n5702), .A3(n5703), .A4(n5704), .ZN(n5700)
         );
  NAND4_X1 U1631 ( .A1(n5732), .A2(n5733), .A3(n5734), .A4(n5735), .ZN(n5701)
         );
  NAND4_X1 U1632 ( .A1(n5723), .A2(n5724), .A3(n5725), .A4(n5726), .ZN(n5702)
         );
  NOR2_X1 U1633 ( .A1(n3280), .A2(n4257), .ZN(N8749) );
  NOR4_X1 U1634 ( .A1(n4258), .A2(n4259), .A3(n4260), .A4(n4261), .ZN(n4257)
         );
  NAND4_X1 U1635 ( .A1(n4289), .A2(n4290), .A3(n4291), .A4(n4292), .ZN(n4258)
         );
  NAND4_X1 U1636 ( .A1(n4280), .A2(n4281), .A3(n4282), .A4(n4283), .ZN(n4259)
         );
  NOR2_X1 U1637 ( .A1(n3269), .A2(n5659), .ZN(N8717) );
  NOR4_X1 U1638 ( .A1(n5660), .A2(n5661), .A3(n5662), .A4(n5663), .ZN(n5659)
         );
  NAND4_X1 U1639 ( .A1(n5691), .A2(n5692), .A3(n5693), .A4(n5694), .ZN(n5660)
         );
  NAND4_X1 U1640 ( .A1(n5682), .A2(n5683), .A3(n5684), .A4(n5685), .ZN(n5661)
         );
  NOR2_X1 U1641 ( .A1(n3280), .A2(n4216), .ZN(N8750) );
  NOR4_X1 U1642 ( .A1(n4217), .A2(n4218), .A3(n4219), .A4(n4220), .ZN(n4216)
         );
  NAND4_X1 U1643 ( .A1(n4248), .A2(n4249), .A3(n4250), .A4(n4251), .ZN(n4217)
         );
  NAND4_X1 U1644 ( .A1(n4239), .A2(n4240), .A3(n4241), .A4(n4242), .ZN(n4218)
         );
  NOR2_X1 U1645 ( .A1(n3269), .A2(n5618), .ZN(N8718) );
  NOR4_X1 U1646 ( .A1(n5619), .A2(n5620), .A3(n5621), .A4(n5622), .ZN(n5618)
         );
  NAND4_X1 U1647 ( .A1(n5650), .A2(n5651), .A3(n5652), .A4(n5653), .ZN(n5619)
         );
  NAND4_X1 U1648 ( .A1(n5641), .A2(n5642), .A3(n5643), .A4(n5644), .ZN(n5620)
         );
  NOR2_X1 U1649 ( .A1(n3281), .A2(n4175), .ZN(N8751) );
  NOR4_X1 U1650 ( .A1(n4176), .A2(n4177), .A3(n4178), .A4(n4179), .ZN(n4175)
         );
  NAND4_X1 U1651 ( .A1(n4207), .A2(n4208), .A3(n4209), .A4(n4210), .ZN(n4176)
         );
  NAND4_X1 U1652 ( .A1(n4198), .A2(n4199), .A3(n4200), .A4(n4201), .ZN(n4177)
         );
  NOR2_X1 U1653 ( .A1(n3270), .A2(n5577), .ZN(N8719) );
  NOR4_X1 U1654 ( .A1(n5578), .A2(n5579), .A3(n5580), .A4(n5581), .ZN(n5577)
         );
  NAND4_X1 U1655 ( .A1(n5609), .A2(n5610), .A3(n5611), .A4(n5612), .ZN(n5578)
         );
  NAND4_X1 U1656 ( .A1(n5600), .A2(n5601), .A3(n5602), .A4(n5603), .ZN(n5579)
         );
  NOR2_X1 U1657 ( .A1(n3281), .A2(n4134), .ZN(N8752) );
  NOR4_X1 U1658 ( .A1(n4135), .A2(n4136), .A3(n4137), .A4(n4138), .ZN(n4134)
         );
  NAND4_X1 U1659 ( .A1(n4166), .A2(n4167), .A3(n4168), .A4(n4169), .ZN(n4135)
         );
  NAND4_X1 U1660 ( .A1(n4157), .A2(n4158), .A3(n4159), .A4(n4160), .ZN(n4136)
         );
  NOR2_X1 U1661 ( .A1(n3270), .A2(n5536), .ZN(N8720) );
  NOR4_X1 U1662 ( .A1(n5537), .A2(n5538), .A3(n5539), .A4(n5540), .ZN(n5536)
         );
  NAND4_X1 U1663 ( .A1(n5568), .A2(n5569), .A3(n5570), .A4(n5571), .ZN(n5537)
         );
  NAND4_X1 U1664 ( .A1(n5559), .A2(n5560), .A3(n5561), .A4(n5562), .ZN(n5538)
         );
  NOR2_X1 U1665 ( .A1(n3281), .A2(n4093), .ZN(N8753) );
  NOR4_X1 U1666 ( .A1(n4094), .A2(n4095), .A3(n4096), .A4(n4097), .ZN(n4093)
         );
  NAND4_X1 U1667 ( .A1(n4125), .A2(n4126), .A3(n4127), .A4(n4128), .ZN(n4094)
         );
  NAND4_X1 U1668 ( .A1(n4116), .A2(n4117), .A3(n4118), .A4(n4119), .ZN(n4095)
         );
  NOR2_X1 U1669 ( .A1(n3270), .A2(n5495), .ZN(N8721) );
  NOR4_X1 U1670 ( .A1(n5496), .A2(n5497), .A3(n5498), .A4(n5499), .ZN(n5495)
         );
  NAND4_X1 U1671 ( .A1(n5527), .A2(n5528), .A3(n5529), .A4(n5530), .ZN(n5496)
         );
  NAND4_X1 U1672 ( .A1(n5518), .A2(n5519), .A3(n5520), .A4(n5521), .ZN(n5497)
         );
  NOR2_X1 U1673 ( .A1(n3281), .A2(n4052), .ZN(N8754) );
  NOR4_X1 U1674 ( .A1(n4053), .A2(n4054), .A3(n4055), .A4(n4056), .ZN(n4052)
         );
  NAND4_X1 U1675 ( .A1(n4084), .A2(n4085), .A3(n4086), .A4(n4087), .ZN(n4053)
         );
  NAND4_X1 U1676 ( .A1(n4075), .A2(n4076), .A3(n4077), .A4(n4078), .ZN(n4054)
         );
  NOR2_X1 U1677 ( .A1(n3270), .A2(n5454), .ZN(N8722) );
  NOR4_X1 U1678 ( .A1(n5455), .A2(n5456), .A3(n5457), .A4(n5458), .ZN(n5454)
         );
  NAND4_X1 U1679 ( .A1(n5486), .A2(n5487), .A3(n5488), .A4(n5489), .ZN(n5455)
         );
  NAND4_X1 U1680 ( .A1(n5477), .A2(n5478), .A3(n5479), .A4(n5480), .ZN(n5456)
         );
  NOR2_X1 U1681 ( .A1(n3282), .A2(n4011), .ZN(N8755) );
  NOR4_X1 U1682 ( .A1(n4012), .A2(n4013), .A3(n4014), .A4(n4015), .ZN(n4011)
         );
  NAND4_X1 U1683 ( .A1(n4043), .A2(n4044), .A3(n4045), .A4(n4046), .ZN(n4012)
         );
  NAND4_X1 U1684 ( .A1(n4034), .A2(n4035), .A3(n4036), .A4(n4037), .ZN(n4013)
         );
  NOR2_X1 U1685 ( .A1(n3272), .A2(n5413), .ZN(N8723) );
  NOR4_X1 U1686 ( .A1(n5414), .A2(n5415), .A3(n5416), .A4(n5417), .ZN(n5413)
         );
  NAND4_X1 U1687 ( .A1(n5445), .A2(n5446), .A3(n5447), .A4(n5448), .ZN(n5414)
         );
  NAND4_X1 U1688 ( .A1(n5436), .A2(n5437), .A3(n5438), .A4(n5439), .ZN(n5415)
         );
  NOR2_X1 U1689 ( .A1(n3282), .A2(n3970), .ZN(N8756) );
  NOR4_X1 U1690 ( .A1(n3971), .A2(n3972), .A3(n3973), .A4(n3974), .ZN(n3970)
         );
  NAND4_X1 U1691 ( .A1(n4002), .A2(n4003), .A3(n4004), .A4(n4005), .ZN(n3971)
         );
  NAND4_X1 U1692 ( .A1(n3993), .A2(n3994), .A3(n3995), .A4(n3996), .ZN(n3972)
         );
  NOR2_X1 U1693 ( .A1(n3272), .A2(n5372), .ZN(N8724) );
  NOR4_X1 U1694 ( .A1(n5373), .A2(n5374), .A3(n5375), .A4(n5376), .ZN(n5372)
         );
  NAND4_X1 U1695 ( .A1(n5404), .A2(n5405), .A3(n5406), .A4(n5407), .ZN(n5373)
         );
  NAND4_X1 U1696 ( .A1(n5395), .A2(n5396), .A3(n5397), .A4(n5398), .ZN(n5374)
         );
  NOR2_X1 U1697 ( .A1(n3282), .A2(n3929), .ZN(N8757) );
  NOR4_X1 U1698 ( .A1(n3930), .A2(n3931), .A3(n3932), .A4(n3933), .ZN(n3929)
         );
  NAND4_X1 U1699 ( .A1(n3961), .A2(n3962), .A3(n3963), .A4(n3964), .ZN(n3930)
         );
  NAND4_X1 U1700 ( .A1(n3952), .A2(n3953), .A3(n3954), .A4(n3955), .ZN(n3931)
         );
  NOR2_X1 U1701 ( .A1(n3272), .A2(n5331), .ZN(N8725) );
  NOR4_X1 U1702 ( .A1(n5332), .A2(n5333), .A3(n5334), .A4(n5335), .ZN(n5331)
         );
  NAND4_X1 U1703 ( .A1(n5363), .A2(n5364), .A3(n5365), .A4(n5366), .ZN(n5332)
         );
  NAND4_X1 U1704 ( .A1(n5354), .A2(n5355), .A3(n5356), .A4(n5357), .ZN(n5333)
         );
  NOR2_X1 U1705 ( .A1(n3282), .A2(n3888), .ZN(N8758) );
  NOR4_X1 U1706 ( .A1(n3889), .A2(n3890), .A3(n3891), .A4(n3892), .ZN(n3888)
         );
  NAND4_X1 U1707 ( .A1(n3920), .A2(n3921), .A3(n3922), .A4(n3923), .ZN(n3889)
         );
  NAND4_X1 U1708 ( .A1(n3911), .A2(n3912), .A3(n3913), .A4(n3914), .ZN(n3890)
         );
  NOR2_X1 U1709 ( .A1(n3272), .A2(n5290), .ZN(N8726) );
  NOR4_X1 U1710 ( .A1(n5291), .A2(n5292), .A3(n5293), .A4(n5294), .ZN(n5290)
         );
  NAND4_X1 U1711 ( .A1(n5322), .A2(n5323), .A3(n5324), .A4(n5325), .ZN(n5291)
         );
  NAND4_X1 U1712 ( .A1(n5313), .A2(n5314), .A3(n5315), .A4(n5316), .ZN(n5292)
         );
  NOR2_X1 U1713 ( .A1(n3284), .A2(n3847), .ZN(N8759) );
  NOR4_X1 U1714 ( .A1(n3848), .A2(n3849), .A3(n3850), .A4(n3851), .ZN(n3847)
         );
  NAND4_X1 U1715 ( .A1(n3879), .A2(n3880), .A3(n3881), .A4(n3882), .ZN(n3848)
         );
  NAND4_X1 U1716 ( .A1(n3870), .A2(n3871), .A3(n3872), .A4(n3873), .ZN(n3849)
         );
  NOR2_X1 U1717 ( .A1(n3273), .A2(n5249), .ZN(N8727) );
  NOR4_X1 U1718 ( .A1(n5250), .A2(n5251), .A3(n5252), .A4(n5253), .ZN(n5249)
         );
  NAND4_X1 U1719 ( .A1(n5281), .A2(n5282), .A3(n5283), .A4(n5284), .ZN(n5250)
         );
  NAND4_X1 U1720 ( .A1(n5272), .A2(n5273), .A3(n5274), .A4(n5275), .ZN(n5251)
         );
  NOR2_X1 U1721 ( .A1(n3284), .A2(n3806), .ZN(N8760) );
  NOR4_X1 U1722 ( .A1(n3807), .A2(n3808), .A3(n3809), .A4(n3810), .ZN(n3806)
         );
  NAND4_X1 U1723 ( .A1(n3838), .A2(n3839), .A3(n3840), .A4(n3841), .ZN(n3807)
         );
  NAND4_X1 U1724 ( .A1(n3829), .A2(n3830), .A3(n3831), .A4(n3832), .ZN(n3808)
         );
  NOR2_X1 U1725 ( .A1(n3273), .A2(n5208), .ZN(N8728) );
  NOR4_X1 U1726 ( .A1(n5209), .A2(n5210), .A3(n5211), .A4(n5212), .ZN(n5208)
         );
  NAND4_X1 U1727 ( .A1(n5240), .A2(n5241), .A3(n5242), .A4(n5243), .ZN(n5209)
         );
  NAND4_X1 U1728 ( .A1(n5231), .A2(n5232), .A3(n5233), .A4(n5234), .ZN(n5210)
         );
  NOR2_X1 U1729 ( .A1(n3284), .A2(n3765), .ZN(N8761) );
  NOR4_X1 U1730 ( .A1(n3766), .A2(n3767), .A3(n3768), .A4(n3769), .ZN(n3765)
         );
  NAND4_X1 U1731 ( .A1(n3797), .A2(n3798), .A3(n3799), .A4(n3800), .ZN(n3766)
         );
  NAND4_X1 U1732 ( .A1(n3788), .A2(n3789), .A3(n3790), .A4(n3791), .ZN(n3767)
         );
  NOR2_X1 U1733 ( .A1(n3273), .A2(n5167), .ZN(N8729) );
  NOR4_X1 U1734 ( .A1(n5168), .A2(n5169), .A3(n5170), .A4(n5171), .ZN(n5167)
         );
  NAND4_X1 U1735 ( .A1(n5199), .A2(n5200), .A3(n5201), .A4(n5202), .ZN(n5168)
         );
  NAND4_X1 U1736 ( .A1(n5190), .A2(n5191), .A3(n5192), .A4(n5193), .ZN(n5169)
         );
  NOR2_X1 U1737 ( .A1(n3284), .A2(n3724), .ZN(N8762) );
  NOR4_X1 U1738 ( .A1(n3725), .A2(n3726), .A3(n3727), .A4(n3728), .ZN(n3724)
         );
  NAND4_X1 U1739 ( .A1(n3756), .A2(n3757), .A3(n3758), .A4(n3759), .ZN(n3725)
         );
  NAND4_X1 U1740 ( .A1(n3747), .A2(n3748), .A3(n3749), .A4(n3750), .ZN(n3726)
         );
  NOR2_X1 U1741 ( .A1(n3273), .A2(n5126), .ZN(N8730) );
  NOR4_X1 U1742 ( .A1(n5127), .A2(n5128), .A3(n5129), .A4(n5130), .ZN(n5126)
         );
  NAND4_X1 U1743 ( .A1(n5158), .A2(n5159), .A3(n5160), .A4(n5161), .ZN(n5127)
         );
  NAND4_X1 U1744 ( .A1(n5149), .A2(n5150), .A3(n5151), .A4(n5152), .ZN(n5128)
         );
  NOR2_X1 U1745 ( .A1(n3285), .A2(n3683), .ZN(N8763) );
  NOR4_X1 U1746 ( .A1(n3684), .A2(n3685), .A3(n3686), .A4(n3687), .ZN(n3683)
         );
  NAND4_X1 U1747 ( .A1(n3715), .A2(n3716), .A3(n3717), .A4(n3718), .ZN(n3684)
         );
  NAND4_X1 U1748 ( .A1(n3706), .A2(n3707), .A3(n3708), .A4(n3709), .ZN(n3685)
         );
  NOR2_X1 U1749 ( .A1(n3274), .A2(n5085), .ZN(N8731) );
  NOR4_X1 U1750 ( .A1(n5086), .A2(n5087), .A3(n5088), .A4(n5089), .ZN(n5085)
         );
  NAND4_X1 U1751 ( .A1(n5117), .A2(n5118), .A3(n5119), .A4(n5120), .ZN(n5086)
         );
  NAND4_X1 U1752 ( .A1(n5108), .A2(n5109), .A3(n5110), .A4(n5111), .ZN(n5087)
         );
  NOR2_X1 U1753 ( .A1(n3285), .A2(n3642), .ZN(N8764) );
  NOR4_X1 U1754 ( .A1(n3643), .A2(n3644), .A3(n3645), .A4(n3646), .ZN(n3642)
         );
  NAND4_X1 U1755 ( .A1(n3674), .A2(n3675), .A3(n3676), .A4(n3677), .ZN(n3643)
         );
  NAND4_X1 U1756 ( .A1(n3665), .A2(n3666), .A3(n3667), .A4(n3668), .ZN(n3644)
         );
  NOR2_X1 U1757 ( .A1(n3274), .A2(n5044), .ZN(N8732) );
  NOR4_X1 U1758 ( .A1(n5045), .A2(n5046), .A3(n5047), .A4(n5048), .ZN(n5044)
         );
  NAND4_X1 U1759 ( .A1(n5076), .A2(n5077), .A3(n5078), .A4(n5079), .ZN(n5045)
         );
  NAND4_X1 U1760 ( .A1(n5067), .A2(n5068), .A3(n5069), .A4(n5070), .ZN(n5046)
         );
  NOR2_X1 U1761 ( .A1(n3285), .A2(n3601), .ZN(N8765) );
  NOR4_X1 U1762 ( .A1(n3602), .A2(n3603), .A3(n3604), .A4(n3605), .ZN(n3601)
         );
  NAND4_X1 U1763 ( .A1(n3633), .A2(n3634), .A3(n3635), .A4(n3636), .ZN(n3602)
         );
  NAND4_X1 U1764 ( .A1(n3624), .A2(n3625), .A3(n3626), .A4(n3627), .ZN(n3603)
         );
  NOR2_X1 U1765 ( .A1(n3274), .A2(n5003), .ZN(N8733) );
  NOR4_X1 U1766 ( .A1(n5004), .A2(n5005), .A3(n5006), .A4(n5007), .ZN(n5003)
         );
  NAND4_X1 U1767 ( .A1(n5035), .A2(n5036), .A3(n5037), .A4(n5038), .ZN(n5004)
         );
  NAND4_X1 U1768 ( .A1(n5026), .A2(n5027), .A3(n5028), .A4(n5029), .ZN(n5005)
         );
  NOR2_X1 U1769 ( .A1(n3285), .A2(n3560), .ZN(N8766) );
  NOR4_X1 U1770 ( .A1(n3561), .A2(n3562), .A3(n3563), .A4(n3564), .ZN(n3560)
         );
  NAND4_X1 U1771 ( .A1(n3592), .A2(n3593), .A3(n3594), .A4(n3595), .ZN(n3561)
         );
  NAND4_X1 U1772 ( .A1(n3583), .A2(n3584), .A3(n3585), .A4(n3586), .ZN(n3562)
         );
  NOR2_X1 U1773 ( .A1(n3274), .A2(n4874), .ZN(N8734) );
  NOR4_X1 U1774 ( .A1(n4875), .A2(n4876), .A3(n4877), .A4(n4878), .ZN(n4874)
         );
  NAND4_X1 U1775 ( .A1(n4972), .A2(n4973), .A3(n4974), .A4(n4975), .ZN(n4875)
         );
  NAND4_X1 U1776 ( .A1(n4941), .A2(n4942), .A3(n4943), .A4(n4944), .ZN(n4876)
         );
  NOR2_X1 U1777 ( .A1(n3276), .A2(n3431), .ZN(N8767) );
  NOR4_X1 U1778 ( .A1(n3432), .A2(n3433), .A3(n3434), .A4(n3435), .ZN(n3431)
         );
  NAND4_X1 U1779 ( .A1(n3529), .A2(n3530), .A3(n3531), .A4(n3532), .ZN(n3432)
         );
  NAND4_X1 U1780 ( .A1(n3498), .A2(n3499), .A3(n3500), .A4(n3501), .ZN(n3433)
         );
  OAI21_X1 U1781 ( .B1(n10920), .B2(n10921), .A(n3415), .ZN(n3416) );
  INV_X1 U1782 ( .A(ENABLE), .ZN(n10920) );
  NAND2_X1 U1783 ( .A1(CALL), .A2(ENABLE), .ZN(n3415) );
  AND3_X1 U1784 ( .A1(n3428), .A2(n10921), .A3(n3416), .ZN(n3420) );
  NAND2_X1 U1785 ( .A1(CWP[6]), .A2(n3429), .ZN(n3428) );
  AND3_X1 U1786 ( .A1(n3416), .A2(n3419), .A3(RETRN), .ZN(n3422) );
  OAI211_X1 U1787 ( .C1(n2898), .C2(n3416), .A(n3417), .B(n3418), .ZN(n9133)
         );
  OAI211_X1 U1788 ( .C1(n3392), .C2(N8834), .A(n3416), .B(RETRN), .ZN(n3418)
         );
  NAND2_X1 U1789 ( .A1(n2), .A2(n3420), .ZN(n3417) );
  XNOR2_X1 U1790 ( .A(CWP[6]), .B(\sub_189/carry[6] ), .ZN(N8834) );
  OAI21_X1 U1791 ( .B1(n3416), .B2(n2916), .A(n3421), .ZN(n9134) );
  AOI22_X1 U1792 ( .A1(N8833), .A2(n3422), .B1(n1), .B2(n3420), .ZN(n3421) );
  XNOR2_X1 U1793 ( .A(CWP[5]), .B(CWP[4]), .ZN(N8833) );
  OAI21_X1 U1794 ( .B1(n3416), .B2(N8791), .A(n3423), .ZN(n9135) );
  AOI22_X1 U1795 ( .A1(N8791), .A2(n3422), .B1(N8791), .B2(n3420), .ZN(n3423)
         );
  OAI21_X1 U1796 ( .B1(n3416), .B2(n2918), .A(n3424), .ZN(n9136) );
  AOI22_X1 U1797 ( .A1(N8790), .A2(n3422), .B1(N8790), .B2(n3420), .ZN(n3424)
         );
  OAI21_X1 U1798 ( .B1(n3416), .B2(n2919), .A(n3425), .ZN(n9137) );
  AOI22_X1 U1799 ( .A1(N8789), .A2(n3422), .B1(N8789), .B2(n3420), .ZN(n3425)
         );
  OAI21_X1 U1800 ( .B1(n3416), .B2(n2920), .A(n3426), .ZN(n9138) );
  AOI22_X1 U1801 ( .A1(N8788), .A2(n3422), .B1(N8788), .B2(n3420), .ZN(n3426)
         );
  OAI21_X1 U1802 ( .B1(n3416), .B2(n2921), .A(n3427), .ZN(n9139) );
  AOI22_X1 U1803 ( .A1(N8787), .A2(n3422), .B1(N8787), .B2(n3420), .ZN(n3427)
         );
  INV_X1 U1804 ( .A(RETRN), .ZN(n10921) );
  NAND2_X1 U1805 ( .A1(n3429), .A2(n2898), .ZN(n3419) );
  OR2_X1 U1806 ( .A1(CWP[5]), .A2(CWP[4]), .ZN(\sub_189/carry[6] ) );
  AND4_X1 U1807 ( .A1(n2920), .A2(n2919), .A3(n2921), .A4(n3430), .ZN(n3429)
         );
  NOR3_X1 U1808 ( .A1(N8790), .A2(CWP[5]), .A3(CWP[4]), .ZN(n3430) );
  XOR2_X1 U1809 ( .A(n2898), .B(n3), .Z(n2) );
  NAND2_X1 U1810 ( .A1(CWP[5]), .A2(CWP[4]), .ZN(n3) );
  AOI22_X1 U1811 ( .A1(N2164), .A2(n3391), .B1(N2157), .B2(N2151), .ZN(n3109)
         );
  XNOR2_X1 U1812 ( .A(ADD_WR[4]), .B(ADD_WR[3]), .ZN(N2164) );
  AOI22_X1 U1813 ( .A1(N8429), .A2(n10918), .B1(N8422), .B2(N8415), .ZN(n6264)
         );
  INV_X1 U1814 ( .A(N8430), .ZN(N8429) );
  AOI22_X1 U1815 ( .A1(N8573), .A2(n10919), .B1(N8566), .B2(N8559), .ZN(n4821)
         );
  INV_X1 U1816 ( .A(N8574), .ZN(N8573) );
  AOI22_X1 U1817 ( .A1(N8426), .A2(n10918), .B1(N8419), .B2(N8415), .ZN(n6315)
         );
  AOI22_X1 U1818 ( .A1(N8570), .A2(n10919), .B1(N8563), .B2(N8559), .ZN(n4872)
         );
  AOI22_X1 U1819 ( .A1(N8428), .A2(n10918), .B1(N8421), .B2(N8415), .ZN(n6265)
         );
  XNOR2_X1 U1820 ( .A(ADD_RD1[4]), .B(ADD_RD1[3]), .ZN(N8428) );
  AOI22_X1 U1821 ( .A1(N8572), .A2(n10919), .B1(N8565), .B2(N8559), .ZN(n4822)
         );
  XNOR2_X1 U1822 ( .A(ADD_RD2[4]), .B(ADD_RD2[3]), .ZN(N8572) );
  AOI22_X1 U1823 ( .A1(N8425), .A2(n10918), .B1(N8418), .B2(N8415), .ZN(n6314)
         );
  AOI22_X1 U1824 ( .A1(N8569), .A2(n10919), .B1(N8562), .B2(N8559), .ZN(n4871)
         );
  AOI22_X1 U1825 ( .A1(N8427), .A2(n10918), .B1(N8420), .B2(N8415), .ZN(n6280)
         );
  INV_X1 U1826 ( .A(ADD_RD1[3]), .ZN(N8427) );
  AOI22_X1 U1827 ( .A1(N8571), .A2(n10919), .B1(N8564), .B2(N8559), .ZN(n4837)
         );
  INV_X1 U1828 ( .A(ADD_RD2[3]), .ZN(N8571) );
  AOI22_X1 U1829 ( .A1(N8424), .A2(n10918), .B1(N8417), .B2(N8415), .ZN(n6278)
         );
  AOI22_X1 U1830 ( .A1(N8568), .A2(n10919), .B1(N8561), .B2(N8559), .ZN(n4835)
         );
  AOI222_X1 U1831 ( .A1(n668), .A2(\REGISTERS[19][0] ), .B1(n667), .B2(
        \REGISTERS[21][0] ), .C1(n664), .C2(\REGISTERS[20][0] ), .ZN(n6239) );
  AOI222_X1 U1832 ( .A1(n602), .A2(\REGISTERS[41][0] ), .B1(n601), .B2(
        \REGISTERS[43][0] ), .C1(n598), .C2(\REGISTERS[42][0] ), .ZN(n6270) );
  AOI222_X1 U1833 ( .A1(n440), .A2(\REGISTERS[52][0] ), .B1(n439), .B2(
        \REGISTERS[54][0] ), .C1(n436), .C2(\REGISTERS[53][0] ), .ZN(n6289) );
  AOI222_X1 U1834 ( .A1(n22), .A2(\REGISTERS[85][0] ), .B1(n21), .B2(
        \REGISTERS[87][0] ), .C1(n18), .C2(\REGISTERS[86][0] ), .ZN(n6302) );
  AOI222_X1 U1835 ( .A1(n1380), .A2(\REGISTERS[19][0] ), .B1(n1379), .B2(
        \REGISTERS[21][0] ), .C1(n1376), .C2(\REGISTERS[20][0] ), .ZN(n4796)
         );
  AOI222_X1 U1836 ( .A1(n1314), .A2(\REGISTERS[41][0] ), .B1(n1313), .B2(
        \REGISTERS[43][0] ), .C1(n1310), .C2(\REGISTERS[42][0] ), .ZN(n4827)
         );
  AOI222_X1 U1837 ( .A1(n1152), .A2(\REGISTERS[52][0] ), .B1(n1151), .B2(
        \REGISTERS[54][0] ), .C1(n1148), .C2(\REGISTERS[53][0] ), .ZN(n4846)
         );
  AOI222_X1 U1838 ( .A1(n734), .A2(\REGISTERS[85][0] ), .B1(n733), .B2(
        \REGISTERS[87][0] ), .C1(n730), .C2(\REGISTERS[86][0] ), .ZN(n4859) );
  AOI222_X1 U1839 ( .A1(n668), .A2(\REGISTERS[19][1] ), .B1(n667), .B2(
        \REGISTERS[21][1] ), .C1(n664), .C2(\REGISTERS[20][1] ), .ZN(n6198) );
  AOI222_X1 U1840 ( .A1(n602), .A2(\REGISTERS[41][1] ), .B1(n601), .B2(
        \REGISTERS[43][1] ), .C1(n598), .C2(\REGISTERS[42][1] ), .ZN(n6207) );
  AOI222_X1 U1841 ( .A1(n440), .A2(\REGISTERS[52][1] ), .B1(n439), .B2(
        \REGISTERS[54][1] ), .C1(n436), .C2(\REGISTERS[53][1] ), .ZN(n6216) );
  AOI222_X1 U1842 ( .A1(n22), .A2(\REGISTERS[85][1] ), .B1(n21), .B2(
        \REGISTERS[87][1] ), .C1(n18), .C2(\REGISTERS[86][1] ), .ZN(n6225) );
  AOI222_X1 U1843 ( .A1(n1380), .A2(\REGISTERS[19][1] ), .B1(n1379), .B2(
        \REGISTERS[21][1] ), .C1(n1376), .C2(\REGISTERS[20][1] ), .ZN(n4755)
         );
  AOI222_X1 U1844 ( .A1(n1314), .A2(\REGISTERS[41][1] ), .B1(n1313), .B2(
        \REGISTERS[43][1] ), .C1(n1310), .C2(\REGISTERS[42][1] ), .ZN(n4764)
         );
  AOI222_X1 U1845 ( .A1(n1152), .A2(\REGISTERS[52][1] ), .B1(n1151), .B2(
        \REGISTERS[54][1] ), .C1(n1148), .C2(\REGISTERS[53][1] ), .ZN(n4773)
         );
  AOI222_X1 U1846 ( .A1(n734), .A2(\REGISTERS[85][1] ), .B1(n733), .B2(
        \REGISTERS[87][1] ), .C1(n730), .C2(\REGISTERS[86][1] ), .ZN(n4782) );
  AOI222_X1 U1847 ( .A1(n668), .A2(\REGISTERS[19][2] ), .B1(n667), .B2(
        \REGISTERS[21][2] ), .C1(n664), .C2(\REGISTERS[20][2] ), .ZN(n6157) );
  AOI222_X1 U1848 ( .A1(n602), .A2(\REGISTERS[41][2] ), .B1(n601), .B2(
        \REGISTERS[43][2] ), .C1(n598), .C2(\REGISTERS[42][2] ), .ZN(n6166) );
  AOI222_X1 U1849 ( .A1(n440), .A2(\REGISTERS[52][2] ), .B1(n439), .B2(
        \REGISTERS[54][2] ), .C1(n436), .C2(\REGISTERS[53][2] ), .ZN(n6175) );
  AOI222_X1 U1850 ( .A1(n22), .A2(\REGISTERS[85][2] ), .B1(n21), .B2(
        \REGISTERS[87][2] ), .C1(n18), .C2(\REGISTERS[86][2] ), .ZN(n6184) );
  AOI222_X1 U1851 ( .A1(n1380), .A2(\REGISTERS[19][2] ), .B1(n1379), .B2(
        \REGISTERS[21][2] ), .C1(n1376), .C2(\REGISTERS[20][2] ), .ZN(n4714)
         );
  AOI222_X1 U1852 ( .A1(n1314), .A2(\REGISTERS[41][2] ), .B1(n1313), .B2(
        \REGISTERS[43][2] ), .C1(n1310), .C2(\REGISTERS[42][2] ), .ZN(n4723)
         );
  AOI222_X1 U1853 ( .A1(n1152), .A2(\REGISTERS[52][2] ), .B1(n1151), .B2(
        \REGISTERS[54][2] ), .C1(n1148), .C2(\REGISTERS[53][2] ), .ZN(n4732)
         );
  AOI222_X1 U1854 ( .A1(n734), .A2(\REGISTERS[85][2] ), .B1(n733), .B2(
        \REGISTERS[87][2] ), .C1(n730), .C2(\REGISTERS[86][2] ), .ZN(n4741) );
  AOI222_X1 U1855 ( .A1(n668), .A2(\REGISTERS[19][3] ), .B1(n667), .B2(
        \REGISTERS[21][3] ), .C1(n664), .C2(\REGISTERS[20][3] ), .ZN(n6116) );
  AOI222_X1 U1856 ( .A1(n602), .A2(\REGISTERS[41][3] ), .B1(n601), .B2(
        \REGISTERS[43][3] ), .C1(n598), .C2(\REGISTERS[42][3] ), .ZN(n6125) );
  AOI222_X1 U1857 ( .A1(n440), .A2(\REGISTERS[52][3] ), .B1(n439), .B2(
        \REGISTERS[54][3] ), .C1(n436), .C2(\REGISTERS[53][3] ), .ZN(n6134) );
  AOI222_X1 U1858 ( .A1(n22), .A2(\REGISTERS[85][3] ), .B1(n21), .B2(
        \REGISTERS[87][3] ), .C1(n18), .C2(\REGISTERS[86][3] ), .ZN(n6143) );
  AOI222_X1 U1859 ( .A1(n1380), .A2(\REGISTERS[19][3] ), .B1(n1379), .B2(
        \REGISTERS[21][3] ), .C1(n1376), .C2(\REGISTERS[20][3] ), .ZN(n4673)
         );
  AOI222_X1 U1860 ( .A1(n1314), .A2(\REGISTERS[41][3] ), .B1(n1313), .B2(
        \REGISTERS[43][3] ), .C1(n1310), .C2(\REGISTERS[42][3] ), .ZN(n4682)
         );
  AOI222_X1 U1861 ( .A1(n1152), .A2(\REGISTERS[52][3] ), .B1(n1151), .B2(
        \REGISTERS[54][3] ), .C1(n1148), .C2(\REGISTERS[53][3] ), .ZN(n4691)
         );
  AOI222_X1 U1862 ( .A1(n734), .A2(\REGISTERS[85][3] ), .B1(n733), .B2(
        \REGISTERS[87][3] ), .C1(n730), .C2(\REGISTERS[86][3] ), .ZN(n4700) );
  AOI222_X1 U1863 ( .A1(n668), .A2(\REGISTERS[19][4] ), .B1(n667), .B2(
        \REGISTERS[21][4] ), .C1(n664), .C2(\REGISTERS[20][4] ), .ZN(n6075) );
  AOI222_X1 U1864 ( .A1(n602), .A2(\REGISTERS[41][4] ), .B1(n601), .B2(
        \REGISTERS[43][4] ), .C1(n598), .C2(\REGISTERS[42][4] ), .ZN(n6084) );
  AOI222_X1 U1865 ( .A1(n440), .A2(\REGISTERS[52][4] ), .B1(n439), .B2(
        \REGISTERS[54][4] ), .C1(n436), .C2(\REGISTERS[53][4] ), .ZN(n6093) );
  AOI222_X1 U1866 ( .A1(n22), .A2(\REGISTERS[85][4] ), .B1(n21), .B2(
        \REGISTERS[87][4] ), .C1(n18), .C2(\REGISTERS[86][4] ), .ZN(n6102) );
  AOI222_X1 U1867 ( .A1(n1380), .A2(\REGISTERS[19][4] ), .B1(n1379), .B2(
        \REGISTERS[21][4] ), .C1(n1376), .C2(\REGISTERS[20][4] ), .ZN(n4632)
         );
  AOI222_X1 U1868 ( .A1(n1314), .A2(\REGISTERS[41][4] ), .B1(n1313), .B2(
        \REGISTERS[43][4] ), .C1(n1310), .C2(\REGISTERS[42][4] ), .ZN(n4641)
         );
  AOI222_X1 U1869 ( .A1(n1152), .A2(\REGISTERS[52][4] ), .B1(n1151), .B2(
        \REGISTERS[54][4] ), .C1(n1148), .C2(\REGISTERS[53][4] ), .ZN(n4650)
         );
  AOI222_X1 U1870 ( .A1(n734), .A2(\REGISTERS[85][4] ), .B1(n733), .B2(
        \REGISTERS[87][4] ), .C1(n730), .C2(\REGISTERS[86][4] ), .ZN(n4659) );
  AOI222_X1 U1871 ( .A1(n668), .A2(\REGISTERS[19][5] ), .B1(n667), .B2(
        \REGISTERS[21][5] ), .C1(n664), .C2(\REGISTERS[20][5] ), .ZN(n6034) );
  AOI222_X1 U1872 ( .A1(n602), .A2(\REGISTERS[41][5] ), .B1(n601), .B2(
        \REGISTERS[43][5] ), .C1(n598), .C2(\REGISTERS[42][5] ), .ZN(n6043) );
  AOI222_X1 U1873 ( .A1(n440), .A2(\REGISTERS[52][5] ), .B1(n439), .B2(
        \REGISTERS[54][5] ), .C1(n436), .C2(\REGISTERS[53][5] ), .ZN(n6052) );
  AOI222_X1 U1874 ( .A1(n22), .A2(\REGISTERS[85][5] ), .B1(n21), .B2(
        \REGISTERS[87][5] ), .C1(n18), .C2(\REGISTERS[86][5] ), .ZN(n6061) );
  AOI222_X1 U1875 ( .A1(n1380), .A2(\REGISTERS[19][5] ), .B1(n1379), .B2(
        \REGISTERS[21][5] ), .C1(n1376), .C2(\REGISTERS[20][5] ), .ZN(n4591)
         );
  AOI222_X1 U1876 ( .A1(n1314), .A2(\REGISTERS[41][5] ), .B1(n1313), .B2(
        \REGISTERS[43][5] ), .C1(n1310), .C2(\REGISTERS[42][5] ), .ZN(n4600)
         );
  AOI222_X1 U1877 ( .A1(n1152), .A2(\REGISTERS[52][5] ), .B1(n1151), .B2(
        \REGISTERS[54][5] ), .C1(n1148), .C2(\REGISTERS[53][5] ), .ZN(n4609)
         );
  AOI222_X1 U1878 ( .A1(n734), .A2(\REGISTERS[85][5] ), .B1(n733), .B2(
        \REGISTERS[87][5] ), .C1(n730), .C2(\REGISTERS[86][5] ), .ZN(n4618) );
  AOI222_X1 U1879 ( .A1(n668), .A2(\REGISTERS[19][6] ), .B1(n667), .B2(
        \REGISTERS[21][6] ), .C1(n664), .C2(\REGISTERS[20][6] ), .ZN(n5993) );
  AOI222_X1 U1880 ( .A1(n602), .A2(\REGISTERS[41][6] ), .B1(n601), .B2(
        \REGISTERS[43][6] ), .C1(n598), .C2(\REGISTERS[42][6] ), .ZN(n6002) );
  AOI222_X1 U1881 ( .A1(n440), .A2(\REGISTERS[52][6] ), .B1(n439), .B2(
        \REGISTERS[54][6] ), .C1(n436), .C2(\REGISTERS[53][6] ), .ZN(n6011) );
  AOI222_X1 U1882 ( .A1(n22), .A2(\REGISTERS[85][6] ), .B1(n21), .B2(
        \REGISTERS[87][6] ), .C1(n18), .C2(\REGISTERS[86][6] ), .ZN(n6020) );
  AOI222_X1 U1883 ( .A1(n1380), .A2(\REGISTERS[19][6] ), .B1(n1379), .B2(
        \REGISTERS[21][6] ), .C1(n1376), .C2(\REGISTERS[20][6] ), .ZN(n4550)
         );
  AOI222_X1 U1884 ( .A1(n1314), .A2(\REGISTERS[41][6] ), .B1(n1313), .B2(
        \REGISTERS[43][6] ), .C1(n1310), .C2(\REGISTERS[42][6] ), .ZN(n4559)
         );
  AOI222_X1 U1885 ( .A1(n1152), .A2(\REGISTERS[52][6] ), .B1(n1151), .B2(
        \REGISTERS[54][6] ), .C1(n1148), .C2(\REGISTERS[53][6] ), .ZN(n4568)
         );
  AOI222_X1 U1886 ( .A1(n734), .A2(\REGISTERS[85][6] ), .B1(n733), .B2(
        \REGISTERS[87][6] ), .C1(n730), .C2(\REGISTERS[86][6] ), .ZN(n4577) );
  AOI222_X1 U1887 ( .A1(n668), .A2(\REGISTERS[19][7] ), .B1(n667), .B2(
        \REGISTERS[21][7] ), .C1(n664), .C2(\REGISTERS[20][7] ), .ZN(n5952) );
  AOI222_X1 U1888 ( .A1(n602), .A2(\REGISTERS[41][7] ), .B1(n601), .B2(
        \REGISTERS[43][7] ), .C1(n598), .C2(\REGISTERS[42][7] ), .ZN(n5961) );
  AOI222_X1 U1889 ( .A1(n440), .A2(\REGISTERS[52][7] ), .B1(n439), .B2(
        \REGISTERS[54][7] ), .C1(n436), .C2(\REGISTERS[53][7] ), .ZN(n5970) );
  AOI222_X1 U1890 ( .A1(n22), .A2(\REGISTERS[85][7] ), .B1(n21), .B2(
        \REGISTERS[87][7] ), .C1(n18), .C2(\REGISTERS[86][7] ), .ZN(n5979) );
  AOI222_X1 U1891 ( .A1(n1380), .A2(\REGISTERS[19][7] ), .B1(n1379), .B2(
        \REGISTERS[21][7] ), .C1(n1376), .C2(\REGISTERS[20][7] ), .ZN(n4509)
         );
  AOI222_X1 U1892 ( .A1(n1314), .A2(\REGISTERS[41][7] ), .B1(n1313), .B2(
        \REGISTERS[43][7] ), .C1(n1310), .C2(\REGISTERS[42][7] ), .ZN(n4518)
         );
  AOI222_X1 U1893 ( .A1(n1152), .A2(\REGISTERS[52][7] ), .B1(n1151), .B2(
        \REGISTERS[54][7] ), .C1(n1148), .C2(\REGISTERS[53][7] ), .ZN(n4527)
         );
  AOI222_X1 U1894 ( .A1(n734), .A2(\REGISTERS[85][7] ), .B1(n733), .B2(
        \REGISTERS[87][7] ), .C1(n730), .C2(\REGISTERS[86][7] ), .ZN(n4536) );
  AOI222_X1 U1895 ( .A1(n668), .A2(\REGISTERS[19][8] ), .B1(n666), .B2(
        \REGISTERS[21][8] ), .C1(n663), .C2(\REGISTERS[20][8] ), .ZN(n5911) );
  AOI222_X1 U1896 ( .A1(n602), .A2(\REGISTERS[41][8] ), .B1(n600), .B2(
        \REGISTERS[43][8] ), .C1(n597), .C2(\REGISTERS[42][8] ), .ZN(n5920) );
  AOI222_X1 U1897 ( .A1(n440), .A2(\REGISTERS[52][8] ), .B1(n438), .B2(
        \REGISTERS[54][8] ), .C1(n435), .C2(\REGISTERS[53][8] ), .ZN(n5929) );
  AOI222_X1 U1898 ( .A1(n22), .A2(\REGISTERS[85][8] ), .B1(n20), .B2(
        \REGISTERS[87][8] ), .C1(n16), .C2(\REGISTERS[86][8] ), .ZN(n5938) );
  AOI222_X1 U1899 ( .A1(n1380), .A2(\REGISTERS[19][8] ), .B1(n1378), .B2(
        \REGISTERS[21][8] ), .C1(n1375), .C2(\REGISTERS[20][8] ), .ZN(n4468)
         );
  AOI222_X1 U1900 ( .A1(n1314), .A2(\REGISTERS[41][8] ), .B1(n1312), .B2(
        \REGISTERS[43][8] ), .C1(n1309), .C2(\REGISTERS[42][8] ), .ZN(n4477)
         );
  AOI222_X1 U1901 ( .A1(n1152), .A2(\REGISTERS[52][8] ), .B1(n1150), .B2(
        \REGISTERS[54][8] ), .C1(n1147), .C2(\REGISTERS[53][8] ), .ZN(n4486)
         );
  AOI222_X1 U1902 ( .A1(n734), .A2(\REGISTERS[85][8] ), .B1(n732), .B2(
        \REGISTERS[87][8] ), .C1(n729), .C2(\REGISTERS[86][8] ), .ZN(n4495) );
  AOI222_X1 U1903 ( .A1(n668), .A2(\REGISTERS[19][9] ), .B1(n666), .B2(
        \REGISTERS[21][9] ), .C1(n663), .C2(\REGISTERS[20][9] ), .ZN(n5870) );
  AOI222_X1 U1904 ( .A1(n602), .A2(\REGISTERS[41][9] ), .B1(n600), .B2(
        \REGISTERS[43][9] ), .C1(n597), .C2(\REGISTERS[42][9] ), .ZN(n5879) );
  AOI222_X1 U1905 ( .A1(n440), .A2(\REGISTERS[52][9] ), .B1(n438), .B2(
        \REGISTERS[54][9] ), .C1(n435), .C2(\REGISTERS[53][9] ), .ZN(n5888) );
  AOI222_X1 U1906 ( .A1(n22), .A2(\REGISTERS[85][9] ), .B1(n20), .B2(
        \REGISTERS[87][9] ), .C1(n16), .C2(\REGISTERS[86][9] ), .ZN(n5897) );
  AOI222_X1 U1907 ( .A1(n1380), .A2(\REGISTERS[19][9] ), .B1(n1378), .B2(
        \REGISTERS[21][9] ), .C1(n1375), .C2(\REGISTERS[20][9] ), .ZN(n4427)
         );
  AOI222_X1 U1908 ( .A1(n1314), .A2(\REGISTERS[41][9] ), .B1(n1312), .B2(
        \REGISTERS[43][9] ), .C1(n1309), .C2(\REGISTERS[42][9] ), .ZN(n4436)
         );
  AOI222_X1 U1909 ( .A1(n1152), .A2(\REGISTERS[52][9] ), .B1(n1150), .B2(
        \REGISTERS[54][9] ), .C1(n1147), .C2(\REGISTERS[53][9] ), .ZN(n4445)
         );
  AOI222_X1 U1910 ( .A1(n734), .A2(\REGISTERS[85][9] ), .B1(n732), .B2(
        \REGISTERS[87][9] ), .C1(n729), .C2(\REGISTERS[86][9] ), .ZN(n4454) );
  AOI222_X1 U1911 ( .A1(n668), .A2(\REGISTERS[19][10] ), .B1(n666), .B2(
        \REGISTERS[21][10] ), .C1(n663), .C2(\REGISTERS[20][10] ), .ZN(n5829)
         );
  AOI222_X1 U1912 ( .A1(n602), .A2(\REGISTERS[41][10] ), .B1(n600), .B2(
        \REGISTERS[43][10] ), .C1(n597), .C2(\REGISTERS[42][10] ), .ZN(n5838)
         );
  AOI222_X1 U1913 ( .A1(n440), .A2(\REGISTERS[52][10] ), .B1(n438), .B2(
        \REGISTERS[54][10] ), .C1(n435), .C2(\REGISTERS[53][10] ), .ZN(n5847)
         );
  AOI222_X1 U1914 ( .A1(n22), .A2(\REGISTERS[85][10] ), .B1(n20), .B2(
        \REGISTERS[87][10] ), .C1(n16), .C2(\REGISTERS[86][10] ), .ZN(n5856)
         );
  AOI222_X1 U1915 ( .A1(n1380), .A2(\REGISTERS[19][10] ), .B1(n1378), .B2(
        \REGISTERS[21][10] ), .C1(n1375), .C2(\REGISTERS[20][10] ), .ZN(n4386)
         );
  AOI222_X1 U1916 ( .A1(n1314), .A2(\REGISTERS[41][10] ), .B1(n1312), .B2(
        \REGISTERS[43][10] ), .C1(n1309), .C2(\REGISTERS[42][10] ), .ZN(n4395)
         );
  AOI222_X1 U1917 ( .A1(n1152), .A2(\REGISTERS[52][10] ), .B1(n1150), .B2(
        \REGISTERS[54][10] ), .C1(n1147), .C2(\REGISTERS[53][10] ), .ZN(n4404)
         );
  AOI222_X1 U1918 ( .A1(n734), .A2(\REGISTERS[85][10] ), .B1(n732), .B2(
        \REGISTERS[87][10] ), .C1(n729), .C2(\REGISTERS[86][10] ), .ZN(n4413)
         );
  AOI222_X1 U1919 ( .A1(n668), .A2(\REGISTERS[19][11] ), .B1(n666), .B2(
        \REGISTERS[21][11] ), .C1(n663), .C2(\REGISTERS[20][11] ), .ZN(n5788)
         );
  AOI222_X1 U1920 ( .A1(n602), .A2(\REGISTERS[41][11] ), .B1(n600), .B2(
        \REGISTERS[43][11] ), .C1(n597), .C2(\REGISTERS[42][11] ), .ZN(n5797)
         );
  AOI222_X1 U1921 ( .A1(n440), .A2(\REGISTERS[52][11] ), .B1(n438), .B2(
        \REGISTERS[54][11] ), .C1(n435), .C2(\REGISTERS[53][11] ), .ZN(n5806)
         );
  AOI222_X1 U1922 ( .A1(n22), .A2(\REGISTERS[85][11] ), .B1(n20), .B2(
        \REGISTERS[87][11] ), .C1(n16), .C2(\REGISTERS[86][11] ), .ZN(n5815)
         );
  AOI222_X1 U1923 ( .A1(n1380), .A2(\REGISTERS[19][11] ), .B1(n1378), .B2(
        \REGISTERS[21][11] ), .C1(n1375), .C2(\REGISTERS[20][11] ), .ZN(n4345)
         );
  AOI222_X1 U1924 ( .A1(n1314), .A2(\REGISTERS[41][11] ), .B1(n1312), .B2(
        \REGISTERS[43][11] ), .C1(n1309), .C2(\REGISTERS[42][11] ), .ZN(n4354)
         );
  AOI222_X1 U1925 ( .A1(n1152), .A2(\REGISTERS[52][11] ), .B1(n1150), .B2(
        \REGISTERS[54][11] ), .C1(n1147), .C2(\REGISTERS[53][11] ), .ZN(n4363)
         );
  AOI222_X1 U1926 ( .A1(n734), .A2(\REGISTERS[85][11] ), .B1(n732), .B2(
        \REGISTERS[87][11] ), .C1(n729), .C2(\REGISTERS[86][11] ), .ZN(n4372)
         );
  AOI222_X1 U1927 ( .A1(n669), .A2(\REGISTERS[19][12] ), .B1(n666), .B2(
        \REGISTERS[21][12] ), .C1(n663), .C2(\REGISTERS[20][12] ), .ZN(n5747)
         );
  AOI222_X1 U1928 ( .A1(n603), .A2(\REGISTERS[41][12] ), .B1(n600), .B2(
        \REGISTERS[43][12] ), .C1(n597), .C2(\REGISTERS[42][12] ), .ZN(n5756)
         );
  AOI222_X1 U1929 ( .A1(n441), .A2(\REGISTERS[52][12] ), .B1(n438), .B2(
        \REGISTERS[54][12] ), .C1(n435), .C2(\REGISTERS[53][12] ), .ZN(n5765)
         );
  AOI222_X1 U1930 ( .A1(n23), .A2(\REGISTERS[85][12] ), .B1(n20), .B2(
        \REGISTERS[87][12] ), .C1(n16), .C2(\REGISTERS[86][12] ), .ZN(n5774)
         );
  AOI222_X1 U1931 ( .A1(n1381), .A2(\REGISTERS[19][12] ), .B1(n1378), .B2(
        \REGISTERS[21][12] ), .C1(n1375), .C2(\REGISTERS[20][12] ), .ZN(n4304)
         );
  AOI222_X1 U1932 ( .A1(n1315), .A2(\REGISTERS[41][12] ), .B1(n1312), .B2(
        \REGISTERS[43][12] ), .C1(n1309), .C2(\REGISTERS[42][12] ), .ZN(n4313)
         );
  AOI222_X1 U1933 ( .A1(n1153), .A2(\REGISTERS[52][12] ), .B1(n1150), .B2(
        \REGISTERS[54][12] ), .C1(n1147), .C2(\REGISTERS[53][12] ), .ZN(n4322)
         );
  AOI222_X1 U1934 ( .A1(n735), .A2(\REGISTERS[85][12] ), .B1(n732), .B2(
        \REGISTERS[87][12] ), .C1(n729), .C2(\REGISTERS[86][12] ), .ZN(n4331)
         );
  AOI222_X1 U1935 ( .A1(n669), .A2(\REGISTERS[19][13] ), .B1(n666), .B2(
        \REGISTERS[21][13] ), .C1(n663), .C2(\REGISTERS[20][13] ), .ZN(n5706)
         );
  AOI222_X1 U1936 ( .A1(n603), .A2(\REGISTERS[41][13] ), .B1(n600), .B2(
        \REGISTERS[43][13] ), .C1(n597), .C2(\REGISTERS[42][13] ), .ZN(n5715)
         );
  AOI222_X1 U1937 ( .A1(n441), .A2(\REGISTERS[52][13] ), .B1(n438), .B2(
        \REGISTERS[54][13] ), .C1(n435), .C2(\REGISTERS[53][13] ), .ZN(n5724)
         );
  AOI222_X1 U1938 ( .A1(n23), .A2(\REGISTERS[85][13] ), .B1(n20), .B2(
        \REGISTERS[87][13] ), .C1(n16), .C2(\REGISTERS[86][13] ), .ZN(n5733)
         );
  AOI222_X1 U1939 ( .A1(n1381), .A2(\REGISTERS[19][13] ), .B1(n1378), .B2(
        \REGISTERS[21][13] ), .C1(n1375), .C2(\REGISTERS[20][13] ), .ZN(n4263)
         );
  AOI222_X1 U1940 ( .A1(n1315), .A2(\REGISTERS[41][13] ), .B1(n1312), .B2(
        \REGISTERS[43][13] ), .C1(n1309), .C2(\REGISTERS[42][13] ), .ZN(n4272)
         );
  AOI222_X1 U1941 ( .A1(n1153), .A2(\REGISTERS[52][13] ), .B1(n1150), .B2(
        \REGISTERS[54][13] ), .C1(n1147), .C2(\REGISTERS[53][13] ), .ZN(n4281)
         );
  AOI222_X1 U1942 ( .A1(n735), .A2(\REGISTERS[85][13] ), .B1(n732), .B2(
        \REGISTERS[87][13] ), .C1(n729), .C2(\REGISTERS[86][13] ), .ZN(n4290)
         );
  AOI222_X1 U1943 ( .A1(n669), .A2(\REGISTERS[19][14] ), .B1(n666), .B2(
        \REGISTERS[21][14] ), .C1(n663), .C2(\REGISTERS[20][14] ), .ZN(n5665)
         );
  AOI222_X1 U1944 ( .A1(n603), .A2(\REGISTERS[41][14] ), .B1(n600), .B2(
        \REGISTERS[43][14] ), .C1(n597), .C2(\REGISTERS[42][14] ), .ZN(n5674)
         );
  AOI222_X1 U1945 ( .A1(n441), .A2(\REGISTERS[52][14] ), .B1(n438), .B2(
        \REGISTERS[54][14] ), .C1(n435), .C2(\REGISTERS[53][14] ), .ZN(n5683)
         );
  AOI222_X1 U1946 ( .A1(n23), .A2(\REGISTERS[85][14] ), .B1(n20), .B2(
        \REGISTERS[87][14] ), .C1(n16), .C2(\REGISTERS[86][14] ), .ZN(n5692)
         );
  AOI222_X1 U1947 ( .A1(n1381), .A2(\REGISTERS[19][14] ), .B1(n1378), .B2(
        \REGISTERS[21][14] ), .C1(n1375), .C2(\REGISTERS[20][14] ), .ZN(n4222)
         );
  AOI222_X1 U1948 ( .A1(n1315), .A2(\REGISTERS[41][14] ), .B1(n1312), .B2(
        \REGISTERS[43][14] ), .C1(n1309), .C2(\REGISTERS[42][14] ), .ZN(n4231)
         );
  AOI222_X1 U1949 ( .A1(n1153), .A2(\REGISTERS[52][14] ), .B1(n1150), .B2(
        \REGISTERS[54][14] ), .C1(n1147), .C2(\REGISTERS[53][14] ), .ZN(n4240)
         );
  AOI222_X1 U1950 ( .A1(n735), .A2(\REGISTERS[85][14] ), .B1(n732), .B2(
        \REGISTERS[87][14] ), .C1(n729), .C2(\REGISTERS[86][14] ), .ZN(n4249)
         );
  AOI222_X1 U1951 ( .A1(n669), .A2(\REGISTERS[19][15] ), .B1(n666), .B2(
        \REGISTERS[21][15] ), .C1(n663), .C2(\REGISTERS[20][15] ), .ZN(n5624)
         );
  AOI222_X1 U1952 ( .A1(n603), .A2(\REGISTERS[41][15] ), .B1(n600), .B2(
        \REGISTERS[43][15] ), .C1(n597), .C2(\REGISTERS[42][15] ), .ZN(n5633)
         );
  AOI222_X1 U1953 ( .A1(n441), .A2(\REGISTERS[52][15] ), .B1(n438), .B2(
        \REGISTERS[54][15] ), .C1(n435), .C2(\REGISTERS[53][15] ), .ZN(n5642)
         );
  AOI222_X1 U1954 ( .A1(n23), .A2(\REGISTERS[85][15] ), .B1(n20), .B2(
        \REGISTERS[87][15] ), .C1(n16), .C2(\REGISTERS[86][15] ), .ZN(n5651)
         );
  AOI222_X1 U1955 ( .A1(n1381), .A2(\REGISTERS[19][15] ), .B1(n1378), .B2(
        \REGISTERS[21][15] ), .C1(n1375), .C2(\REGISTERS[20][15] ), .ZN(n4181)
         );
  AOI222_X1 U1956 ( .A1(n1315), .A2(\REGISTERS[41][15] ), .B1(n1312), .B2(
        \REGISTERS[43][15] ), .C1(n1309), .C2(\REGISTERS[42][15] ), .ZN(n4190)
         );
  AOI222_X1 U1957 ( .A1(n1153), .A2(\REGISTERS[52][15] ), .B1(n1150), .B2(
        \REGISTERS[54][15] ), .C1(n1147), .C2(\REGISTERS[53][15] ), .ZN(n4199)
         );
  AOI222_X1 U1958 ( .A1(n735), .A2(\REGISTERS[85][15] ), .B1(n732), .B2(
        \REGISTERS[87][15] ), .C1(n729), .C2(\REGISTERS[86][15] ), .ZN(n4208)
         );
  AOI222_X1 U1959 ( .A1(n669), .A2(\REGISTERS[19][16] ), .B1(n666), .B2(
        \REGISTERS[21][16] ), .C1(n663), .C2(\REGISTERS[20][16] ), .ZN(n5583)
         );
  AOI222_X1 U1960 ( .A1(n603), .A2(\REGISTERS[41][16] ), .B1(n600), .B2(
        \REGISTERS[43][16] ), .C1(n597), .C2(\REGISTERS[42][16] ), .ZN(n5592)
         );
  AOI222_X1 U1961 ( .A1(n441), .A2(\REGISTERS[52][16] ), .B1(n438), .B2(
        \REGISTERS[54][16] ), .C1(n435), .C2(\REGISTERS[53][16] ), .ZN(n5601)
         );
  AOI222_X1 U1962 ( .A1(n23), .A2(\REGISTERS[85][16] ), .B1(n20), .B2(
        \REGISTERS[87][16] ), .C1(n16), .C2(\REGISTERS[86][16] ), .ZN(n5610)
         );
  AOI222_X1 U1963 ( .A1(n1381), .A2(\REGISTERS[19][16] ), .B1(n1378), .B2(
        \REGISTERS[21][16] ), .C1(n1375), .C2(\REGISTERS[20][16] ), .ZN(n4140)
         );
  AOI222_X1 U1964 ( .A1(n1315), .A2(\REGISTERS[41][16] ), .B1(n1312), .B2(
        \REGISTERS[43][16] ), .C1(n1309), .C2(\REGISTERS[42][16] ), .ZN(n4149)
         );
  AOI222_X1 U1965 ( .A1(n1153), .A2(\REGISTERS[52][16] ), .B1(n1150), .B2(
        \REGISTERS[54][16] ), .C1(n1147), .C2(\REGISTERS[53][16] ), .ZN(n4158)
         );
  AOI222_X1 U1966 ( .A1(n735), .A2(\REGISTERS[85][16] ), .B1(n732), .B2(
        \REGISTERS[87][16] ), .C1(n729), .C2(\REGISTERS[86][16] ), .ZN(n4167)
         );
  AOI222_X1 U1967 ( .A1(n669), .A2(\REGISTERS[19][17] ), .B1(n666), .B2(
        \REGISTERS[21][17] ), .C1(n663), .C2(\REGISTERS[20][17] ), .ZN(n5542)
         );
  AOI222_X1 U1968 ( .A1(n603), .A2(\REGISTERS[41][17] ), .B1(n600), .B2(
        \REGISTERS[43][17] ), .C1(n597), .C2(\REGISTERS[42][17] ), .ZN(n5551)
         );
  AOI222_X1 U1969 ( .A1(n441), .A2(\REGISTERS[52][17] ), .B1(n438), .B2(
        \REGISTERS[54][17] ), .C1(n435), .C2(\REGISTERS[53][17] ), .ZN(n5560)
         );
  AOI222_X1 U1970 ( .A1(n23), .A2(\REGISTERS[85][17] ), .B1(n20), .B2(
        \REGISTERS[87][17] ), .C1(n16), .C2(\REGISTERS[86][17] ), .ZN(n5569)
         );
  AOI222_X1 U1971 ( .A1(n1381), .A2(\REGISTERS[19][17] ), .B1(n1378), .B2(
        \REGISTERS[21][17] ), .C1(n1375), .C2(\REGISTERS[20][17] ), .ZN(n4099)
         );
  AOI222_X1 U1972 ( .A1(n1315), .A2(\REGISTERS[41][17] ), .B1(n1312), .B2(
        \REGISTERS[43][17] ), .C1(n1309), .C2(\REGISTERS[42][17] ), .ZN(n4108)
         );
  AOI222_X1 U1973 ( .A1(n1153), .A2(\REGISTERS[52][17] ), .B1(n1150), .B2(
        \REGISTERS[54][17] ), .C1(n1147), .C2(\REGISTERS[53][17] ), .ZN(n4117)
         );
  AOI222_X1 U1974 ( .A1(n735), .A2(\REGISTERS[85][17] ), .B1(n732), .B2(
        \REGISTERS[87][17] ), .C1(n729), .C2(\REGISTERS[86][17] ), .ZN(n4126)
         );
  AOI222_X1 U1975 ( .A1(n669), .A2(\REGISTERS[19][18] ), .B1(n666), .B2(
        \REGISTERS[21][18] ), .C1(n663), .C2(\REGISTERS[20][18] ), .ZN(n5501)
         );
  AOI222_X1 U1976 ( .A1(n603), .A2(\REGISTERS[41][18] ), .B1(n600), .B2(
        \REGISTERS[43][18] ), .C1(n597), .C2(\REGISTERS[42][18] ), .ZN(n5510)
         );
  AOI222_X1 U1977 ( .A1(n441), .A2(\REGISTERS[52][18] ), .B1(n438), .B2(
        \REGISTERS[54][18] ), .C1(n435), .C2(\REGISTERS[53][18] ), .ZN(n5519)
         );
  AOI222_X1 U1978 ( .A1(n23), .A2(\REGISTERS[85][18] ), .B1(n20), .B2(
        \REGISTERS[87][18] ), .C1(n16), .C2(\REGISTERS[86][18] ), .ZN(n5528)
         );
  AOI222_X1 U1979 ( .A1(n1381), .A2(\REGISTERS[19][18] ), .B1(n1378), .B2(
        \REGISTERS[21][18] ), .C1(n1375), .C2(\REGISTERS[20][18] ), .ZN(n4058)
         );
  AOI222_X1 U1980 ( .A1(n1315), .A2(\REGISTERS[41][18] ), .B1(n1312), .B2(
        \REGISTERS[43][18] ), .C1(n1309), .C2(\REGISTERS[42][18] ), .ZN(n4067)
         );
  AOI222_X1 U1981 ( .A1(n1153), .A2(\REGISTERS[52][18] ), .B1(n1150), .B2(
        \REGISTERS[54][18] ), .C1(n1147), .C2(\REGISTERS[53][18] ), .ZN(n4076)
         );
  AOI222_X1 U1982 ( .A1(n735), .A2(\REGISTERS[85][18] ), .B1(n732), .B2(
        \REGISTERS[87][18] ), .C1(n729), .C2(\REGISTERS[86][18] ), .ZN(n4085)
         );
  AOI222_X1 U1983 ( .A1(n669), .A2(\REGISTERS[19][19] ), .B1(n666), .B2(
        \REGISTERS[21][19] ), .C1(n663), .C2(\REGISTERS[20][19] ), .ZN(n5460)
         );
  AOI222_X1 U1984 ( .A1(n603), .A2(\REGISTERS[41][19] ), .B1(n600), .B2(
        \REGISTERS[43][19] ), .C1(n597), .C2(\REGISTERS[42][19] ), .ZN(n5469)
         );
  AOI222_X1 U1985 ( .A1(n441), .A2(\REGISTERS[52][19] ), .B1(n438), .B2(
        \REGISTERS[54][19] ), .C1(n435), .C2(\REGISTERS[53][19] ), .ZN(n5478)
         );
  AOI222_X1 U1986 ( .A1(n23), .A2(\REGISTERS[85][19] ), .B1(n20), .B2(
        \REGISTERS[87][19] ), .C1(n16), .C2(\REGISTERS[86][19] ), .ZN(n5487)
         );
  AOI222_X1 U1987 ( .A1(n1381), .A2(\REGISTERS[19][19] ), .B1(n1378), .B2(
        \REGISTERS[21][19] ), .C1(n1375), .C2(\REGISTERS[20][19] ), .ZN(n4017)
         );
  AOI222_X1 U1988 ( .A1(n1315), .A2(\REGISTERS[41][19] ), .B1(n1312), .B2(
        \REGISTERS[43][19] ), .C1(n1309), .C2(\REGISTERS[42][19] ), .ZN(n4026)
         );
  AOI222_X1 U1989 ( .A1(n1153), .A2(\REGISTERS[52][19] ), .B1(n1150), .B2(
        \REGISTERS[54][19] ), .C1(n1147), .C2(\REGISTERS[53][19] ), .ZN(n4035)
         );
  AOI222_X1 U1990 ( .A1(n735), .A2(\REGISTERS[85][19] ), .B1(n732), .B2(
        \REGISTERS[87][19] ), .C1(n729), .C2(\REGISTERS[86][19] ), .ZN(n4044)
         );
  AOI222_X1 U1991 ( .A1(n669), .A2(\REGISTERS[19][20] ), .B1(n665), .B2(
        \REGISTERS[21][20] ), .C1(n662), .C2(\REGISTERS[20][20] ), .ZN(n5419)
         );
  AOI222_X1 U1992 ( .A1(n603), .A2(\REGISTERS[41][20] ), .B1(n599), .B2(
        \REGISTERS[43][20] ), .C1(n596), .C2(\REGISTERS[42][20] ), .ZN(n5428)
         );
  AOI222_X1 U1993 ( .A1(n441), .A2(\REGISTERS[52][20] ), .B1(n437), .B2(
        \REGISTERS[54][20] ), .C1(n434), .C2(\REGISTERS[53][20] ), .ZN(n5437)
         );
  AOI222_X1 U1994 ( .A1(n23), .A2(\REGISTERS[85][20] ), .B1(n19), .B2(
        \REGISTERS[87][20] ), .C1(n15), .C2(\REGISTERS[86][20] ), .ZN(n5446)
         );
  AOI222_X1 U1995 ( .A1(n1381), .A2(\REGISTERS[19][20] ), .B1(n1377), .B2(
        \REGISTERS[21][20] ), .C1(n1374), .C2(\REGISTERS[20][20] ), .ZN(n3976)
         );
  AOI222_X1 U1996 ( .A1(n1315), .A2(\REGISTERS[41][20] ), .B1(n1311), .B2(
        \REGISTERS[43][20] ), .C1(n1308), .C2(\REGISTERS[42][20] ), .ZN(n3985)
         );
  AOI222_X1 U1997 ( .A1(n1153), .A2(\REGISTERS[52][20] ), .B1(n1149), .B2(
        \REGISTERS[54][20] ), .C1(n1146), .C2(\REGISTERS[53][20] ), .ZN(n3994)
         );
  AOI222_X1 U1998 ( .A1(n735), .A2(\REGISTERS[85][20] ), .B1(n731), .B2(
        \REGISTERS[87][20] ), .C1(n728), .C2(\REGISTERS[86][20] ), .ZN(n4003)
         );
  AOI222_X1 U1999 ( .A1(n669), .A2(\REGISTERS[19][21] ), .B1(n665), .B2(
        \REGISTERS[21][21] ), .C1(n662), .C2(\REGISTERS[20][21] ), .ZN(n5378)
         );
  AOI222_X1 U2000 ( .A1(n603), .A2(\REGISTERS[41][21] ), .B1(n599), .B2(
        \REGISTERS[43][21] ), .C1(n596), .C2(\REGISTERS[42][21] ), .ZN(n5387)
         );
  AOI222_X1 U2001 ( .A1(n441), .A2(\REGISTERS[52][21] ), .B1(n437), .B2(
        \REGISTERS[54][21] ), .C1(n434), .C2(\REGISTERS[53][21] ), .ZN(n5396)
         );
  AOI222_X1 U2002 ( .A1(n23), .A2(\REGISTERS[85][21] ), .B1(n19), .B2(
        \REGISTERS[87][21] ), .C1(n15), .C2(\REGISTERS[86][21] ), .ZN(n5405)
         );
  AOI222_X1 U2003 ( .A1(n1381), .A2(\REGISTERS[19][21] ), .B1(n1377), .B2(
        \REGISTERS[21][21] ), .C1(n1374), .C2(\REGISTERS[20][21] ), .ZN(n3935)
         );
  AOI222_X1 U2004 ( .A1(n1315), .A2(\REGISTERS[41][21] ), .B1(n1311), .B2(
        \REGISTERS[43][21] ), .C1(n1308), .C2(\REGISTERS[42][21] ), .ZN(n3944)
         );
  AOI222_X1 U2005 ( .A1(n1153), .A2(\REGISTERS[52][21] ), .B1(n1149), .B2(
        \REGISTERS[54][21] ), .C1(n1146), .C2(\REGISTERS[53][21] ), .ZN(n3953)
         );
  AOI222_X1 U2006 ( .A1(n735), .A2(\REGISTERS[85][21] ), .B1(n731), .B2(
        \REGISTERS[87][21] ), .C1(n728), .C2(\REGISTERS[86][21] ), .ZN(n3962)
         );
  AOI222_X1 U2007 ( .A1(n669), .A2(\REGISTERS[19][22] ), .B1(n665), .B2(
        \REGISTERS[21][22] ), .C1(n662), .C2(\REGISTERS[20][22] ), .ZN(n5337)
         );
  AOI222_X1 U2008 ( .A1(n603), .A2(\REGISTERS[41][22] ), .B1(n599), .B2(
        \REGISTERS[43][22] ), .C1(n596), .C2(\REGISTERS[42][22] ), .ZN(n5346)
         );
  AOI222_X1 U2009 ( .A1(n441), .A2(\REGISTERS[52][22] ), .B1(n437), .B2(
        \REGISTERS[54][22] ), .C1(n434), .C2(\REGISTERS[53][22] ), .ZN(n5355)
         );
  AOI222_X1 U2010 ( .A1(n23), .A2(\REGISTERS[85][22] ), .B1(n19), .B2(
        \REGISTERS[87][22] ), .C1(n15), .C2(\REGISTERS[86][22] ), .ZN(n5364)
         );
  AOI222_X1 U2011 ( .A1(n1381), .A2(\REGISTERS[19][22] ), .B1(n1377), .B2(
        \REGISTERS[21][22] ), .C1(n1374), .C2(\REGISTERS[20][22] ), .ZN(n3894)
         );
  AOI222_X1 U2012 ( .A1(n1315), .A2(\REGISTERS[41][22] ), .B1(n1311), .B2(
        \REGISTERS[43][22] ), .C1(n1308), .C2(\REGISTERS[42][22] ), .ZN(n3903)
         );
  AOI222_X1 U2013 ( .A1(n1153), .A2(\REGISTERS[52][22] ), .B1(n1149), .B2(
        \REGISTERS[54][22] ), .C1(n1146), .C2(\REGISTERS[53][22] ), .ZN(n3912)
         );
  AOI222_X1 U2014 ( .A1(n735), .A2(\REGISTERS[85][22] ), .B1(n731), .B2(
        \REGISTERS[87][22] ), .C1(n728), .C2(\REGISTERS[86][22] ), .ZN(n3921)
         );
  AOI222_X1 U2015 ( .A1(n669), .A2(\REGISTERS[19][23] ), .B1(n665), .B2(
        \REGISTERS[21][23] ), .C1(n662), .C2(\REGISTERS[20][23] ), .ZN(n5296)
         );
  AOI222_X1 U2016 ( .A1(n603), .A2(\REGISTERS[41][23] ), .B1(n599), .B2(
        \REGISTERS[43][23] ), .C1(n596), .C2(\REGISTERS[42][23] ), .ZN(n5305)
         );
  AOI222_X1 U2017 ( .A1(n441), .A2(\REGISTERS[52][23] ), .B1(n437), .B2(
        \REGISTERS[54][23] ), .C1(n434), .C2(\REGISTERS[53][23] ), .ZN(n5314)
         );
  AOI222_X1 U2018 ( .A1(n23), .A2(\REGISTERS[85][23] ), .B1(n19), .B2(
        \REGISTERS[87][23] ), .C1(n15), .C2(\REGISTERS[86][23] ), .ZN(n5323)
         );
  AOI222_X1 U2019 ( .A1(n1381), .A2(\REGISTERS[19][23] ), .B1(n1377), .B2(
        \REGISTERS[21][23] ), .C1(n1374), .C2(\REGISTERS[20][23] ), .ZN(n3853)
         );
  AOI222_X1 U2020 ( .A1(n1315), .A2(\REGISTERS[41][23] ), .B1(n1311), .B2(
        \REGISTERS[43][23] ), .C1(n1308), .C2(\REGISTERS[42][23] ), .ZN(n3862)
         );
  AOI222_X1 U2021 ( .A1(n1153), .A2(\REGISTERS[52][23] ), .B1(n1149), .B2(
        \REGISTERS[54][23] ), .C1(n1146), .C2(\REGISTERS[53][23] ), .ZN(n3871)
         );
  AOI222_X1 U2022 ( .A1(n735), .A2(\REGISTERS[85][23] ), .B1(n731), .B2(
        \REGISTERS[87][23] ), .C1(n728), .C2(\REGISTERS[86][23] ), .ZN(n3880)
         );
  AOI222_X1 U2023 ( .A1(n670), .A2(\REGISTERS[19][24] ), .B1(n665), .B2(
        \REGISTERS[21][24] ), .C1(n662), .C2(\REGISTERS[20][24] ), .ZN(n5255)
         );
  AOI222_X1 U2024 ( .A1(n604), .A2(\REGISTERS[41][24] ), .B1(n599), .B2(
        \REGISTERS[43][24] ), .C1(n596), .C2(\REGISTERS[42][24] ), .ZN(n5264)
         );
  AOI222_X1 U2025 ( .A1(n442), .A2(\REGISTERS[52][24] ), .B1(n437), .B2(
        \REGISTERS[54][24] ), .C1(n434), .C2(\REGISTERS[53][24] ), .ZN(n5273)
         );
  AOI222_X1 U2026 ( .A1(n24), .A2(\REGISTERS[85][24] ), .B1(n19), .B2(
        \REGISTERS[87][24] ), .C1(n15), .C2(\REGISTERS[86][24] ), .ZN(n5282)
         );
  AOI222_X1 U2027 ( .A1(n1382), .A2(\REGISTERS[19][24] ), .B1(n1377), .B2(
        \REGISTERS[21][24] ), .C1(n1374), .C2(\REGISTERS[20][24] ), .ZN(n3812)
         );
  AOI222_X1 U2028 ( .A1(n1316), .A2(\REGISTERS[41][24] ), .B1(n1311), .B2(
        \REGISTERS[43][24] ), .C1(n1308), .C2(\REGISTERS[42][24] ), .ZN(n3821)
         );
  AOI222_X1 U2029 ( .A1(n1154), .A2(\REGISTERS[52][24] ), .B1(n1149), .B2(
        \REGISTERS[54][24] ), .C1(n1146), .C2(\REGISTERS[53][24] ), .ZN(n3830)
         );
  AOI222_X1 U2030 ( .A1(n736), .A2(\REGISTERS[85][24] ), .B1(n731), .B2(
        \REGISTERS[87][24] ), .C1(n728), .C2(\REGISTERS[86][24] ), .ZN(n3839)
         );
  AOI222_X1 U2031 ( .A1(n670), .A2(\REGISTERS[19][25] ), .B1(n665), .B2(
        \REGISTERS[21][25] ), .C1(n662), .C2(\REGISTERS[20][25] ), .ZN(n5214)
         );
  AOI222_X1 U2032 ( .A1(n604), .A2(\REGISTERS[41][25] ), .B1(n599), .B2(
        \REGISTERS[43][25] ), .C1(n596), .C2(\REGISTERS[42][25] ), .ZN(n5223)
         );
  AOI222_X1 U2033 ( .A1(n442), .A2(\REGISTERS[52][25] ), .B1(n437), .B2(
        \REGISTERS[54][25] ), .C1(n434), .C2(\REGISTERS[53][25] ), .ZN(n5232)
         );
  AOI222_X1 U2034 ( .A1(n24), .A2(\REGISTERS[85][25] ), .B1(n19), .B2(
        \REGISTERS[87][25] ), .C1(n15), .C2(\REGISTERS[86][25] ), .ZN(n5241)
         );
  AOI222_X1 U2035 ( .A1(n1382), .A2(\REGISTERS[19][25] ), .B1(n1377), .B2(
        \REGISTERS[21][25] ), .C1(n1374), .C2(\REGISTERS[20][25] ), .ZN(n3771)
         );
  AOI222_X1 U2036 ( .A1(n1316), .A2(\REGISTERS[41][25] ), .B1(n1311), .B2(
        \REGISTERS[43][25] ), .C1(n1308), .C2(\REGISTERS[42][25] ), .ZN(n3780)
         );
  AOI222_X1 U2037 ( .A1(n1154), .A2(\REGISTERS[52][25] ), .B1(n1149), .B2(
        \REGISTERS[54][25] ), .C1(n1146), .C2(\REGISTERS[53][25] ), .ZN(n3789)
         );
  AOI222_X1 U2038 ( .A1(n736), .A2(\REGISTERS[85][25] ), .B1(n731), .B2(
        \REGISTERS[87][25] ), .C1(n728), .C2(\REGISTERS[86][25] ), .ZN(n3798)
         );
  AOI222_X1 U2039 ( .A1(n670), .A2(\REGISTERS[19][26] ), .B1(n665), .B2(
        \REGISTERS[21][26] ), .C1(n662), .C2(\REGISTERS[20][26] ), .ZN(n5173)
         );
  AOI222_X1 U2040 ( .A1(n604), .A2(\REGISTERS[41][26] ), .B1(n599), .B2(
        \REGISTERS[43][26] ), .C1(n596), .C2(\REGISTERS[42][26] ), .ZN(n5182)
         );
  AOI222_X1 U2041 ( .A1(n442), .A2(\REGISTERS[52][26] ), .B1(n437), .B2(
        \REGISTERS[54][26] ), .C1(n434), .C2(\REGISTERS[53][26] ), .ZN(n5191)
         );
  AOI222_X1 U2042 ( .A1(n24), .A2(\REGISTERS[85][26] ), .B1(n19), .B2(
        \REGISTERS[87][26] ), .C1(n15), .C2(\REGISTERS[86][26] ), .ZN(n5200)
         );
  AOI222_X1 U2043 ( .A1(n1382), .A2(\REGISTERS[19][26] ), .B1(n1377), .B2(
        \REGISTERS[21][26] ), .C1(n1374), .C2(\REGISTERS[20][26] ), .ZN(n3730)
         );
  AOI222_X1 U2044 ( .A1(n1316), .A2(\REGISTERS[41][26] ), .B1(n1311), .B2(
        \REGISTERS[43][26] ), .C1(n1308), .C2(\REGISTERS[42][26] ), .ZN(n3739)
         );
  AOI222_X1 U2045 ( .A1(n1154), .A2(\REGISTERS[52][26] ), .B1(n1149), .B2(
        \REGISTERS[54][26] ), .C1(n1146), .C2(\REGISTERS[53][26] ), .ZN(n3748)
         );
  AOI222_X1 U2046 ( .A1(n736), .A2(\REGISTERS[85][26] ), .B1(n731), .B2(
        \REGISTERS[87][26] ), .C1(n728), .C2(\REGISTERS[86][26] ), .ZN(n3757)
         );
  AOI222_X1 U2047 ( .A1(n670), .A2(\REGISTERS[19][27] ), .B1(n665), .B2(
        \REGISTERS[21][27] ), .C1(n662), .C2(\REGISTERS[20][27] ), .ZN(n5132)
         );
  AOI222_X1 U2048 ( .A1(n604), .A2(\REGISTERS[41][27] ), .B1(n599), .B2(
        \REGISTERS[43][27] ), .C1(n596), .C2(\REGISTERS[42][27] ), .ZN(n5141)
         );
  AOI222_X1 U2049 ( .A1(n442), .A2(\REGISTERS[52][27] ), .B1(n437), .B2(
        \REGISTERS[54][27] ), .C1(n434), .C2(\REGISTERS[53][27] ), .ZN(n5150)
         );
  AOI222_X1 U2050 ( .A1(n24), .A2(\REGISTERS[85][27] ), .B1(n19), .B2(
        \REGISTERS[87][27] ), .C1(n15), .C2(\REGISTERS[86][27] ), .ZN(n5159)
         );
  AOI222_X1 U2051 ( .A1(n1382), .A2(\REGISTERS[19][27] ), .B1(n1377), .B2(
        \REGISTERS[21][27] ), .C1(n1374), .C2(\REGISTERS[20][27] ), .ZN(n3689)
         );
  AOI222_X1 U2052 ( .A1(n1316), .A2(\REGISTERS[41][27] ), .B1(n1311), .B2(
        \REGISTERS[43][27] ), .C1(n1308), .C2(\REGISTERS[42][27] ), .ZN(n3698)
         );
  AOI222_X1 U2053 ( .A1(n1154), .A2(\REGISTERS[52][27] ), .B1(n1149), .B2(
        \REGISTERS[54][27] ), .C1(n1146), .C2(\REGISTERS[53][27] ), .ZN(n3707)
         );
  AOI222_X1 U2054 ( .A1(n736), .A2(\REGISTERS[85][27] ), .B1(n731), .B2(
        \REGISTERS[87][27] ), .C1(n728), .C2(\REGISTERS[86][27] ), .ZN(n3716)
         );
  AOI222_X1 U2055 ( .A1(n670), .A2(\REGISTERS[19][28] ), .B1(n665), .B2(
        \REGISTERS[21][28] ), .C1(n662), .C2(\REGISTERS[20][28] ), .ZN(n5091)
         );
  AOI222_X1 U2056 ( .A1(n604), .A2(\REGISTERS[41][28] ), .B1(n599), .B2(
        \REGISTERS[43][28] ), .C1(n596), .C2(\REGISTERS[42][28] ), .ZN(n5100)
         );
  AOI222_X1 U2057 ( .A1(n442), .A2(\REGISTERS[52][28] ), .B1(n437), .B2(
        \REGISTERS[54][28] ), .C1(n434), .C2(\REGISTERS[53][28] ), .ZN(n5109)
         );
  AOI222_X1 U2058 ( .A1(n24), .A2(\REGISTERS[85][28] ), .B1(n19), .B2(
        \REGISTERS[87][28] ), .C1(n15), .C2(\REGISTERS[86][28] ), .ZN(n5118)
         );
  AOI222_X1 U2059 ( .A1(n1382), .A2(\REGISTERS[19][28] ), .B1(n1377), .B2(
        \REGISTERS[21][28] ), .C1(n1374), .C2(\REGISTERS[20][28] ), .ZN(n3648)
         );
  AOI222_X1 U2060 ( .A1(n1316), .A2(\REGISTERS[41][28] ), .B1(n1311), .B2(
        \REGISTERS[43][28] ), .C1(n1308), .C2(\REGISTERS[42][28] ), .ZN(n3657)
         );
  AOI222_X1 U2061 ( .A1(n1154), .A2(\REGISTERS[52][28] ), .B1(n1149), .B2(
        \REGISTERS[54][28] ), .C1(n1146), .C2(\REGISTERS[53][28] ), .ZN(n3666)
         );
  AOI222_X1 U2062 ( .A1(n736), .A2(\REGISTERS[85][28] ), .B1(n731), .B2(
        \REGISTERS[87][28] ), .C1(n728), .C2(\REGISTERS[86][28] ), .ZN(n3675)
         );
  AOI222_X1 U2063 ( .A1(n670), .A2(\REGISTERS[19][29] ), .B1(n665), .B2(
        \REGISTERS[21][29] ), .C1(n662), .C2(\REGISTERS[20][29] ), .ZN(n5050)
         );
  AOI222_X1 U2064 ( .A1(n604), .A2(\REGISTERS[41][29] ), .B1(n599), .B2(
        \REGISTERS[43][29] ), .C1(n596), .C2(\REGISTERS[42][29] ), .ZN(n5059)
         );
  AOI222_X1 U2065 ( .A1(n442), .A2(\REGISTERS[52][29] ), .B1(n437), .B2(
        \REGISTERS[54][29] ), .C1(n434), .C2(\REGISTERS[53][29] ), .ZN(n5068)
         );
  AOI222_X1 U2066 ( .A1(n24), .A2(\REGISTERS[85][29] ), .B1(n19), .B2(
        \REGISTERS[87][29] ), .C1(n15), .C2(\REGISTERS[86][29] ), .ZN(n5077)
         );
  AOI222_X1 U2067 ( .A1(n1382), .A2(\REGISTERS[19][29] ), .B1(n1377), .B2(
        \REGISTERS[21][29] ), .C1(n1374), .C2(\REGISTERS[20][29] ), .ZN(n3607)
         );
  AOI222_X1 U2068 ( .A1(n1316), .A2(\REGISTERS[41][29] ), .B1(n1311), .B2(
        \REGISTERS[43][29] ), .C1(n1308), .C2(\REGISTERS[42][29] ), .ZN(n3616)
         );
  AOI222_X1 U2069 ( .A1(n1154), .A2(\REGISTERS[52][29] ), .B1(n1149), .B2(
        \REGISTERS[54][29] ), .C1(n1146), .C2(\REGISTERS[53][29] ), .ZN(n3625)
         );
  AOI222_X1 U2070 ( .A1(n736), .A2(\REGISTERS[85][29] ), .B1(n731), .B2(
        \REGISTERS[87][29] ), .C1(n728), .C2(\REGISTERS[86][29] ), .ZN(n3634)
         );
  AOI222_X1 U2071 ( .A1(n670), .A2(\REGISTERS[19][30] ), .B1(n665), .B2(
        \REGISTERS[21][30] ), .C1(n662), .C2(\REGISTERS[20][30] ), .ZN(n5009)
         );
  AOI222_X1 U2072 ( .A1(n604), .A2(\REGISTERS[41][30] ), .B1(n599), .B2(
        \REGISTERS[43][30] ), .C1(n596), .C2(\REGISTERS[42][30] ), .ZN(n5018)
         );
  AOI222_X1 U2073 ( .A1(n442), .A2(\REGISTERS[52][30] ), .B1(n437), .B2(
        \REGISTERS[54][30] ), .C1(n434), .C2(\REGISTERS[53][30] ), .ZN(n5027)
         );
  AOI222_X1 U2074 ( .A1(n24), .A2(\REGISTERS[85][30] ), .B1(n19), .B2(
        \REGISTERS[87][30] ), .C1(n15), .C2(\REGISTERS[86][30] ), .ZN(n5036)
         );
  AOI222_X1 U2075 ( .A1(n1382), .A2(\REGISTERS[19][30] ), .B1(n1377), .B2(
        \REGISTERS[21][30] ), .C1(n1374), .C2(\REGISTERS[20][30] ), .ZN(n3566)
         );
  AOI222_X1 U2076 ( .A1(n1316), .A2(\REGISTERS[41][30] ), .B1(n1311), .B2(
        \REGISTERS[43][30] ), .C1(n1308), .C2(\REGISTERS[42][30] ), .ZN(n3575)
         );
  AOI222_X1 U2077 ( .A1(n1154), .A2(\REGISTERS[52][30] ), .B1(n1149), .B2(
        \REGISTERS[54][30] ), .C1(n1146), .C2(\REGISTERS[53][30] ), .ZN(n3584)
         );
  AOI222_X1 U2078 ( .A1(n736), .A2(\REGISTERS[85][30] ), .B1(n731), .B2(
        \REGISTERS[87][30] ), .C1(n728), .C2(\REGISTERS[86][30] ), .ZN(n3593)
         );
  AOI222_X1 U2079 ( .A1(n670), .A2(\REGISTERS[19][31] ), .B1(n665), .B2(
        \REGISTERS[21][31] ), .C1(n662), .C2(\REGISTERS[20][31] ), .ZN(n4880)
         );
  AOI222_X1 U2080 ( .A1(n604), .A2(\REGISTERS[41][31] ), .B1(n599), .B2(
        \REGISTERS[43][31] ), .C1(n596), .C2(\REGISTERS[42][31] ), .ZN(n4911)
         );
  AOI222_X1 U2081 ( .A1(n442), .A2(\REGISTERS[52][31] ), .B1(n437), .B2(
        \REGISTERS[54][31] ), .C1(n434), .C2(\REGISTERS[53][31] ), .ZN(n4942)
         );
  AOI222_X1 U2082 ( .A1(n24), .A2(\REGISTERS[85][31] ), .B1(n19), .B2(
        \REGISTERS[87][31] ), .C1(n15), .C2(\REGISTERS[86][31] ), .ZN(n4973)
         );
  AOI222_X1 U2083 ( .A1(n1382), .A2(\REGISTERS[19][31] ), .B1(n1377), .B2(
        \REGISTERS[21][31] ), .C1(n1374), .C2(\REGISTERS[20][31] ), .ZN(n3437)
         );
  AOI222_X1 U2084 ( .A1(n1316), .A2(\REGISTERS[41][31] ), .B1(n1311), .B2(
        \REGISTERS[43][31] ), .C1(n1308), .C2(\REGISTERS[42][31] ), .ZN(n3468)
         );
  AOI222_X1 U2085 ( .A1(n1154), .A2(\REGISTERS[52][31] ), .B1(n1149), .B2(
        \REGISTERS[54][31] ), .C1(n1146), .C2(\REGISTERS[53][31] ), .ZN(n3499)
         );
  AOI222_X1 U2086 ( .A1(n736), .A2(\REGISTERS[85][31] ), .B1(n731), .B2(
        \REGISTERS[87][31] ), .C1(n728), .C2(\REGISTERS[86][31] ), .ZN(n3530)
         );
  OAI222_X1 U2087 ( .A1(n207), .A2(n710), .B1(n239), .B2(n707), .C1(n175), 
        .C2(n704), .ZN(n6244) );
  OAI222_X1 U2088 ( .A1(n911), .A2(n644), .B1(n943), .B2(n641), .C1(n879), 
        .C2(n638), .ZN(n6275) );
  OAI222_X1 U2089 ( .A1(n1967), .A2(n482), .B1(n1999), .B2(n479), .C1(n1935), 
        .C2(n476), .ZN(n6294) );
  OAI222_X1 U2090 ( .A1(n2319), .A2(n64), .B1(n2351), .B2(n61), .C1(n2287), 
        .C2(n58), .ZN(n6307) );
  OAI222_X1 U2091 ( .A1(n207), .A2(n1422), .B1(n239), .B2(n1419), .C1(n175), 
        .C2(n1416), .ZN(n4801) );
  OAI222_X1 U2092 ( .A1(n911), .A2(n1356), .B1(n943), .B2(n1353), .C1(n879), 
        .C2(n1350), .ZN(n4832) );
  OAI222_X1 U2093 ( .A1(n1967), .A2(n1194), .B1(n1999), .B2(n1191), .C1(n1935), 
        .C2(n1188), .ZN(n4851) );
  OAI222_X1 U2094 ( .A1(n2319), .A2(n776), .B1(n2351), .B2(n773), .C1(n2287), 
        .C2(n770), .ZN(n4864) );
  OAI222_X1 U2095 ( .A1(n206), .A2(n710), .B1(n238), .B2(n707), .C1(n174), 
        .C2(n704), .ZN(n6203) );
  OAI222_X1 U2096 ( .A1(n910), .A2(n644), .B1(n942), .B2(n641), .C1(n878), 
        .C2(n638), .ZN(n6212) );
  OAI222_X1 U2097 ( .A1(n1966), .A2(n482), .B1(n1998), .B2(n479), .C1(n1934), 
        .C2(n476), .ZN(n6221) );
  OAI222_X1 U2098 ( .A1(n2318), .A2(n64), .B1(n2350), .B2(n61), .C1(n2286), 
        .C2(n58), .ZN(n6230) );
  OAI222_X1 U2099 ( .A1(n206), .A2(n1422), .B1(n238), .B2(n1419), .C1(n174), 
        .C2(n1416), .ZN(n4760) );
  OAI222_X1 U2100 ( .A1(n910), .A2(n1356), .B1(n942), .B2(n1353), .C1(n878), 
        .C2(n1350), .ZN(n4769) );
  OAI222_X1 U2101 ( .A1(n1966), .A2(n1194), .B1(n1998), .B2(n1191), .C1(n1934), 
        .C2(n1188), .ZN(n4778) );
  OAI222_X1 U2102 ( .A1(n2318), .A2(n776), .B1(n2350), .B2(n773), .C1(n2286), 
        .C2(n770), .ZN(n4787) );
  OAI222_X1 U2103 ( .A1(n205), .A2(n710), .B1(n237), .B2(n707), .C1(n173), 
        .C2(n704), .ZN(n6162) );
  OAI222_X1 U2104 ( .A1(n909), .A2(n644), .B1(n941), .B2(n641), .C1(n877), 
        .C2(n638), .ZN(n6171) );
  OAI222_X1 U2105 ( .A1(n1965), .A2(n482), .B1(n1997), .B2(n479), .C1(n1933), 
        .C2(n476), .ZN(n6180) );
  OAI222_X1 U2106 ( .A1(n2317), .A2(n64), .B1(n2349), .B2(n61), .C1(n2285), 
        .C2(n58), .ZN(n6189) );
  OAI222_X1 U2107 ( .A1(n205), .A2(n1422), .B1(n237), .B2(n1419), .C1(n173), 
        .C2(n1416), .ZN(n4719) );
  OAI222_X1 U2108 ( .A1(n909), .A2(n1356), .B1(n941), .B2(n1353), .C1(n877), 
        .C2(n1350), .ZN(n4728) );
  OAI222_X1 U2109 ( .A1(n1965), .A2(n1194), .B1(n1997), .B2(n1191), .C1(n1933), 
        .C2(n1188), .ZN(n4737) );
  OAI222_X1 U2110 ( .A1(n2317), .A2(n776), .B1(n2349), .B2(n773), .C1(n2285), 
        .C2(n770), .ZN(n4746) );
  OAI222_X1 U2111 ( .A1(n204), .A2(n710), .B1(n236), .B2(n707), .C1(n172), 
        .C2(n704), .ZN(n6121) );
  OAI222_X1 U2112 ( .A1(n908), .A2(n644), .B1(n940), .B2(n641), .C1(n876), 
        .C2(n638), .ZN(n6130) );
  OAI222_X1 U2113 ( .A1(n1964), .A2(n482), .B1(n1996), .B2(n479), .C1(n1932), 
        .C2(n476), .ZN(n6139) );
  OAI222_X1 U2114 ( .A1(n2316), .A2(n64), .B1(n2348), .B2(n61), .C1(n2284), 
        .C2(n58), .ZN(n6148) );
  OAI222_X1 U2115 ( .A1(n204), .A2(n1422), .B1(n236), .B2(n1419), .C1(n172), 
        .C2(n1416), .ZN(n4678) );
  OAI222_X1 U2116 ( .A1(n908), .A2(n1356), .B1(n940), .B2(n1353), .C1(n876), 
        .C2(n1350), .ZN(n4687) );
  OAI222_X1 U2117 ( .A1(n1964), .A2(n1194), .B1(n1996), .B2(n1191), .C1(n1932), 
        .C2(n1188), .ZN(n4696) );
  OAI222_X1 U2118 ( .A1(n2316), .A2(n776), .B1(n2348), .B2(n773), .C1(n2284), 
        .C2(n770), .ZN(n4705) );
  OAI222_X1 U2119 ( .A1(n203), .A2(n710), .B1(n235), .B2(n707), .C1(n171), 
        .C2(n704), .ZN(n6080) );
  OAI222_X1 U2120 ( .A1(n907), .A2(n644), .B1(n939), .B2(n641), .C1(n875), 
        .C2(n638), .ZN(n6089) );
  OAI222_X1 U2121 ( .A1(n1963), .A2(n482), .B1(n1995), .B2(n479), .C1(n1931), 
        .C2(n476), .ZN(n6098) );
  OAI222_X1 U2122 ( .A1(n2315), .A2(n64), .B1(n2347), .B2(n61), .C1(n2283), 
        .C2(n58), .ZN(n6107) );
  OAI222_X1 U2123 ( .A1(n203), .A2(n1422), .B1(n235), .B2(n1419), .C1(n171), 
        .C2(n1416), .ZN(n4637) );
  OAI222_X1 U2124 ( .A1(n907), .A2(n1356), .B1(n939), .B2(n1353), .C1(n875), 
        .C2(n1350), .ZN(n4646) );
  OAI222_X1 U2125 ( .A1(n1963), .A2(n1194), .B1(n1995), .B2(n1191), .C1(n1931), 
        .C2(n1188), .ZN(n4655) );
  OAI222_X1 U2126 ( .A1(n2315), .A2(n776), .B1(n2347), .B2(n773), .C1(n2283), 
        .C2(n770), .ZN(n4664) );
  OAI222_X1 U2127 ( .A1(n202), .A2(n710), .B1(n234), .B2(n707), .C1(n170), 
        .C2(n704), .ZN(n6039) );
  OAI222_X1 U2128 ( .A1(n906), .A2(n644), .B1(n938), .B2(n641), .C1(n874), 
        .C2(n638), .ZN(n6048) );
  OAI222_X1 U2129 ( .A1(n1962), .A2(n482), .B1(n1994), .B2(n479), .C1(n1930), 
        .C2(n476), .ZN(n6057) );
  OAI222_X1 U2130 ( .A1(n2314), .A2(n64), .B1(n2346), .B2(n61), .C1(n2282), 
        .C2(n58), .ZN(n6066) );
  OAI222_X1 U2131 ( .A1(n202), .A2(n1422), .B1(n234), .B2(n1419), .C1(n170), 
        .C2(n1416), .ZN(n4596) );
  OAI222_X1 U2132 ( .A1(n906), .A2(n1356), .B1(n938), .B2(n1353), .C1(n874), 
        .C2(n1350), .ZN(n4605) );
  OAI222_X1 U2133 ( .A1(n1962), .A2(n1194), .B1(n1994), .B2(n1191), .C1(n1930), 
        .C2(n1188), .ZN(n4614) );
  OAI222_X1 U2134 ( .A1(n2314), .A2(n776), .B1(n2346), .B2(n773), .C1(n2282), 
        .C2(n770), .ZN(n4623) );
  OAI222_X1 U2135 ( .A1(n201), .A2(n710), .B1(n233), .B2(n707), .C1(n169), 
        .C2(n704), .ZN(n5998) );
  OAI222_X1 U2136 ( .A1(n905), .A2(n644), .B1(n937), .B2(n641), .C1(n873), 
        .C2(n638), .ZN(n6007) );
  OAI222_X1 U2137 ( .A1(n1961), .A2(n482), .B1(n1993), .B2(n479), .C1(n1929), 
        .C2(n476), .ZN(n6016) );
  OAI222_X1 U2138 ( .A1(n2313), .A2(n64), .B1(n2345), .B2(n61), .C1(n2281), 
        .C2(n58), .ZN(n6025) );
  OAI222_X1 U2139 ( .A1(n201), .A2(n1422), .B1(n233), .B2(n1419), .C1(n169), 
        .C2(n1416), .ZN(n4555) );
  OAI222_X1 U2140 ( .A1(n905), .A2(n1356), .B1(n937), .B2(n1353), .C1(n873), 
        .C2(n1350), .ZN(n4564) );
  OAI222_X1 U2141 ( .A1(n1961), .A2(n1194), .B1(n1993), .B2(n1191), .C1(n1929), 
        .C2(n1188), .ZN(n4573) );
  OAI222_X1 U2142 ( .A1(n2313), .A2(n776), .B1(n2345), .B2(n773), .C1(n2281), 
        .C2(n770), .ZN(n4582) );
  OAI222_X1 U2143 ( .A1(n200), .A2(n710), .B1(n232), .B2(n707), .C1(n168), 
        .C2(n704), .ZN(n5957) );
  OAI222_X1 U2144 ( .A1(n904), .A2(n644), .B1(n936), .B2(n641), .C1(n872), 
        .C2(n638), .ZN(n5966) );
  OAI222_X1 U2145 ( .A1(n1960), .A2(n482), .B1(n1992), .B2(n479), .C1(n1928), 
        .C2(n476), .ZN(n5975) );
  OAI222_X1 U2146 ( .A1(n2312), .A2(n64), .B1(n2344), .B2(n61), .C1(n2280), 
        .C2(n58), .ZN(n5984) );
  OAI222_X1 U2147 ( .A1(n200), .A2(n1422), .B1(n232), .B2(n1419), .C1(n168), 
        .C2(n1416), .ZN(n4514) );
  OAI222_X1 U2148 ( .A1(n904), .A2(n1356), .B1(n936), .B2(n1353), .C1(n872), 
        .C2(n1350), .ZN(n4523) );
  OAI222_X1 U2149 ( .A1(n1960), .A2(n1194), .B1(n1992), .B2(n1191), .C1(n1928), 
        .C2(n1188), .ZN(n4532) );
  OAI222_X1 U2150 ( .A1(n2312), .A2(n776), .B1(n2344), .B2(n773), .C1(n2280), 
        .C2(n770), .ZN(n4541) );
  OAI222_X1 U2151 ( .A1(n199), .A2(n710), .B1(n231), .B2(n707), .C1(n167), 
        .C2(n704), .ZN(n5916) );
  OAI222_X1 U2152 ( .A1(n903), .A2(n644), .B1(n935), .B2(n641), .C1(n871), 
        .C2(n638), .ZN(n5925) );
  OAI222_X1 U2153 ( .A1(n1959), .A2(n482), .B1(n1991), .B2(n479), .C1(n1927), 
        .C2(n476), .ZN(n5934) );
  OAI222_X1 U2154 ( .A1(n2311), .A2(n64), .B1(n2343), .B2(n61), .C1(n2279), 
        .C2(n58), .ZN(n5943) );
  OAI222_X1 U2155 ( .A1(n199), .A2(n1422), .B1(n231), .B2(n1419), .C1(n167), 
        .C2(n1416), .ZN(n4473) );
  OAI222_X1 U2156 ( .A1(n903), .A2(n1356), .B1(n935), .B2(n1353), .C1(n871), 
        .C2(n1350), .ZN(n4482) );
  OAI222_X1 U2157 ( .A1(n1959), .A2(n1194), .B1(n1991), .B2(n1191), .C1(n1927), 
        .C2(n1188), .ZN(n4491) );
  OAI222_X1 U2158 ( .A1(n2311), .A2(n776), .B1(n2343), .B2(n773), .C1(n2279), 
        .C2(n770), .ZN(n4500) );
  OAI222_X1 U2159 ( .A1(n198), .A2(n710), .B1(n230), .B2(n707), .C1(n166), 
        .C2(n704), .ZN(n5875) );
  OAI222_X1 U2160 ( .A1(n902), .A2(n644), .B1(n934), .B2(n641), .C1(n870), 
        .C2(n638), .ZN(n5884) );
  OAI222_X1 U2161 ( .A1(n1958), .A2(n482), .B1(n1990), .B2(n479), .C1(n1926), 
        .C2(n476), .ZN(n5893) );
  OAI222_X1 U2162 ( .A1(n2310), .A2(n64), .B1(n2342), .B2(n61), .C1(n2278), 
        .C2(n58), .ZN(n5902) );
  OAI222_X1 U2163 ( .A1(n198), .A2(n1422), .B1(n230), .B2(n1419), .C1(n166), 
        .C2(n1416), .ZN(n4432) );
  OAI222_X1 U2164 ( .A1(n902), .A2(n1356), .B1(n934), .B2(n1353), .C1(n870), 
        .C2(n1350), .ZN(n4441) );
  OAI222_X1 U2165 ( .A1(n1958), .A2(n1194), .B1(n1990), .B2(n1191), .C1(n1926), 
        .C2(n1188), .ZN(n4450) );
  OAI222_X1 U2166 ( .A1(n2310), .A2(n776), .B1(n2342), .B2(n773), .C1(n2278), 
        .C2(n770), .ZN(n4459) );
  OAI222_X1 U2167 ( .A1(n197), .A2(n710), .B1(n229), .B2(n707), .C1(n165), 
        .C2(n704), .ZN(n5834) );
  OAI222_X1 U2168 ( .A1(n901), .A2(n644), .B1(n933), .B2(n641), .C1(n869), 
        .C2(n638), .ZN(n5843) );
  OAI222_X1 U2169 ( .A1(n1957), .A2(n482), .B1(n1989), .B2(n479), .C1(n1925), 
        .C2(n476), .ZN(n5852) );
  OAI222_X1 U2170 ( .A1(n2309), .A2(n64), .B1(n2341), .B2(n61), .C1(n2277), 
        .C2(n58), .ZN(n5861) );
  OAI222_X1 U2171 ( .A1(n197), .A2(n1422), .B1(n229), .B2(n1419), .C1(n165), 
        .C2(n1416), .ZN(n4391) );
  OAI222_X1 U2172 ( .A1(n901), .A2(n1356), .B1(n933), .B2(n1353), .C1(n869), 
        .C2(n1350), .ZN(n4400) );
  OAI222_X1 U2173 ( .A1(n1957), .A2(n1194), .B1(n1989), .B2(n1191), .C1(n1925), 
        .C2(n1188), .ZN(n4409) );
  OAI222_X1 U2174 ( .A1(n2309), .A2(n776), .B1(n2341), .B2(n773), .C1(n2277), 
        .C2(n770), .ZN(n4418) );
  OAI222_X1 U2175 ( .A1(n196), .A2(n710), .B1(n228), .B2(n707), .C1(n164), 
        .C2(n704), .ZN(n5793) );
  OAI222_X1 U2176 ( .A1(n900), .A2(n644), .B1(n932), .B2(n641), .C1(n868), 
        .C2(n638), .ZN(n5802) );
  OAI222_X1 U2177 ( .A1(n1956), .A2(n482), .B1(n1988), .B2(n479), .C1(n1924), 
        .C2(n476), .ZN(n5811) );
  OAI222_X1 U2178 ( .A1(n2308), .A2(n64), .B1(n2340), .B2(n61), .C1(n2276), 
        .C2(n58), .ZN(n5820) );
  OAI222_X1 U2179 ( .A1(n196), .A2(n1422), .B1(n228), .B2(n1419), .C1(n164), 
        .C2(n1416), .ZN(n4350) );
  OAI222_X1 U2180 ( .A1(n900), .A2(n1356), .B1(n932), .B2(n1353), .C1(n868), 
        .C2(n1350), .ZN(n4359) );
  OAI222_X1 U2181 ( .A1(n1956), .A2(n1194), .B1(n1988), .B2(n1191), .C1(n1924), 
        .C2(n1188), .ZN(n4368) );
  OAI222_X1 U2182 ( .A1(n2308), .A2(n776), .B1(n2340), .B2(n773), .C1(n2276), 
        .C2(n770), .ZN(n4377) );
  OAI222_X1 U2183 ( .A1(n195), .A2(n711), .B1(n227), .B2(n708), .C1(n163), 
        .C2(n705), .ZN(n5752) );
  OAI222_X1 U2184 ( .A1(n899), .A2(n645), .B1(n931), .B2(n642), .C1(n867), 
        .C2(n639), .ZN(n5761) );
  OAI222_X1 U2185 ( .A1(n1955), .A2(n483), .B1(n1987), .B2(n480), .C1(n1923), 
        .C2(n477), .ZN(n5770) );
  OAI222_X1 U2186 ( .A1(n2307), .A2(n65), .B1(n2339), .B2(n62), .C1(n2275), 
        .C2(n59), .ZN(n5779) );
  OAI222_X1 U2187 ( .A1(n195), .A2(n1423), .B1(n227), .B2(n1420), .C1(n163), 
        .C2(n1417), .ZN(n4309) );
  OAI222_X1 U2188 ( .A1(n899), .A2(n1357), .B1(n931), .B2(n1354), .C1(n867), 
        .C2(n1351), .ZN(n4318) );
  OAI222_X1 U2189 ( .A1(n1955), .A2(n1195), .B1(n1987), .B2(n1192), .C1(n1923), 
        .C2(n1189), .ZN(n4327) );
  OAI222_X1 U2190 ( .A1(n2307), .A2(n777), .B1(n2339), .B2(n774), .C1(n2275), 
        .C2(n771), .ZN(n4336) );
  OAI222_X1 U2191 ( .A1(n194), .A2(n711), .B1(n226), .B2(n708), .C1(n162), 
        .C2(n705), .ZN(n5711) );
  OAI222_X1 U2192 ( .A1(n898), .A2(n645), .B1(n930), .B2(n642), .C1(n866), 
        .C2(n639), .ZN(n5720) );
  OAI222_X1 U2193 ( .A1(n1954), .A2(n483), .B1(n1986), .B2(n480), .C1(n1922), 
        .C2(n477), .ZN(n5729) );
  OAI222_X1 U2194 ( .A1(n2306), .A2(n65), .B1(n2338), .B2(n62), .C1(n2274), 
        .C2(n59), .ZN(n5738) );
  OAI222_X1 U2195 ( .A1(n194), .A2(n1423), .B1(n226), .B2(n1420), .C1(n162), 
        .C2(n1417), .ZN(n4268) );
  OAI222_X1 U2196 ( .A1(n898), .A2(n1357), .B1(n930), .B2(n1354), .C1(n866), 
        .C2(n1351), .ZN(n4277) );
  OAI222_X1 U2197 ( .A1(n1954), .A2(n1195), .B1(n1986), .B2(n1192), .C1(n1922), 
        .C2(n1189), .ZN(n4286) );
  OAI222_X1 U2198 ( .A1(n2306), .A2(n777), .B1(n2338), .B2(n774), .C1(n2274), 
        .C2(n771), .ZN(n4295) );
  OAI222_X1 U2199 ( .A1(n193), .A2(n711), .B1(n225), .B2(n708), .C1(n161), 
        .C2(n705), .ZN(n5670) );
  OAI222_X1 U2200 ( .A1(n897), .A2(n645), .B1(n929), .B2(n642), .C1(n865), 
        .C2(n639), .ZN(n5679) );
  OAI222_X1 U2201 ( .A1(n1953), .A2(n483), .B1(n1985), .B2(n480), .C1(n1921), 
        .C2(n477), .ZN(n5688) );
  OAI222_X1 U2202 ( .A1(n2305), .A2(n65), .B1(n2337), .B2(n62), .C1(n2273), 
        .C2(n59), .ZN(n5697) );
  OAI222_X1 U2203 ( .A1(n193), .A2(n1423), .B1(n225), .B2(n1420), .C1(n161), 
        .C2(n1417), .ZN(n4227) );
  OAI222_X1 U2204 ( .A1(n897), .A2(n1357), .B1(n929), .B2(n1354), .C1(n865), 
        .C2(n1351), .ZN(n4236) );
  OAI222_X1 U2205 ( .A1(n1953), .A2(n1195), .B1(n1985), .B2(n1192), .C1(n1921), 
        .C2(n1189), .ZN(n4245) );
  OAI222_X1 U2206 ( .A1(n2305), .A2(n777), .B1(n2337), .B2(n774), .C1(n2273), 
        .C2(n771), .ZN(n4254) );
  OAI222_X1 U2207 ( .A1(n192), .A2(n711), .B1(n224), .B2(n708), .C1(n160), 
        .C2(n705), .ZN(n5629) );
  OAI222_X1 U2208 ( .A1(n896), .A2(n645), .B1(n928), .B2(n642), .C1(n864), 
        .C2(n639), .ZN(n5638) );
  OAI222_X1 U2209 ( .A1(n1952), .A2(n483), .B1(n1984), .B2(n480), .C1(n1920), 
        .C2(n477), .ZN(n5647) );
  OAI222_X1 U2210 ( .A1(n2304), .A2(n65), .B1(n2336), .B2(n62), .C1(n2272), 
        .C2(n59), .ZN(n5656) );
  OAI222_X1 U2211 ( .A1(n192), .A2(n1423), .B1(n224), .B2(n1420), .C1(n160), 
        .C2(n1417), .ZN(n4186) );
  OAI222_X1 U2212 ( .A1(n896), .A2(n1357), .B1(n928), .B2(n1354), .C1(n864), 
        .C2(n1351), .ZN(n4195) );
  OAI222_X1 U2213 ( .A1(n1952), .A2(n1195), .B1(n1984), .B2(n1192), .C1(n1920), 
        .C2(n1189), .ZN(n4204) );
  OAI222_X1 U2214 ( .A1(n2304), .A2(n777), .B1(n2336), .B2(n774), .C1(n2272), 
        .C2(n771), .ZN(n4213) );
  OAI222_X1 U2215 ( .A1(n191), .A2(n711), .B1(n223), .B2(n708), .C1(n159), 
        .C2(n705), .ZN(n5588) );
  OAI222_X1 U2216 ( .A1(n895), .A2(n645), .B1(n927), .B2(n642), .C1(n863), 
        .C2(n639), .ZN(n5597) );
  OAI222_X1 U2217 ( .A1(n1951), .A2(n483), .B1(n1983), .B2(n480), .C1(n1919), 
        .C2(n477), .ZN(n5606) );
  OAI222_X1 U2218 ( .A1(n2303), .A2(n65), .B1(n2335), .B2(n62), .C1(n2271), 
        .C2(n59), .ZN(n5615) );
  OAI222_X1 U2219 ( .A1(n191), .A2(n1423), .B1(n223), .B2(n1420), .C1(n159), 
        .C2(n1417), .ZN(n4145) );
  OAI222_X1 U2220 ( .A1(n895), .A2(n1357), .B1(n927), .B2(n1354), .C1(n863), 
        .C2(n1351), .ZN(n4154) );
  OAI222_X1 U2221 ( .A1(n1951), .A2(n1195), .B1(n1983), .B2(n1192), .C1(n1919), 
        .C2(n1189), .ZN(n4163) );
  OAI222_X1 U2222 ( .A1(n2303), .A2(n777), .B1(n2335), .B2(n774), .C1(n2271), 
        .C2(n771), .ZN(n4172) );
  OAI222_X1 U2223 ( .A1(n190), .A2(n711), .B1(n222), .B2(n708), .C1(n158), 
        .C2(n705), .ZN(n5547) );
  OAI222_X1 U2224 ( .A1(n894), .A2(n645), .B1(n926), .B2(n642), .C1(n862), 
        .C2(n639), .ZN(n5556) );
  OAI222_X1 U2225 ( .A1(n1950), .A2(n483), .B1(n1982), .B2(n480), .C1(n1918), 
        .C2(n477), .ZN(n5565) );
  OAI222_X1 U2226 ( .A1(n2302), .A2(n65), .B1(n2334), .B2(n62), .C1(n2270), 
        .C2(n59), .ZN(n5574) );
  OAI222_X1 U2227 ( .A1(n190), .A2(n1423), .B1(n222), .B2(n1420), .C1(n158), 
        .C2(n1417), .ZN(n4104) );
  OAI222_X1 U2228 ( .A1(n894), .A2(n1357), .B1(n926), .B2(n1354), .C1(n862), 
        .C2(n1351), .ZN(n4113) );
  OAI222_X1 U2229 ( .A1(n1950), .A2(n1195), .B1(n1982), .B2(n1192), .C1(n1918), 
        .C2(n1189), .ZN(n4122) );
  OAI222_X1 U2230 ( .A1(n2302), .A2(n777), .B1(n2334), .B2(n774), .C1(n2270), 
        .C2(n771), .ZN(n4131) );
  OAI222_X1 U2231 ( .A1(n189), .A2(n711), .B1(n221), .B2(n708), .C1(n157), 
        .C2(n705), .ZN(n5506) );
  OAI222_X1 U2232 ( .A1(n893), .A2(n645), .B1(n925), .B2(n642), .C1(n861), 
        .C2(n639), .ZN(n5515) );
  OAI222_X1 U2233 ( .A1(n1949), .A2(n483), .B1(n1981), .B2(n480), .C1(n1917), 
        .C2(n477), .ZN(n5524) );
  OAI222_X1 U2234 ( .A1(n2301), .A2(n65), .B1(n2333), .B2(n62), .C1(n2269), 
        .C2(n59), .ZN(n5533) );
  OAI222_X1 U2235 ( .A1(n189), .A2(n1423), .B1(n221), .B2(n1420), .C1(n157), 
        .C2(n1417), .ZN(n4063) );
  OAI222_X1 U2236 ( .A1(n893), .A2(n1357), .B1(n925), .B2(n1354), .C1(n861), 
        .C2(n1351), .ZN(n4072) );
  OAI222_X1 U2237 ( .A1(n1949), .A2(n1195), .B1(n1981), .B2(n1192), .C1(n1917), 
        .C2(n1189), .ZN(n4081) );
  OAI222_X1 U2238 ( .A1(n2301), .A2(n777), .B1(n2333), .B2(n774), .C1(n2269), 
        .C2(n771), .ZN(n4090) );
  OAI222_X1 U2239 ( .A1(n188), .A2(n711), .B1(n220), .B2(n708), .C1(n156), 
        .C2(n705), .ZN(n5465) );
  OAI222_X1 U2240 ( .A1(n892), .A2(n645), .B1(n924), .B2(n642), .C1(n860), 
        .C2(n639), .ZN(n5474) );
  OAI222_X1 U2241 ( .A1(n1948), .A2(n483), .B1(n1980), .B2(n480), .C1(n1916), 
        .C2(n477), .ZN(n5483) );
  OAI222_X1 U2242 ( .A1(n2300), .A2(n65), .B1(n2332), .B2(n62), .C1(n2268), 
        .C2(n59), .ZN(n5492) );
  OAI222_X1 U2243 ( .A1(n188), .A2(n1423), .B1(n220), .B2(n1420), .C1(n156), 
        .C2(n1417), .ZN(n4022) );
  OAI222_X1 U2244 ( .A1(n892), .A2(n1357), .B1(n924), .B2(n1354), .C1(n860), 
        .C2(n1351), .ZN(n4031) );
  OAI222_X1 U2245 ( .A1(n1948), .A2(n1195), .B1(n1980), .B2(n1192), .C1(n1916), 
        .C2(n1189), .ZN(n4040) );
  OAI222_X1 U2246 ( .A1(n2300), .A2(n777), .B1(n2332), .B2(n774), .C1(n2268), 
        .C2(n771), .ZN(n4049) );
  OAI222_X1 U2247 ( .A1(n187), .A2(n711), .B1(n219), .B2(n708), .C1(n155), 
        .C2(n705), .ZN(n5424) );
  OAI222_X1 U2248 ( .A1(n891), .A2(n645), .B1(n923), .B2(n642), .C1(n859), 
        .C2(n639), .ZN(n5433) );
  OAI222_X1 U2249 ( .A1(n1947), .A2(n483), .B1(n1979), .B2(n480), .C1(n1915), 
        .C2(n477), .ZN(n5442) );
  OAI222_X1 U2250 ( .A1(n2299), .A2(n65), .B1(n2331), .B2(n62), .C1(n2267), 
        .C2(n59), .ZN(n5451) );
  OAI222_X1 U2251 ( .A1(n187), .A2(n1423), .B1(n219), .B2(n1420), .C1(n155), 
        .C2(n1417), .ZN(n3981) );
  OAI222_X1 U2252 ( .A1(n891), .A2(n1357), .B1(n923), .B2(n1354), .C1(n859), 
        .C2(n1351), .ZN(n3990) );
  OAI222_X1 U2253 ( .A1(n1947), .A2(n1195), .B1(n1979), .B2(n1192), .C1(n1915), 
        .C2(n1189), .ZN(n3999) );
  OAI222_X1 U2254 ( .A1(n2299), .A2(n777), .B1(n2331), .B2(n774), .C1(n2267), 
        .C2(n771), .ZN(n4008) );
  OAI222_X1 U2255 ( .A1(n186), .A2(n711), .B1(n218), .B2(n708), .C1(n154), 
        .C2(n705), .ZN(n5383) );
  OAI222_X1 U2256 ( .A1(n890), .A2(n645), .B1(n922), .B2(n642), .C1(n858), 
        .C2(n639), .ZN(n5392) );
  OAI222_X1 U2257 ( .A1(n1946), .A2(n483), .B1(n1978), .B2(n480), .C1(n1914), 
        .C2(n477), .ZN(n5401) );
  OAI222_X1 U2258 ( .A1(n2298), .A2(n65), .B1(n2330), .B2(n62), .C1(n2266), 
        .C2(n59), .ZN(n5410) );
  OAI222_X1 U2259 ( .A1(n186), .A2(n1423), .B1(n218), .B2(n1420), .C1(n154), 
        .C2(n1417), .ZN(n3940) );
  OAI222_X1 U2260 ( .A1(n890), .A2(n1357), .B1(n922), .B2(n1354), .C1(n858), 
        .C2(n1351), .ZN(n3949) );
  OAI222_X1 U2261 ( .A1(n1946), .A2(n1195), .B1(n1978), .B2(n1192), .C1(n1914), 
        .C2(n1189), .ZN(n3958) );
  OAI222_X1 U2262 ( .A1(n2298), .A2(n777), .B1(n2330), .B2(n774), .C1(n2266), 
        .C2(n771), .ZN(n3967) );
  OAI222_X1 U2263 ( .A1(n185), .A2(n711), .B1(n217), .B2(n708), .C1(n153), 
        .C2(n705), .ZN(n5342) );
  OAI222_X1 U2264 ( .A1(n889), .A2(n645), .B1(n921), .B2(n642), .C1(n857), 
        .C2(n639), .ZN(n5351) );
  OAI222_X1 U2265 ( .A1(n1945), .A2(n483), .B1(n1977), .B2(n480), .C1(n1913), 
        .C2(n477), .ZN(n5360) );
  OAI222_X1 U2266 ( .A1(n2297), .A2(n65), .B1(n2329), .B2(n62), .C1(n2265), 
        .C2(n59), .ZN(n5369) );
  OAI222_X1 U2267 ( .A1(n185), .A2(n1423), .B1(n217), .B2(n1420), .C1(n153), 
        .C2(n1417), .ZN(n3899) );
  OAI222_X1 U2268 ( .A1(n889), .A2(n1357), .B1(n921), .B2(n1354), .C1(n857), 
        .C2(n1351), .ZN(n3908) );
  OAI222_X1 U2269 ( .A1(n1945), .A2(n1195), .B1(n1977), .B2(n1192), .C1(n1913), 
        .C2(n1189), .ZN(n3917) );
  OAI222_X1 U2270 ( .A1(n2297), .A2(n777), .B1(n2329), .B2(n774), .C1(n2265), 
        .C2(n771), .ZN(n3926) );
  OAI222_X1 U2271 ( .A1(n184), .A2(n711), .B1(n216), .B2(n708), .C1(n152), 
        .C2(n705), .ZN(n5301) );
  OAI222_X1 U2272 ( .A1(n888), .A2(n645), .B1(n920), .B2(n642), .C1(n856), 
        .C2(n639), .ZN(n5310) );
  OAI222_X1 U2273 ( .A1(n1944), .A2(n483), .B1(n1976), .B2(n480), .C1(n1912), 
        .C2(n477), .ZN(n5319) );
  OAI222_X1 U2274 ( .A1(n2296), .A2(n65), .B1(n2328), .B2(n62), .C1(n2264), 
        .C2(n59), .ZN(n5328) );
  OAI222_X1 U2275 ( .A1(n184), .A2(n1423), .B1(n216), .B2(n1420), .C1(n152), 
        .C2(n1417), .ZN(n3858) );
  OAI222_X1 U2276 ( .A1(n888), .A2(n1357), .B1(n920), .B2(n1354), .C1(n856), 
        .C2(n1351), .ZN(n3867) );
  OAI222_X1 U2277 ( .A1(n1944), .A2(n1195), .B1(n1976), .B2(n1192), .C1(n1912), 
        .C2(n1189), .ZN(n3876) );
  OAI222_X1 U2278 ( .A1(n2296), .A2(n777), .B1(n2328), .B2(n774), .C1(n2264), 
        .C2(n771), .ZN(n3885) );
  OAI222_X1 U2279 ( .A1(n183), .A2(n712), .B1(n215), .B2(n709), .C1(n151), 
        .C2(n706), .ZN(n5260) );
  OAI222_X1 U2280 ( .A1(n887), .A2(n646), .B1(n919), .B2(n643), .C1(n855), 
        .C2(n640), .ZN(n5269) );
  OAI222_X1 U2281 ( .A1(n1943), .A2(n484), .B1(n1975), .B2(n481), .C1(n1911), 
        .C2(n478), .ZN(n5278) );
  OAI222_X1 U2282 ( .A1(n2295), .A2(n66), .B1(n2327), .B2(n63), .C1(n2263), 
        .C2(n60), .ZN(n5287) );
  OAI222_X1 U2283 ( .A1(n183), .A2(n1424), .B1(n215), .B2(n1421), .C1(n151), 
        .C2(n1418), .ZN(n3817) );
  OAI222_X1 U2284 ( .A1(n887), .A2(n1358), .B1(n919), .B2(n1355), .C1(n855), 
        .C2(n1352), .ZN(n3826) );
  OAI222_X1 U2285 ( .A1(n1943), .A2(n1196), .B1(n1975), .B2(n1193), .C1(n1911), 
        .C2(n1190), .ZN(n3835) );
  OAI222_X1 U2286 ( .A1(n2295), .A2(n778), .B1(n2327), .B2(n775), .C1(n2263), 
        .C2(n772), .ZN(n3844) );
  OAI222_X1 U2287 ( .A1(n182), .A2(n712), .B1(n214), .B2(n709), .C1(n150), 
        .C2(n706), .ZN(n5219) );
  OAI222_X1 U2288 ( .A1(n886), .A2(n646), .B1(n918), .B2(n643), .C1(n854), 
        .C2(n640), .ZN(n5228) );
  OAI222_X1 U2289 ( .A1(n1942), .A2(n484), .B1(n1974), .B2(n481), .C1(n1910), 
        .C2(n478), .ZN(n5237) );
  OAI222_X1 U2290 ( .A1(n2294), .A2(n66), .B1(n2326), .B2(n63), .C1(n2262), 
        .C2(n60), .ZN(n5246) );
  OAI222_X1 U2291 ( .A1(n182), .A2(n1424), .B1(n214), .B2(n1421), .C1(n150), 
        .C2(n1418), .ZN(n3776) );
  OAI222_X1 U2292 ( .A1(n886), .A2(n1358), .B1(n918), .B2(n1355), .C1(n854), 
        .C2(n1352), .ZN(n3785) );
  OAI222_X1 U2293 ( .A1(n1942), .A2(n1196), .B1(n1974), .B2(n1193), .C1(n1910), 
        .C2(n1190), .ZN(n3794) );
  OAI222_X1 U2294 ( .A1(n2294), .A2(n778), .B1(n2326), .B2(n775), .C1(n2262), 
        .C2(n772), .ZN(n3803) );
  OAI222_X1 U2295 ( .A1(n181), .A2(n712), .B1(n213), .B2(n709), .C1(n149), 
        .C2(n706), .ZN(n5178) );
  OAI222_X1 U2296 ( .A1(n885), .A2(n646), .B1(n917), .B2(n643), .C1(n853), 
        .C2(n640), .ZN(n5187) );
  OAI222_X1 U2297 ( .A1(n1941), .A2(n484), .B1(n1973), .B2(n481), .C1(n1909), 
        .C2(n478), .ZN(n5196) );
  OAI222_X1 U2298 ( .A1(n2293), .A2(n66), .B1(n2325), .B2(n63), .C1(n2261), 
        .C2(n60), .ZN(n5205) );
  OAI222_X1 U2299 ( .A1(n181), .A2(n1424), .B1(n213), .B2(n1421), .C1(n149), 
        .C2(n1418), .ZN(n3735) );
  OAI222_X1 U2300 ( .A1(n885), .A2(n1358), .B1(n917), .B2(n1355), .C1(n853), 
        .C2(n1352), .ZN(n3744) );
  OAI222_X1 U2301 ( .A1(n1941), .A2(n1196), .B1(n1973), .B2(n1193), .C1(n1909), 
        .C2(n1190), .ZN(n3753) );
  OAI222_X1 U2302 ( .A1(n2293), .A2(n778), .B1(n2325), .B2(n775), .C1(n2261), 
        .C2(n772), .ZN(n3762) );
  OAI222_X1 U2303 ( .A1(n180), .A2(n712), .B1(n212), .B2(n709), .C1(n148), 
        .C2(n706), .ZN(n5137) );
  OAI222_X1 U2304 ( .A1(n884), .A2(n646), .B1(n916), .B2(n643), .C1(n852), 
        .C2(n640), .ZN(n5146) );
  OAI222_X1 U2305 ( .A1(n1940), .A2(n484), .B1(n1972), .B2(n481), .C1(n1908), 
        .C2(n478), .ZN(n5155) );
  OAI222_X1 U2306 ( .A1(n2292), .A2(n66), .B1(n2324), .B2(n63), .C1(n2260), 
        .C2(n60), .ZN(n5164) );
  OAI222_X1 U2307 ( .A1(n180), .A2(n1424), .B1(n212), .B2(n1421), .C1(n148), 
        .C2(n1418), .ZN(n3694) );
  OAI222_X1 U2308 ( .A1(n884), .A2(n1358), .B1(n916), .B2(n1355), .C1(n852), 
        .C2(n1352), .ZN(n3703) );
  OAI222_X1 U2309 ( .A1(n1940), .A2(n1196), .B1(n1972), .B2(n1193), .C1(n1908), 
        .C2(n1190), .ZN(n3712) );
  OAI222_X1 U2310 ( .A1(n2292), .A2(n778), .B1(n2324), .B2(n775), .C1(n2260), 
        .C2(n772), .ZN(n3721) );
  OAI222_X1 U2311 ( .A1(n179), .A2(n712), .B1(n211), .B2(n709), .C1(n147), 
        .C2(n706), .ZN(n5096) );
  OAI222_X1 U2312 ( .A1(n883), .A2(n646), .B1(n915), .B2(n643), .C1(n851), 
        .C2(n640), .ZN(n5105) );
  OAI222_X1 U2313 ( .A1(n1939), .A2(n484), .B1(n1971), .B2(n481), .C1(n1907), 
        .C2(n478), .ZN(n5114) );
  OAI222_X1 U2314 ( .A1(n2291), .A2(n66), .B1(n2323), .B2(n63), .C1(n2259), 
        .C2(n60), .ZN(n5123) );
  OAI222_X1 U2315 ( .A1(n179), .A2(n1424), .B1(n211), .B2(n1421), .C1(n147), 
        .C2(n1418), .ZN(n3653) );
  OAI222_X1 U2316 ( .A1(n883), .A2(n1358), .B1(n915), .B2(n1355), .C1(n851), 
        .C2(n1352), .ZN(n3662) );
  OAI222_X1 U2317 ( .A1(n1939), .A2(n1196), .B1(n1971), .B2(n1193), .C1(n1907), 
        .C2(n1190), .ZN(n3671) );
  OAI222_X1 U2318 ( .A1(n2291), .A2(n778), .B1(n2323), .B2(n775), .C1(n2259), 
        .C2(n772), .ZN(n3680) );
  OAI222_X1 U2319 ( .A1(n178), .A2(n712), .B1(n210), .B2(n709), .C1(n146), 
        .C2(n706), .ZN(n5055) );
  OAI222_X1 U2320 ( .A1(n882), .A2(n646), .B1(n914), .B2(n643), .C1(n850), 
        .C2(n640), .ZN(n5064) );
  OAI222_X1 U2321 ( .A1(n1938), .A2(n484), .B1(n1970), .B2(n481), .C1(n1906), 
        .C2(n478), .ZN(n5073) );
  OAI222_X1 U2322 ( .A1(n2290), .A2(n66), .B1(n2322), .B2(n63), .C1(n2258), 
        .C2(n60), .ZN(n5082) );
  OAI222_X1 U2323 ( .A1(n178), .A2(n1424), .B1(n210), .B2(n1421), .C1(n146), 
        .C2(n1418), .ZN(n3612) );
  OAI222_X1 U2324 ( .A1(n882), .A2(n1358), .B1(n914), .B2(n1355), .C1(n850), 
        .C2(n1352), .ZN(n3621) );
  OAI222_X1 U2325 ( .A1(n1938), .A2(n1196), .B1(n1970), .B2(n1193), .C1(n1906), 
        .C2(n1190), .ZN(n3630) );
  OAI222_X1 U2326 ( .A1(n2290), .A2(n778), .B1(n2322), .B2(n775), .C1(n2258), 
        .C2(n772), .ZN(n3639) );
  OAI222_X1 U2327 ( .A1(n177), .A2(n712), .B1(n209), .B2(n709), .C1(n145), 
        .C2(n706), .ZN(n5014) );
  OAI222_X1 U2328 ( .A1(n881), .A2(n646), .B1(n913), .B2(n643), .C1(n849), 
        .C2(n640), .ZN(n5023) );
  OAI222_X1 U2329 ( .A1(n1937), .A2(n484), .B1(n1969), .B2(n481), .C1(n1905), 
        .C2(n478), .ZN(n5032) );
  OAI222_X1 U2330 ( .A1(n2289), .A2(n66), .B1(n2321), .B2(n63), .C1(n2257), 
        .C2(n60), .ZN(n5041) );
  OAI222_X1 U2331 ( .A1(n177), .A2(n1424), .B1(n209), .B2(n1421), .C1(n145), 
        .C2(n1418), .ZN(n3571) );
  OAI222_X1 U2332 ( .A1(n881), .A2(n1358), .B1(n913), .B2(n1355), .C1(n849), 
        .C2(n1352), .ZN(n3580) );
  OAI222_X1 U2333 ( .A1(n1937), .A2(n1196), .B1(n1969), .B2(n1193), .C1(n1905), 
        .C2(n1190), .ZN(n3589) );
  OAI222_X1 U2334 ( .A1(n2289), .A2(n778), .B1(n2321), .B2(n775), .C1(n2257), 
        .C2(n772), .ZN(n3598) );
  OAI222_X1 U2335 ( .A1(n176), .A2(n712), .B1(n208), .B2(n709), .C1(n144), 
        .C2(n706), .ZN(n4885) );
  OAI222_X1 U2336 ( .A1(n880), .A2(n646), .B1(n912), .B2(n643), .C1(n848), 
        .C2(n640), .ZN(n4916) );
  OAI222_X1 U2337 ( .A1(n1936), .A2(n484), .B1(n1968), .B2(n481), .C1(n1904), 
        .C2(n478), .ZN(n4947) );
  OAI222_X1 U2338 ( .A1(n2288), .A2(n66), .B1(n2320), .B2(n63), .C1(n2256), 
        .C2(n60), .ZN(n4978) );
  OAI222_X1 U2339 ( .A1(n176), .A2(n1424), .B1(n208), .B2(n1421), .C1(n144), 
        .C2(n1418), .ZN(n3442) );
  OAI222_X1 U2340 ( .A1(n880), .A2(n1358), .B1(n912), .B2(n1355), .C1(n848), 
        .C2(n1352), .ZN(n3473) );
  OAI222_X1 U2341 ( .A1(n1936), .A2(n1196), .B1(n1968), .B2(n1193), .C1(n1904), 
        .C2(n1190), .ZN(n3504) );
  OAI222_X1 U2342 ( .A1(n2288), .A2(n778), .B1(n2320), .B2(n775), .C1(n2256), 
        .C2(n772), .ZN(n3535) );
  OAI222_X1 U2343 ( .A1(n559), .A2(n677), .B1(n591), .B2(n674), .C1(n527), 
        .C2(n671), .ZN(n6258) );
  OAI222_X1 U2344 ( .A1(n1263), .A2(n611), .B1(n1295), .B2(n608), .C1(n1231), 
        .C2(n605), .ZN(n6282) );
  OAI222_X1 U2345 ( .A1(n559), .A2(n1389), .B1(n591), .B2(n1386), .C1(n527), 
        .C2(n1383), .ZN(n4815) );
  OAI222_X1 U2346 ( .A1(n1263), .A2(n1323), .B1(n1295), .B2(n1320), .C1(n1231), 
        .C2(n1317), .ZN(n4839) );
  OAI222_X1 U2347 ( .A1(n558), .A2(n677), .B1(n590), .B2(n674), .C1(n526), 
        .C2(n671), .ZN(n6205) );
  OAI222_X1 U2348 ( .A1(n1262), .A2(n611), .B1(n1294), .B2(n608), .C1(n1230), 
        .C2(n605), .ZN(n6214) );
  OAI222_X1 U2349 ( .A1(n558), .A2(n1389), .B1(n590), .B2(n1386), .C1(n526), 
        .C2(n1383), .ZN(n4762) );
  OAI222_X1 U2350 ( .A1(n1262), .A2(n1323), .B1(n1294), .B2(n1320), .C1(n1230), 
        .C2(n1317), .ZN(n4771) );
  OAI222_X1 U2351 ( .A1(n557), .A2(n677), .B1(n589), .B2(n674), .C1(n525), 
        .C2(n671), .ZN(n6164) );
  OAI222_X1 U2352 ( .A1(n1261), .A2(n611), .B1(n1293), .B2(n608), .C1(n1229), 
        .C2(n605), .ZN(n6173) );
  OAI222_X1 U2353 ( .A1(n557), .A2(n1389), .B1(n589), .B2(n1386), .C1(n525), 
        .C2(n1383), .ZN(n4721) );
  OAI222_X1 U2354 ( .A1(n1261), .A2(n1323), .B1(n1293), .B2(n1320), .C1(n1229), 
        .C2(n1317), .ZN(n4730) );
  OAI222_X1 U2355 ( .A1(n556), .A2(n677), .B1(n588), .B2(n674), .C1(n524), 
        .C2(n671), .ZN(n6123) );
  OAI222_X1 U2356 ( .A1(n1260), .A2(n611), .B1(n1292), .B2(n608), .C1(n1228), 
        .C2(n605), .ZN(n6132) );
  OAI222_X1 U2357 ( .A1(n556), .A2(n1389), .B1(n588), .B2(n1386), .C1(n524), 
        .C2(n1383), .ZN(n4680) );
  OAI222_X1 U2358 ( .A1(n1260), .A2(n1323), .B1(n1292), .B2(n1320), .C1(n1228), 
        .C2(n1317), .ZN(n4689) );
  OAI222_X1 U2359 ( .A1(n555), .A2(n677), .B1(n587), .B2(n674), .C1(n523), 
        .C2(n671), .ZN(n6082) );
  OAI222_X1 U2360 ( .A1(n1259), .A2(n611), .B1(n1291), .B2(n608), .C1(n1227), 
        .C2(n605), .ZN(n6091) );
  OAI222_X1 U2361 ( .A1(n555), .A2(n1389), .B1(n587), .B2(n1386), .C1(n523), 
        .C2(n1383), .ZN(n4639) );
  OAI222_X1 U2362 ( .A1(n1259), .A2(n1323), .B1(n1291), .B2(n1320), .C1(n1227), 
        .C2(n1317), .ZN(n4648) );
  OAI222_X1 U2363 ( .A1(n554), .A2(n677), .B1(n586), .B2(n674), .C1(n522), 
        .C2(n671), .ZN(n6041) );
  OAI222_X1 U2364 ( .A1(n1258), .A2(n611), .B1(n1290), .B2(n608), .C1(n1226), 
        .C2(n605), .ZN(n6050) );
  OAI222_X1 U2365 ( .A1(n554), .A2(n1389), .B1(n586), .B2(n1386), .C1(n522), 
        .C2(n1383), .ZN(n4598) );
  OAI222_X1 U2366 ( .A1(n1258), .A2(n1323), .B1(n1290), .B2(n1320), .C1(n1226), 
        .C2(n1317), .ZN(n4607) );
  OAI222_X1 U2367 ( .A1(n553), .A2(n677), .B1(n585), .B2(n674), .C1(n521), 
        .C2(n671), .ZN(n6000) );
  OAI222_X1 U2368 ( .A1(n1257), .A2(n611), .B1(n1289), .B2(n608), .C1(n1225), 
        .C2(n605), .ZN(n6009) );
  OAI222_X1 U2369 ( .A1(n553), .A2(n1389), .B1(n585), .B2(n1386), .C1(n521), 
        .C2(n1383), .ZN(n4557) );
  OAI222_X1 U2370 ( .A1(n1257), .A2(n1323), .B1(n1289), .B2(n1320), .C1(n1225), 
        .C2(n1317), .ZN(n4566) );
  OAI222_X1 U2371 ( .A1(n552), .A2(n677), .B1(n584), .B2(n674), .C1(n520), 
        .C2(n671), .ZN(n5959) );
  OAI222_X1 U2372 ( .A1(n1256), .A2(n611), .B1(n1288), .B2(n608), .C1(n1224), 
        .C2(n605), .ZN(n5968) );
  OAI222_X1 U2373 ( .A1(n552), .A2(n1389), .B1(n584), .B2(n1386), .C1(n520), 
        .C2(n1383), .ZN(n4516) );
  OAI222_X1 U2374 ( .A1(n1256), .A2(n1323), .B1(n1288), .B2(n1320), .C1(n1224), 
        .C2(n1317), .ZN(n4525) );
  OAI222_X1 U2375 ( .A1(n551), .A2(n677), .B1(n583), .B2(n674), .C1(n519), 
        .C2(n671), .ZN(n5918) );
  OAI222_X1 U2376 ( .A1(n1255), .A2(n611), .B1(n1287), .B2(n608), .C1(n1223), 
        .C2(n605), .ZN(n5927) );
  OAI222_X1 U2377 ( .A1(n551), .A2(n1389), .B1(n583), .B2(n1386), .C1(n519), 
        .C2(n1383), .ZN(n4475) );
  OAI222_X1 U2378 ( .A1(n1255), .A2(n1323), .B1(n1287), .B2(n1320), .C1(n1223), 
        .C2(n1317), .ZN(n4484) );
  OAI222_X1 U2379 ( .A1(n550), .A2(n677), .B1(n582), .B2(n674), .C1(n518), 
        .C2(n671), .ZN(n5877) );
  OAI222_X1 U2380 ( .A1(n1254), .A2(n611), .B1(n1286), .B2(n608), .C1(n1222), 
        .C2(n605), .ZN(n5886) );
  OAI222_X1 U2381 ( .A1(n550), .A2(n1389), .B1(n582), .B2(n1386), .C1(n518), 
        .C2(n1383), .ZN(n4434) );
  OAI222_X1 U2382 ( .A1(n1254), .A2(n1323), .B1(n1286), .B2(n1320), .C1(n1222), 
        .C2(n1317), .ZN(n4443) );
  OAI222_X1 U2383 ( .A1(n549), .A2(n677), .B1(n581), .B2(n674), .C1(n517), 
        .C2(n671), .ZN(n5836) );
  OAI222_X1 U2384 ( .A1(n1253), .A2(n611), .B1(n1285), .B2(n608), .C1(n1221), 
        .C2(n605), .ZN(n5845) );
  OAI222_X1 U2385 ( .A1(n549), .A2(n1389), .B1(n581), .B2(n1386), .C1(n517), 
        .C2(n1383), .ZN(n4393) );
  OAI222_X1 U2386 ( .A1(n1253), .A2(n1323), .B1(n1285), .B2(n1320), .C1(n1221), 
        .C2(n1317), .ZN(n4402) );
  OAI222_X1 U2387 ( .A1(n548), .A2(n677), .B1(n580), .B2(n674), .C1(n516), 
        .C2(n671), .ZN(n5795) );
  OAI222_X1 U2388 ( .A1(n1252), .A2(n611), .B1(n1284), .B2(n608), .C1(n1220), 
        .C2(n605), .ZN(n5804) );
  OAI222_X1 U2389 ( .A1(n548), .A2(n1389), .B1(n580), .B2(n1386), .C1(n516), 
        .C2(n1383), .ZN(n4352) );
  OAI222_X1 U2390 ( .A1(n1252), .A2(n1323), .B1(n1284), .B2(n1320), .C1(n1220), 
        .C2(n1317), .ZN(n4361) );
  OAI222_X1 U2391 ( .A1(n547), .A2(n678), .B1(n579), .B2(n675), .C1(n515), 
        .C2(n672), .ZN(n5754) );
  OAI222_X1 U2392 ( .A1(n1251), .A2(n612), .B1(n1283), .B2(n609), .C1(n1219), 
        .C2(n606), .ZN(n5763) );
  OAI222_X1 U2393 ( .A1(n547), .A2(n1390), .B1(n579), .B2(n1387), .C1(n515), 
        .C2(n1384), .ZN(n4311) );
  OAI222_X1 U2394 ( .A1(n1251), .A2(n1324), .B1(n1283), .B2(n1321), .C1(n1219), 
        .C2(n1318), .ZN(n4320) );
  OAI222_X1 U2395 ( .A1(n546), .A2(n678), .B1(n578), .B2(n675), .C1(n514), 
        .C2(n672), .ZN(n5713) );
  OAI222_X1 U2396 ( .A1(n1250), .A2(n612), .B1(n1282), .B2(n609), .C1(n1218), 
        .C2(n606), .ZN(n5722) );
  OAI222_X1 U2397 ( .A1(n546), .A2(n1390), .B1(n578), .B2(n1387), .C1(n514), 
        .C2(n1384), .ZN(n4270) );
  OAI222_X1 U2398 ( .A1(n1250), .A2(n1324), .B1(n1282), .B2(n1321), .C1(n1218), 
        .C2(n1318), .ZN(n4279) );
  OAI222_X1 U2399 ( .A1(n545), .A2(n678), .B1(n577), .B2(n675), .C1(n513), 
        .C2(n672), .ZN(n5672) );
  OAI222_X1 U2400 ( .A1(n1249), .A2(n612), .B1(n1281), .B2(n609), .C1(n1217), 
        .C2(n606), .ZN(n5681) );
  OAI222_X1 U2401 ( .A1(n545), .A2(n1390), .B1(n577), .B2(n1387), .C1(n513), 
        .C2(n1384), .ZN(n4229) );
  OAI222_X1 U2402 ( .A1(n1249), .A2(n1324), .B1(n1281), .B2(n1321), .C1(n1217), 
        .C2(n1318), .ZN(n4238) );
  OAI222_X1 U2403 ( .A1(n544), .A2(n678), .B1(n576), .B2(n675), .C1(n512), 
        .C2(n672), .ZN(n5631) );
  OAI222_X1 U2404 ( .A1(n1248), .A2(n612), .B1(n1280), .B2(n609), .C1(n1216), 
        .C2(n606), .ZN(n5640) );
  OAI222_X1 U2405 ( .A1(n544), .A2(n1390), .B1(n576), .B2(n1387), .C1(n512), 
        .C2(n1384), .ZN(n4188) );
  OAI222_X1 U2406 ( .A1(n1248), .A2(n1324), .B1(n1280), .B2(n1321), .C1(n1216), 
        .C2(n1318), .ZN(n4197) );
  OAI222_X1 U2407 ( .A1(n543), .A2(n678), .B1(n575), .B2(n675), .C1(n511), 
        .C2(n672), .ZN(n5590) );
  OAI222_X1 U2408 ( .A1(n1247), .A2(n612), .B1(n1279), .B2(n609), .C1(n1215), 
        .C2(n606), .ZN(n5599) );
  OAI222_X1 U2409 ( .A1(n543), .A2(n1390), .B1(n575), .B2(n1387), .C1(n511), 
        .C2(n1384), .ZN(n4147) );
  OAI222_X1 U2410 ( .A1(n1247), .A2(n1324), .B1(n1279), .B2(n1321), .C1(n1215), 
        .C2(n1318), .ZN(n4156) );
  OAI222_X1 U2411 ( .A1(n542), .A2(n678), .B1(n574), .B2(n675), .C1(n510), 
        .C2(n672), .ZN(n5549) );
  OAI222_X1 U2412 ( .A1(n1246), .A2(n612), .B1(n1278), .B2(n609), .C1(n1214), 
        .C2(n606), .ZN(n5558) );
  OAI222_X1 U2413 ( .A1(n542), .A2(n1390), .B1(n574), .B2(n1387), .C1(n510), 
        .C2(n1384), .ZN(n4106) );
  OAI222_X1 U2414 ( .A1(n1246), .A2(n1324), .B1(n1278), .B2(n1321), .C1(n1214), 
        .C2(n1318), .ZN(n4115) );
  OAI222_X1 U2415 ( .A1(n541), .A2(n678), .B1(n573), .B2(n675), .C1(n509), 
        .C2(n672), .ZN(n5508) );
  OAI222_X1 U2416 ( .A1(n1245), .A2(n612), .B1(n1277), .B2(n609), .C1(n1213), 
        .C2(n606), .ZN(n5517) );
  OAI222_X1 U2417 ( .A1(n541), .A2(n1390), .B1(n573), .B2(n1387), .C1(n509), 
        .C2(n1384), .ZN(n4065) );
  OAI222_X1 U2418 ( .A1(n1245), .A2(n1324), .B1(n1277), .B2(n1321), .C1(n1213), 
        .C2(n1318), .ZN(n4074) );
  OAI222_X1 U2419 ( .A1(n540), .A2(n678), .B1(n572), .B2(n675), .C1(n508), 
        .C2(n672), .ZN(n5467) );
  OAI222_X1 U2420 ( .A1(n1244), .A2(n612), .B1(n1276), .B2(n609), .C1(n1212), 
        .C2(n606), .ZN(n5476) );
  OAI222_X1 U2421 ( .A1(n540), .A2(n1390), .B1(n572), .B2(n1387), .C1(n508), 
        .C2(n1384), .ZN(n4024) );
  OAI222_X1 U2422 ( .A1(n1244), .A2(n1324), .B1(n1276), .B2(n1321), .C1(n1212), 
        .C2(n1318), .ZN(n4033) );
  OAI222_X1 U2423 ( .A1(n539), .A2(n678), .B1(n571), .B2(n675), .C1(n507), 
        .C2(n672), .ZN(n5426) );
  OAI222_X1 U2424 ( .A1(n1243), .A2(n612), .B1(n1275), .B2(n609), .C1(n1211), 
        .C2(n606), .ZN(n5435) );
  OAI222_X1 U2425 ( .A1(n539), .A2(n1390), .B1(n571), .B2(n1387), .C1(n507), 
        .C2(n1384), .ZN(n3983) );
  OAI222_X1 U2426 ( .A1(n1243), .A2(n1324), .B1(n1275), .B2(n1321), .C1(n1211), 
        .C2(n1318), .ZN(n3992) );
  OAI222_X1 U2427 ( .A1(n538), .A2(n678), .B1(n570), .B2(n675), .C1(n506), 
        .C2(n672), .ZN(n5385) );
  OAI222_X1 U2428 ( .A1(n1242), .A2(n612), .B1(n1274), .B2(n609), .C1(n1210), 
        .C2(n606), .ZN(n5394) );
  OAI222_X1 U2429 ( .A1(n538), .A2(n1390), .B1(n570), .B2(n1387), .C1(n506), 
        .C2(n1384), .ZN(n3942) );
  OAI222_X1 U2430 ( .A1(n1242), .A2(n1324), .B1(n1274), .B2(n1321), .C1(n1210), 
        .C2(n1318), .ZN(n3951) );
  OAI222_X1 U2431 ( .A1(n537), .A2(n678), .B1(n569), .B2(n675), .C1(n505), 
        .C2(n672), .ZN(n5344) );
  OAI222_X1 U2432 ( .A1(n1241), .A2(n612), .B1(n1273), .B2(n609), .C1(n1209), 
        .C2(n606), .ZN(n5353) );
  OAI222_X1 U2433 ( .A1(n537), .A2(n1390), .B1(n569), .B2(n1387), .C1(n505), 
        .C2(n1384), .ZN(n3901) );
  OAI222_X1 U2434 ( .A1(n1241), .A2(n1324), .B1(n1273), .B2(n1321), .C1(n1209), 
        .C2(n1318), .ZN(n3910) );
  OAI222_X1 U2435 ( .A1(n536), .A2(n678), .B1(n568), .B2(n675), .C1(n504), 
        .C2(n672), .ZN(n5303) );
  OAI222_X1 U2436 ( .A1(n1240), .A2(n612), .B1(n1272), .B2(n609), .C1(n1208), 
        .C2(n606), .ZN(n5312) );
  OAI222_X1 U2437 ( .A1(n536), .A2(n1390), .B1(n568), .B2(n1387), .C1(n504), 
        .C2(n1384), .ZN(n3860) );
  OAI222_X1 U2438 ( .A1(n1240), .A2(n1324), .B1(n1272), .B2(n1321), .C1(n1208), 
        .C2(n1318), .ZN(n3869) );
  OAI222_X1 U2439 ( .A1(n535), .A2(n679), .B1(n567), .B2(n676), .C1(n503), 
        .C2(n673), .ZN(n5262) );
  OAI222_X1 U2440 ( .A1(n1239), .A2(n613), .B1(n1271), .B2(n610), .C1(n1207), 
        .C2(n607), .ZN(n5271) );
  OAI222_X1 U2441 ( .A1(n535), .A2(n1391), .B1(n567), .B2(n1388), .C1(n503), 
        .C2(n1385), .ZN(n3819) );
  OAI222_X1 U2442 ( .A1(n1239), .A2(n1325), .B1(n1271), .B2(n1322), .C1(n1207), 
        .C2(n1319), .ZN(n3828) );
  OAI222_X1 U2443 ( .A1(n534), .A2(n679), .B1(n566), .B2(n676), .C1(n502), 
        .C2(n673), .ZN(n5221) );
  OAI222_X1 U2444 ( .A1(n1238), .A2(n613), .B1(n1270), .B2(n610), .C1(n1206), 
        .C2(n607), .ZN(n5230) );
  OAI222_X1 U2445 ( .A1(n534), .A2(n1391), .B1(n566), .B2(n1388), .C1(n502), 
        .C2(n1385), .ZN(n3778) );
  OAI222_X1 U2446 ( .A1(n1238), .A2(n1325), .B1(n1270), .B2(n1322), .C1(n1206), 
        .C2(n1319), .ZN(n3787) );
  OAI222_X1 U2447 ( .A1(n533), .A2(n679), .B1(n565), .B2(n676), .C1(n501), 
        .C2(n673), .ZN(n5180) );
  OAI222_X1 U2448 ( .A1(n1237), .A2(n613), .B1(n1269), .B2(n610), .C1(n1205), 
        .C2(n607), .ZN(n5189) );
  OAI222_X1 U2449 ( .A1(n533), .A2(n1391), .B1(n565), .B2(n1388), .C1(n501), 
        .C2(n1385), .ZN(n3737) );
  OAI222_X1 U2450 ( .A1(n1237), .A2(n1325), .B1(n1269), .B2(n1322), .C1(n1205), 
        .C2(n1319), .ZN(n3746) );
  OAI222_X1 U2451 ( .A1(n532), .A2(n679), .B1(n564), .B2(n676), .C1(n500), 
        .C2(n673), .ZN(n5139) );
  OAI222_X1 U2452 ( .A1(n1236), .A2(n613), .B1(n1268), .B2(n610), .C1(n1204), 
        .C2(n607), .ZN(n5148) );
  OAI222_X1 U2453 ( .A1(n532), .A2(n1391), .B1(n564), .B2(n1388), .C1(n500), 
        .C2(n1385), .ZN(n3696) );
  OAI222_X1 U2454 ( .A1(n1236), .A2(n1325), .B1(n1268), .B2(n1322), .C1(n1204), 
        .C2(n1319), .ZN(n3705) );
  OAI222_X1 U2455 ( .A1(n531), .A2(n679), .B1(n563), .B2(n676), .C1(n499), 
        .C2(n673), .ZN(n5098) );
  OAI222_X1 U2456 ( .A1(n1235), .A2(n613), .B1(n1267), .B2(n610), .C1(n1203), 
        .C2(n607), .ZN(n5107) );
  OAI222_X1 U2457 ( .A1(n531), .A2(n1391), .B1(n563), .B2(n1388), .C1(n499), 
        .C2(n1385), .ZN(n3655) );
  OAI222_X1 U2458 ( .A1(n1235), .A2(n1325), .B1(n1267), .B2(n1322), .C1(n1203), 
        .C2(n1319), .ZN(n3664) );
  OAI222_X1 U2459 ( .A1(n530), .A2(n679), .B1(n562), .B2(n676), .C1(n498), 
        .C2(n673), .ZN(n5057) );
  OAI222_X1 U2460 ( .A1(n1234), .A2(n613), .B1(n1266), .B2(n610), .C1(n1202), 
        .C2(n607), .ZN(n5066) );
  OAI222_X1 U2461 ( .A1(n530), .A2(n1391), .B1(n562), .B2(n1388), .C1(n498), 
        .C2(n1385), .ZN(n3614) );
  OAI222_X1 U2462 ( .A1(n1234), .A2(n1325), .B1(n1266), .B2(n1322), .C1(n1202), 
        .C2(n1319), .ZN(n3623) );
  OAI222_X1 U2463 ( .A1(n529), .A2(n679), .B1(n561), .B2(n676), .C1(n497), 
        .C2(n673), .ZN(n5016) );
  OAI222_X1 U2464 ( .A1(n1233), .A2(n613), .B1(n1265), .B2(n610), .C1(n1201), 
        .C2(n607), .ZN(n5025) );
  OAI222_X1 U2465 ( .A1(n529), .A2(n1391), .B1(n561), .B2(n1388), .C1(n497), 
        .C2(n1385), .ZN(n3573) );
  OAI222_X1 U2466 ( .A1(n1233), .A2(n1325), .B1(n1265), .B2(n1322), .C1(n1201), 
        .C2(n1319), .ZN(n3582) );
  OAI222_X1 U2467 ( .A1(n528), .A2(n679), .B1(n560), .B2(n676), .C1(n496), 
        .C2(n673), .ZN(n4900) );
  OAI222_X1 U2468 ( .A1(n1232), .A2(n613), .B1(n1264), .B2(n610), .C1(n1200), 
        .C2(n607), .ZN(n4931) );
  OAI222_X1 U2469 ( .A1(n528), .A2(n1391), .B1(n560), .B2(n1388), .C1(n496), 
        .C2(n1385), .ZN(n3457) );
  OAI222_X1 U2470 ( .A1(n1232), .A2(n1325), .B1(n1264), .B2(n1322), .C1(n1200), 
        .C2(n1319), .ZN(n3488) );
  OAI222_X1 U2471 ( .A1(n303), .A2(n701), .B1(n335), .B2(n698), .C1(n271), 
        .C2(n695), .ZN(n6243) );
  OAI222_X1 U2472 ( .A1(n1007), .A2(n635), .B1(n1039), .B2(n632), .C1(n975), 
        .C2(n629), .ZN(n6274) );
  OAI222_X1 U2473 ( .A1(n303), .A2(n1413), .B1(n335), .B2(n1410), .C1(n271), 
        .C2(n1407), .ZN(n4800) );
  OAI222_X1 U2474 ( .A1(n1007), .A2(n1347), .B1(n1039), .B2(n1344), .C1(n975), 
        .C2(n1341), .ZN(n4831) );
  OAI222_X1 U2475 ( .A1(n302), .A2(n701), .B1(n334), .B2(n698), .C1(n270), 
        .C2(n695), .ZN(n6202) );
  OAI222_X1 U2476 ( .A1(n1006), .A2(n635), .B1(n1038), .B2(n632), .C1(n974), 
        .C2(n629), .ZN(n6211) );
  OAI222_X1 U2477 ( .A1(n302), .A2(n1413), .B1(n334), .B2(n1410), .C1(n270), 
        .C2(n1407), .ZN(n4759) );
  OAI222_X1 U2478 ( .A1(n1006), .A2(n1347), .B1(n1038), .B2(n1344), .C1(n974), 
        .C2(n1341), .ZN(n4768) );
  OAI222_X1 U2479 ( .A1(n301), .A2(n701), .B1(n333), .B2(n698), .C1(n269), 
        .C2(n695), .ZN(n6161) );
  OAI222_X1 U2480 ( .A1(n1005), .A2(n635), .B1(n1037), .B2(n632), .C1(n973), 
        .C2(n629), .ZN(n6170) );
  OAI222_X1 U2481 ( .A1(n301), .A2(n1413), .B1(n333), .B2(n1410), .C1(n269), 
        .C2(n1407), .ZN(n4718) );
  OAI222_X1 U2482 ( .A1(n1005), .A2(n1347), .B1(n1037), .B2(n1344), .C1(n973), 
        .C2(n1341), .ZN(n4727) );
  OAI222_X1 U2483 ( .A1(n300), .A2(n701), .B1(n332), .B2(n698), .C1(n268), 
        .C2(n695), .ZN(n6120) );
  OAI222_X1 U2484 ( .A1(n1004), .A2(n635), .B1(n1036), .B2(n632), .C1(n972), 
        .C2(n629), .ZN(n6129) );
  OAI222_X1 U2485 ( .A1(n300), .A2(n1413), .B1(n332), .B2(n1410), .C1(n268), 
        .C2(n1407), .ZN(n4677) );
  OAI222_X1 U2486 ( .A1(n1004), .A2(n1347), .B1(n1036), .B2(n1344), .C1(n972), 
        .C2(n1341), .ZN(n4686) );
  OAI222_X1 U2487 ( .A1(n299), .A2(n701), .B1(n331), .B2(n698), .C1(n267), 
        .C2(n695), .ZN(n6079) );
  OAI222_X1 U2488 ( .A1(n1003), .A2(n635), .B1(n1035), .B2(n632), .C1(n971), 
        .C2(n629), .ZN(n6088) );
  OAI222_X1 U2489 ( .A1(n299), .A2(n1413), .B1(n331), .B2(n1410), .C1(n267), 
        .C2(n1407), .ZN(n4636) );
  OAI222_X1 U2490 ( .A1(n1003), .A2(n1347), .B1(n1035), .B2(n1344), .C1(n971), 
        .C2(n1341), .ZN(n4645) );
  OAI222_X1 U2491 ( .A1(n298), .A2(n701), .B1(n330), .B2(n698), .C1(n266), 
        .C2(n695), .ZN(n6038) );
  OAI222_X1 U2492 ( .A1(n1002), .A2(n635), .B1(n1034), .B2(n632), .C1(n970), 
        .C2(n629), .ZN(n6047) );
  OAI222_X1 U2493 ( .A1(n298), .A2(n1413), .B1(n330), .B2(n1410), .C1(n266), 
        .C2(n1407), .ZN(n4595) );
  OAI222_X1 U2494 ( .A1(n1002), .A2(n1347), .B1(n1034), .B2(n1344), .C1(n970), 
        .C2(n1341), .ZN(n4604) );
  OAI222_X1 U2495 ( .A1(n297), .A2(n701), .B1(n329), .B2(n698), .C1(n265), 
        .C2(n695), .ZN(n5997) );
  OAI222_X1 U2496 ( .A1(n1001), .A2(n635), .B1(n1033), .B2(n632), .C1(n969), 
        .C2(n629), .ZN(n6006) );
  OAI222_X1 U2497 ( .A1(n297), .A2(n1413), .B1(n329), .B2(n1410), .C1(n265), 
        .C2(n1407), .ZN(n4554) );
  OAI222_X1 U2498 ( .A1(n1001), .A2(n1347), .B1(n1033), .B2(n1344), .C1(n969), 
        .C2(n1341), .ZN(n4563) );
  OAI222_X1 U2499 ( .A1(n296), .A2(n701), .B1(n328), .B2(n698), .C1(n264), 
        .C2(n695), .ZN(n5956) );
  OAI222_X1 U2500 ( .A1(n1000), .A2(n635), .B1(n1032), .B2(n632), .C1(n968), 
        .C2(n629), .ZN(n5965) );
  OAI222_X1 U2501 ( .A1(n296), .A2(n1413), .B1(n328), .B2(n1410), .C1(n264), 
        .C2(n1407), .ZN(n4513) );
  OAI222_X1 U2502 ( .A1(n1000), .A2(n1347), .B1(n1032), .B2(n1344), .C1(n968), 
        .C2(n1341), .ZN(n4522) );
  OAI222_X1 U2503 ( .A1(n295), .A2(n701), .B1(n327), .B2(n698), .C1(n263), 
        .C2(n695), .ZN(n5915) );
  OAI222_X1 U2504 ( .A1(n999), .A2(n635), .B1(n1031), .B2(n632), .C1(n967), 
        .C2(n629), .ZN(n5924) );
  OAI222_X1 U2505 ( .A1(n295), .A2(n1413), .B1(n327), .B2(n1410), .C1(n263), 
        .C2(n1407), .ZN(n4472) );
  OAI222_X1 U2506 ( .A1(n999), .A2(n1347), .B1(n1031), .B2(n1344), .C1(n967), 
        .C2(n1341), .ZN(n4481) );
  OAI222_X1 U2507 ( .A1(n294), .A2(n701), .B1(n326), .B2(n698), .C1(n262), 
        .C2(n695), .ZN(n5874) );
  OAI222_X1 U2508 ( .A1(n998), .A2(n635), .B1(n1030), .B2(n632), .C1(n966), 
        .C2(n629), .ZN(n5883) );
  OAI222_X1 U2509 ( .A1(n294), .A2(n1413), .B1(n326), .B2(n1410), .C1(n262), 
        .C2(n1407), .ZN(n4431) );
  OAI222_X1 U2510 ( .A1(n998), .A2(n1347), .B1(n1030), .B2(n1344), .C1(n966), 
        .C2(n1341), .ZN(n4440) );
  OAI222_X1 U2511 ( .A1(n293), .A2(n701), .B1(n325), .B2(n698), .C1(n261), 
        .C2(n695), .ZN(n5833) );
  OAI222_X1 U2512 ( .A1(n997), .A2(n635), .B1(n1029), .B2(n632), .C1(n965), 
        .C2(n629), .ZN(n5842) );
  OAI222_X1 U2513 ( .A1(n293), .A2(n1413), .B1(n325), .B2(n1410), .C1(n261), 
        .C2(n1407), .ZN(n4390) );
  OAI222_X1 U2514 ( .A1(n997), .A2(n1347), .B1(n1029), .B2(n1344), .C1(n965), 
        .C2(n1341), .ZN(n4399) );
  OAI222_X1 U2515 ( .A1(n292), .A2(n701), .B1(n324), .B2(n698), .C1(n260), 
        .C2(n695), .ZN(n5792) );
  OAI222_X1 U2516 ( .A1(n996), .A2(n635), .B1(n1028), .B2(n632), .C1(n964), 
        .C2(n629), .ZN(n5801) );
  OAI222_X1 U2517 ( .A1(n292), .A2(n1413), .B1(n324), .B2(n1410), .C1(n260), 
        .C2(n1407), .ZN(n4349) );
  OAI222_X1 U2518 ( .A1(n996), .A2(n1347), .B1(n1028), .B2(n1344), .C1(n964), 
        .C2(n1341), .ZN(n4358) );
  OAI222_X1 U2519 ( .A1(n291), .A2(n702), .B1(n323), .B2(n699), .C1(n259), 
        .C2(n696), .ZN(n5751) );
  OAI222_X1 U2520 ( .A1(n995), .A2(n636), .B1(n1027), .B2(n633), .C1(n963), 
        .C2(n630), .ZN(n5760) );
  OAI222_X1 U2521 ( .A1(n291), .A2(n1414), .B1(n323), .B2(n1411), .C1(n259), 
        .C2(n1408), .ZN(n4308) );
  OAI222_X1 U2522 ( .A1(n995), .A2(n1348), .B1(n1027), .B2(n1345), .C1(n963), 
        .C2(n1342), .ZN(n4317) );
  OAI222_X1 U2523 ( .A1(n290), .A2(n702), .B1(n322), .B2(n699), .C1(n258), 
        .C2(n696), .ZN(n5710) );
  OAI222_X1 U2524 ( .A1(n994), .A2(n636), .B1(n1026), .B2(n633), .C1(n962), 
        .C2(n630), .ZN(n5719) );
  OAI222_X1 U2525 ( .A1(n290), .A2(n1414), .B1(n322), .B2(n1411), .C1(n258), 
        .C2(n1408), .ZN(n4267) );
  OAI222_X1 U2526 ( .A1(n994), .A2(n1348), .B1(n1026), .B2(n1345), .C1(n962), 
        .C2(n1342), .ZN(n4276) );
  OAI222_X1 U2527 ( .A1(n289), .A2(n702), .B1(n321), .B2(n699), .C1(n257), 
        .C2(n696), .ZN(n5669) );
  OAI222_X1 U2528 ( .A1(n993), .A2(n636), .B1(n1025), .B2(n633), .C1(n961), 
        .C2(n630), .ZN(n5678) );
  OAI222_X1 U2529 ( .A1(n289), .A2(n1414), .B1(n321), .B2(n1411), .C1(n257), 
        .C2(n1408), .ZN(n4226) );
  OAI222_X1 U2530 ( .A1(n993), .A2(n1348), .B1(n1025), .B2(n1345), .C1(n961), 
        .C2(n1342), .ZN(n4235) );
  OAI222_X1 U2531 ( .A1(n288), .A2(n702), .B1(n320), .B2(n699), .C1(n256), 
        .C2(n696), .ZN(n5628) );
  OAI222_X1 U2532 ( .A1(n992), .A2(n636), .B1(n1024), .B2(n633), .C1(n960), 
        .C2(n630), .ZN(n5637) );
  OAI222_X1 U2533 ( .A1(n288), .A2(n1414), .B1(n320), .B2(n1411), .C1(n256), 
        .C2(n1408), .ZN(n4185) );
  OAI222_X1 U2534 ( .A1(n992), .A2(n1348), .B1(n1024), .B2(n1345), .C1(n960), 
        .C2(n1342), .ZN(n4194) );
  OAI222_X1 U2535 ( .A1(n287), .A2(n702), .B1(n319), .B2(n699), .C1(n255), 
        .C2(n696), .ZN(n5587) );
  OAI222_X1 U2536 ( .A1(n991), .A2(n636), .B1(n1023), .B2(n633), .C1(n959), 
        .C2(n630), .ZN(n5596) );
  OAI222_X1 U2537 ( .A1(n287), .A2(n1414), .B1(n319), .B2(n1411), .C1(n255), 
        .C2(n1408), .ZN(n4144) );
  OAI222_X1 U2538 ( .A1(n991), .A2(n1348), .B1(n1023), .B2(n1345), .C1(n959), 
        .C2(n1342), .ZN(n4153) );
  OAI222_X1 U2539 ( .A1(n286), .A2(n702), .B1(n318), .B2(n699), .C1(n254), 
        .C2(n696), .ZN(n5546) );
  OAI222_X1 U2540 ( .A1(n990), .A2(n636), .B1(n1022), .B2(n633), .C1(n958), 
        .C2(n630), .ZN(n5555) );
  OAI222_X1 U2541 ( .A1(n286), .A2(n1414), .B1(n318), .B2(n1411), .C1(n254), 
        .C2(n1408), .ZN(n4103) );
  OAI222_X1 U2542 ( .A1(n990), .A2(n1348), .B1(n1022), .B2(n1345), .C1(n958), 
        .C2(n1342), .ZN(n4112) );
  OAI222_X1 U2543 ( .A1(n285), .A2(n702), .B1(n317), .B2(n699), .C1(n253), 
        .C2(n696), .ZN(n5505) );
  OAI222_X1 U2544 ( .A1(n989), .A2(n636), .B1(n1021), .B2(n633), .C1(n957), 
        .C2(n630), .ZN(n5514) );
  OAI222_X1 U2545 ( .A1(n285), .A2(n1414), .B1(n317), .B2(n1411), .C1(n253), 
        .C2(n1408), .ZN(n4062) );
  OAI222_X1 U2546 ( .A1(n989), .A2(n1348), .B1(n1021), .B2(n1345), .C1(n957), 
        .C2(n1342), .ZN(n4071) );
  OAI222_X1 U2547 ( .A1(n284), .A2(n702), .B1(n316), .B2(n699), .C1(n252), 
        .C2(n696), .ZN(n5464) );
  OAI222_X1 U2548 ( .A1(n988), .A2(n636), .B1(n1020), .B2(n633), .C1(n956), 
        .C2(n630), .ZN(n5473) );
  OAI222_X1 U2549 ( .A1(n284), .A2(n1414), .B1(n316), .B2(n1411), .C1(n252), 
        .C2(n1408), .ZN(n4021) );
  OAI222_X1 U2550 ( .A1(n988), .A2(n1348), .B1(n1020), .B2(n1345), .C1(n956), 
        .C2(n1342), .ZN(n4030) );
  OAI222_X1 U2551 ( .A1(n283), .A2(n702), .B1(n315), .B2(n699), .C1(n251), 
        .C2(n696), .ZN(n5423) );
  OAI222_X1 U2552 ( .A1(n987), .A2(n636), .B1(n1019), .B2(n633), .C1(n955), 
        .C2(n630), .ZN(n5432) );
  OAI222_X1 U2553 ( .A1(n283), .A2(n1414), .B1(n315), .B2(n1411), .C1(n251), 
        .C2(n1408), .ZN(n3980) );
  OAI222_X1 U2554 ( .A1(n987), .A2(n1348), .B1(n1019), .B2(n1345), .C1(n955), 
        .C2(n1342), .ZN(n3989) );
  OAI222_X1 U2555 ( .A1(n282), .A2(n702), .B1(n314), .B2(n699), .C1(n250), 
        .C2(n696), .ZN(n5382) );
  OAI222_X1 U2556 ( .A1(n986), .A2(n636), .B1(n1018), .B2(n633), .C1(n954), 
        .C2(n630), .ZN(n5391) );
  OAI222_X1 U2557 ( .A1(n282), .A2(n1414), .B1(n314), .B2(n1411), .C1(n250), 
        .C2(n1408), .ZN(n3939) );
  OAI222_X1 U2558 ( .A1(n986), .A2(n1348), .B1(n1018), .B2(n1345), .C1(n954), 
        .C2(n1342), .ZN(n3948) );
  OAI222_X1 U2559 ( .A1(n281), .A2(n702), .B1(n313), .B2(n699), .C1(n249), 
        .C2(n696), .ZN(n5341) );
  OAI222_X1 U2560 ( .A1(n985), .A2(n636), .B1(n1017), .B2(n633), .C1(n953), 
        .C2(n630), .ZN(n5350) );
  OAI222_X1 U2561 ( .A1(n281), .A2(n1414), .B1(n313), .B2(n1411), .C1(n249), 
        .C2(n1408), .ZN(n3898) );
  OAI222_X1 U2562 ( .A1(n985), .A2(n1348), .B1(n1017), .B2(n1345), .C1(n953), 
        .C2(n1342), .ZN(n3907) );
  OAI222_X1 U2563 ( .A1(n280), .A2(n702), .B1(n312), .B2(n699), .C1(n248), 
        .C2(n696), .ZN(n5300) );
  OAI222_X1 U2564 ( .A1(n984), .A2(n636), .B1(n1016), .B2(n633), .C1(n952), 
        .C2(n630), .ZN(n5309) );
  OAI222_X1 U2565 ( .A1(n280), .A2(n1414), .B1(n312), .B2(n1411), .C1(n248), 
        .C2(n1408), .ZN(n3857) );
  OAI222_X1 U2566 ( .A1(n984), .A2(n1348), .B1(n1016), .B2(n1345), .C1(n952), 
        .C2(n1342), .ZN(n3866) );
  OAI222_X1 U2567 ( .A1(n279), .A2(n703), .B1(n311), .B2(n700), .C1(n247), 
        .C2(n697), .ZN(n5259) );
  OAI222_X1 U2568 ( .A1(n983), .A2(n637), .B1(n1015), .B2(n634), .C1(n951), 
        .C2(n631), .ZN(n5268) );
  OAI222_X1 U2569 ( .A1(n279), .A2(n1415), .B1(n311), .B2(n1412), .C1(n247), 
        .C2(n1409), .ZN(n3816) );
  OAI222_X1 U2570 ( .A1(n983), .A2(n1349), .B1(n1015), .B2(n1346), .C1(n951), 
        .C2(n1343), .ZN(n3825) );
  OAI222_X1 U2571 ( .A1(n278), .A2(n703), .B1(n310), .B2(n700), .C1(n246), 
        .C2(n697), .ZN(n5218) );
  OAI222_X1 U2572 ( .A1(n982), .A2(n637), .B1(n1014), .B2(n634), .C1(n950), 
        .C2(n631), .ZN(n5227) );
  OAI222_X1 U2573 ( .A1(n278), .A2(n1415), .B1(n310), .B2(n1412), .C1(n246), 
        .C2(n1409), .ZN(n3775) );
  OAI222_X1 U2574 ( .A1(n982), .A2(n1349), .B1(n1014), .B2(n1346), .C1(n950), 
        .C2(n1343), .ZN(n3784) );
  OAI222_X1 U2575 ( .A1(n277), .A2(n703), .B1(n309), .B2(n700), .C1(n245), 
        .C2(n697), .ZN(n5177) );
  OAI222_X1 U2576 ( .A1(n981), .A2(n637), .B1(n1013), .B2(n634), .C1(n949), 
        .C2(n631), .ZN(n5186) );
  OAI222_X1 U2577 ( .A1(n277), .A2(n1415), .B1(n309), .B2(n1412), .C1(n245), 
        .C2(n1409), .ZN(n3734) );
  OAI222_X1 U2578 ( .A1(n981), .A2(n1349), .B1(n1013), .B2(n1346), .C1(n949), 
        .C2(n1343), .ZN(n3743) );
  OAI222_X1 U2579 ( .A1(n276), .A2(n703), .B1(n308), .B2(n700), .C1(n244), 
        .C2(n697), .ZN(n5136) );
  OAI222_X1 U2580 ( .A1(n980), .A2(n637), .B1(n1012), .B2(n634), .C1(n948), 
        .C2(n631), .ZN(n5145) );
  OAI222_X1 U2581 ( .A1(n276), .A2(n1415), .B1(n308), .B2(n1412), .C1(n244), 
        .C2(n1409), .ZN(n3693) );
  OAI222_X1 U2582 ( .A1(n980), .A2(n1349), .B1(n1012), .B2(n1346), .C1(n948), 
        .C2(n1343), .ZN(n3702) );
  OAI222_X1 U2583 ( .A1(n275), .A2(n703), .B1(n307), .B2(n700), .C1(n243), 
        .C2(n697), .ZN(n5095) );
  OAI222_X1 U2584 ( .A1(n979), .A2(n637), .B1(n1011), .B2(n634), .C1(n947), 
        .C2(n631), .ZN(n5104) );
  OAI222_X1 U2585 ( .A1(n275), .A2(n1415), .B1(n307), .B2(n1412), .C1(n243), 
        .C2(n1409), .ZN(n3652) );
  OAI222_X1 U2586 ( .A1(n979), .A2(n1349), .B1(n1011), .B2(n1346), .C1(n947), 
        .C2(n1343), .ZN(n3661) );
  OAI222_X1 U2587 ( .A1(n274), .A2(n703), .B1(n306), .B2(n700), .C1(n242), 
        .C2(n697), .ZN(n5054) );
  OAI222_X1 U2588 ( .A1(n978), .A2(n637), .B1(n1010), .B2(n634), .C1(n946), 
        .C2(n631), .ZN(n5063) );
  OAI222_X1 U2589 ( .A1(n274), .A2(n1415), .B1(n306), .B2(n1412), .C1(n242), 
        .C2(n1409), .ZN(n3611) );
  OAI222_X1 U2590 ( .A1(n978), .A2(n1349), .B1(n1010), .B2(n1346), .C1(n946), 
        .C2(n1343), .ZN(n3620) );
  OAI222_X1 U2591 ( .A1(n273), .A2(n703), .B1(n305), .B2(n700), .C1(n241), 
        .C2(n697), .ZN(n5013) );
  OAI222_X1 U2592 ( .A1(n977), .A2(n637), .B1(n1009), .B2(n634), .C1(n945), 
        .C2(n631), .ZN(n5022) );
  OAI222_X1 U2593 ( .A1(n273), .A2(n1415), .B1(n305), .B2(n1412), .C1(n241), 
        .C2(n1409), .ZN(n3570) );
  OAI222_X1 U2594 ( .A1(n977), .A2(n1349), .B1(n1009), .B2(n1346), .C1(n945), 
        .C2(n1343), .ZN(n3579) );
  OAI222_X1 U2595 ( .A1(n272), .A2(n703), .B1(n304), .B2(n700), .C1(n240), 
        .C2(n697), .ZN(n4884) );
  OAI222_X1 U2596 ( .A1(n976), .A2(n637), .B1(n1008), .B2(n634), .C1(n944), 
        .C2(n631), .ZN(n4915) );
  OAI222_X1 U2597 ( .A1(n272), .A2(n1415), .B1(n304), .B2(n1412), .C1(n240), 
        .C2(n1409), .ZN(n3441) );
  OAI222_X1 U2598 ( .A1(n976), .A2(n1349), .B1(n1008), .B2(n1346), .C1(n944), 
        .C2(n1343), .ZN(n3472) );
  OAI222_X1 U2599 ( .A1(n399), .A2(n692), .B1(n431), .B2(n689), .C1(n367), 
        .C2(n686), .ZN(n6242) );
  OAI222_X1 U2600 ( .A1(n1103), .A2(n626), .B1(n1135), .B2(n623), .C1(n1071), 
        .C2(n620), .ZN(n6273) );
  OAI222_X1 U2601 ( .A1(n399), .A2(n1404), .B1(n431), .B2(n1401), .C1(n367), 
        .C2(n1398), .ZN(n4799) );
  OAI222_X1 U2602 ( .A1(n1103), .A2(n1338), .B1(n1135), .B2(n1335), .C1(n1071), 
        .C2(n1332), .ZN(n4830) );
  OAI222_X1 U2603 ( .A1(n398), .A2(n692), .B1(n430), .B2(n689), .C1(n366), 
        .C2(n686), .ZN(n6201) );
  OAI222_X1 U2604 ( .A1(n1102), .A2(n626), .B1(n1134), .B2(n623), .C1(n1070), 
        .C2(n620), .ZN(n6210) );
  OAI222_X1 U2605 ( .A1(n398), .A2(n1404), .B1(n430), .B2(n1401), .C1(n366), 
        .C2(n1398), .ZN(n4758) );
  OAI222_X1 U2606 ( .A1(n1102), .A2(n1338), .B1(n1134), .B2(n1335), .C1(n1070), 
        .C2(n1332), .ZN(n4767) );
  OAI222_X1 U2607 ( .A1(n397), .A2(n692), .B1(n429), .B2(n689), .C1(n365), 
        .C2(n686), .ZN(n6160) );
  OAI222_X1 U2608 ( .A1(n1101), .A2(n626), .B1(n1133), .B2(n623), .C1(n1069), 
        .C2(n620), .ZN(n6169) );
  OAI222_X1 U2609 ( .A1(n397), .A2(n1404), .B1(n429), .B2(n1401), .C1(n365), 
        .C2(n1398), .ZN(n4717) );
  OAI222_X1 U2610 ( .A1(n1101), .A2(n1338), .B1(n1133), .B2(n1335), .C1(n1069), 
        .C2(n1332), .ZN(n4726) );
  OAI222_X1 U2611 ( .A1(n396), .A2(n692), .B1(n428), .B2(n689), .C1(n364), 
        .C2(n686), .ZN(n6119) );
  OAI222_X1 U2612 ( .A1(n1100), .A2(n626), .B1(n1132), .B2(n623), .C1(n1068), 
        .C2(n620), .ZN(n6128) );
  OAI222_X1 U2613 ( .A1(n396), .A2(n1404), .B1(n428), .B2(n1401), .C1(n364), 
        .C2(n1398), .ZN(n4676) );
  OAI222_X1 U2614 ( .A1(n1100), .A2(n1338), .B1(n1132), .B2(n1335), .C1(n1068), 
        .C2(n1332), .ZN(n4685) );
  OAI222_X1 U2615 ( .A1(n395), .A2(n692), .B1(n427), .B2(n689), .C1(n363), 
        .C2(n686), .ZN(n6078) );
  OAI222_X1 U2616 ( .A1(n1099), .A2(n626), .B1(n1131), .B2(n623), .C1(n1067), 
        .C2(n620), .ZN(n6087) );
  OAI222_X1 U2617 ( .A1(n395), .A2(n1404), .B1(n427), .B2(n1401), .C1(n363), 
        .C2(n1398), .ZN(n4635) );
  OAI222_X1 U2618 ( .A1(n1099), .A2(n1338), .B1(n1131), .B2(n1335), .C1(n1067), 
        .C2(n1332), .ZN(n4644) );
  OAI222_X1 U2619 ( .A1(n394), .A2(n692), .B1(n426), .B2(n689), .C1(n362), 
        .C2(n686), .ZN(n6037) );
  OAI222_X1 U2620 ( .A1(n1098), .A2(n626), .B1(n1130), .B2(n623), .C1(n1066), 
        .C2(n620), .ZN(n6046) );
  OAI222_X1 U2621 ( .A1(n394), .A2(n1404), .B1(n426), .B2(n1401), .C1(n362), 
        .C2(n1398), .ZN(n4594) );
  OAI222_X1 U2622 ( .A1(n1098), .A2(n1338), .B1(n1130), .B2(n1335), .C1(n1066), 
        .C2(n1332), .ZN(n4603) );
  OAI222_X1 U2623 ( .A1(n393), .A2(n692), .B1(n425), .B2(n689), .C1(n361), 
        .C2(n686), .ZN(n5996) );
  OAI222_X1 U2624 ( .A1(n1097), .A2(n626), .B1(n1129), .B2(n623), .C1(n1065), 
        .C2(n620), .ZN(n6005) );
  OAI222_X1 U2625 ( .A1(n393), .A2(n1404), .B1(n425), .B2(n1401), .C1(n361), 
        .C2(n1398), .ZN(n4553) );
  OAI222_X1 U2626 ( .A1(n1097), .A2(n1338), .B1(n1129), .B2(n1335), .C1(n1065), 
        .C2(n1332), .ZN(n4562) );
  OAI222_X1 U2627 ( .A1(n392), .A2(n692), .B1(n424), .B2(n689), .C1(n360), 
        .C2(n686), .ZN(n5955) );
  OAI222_X1 U2628 ( .A1(n1096), .A2(n626), .B1(n1128), .B2(n623), .C1(n1064), 
        .C2(n620), .ZN(n5964) );
  OAI222_X1 U2629 ( .A1(n392), .A2(n1404), .B1(n424), .B2(n1401), .C1(n360), 
        .C2(n1398), .ZN(n4512) );
  OAI222_X1 U2630 ( .A1(n1096), .A2(n1338), .B1(n1128), .B2(n1335), .C1(n1064), 
        .C2(n1332), .ZN(n4521) );
  OAI222_X1 U2631 ( .A1(n391), .A2(n692), .B1(n423), .B2(n689), .C1(n359), 
        .C2(n686), .ZN(n5914) );
  OAI222_X1 U2632 ( .A1(n1095), .A2(n626), .B1(n1127), .B2(n623), .C1(n1063), 
        .C2(n620), .ZN(n5923) );
  OAI222_X1 U2633 ( .A1(n391), .A2(n1404), .B1(n423), .B2(n1401), .C1(n359), 
        .C2(n1398), .ZN(n4471) );
  OAI222_X1 U2634 ( .A1(n1095), .A2(n1338), .B1(n1127), .B2(n1335), .C1(n1063), 
        .C2(n1332), .ZN(n4480) );
  OAI222_X1 U2635 ( .A1(n390), .A2(n692), .B1(n422), .B2(n689), .C1(n358), 
        .C2(n686), .ZN(n5873) );
  OAI222_X1 U2636 ( .A1(n1094), .A2(n626), .B1(n1126), .B2(n623), .C1(n1062), 
        .C2(n620), .ZN(n5882) );
  OAI222_X1 U2637 ( .A1(n390), .A2(n1404), .B1(n422), .B2(n1401), .C1(n358), 
        .C2(n1398), .ZN(n4430) );
  OAI222_X1 U2638 ( .A1(n1094), .A2(n1338), .B1(n1126), .B2(n1335), .C1(n1062), 
        .C2(n1332), .ZN(n4439) );
  OAI222_X1 U2639 ( .A1(n389), .A2(n692), .B1(n421), .B2(n689), .C1(n357), 
        .C2(n686), .ZN(n5832) );
  OAI222_X1 U2640 ( .A1(n1093), .A2(n626), .B1(n1125), .B2(n623), .C1(n1061), 
        .C2(n620), .ZN(n5841) );
  OAI222_X1 U2641 ( .A1(n389), .A2(n1404), .B1(n421), .B2(n1401), .C1(n357), 
        .C2(n1398), .ZN(n4389) );
  OAI222_X1 U2642 ( .A1(n1093), .A2(n1338), .B1(n1125), .B2(n1335), .C1(n1061), 
        .C2(n1332), .ZN(n4398) );
  OAI222_X1 U2643 ( .A1(n388), .A2(n692), .B1(n420), .B2(n689), .C1(n356), 
        .C2(n686), .ZN(n5791) );
  OAI222_X1 U2644 ( .A1(n1092), .A2(n626), .B1(n1124), .B2(n623), .C1(n1060), 
        .C2(n620), .ZN(n5800) );
  OAI222_X1 U2645 ( .A1(n388), .A2(n1404), .B1(n420), .B2(n1401), .C1(n356), 
        .C2(n1398), .ZN(n4348) );
  OAI222_X1 U2646 ( .A1(n1092), .A2(n1338), .B1(n1124), .B2(n1335), .C1(n1060), 
        .C2(n1332), .ZN(n4357) );
  OAI222_X1 U2647 ( .A1(n387), .A2(n693), .B1(n419), .B2(n690), .C1(n355), 
        .C2(n687), .ZN(n5750) );
  OAI222_X1 U2648 ( .A1(n1091), .A2(n627), .B1(n1123), .B2(n624), .C1(n1059), 
        .C2(n621), .ZN(n5759) );
  OAI222_X1 U2649 ( .A1(n387), .A2(n1405), .B1(n419), .B2(n1402), .C1(n355), 
        .C2(n1399), .ZN(n4307) );
  OAI222_X1 U2650 ( .A1(n1091), .A2(n1339), .B1(n1123), .B2(n1336), .C1(n1059), 
        .C2(n1333), .ZN(n4316) );
  OAI222_X1 U2651 ( .A1(n386), .A2(n693), .B1(n418), .B2(n690), .C1(n354), 
        .C2(n687), .ZN(n5709) );
  OAI222_X1 U2652 ( .A1(n1090), .A2(n627), .B1(n1122), .B2(n624), .C1(n1058), 
        .C2(n621), .ZN(n5718) );
  OAI222_X1 U2653 ( .A1(n386), .A2(n1405), .B1(n418), .B2(n1402), .C1(n354), 
        .C2(n1399), .ZN(n4266) );
  OAI222_X1 U2654 ( .A1(n1090), .A2(n1339), .B1(n1122), .B2(n1336), .C1(n1058), 
        .C2(n1333), .ZN(n4275) );
  OAI222_X1 U2655 ( .A1(n385), .A2(n693), .B1(n417), .B2(n690), .C1(n353), 
        .C2(n687), .ZN(n5668) );
  OAI222_X1 U2656 ( .A1(n1089), .A2(n627), .B1(n1121), .B2(n624), .C1(n1057), 
        .C2(n621), .ZN(n5677) );
  OAI222_X1 U2657 ( .A1(n385), .A2(n1405), .B1(n417), .B2(n1402), .C1(n353), 
        .C2(n1399), .ZN(n4225) );
  OAI222_X1 U2658 ( .A1(n1089), .A2(n1339), .B1(n1121), .B2(n1336), .C1(n1057), 
        .C2(n1333), .ZN(n4234) );
  OAI222_X1 U2659 ( .A1(n384), .A2(n693), .B1(n416), .B2(n690), .C1(n352), 
        .C2(n687), .ZN(n5627) );
  OAI222_X1 U2660 ( .A1(n1088), .A2(n627), .B1(n1120), .B2(n624), .C1(n1056), 
        .C2(n621), .ZN(n5636) );
  OAI222_X1 U2661 ( .A1(n384), .A2(n1405), .B1(n416), .B2(n1402), .C1(n352), 
        .C2(n1399), .ZN(n4184) );
  OAI222_X1 U2662 ( .A1(n1088), .A2(n1339), .B1(n1120), .B2(n1336), .C1(n1056), 
        .C2(n1333), .ZN(n4193) );
  OAI222_X1 U2663 ( .A1(n383), .A2(n693), .B1(n415), .B2(n690), .C1(n351), 
        .C2(n687), .ZN(n5586) );
  OAI222_X1 U2664 ( .A1(n1087), .A2(n627), .B1(n1119), .B2(n624), .C1(n1055), 
        .C2(n621), .ZN(n5595) );
  OAI222_X1 U2665 ( .A1(n383), .A2(n1405), .B1(n415), .B2(n1402), .C1(n351), 
        .C2(n1399), .ZN(n4143) );
  OAI222_X1 U2666 ( .A1(n1087), .A2(n1339), .B1(n1119), .B2(n1336), .C1(n1055), 
        .C2(n1333), .ZN(n4152) );
  OAI222_X1 U2667 ( .A1(n382), .A2(n693), .B1(n414), .B2(n690), .C1(n350), 
        .C2(n687), .ZN(n5545) );
  OAI222_X1 U2668 ( .A1(n1086), .A2(n627), .B1(n1118), .B2(n624), .C1(n1054), 
        .C2(n621), .ZN(n5554) );
  OAI222_X1 U2669 ( .A1(n382), .A2(n1405), .B1(n414), .B2(n1402), .C1(n350), 
        .C2(n1399), .ZN(n4102) );
  OAI222_X1 U2670 ( .A1(n1086), .A2(n1339), .B1(n1118), .B2(n1336), .C1(n1054), 
        .C2(n1333), .ZN(n4111) );
  OAI222_X1 U2671 ( .A1(n381), .A2(n693), .B1(n413), .B2(n690), .C1(n349), 
        .C2(n687), .ZN(n5504) );
  OAI222_X1 U2672 ( .A1(n1085), .A2(n627), .B1(n1117), .B2(n624), .C1(n1053), 
        .C2(n621), .ZN(n5513) );
  OAI222_X1 U2673 ( .A1(n381), .A2(n1405), .B1(n413), .B2(n1402), .C1(n349), 
        .C2(n1399), .ZN(n4061) );
  OAI222_X1 U2674 ( .A1(n1085), .A2(n1339), .B1(n1117), .B2(n1336), .C1(n1053), 
        .C2(n1333), .ZN(n4070) );
  OAI222_X1 U2675 ( .A1(n380), .A2(n693), .B1(n412), .B2(n690), .C1(n348), 
        .C2(n687), .ZN(n5463) );
  OAI222_X1 U2676 ( .A1(n1084), .A2(n627), .B1(n1116), .B2(n624), .C1(n1052), 
        .C2(n621), .ZN(n5472) );
  OAI222_X1 U2677 ( .A1(n380), .A2(n1405), .B1(n412), .B2(n1402), .C1(n348), 
        .C2(n1399), .ZN(n4020) );
  OAI222_X1 U2678 ( .A1(n1084), .A2(n1339), .B1(n1116), .B2(n1336), .C1(n1052), 
        .C2(n1333), .ZN(n4029) );
  OAI222_X1 U2679 ( .A1(n379), .A2(n693), .B1(n411), .B2(n690), .C1(n347), 
        .C2(n687), .ZN(n5422) );
  OAI222_X1 U2680 ( .A1(n1083), .A2(n627), .B1(n1115), .B2(n624), .C1(n1051), 
        .C2(n621), .ZN(n5431) );
  OAI222_X1 U2681 ( .A1(n379), .A2(n1405), .B1(n411), .B2(n1402), .C1(n347), 
        .C2(n1399), .ZN(n3979) );
  OAI222_X1 U2682 ( .A1(n1083), .A2(n1339), .B1(n1115), .B2(n1336), .C1(n1051), 
        .C2(n1333), .ZN(n3988) );
  OAI222_X1 U2683 ( .A1(n378), .A2(n693), .B1(n410), .B2(n690), .C1(n346), 
        .C2(n687), .ZN(n5381) );
  OAI222_X1 U2684 ( .A1(n1082), .A2(n627), .B1(n1114), .B2(n624), .C1(n1050), 
        .C2(n621), .ZN(n5390) );
  OAI222_X1 U2685 ( .A1(n378), .A2(n1405), .B1(n410), .B2(n1402), .C1(n346), 
        .C2(n1399), .ZN(n3938) );
  OAI222_X1 U2686 ( .A1(n1082), .A2(n1339), .B1(n1114), .B2(n1336), .C1(n1050), 
        .C2(n1333), .ZN(n3947) );
  OAI222_X1 U2687 ( .A1(n377), .A2(n693), .B1(n409), .B2(n690), .C1(n345), 
        .C2(n687), .ZN(n5340) );
  OAI222_X1 U2688 ( .A1(n1081), .A2(n627), .B1(n1113), .B2(n624), .C1(n1049), 
        .C2(n621), .ZN(n5349) );
  OAI222_X1 U2689 ( .A1(n377), .A2(n1405), .B1(n409), .B2(n1402), .C1(n345), 
        .C2(n1399), .ZN(n3897) );
  OAI222_X1 U2690 ( .A1(n1081), .A2(n1339), .B1(n1113), .B2(n1336), .C1(n1049), 
        .C2(n1333), .ZN(n3906) );
  OAI222_X1 U2691 ( .A1(n376), .A2(n693), .B1(n408), .B2(n690), .C1(n344), 
        .C2(n687), .ZN(n5299) );
  OAI222_X1 U2692 ( .A1(n1080), .A2(n627), .B1(n1112), .B2(n624), .C1(n1048), 
        .C2(n621), .ZN(n5308) );
  OAI222_X1 U2693 ( .A1(n376), .A2(n1405), .B1(n408), .B2(n1402), .C1(n344), 
        .C2(n1399), .ZN(n3856) );
  OAI222_X1 U2694 ( .A1(n1080), .A2(n1339), .B1(n1112), .B2(n1336), .C1(n1048), 
        .C2(n1333), .ZN(n3865) );
  OAI222_X1 U2695 ( .A1(n375), .A2(n694), .B1(n407), .B2(n691), .C1(n343), 
        .C2(n688), .ZN(n5258) );
  OAI222_X1 U2696 ( .A1(n1079), .A2(n628), .B1(n1111), .B2(n625), .C1(n1047), 
        .C2(n622), .ZN(n5267) );
  OAI222_X1 U2697 ( .A1(n375), .A2(n1406), .B1(n407), .B2(n1403), .C1(n343), 
        .C2(n1400), .ZN(n3815) );
  OAI222_X1 U2698 ( .A1(n1079), .A2(n1340), .B1(n1111), .B2(n1337), .C1(n1047), 
        .C2(n1334), .ZN(n3824) );
  OAI222_X1 U2699 ( .A1(n374), .A2(n694), .B1(n406), .B2(n691), .C1(n342), 
        .C2(n688), .ZN(n5217) );
  OAI222_X1 U2700 ( .A1(n1078), .A2(n628), .B1(n1110), .B2(n625), .C1(n1046), 
        .C2(n622), .ZN(n5226) );
  OAI222_X1 U2701 ( .A1(n374), .A2(n1406), .B1(n406), .B2(n1403), .C1(n342), 
        .C2(n1400), .ZN(n3774) );
  OAI222_X1 U2702 ( .A1(n1078), .A2(n1340), .B1(n1110), .B2(n1337), .C1(n1046), 
        .C2(n1334), .ZN(n3783) );
  OAI222_X1 U2703 ( .A1(n373), .A2(n694), .B1(n405), .B2(n691), .C1(n341), 
        .C2(n688), .ZN(n5176) );
  OAI222_X1 U2704 ( .A1(n1077), .A2(n628), .B1(n1109), .B2(n625), .C1(n1045), 
        .C2(n622), .ZN(n5185) );
  OAI222_X1 U2705 ( .A1(n373), .A2(n1406), .B1(n405), .B2(n1403), .C1(n341), 
        .C2(n1400), .ZN(n3733) );
  OAI222_X1 U2706 ( .A1(n1077), .A2(n1340), .B1(n1109), .B2(n1337), .C1(n1045), 
        .C2(n1334), .ZN(n3742) );
  OAI222_X1 U2707 ( .A1(n372), .A2(n694), .B1(n404), .B2(n691), .C1(n340), 
        .C2(n688), .ZN(n5135) );
  OAI222_X1 U2708 ( .A1(n1076), .A2(n628), .B1(n1108), .B2(n625), .C1(n1044), 
        .C2(n622), .ZN(n5144) );
  OAI222_X1 U2709 ( .A1(n372), .A2(n1406), .B1(n404), .B2(n1403), .C1(n340), 
        .C2(n1400), .ZN(n3692) );
  OAI222_X1 U2710 ( .A1(n1076), .A2(n1340), .B1(n1108), .B2(n1337), .C1(n1044), 
        .C2(n1334), .ZN(n3701) );
  OAI222_X1 U2711 ( .A1(n371), .A2(n694), .B1(n403), .B2(n691), .C1(n339), 
        .C2(n688), .ZN(n5094) );
  OAI222_X1 U2712 ( .A1(n1075), .A2(n628), .B1(n1107), .B2(n625), .C1(n1043), 
        .C2(n622), .ZN(n5103) );
  OAI222_X1 U2713 ( .A1(n371), .A2(n1406), .B1(n403), .B2(n1403), .C1(n339), 
        .C2(n1400), .ZN(n3651) );
  OAI222_X1 U2714 ( .A1(n1075), .A2(n1340), .B1(n1107), .B2(n1337), .C1(n1043), 
        .C2(n1334), .ZN(n3660) );
  OAI222_X1 U2715 ( .A1(n370), .A2(n694), .B1(n402), .B2(n691), .C1(n338), 
        .C2(n688), .ZN(n5053) );
  OAI222_X1 U2716 ( .A1(n1074), .A2(n628), .B1(n1106), .B2(n625), .C1(n1042), 
        .C2(n622), .ZN(n5062) );
  OAI222_X1 U2717 ( .A1(n370), .A2(n1406), .B1(n402), .B2(n1403), .C1(n338), 
        .C2(n1400), .ZN(n3610) );
  OAI222_X1 U2718 ( .A1(n1074), .A2(n1340), .B1(n1106), .B2(n1337), .C1(n1042), 
        .C2(n1334), .ZN(n3619) );
  OAI222_X1 U2719 ( .A1(n369), .A2(n694), .B1(n401), .B2(n691), .C1(n337), 
        .C2(n688), .ZN(n5012) );
  OAI222_X1 U2720 ( .A1(n1073), .A2(n628), .B1(n1105), .B2(n625), .C1(n1041), 
        .C2(n622), .ZN(n5021) );
  OAI222_X1 U2721 ( .A1(n369), .A2(n1406), .B1(n401), .B2(n1403), .C1(n337), 
        .C2(n1400), .ZN(n3569) );
  OAI222_X1 U2722 ( .A1(n1073), .A2(n1340), .B1(n1105), .B2(n1337), .C1(n1041), 
        .C2(n1334), .ZN(n3578) );
  OAI222_X1 U2723 ( .A1(n368), .A2(n694), .B1(n400), .B2(n691), .C1(n336), 
        .C2(n688), .ZN(n4883) );
  OAI222_X1 U2724 ( .A1(n1072), .A2(n628), .B1(n1104), .B2(n625), .C1(n1040), 
        .C2(n622), .ZN(n4914) );
  OAI222_X1 U2725 ( .A1(n368), .A2(n1406), .B1(n400), .B2(n1403), .C1(n336), 
        .C2(n1400), .ZN(n3440) );
  OAI222_X1 U2726 ( .A1(n1072), .A2(n1340), .B1(n1104), .B2(n1337), .C1(n1040), 
        .C2(n1334), .ZN(n3471) );
  AOI222_X1 U2727 ( .A1(n79), .A2(\REGISTERS[49][0] ), .B1(n78), .B2(
        \REGISTERS[51][0] ), .C1(n75), .C2(\REGISTERS[50][0] ), .ZN(n6288) );
  AOI222_X1 U2728 ( .A1(n12), .A2(\REGISTERS[82][0] ), .B1(n10), .B2(
        \REGISTERS[84][0] ), .C1(n6), .C2(\REGISTERS[83][0] ), .ZN(n6301) );
  AOI222_X1 U2729 ( .A1(n1143), .A2(\REGISTERS[49][0] ), .B1(n1142), .B2(
        \REGISTERS[51][0] ), .C1(n1139), .C2(\REGISTERS[50][0] ), .ZN(n4845)
         );
  AOI222_X1 U2730 ( .A1(n725), .A2(\REGISTERS[82][0] ), .B1(n724), .B2(
        \REGISTERS[84][0] ), .C1(n721), .C2(\REGISTERS[83][0] ), .ZN(n4858) );
  AOI222_X1 U2731 ( .A1(n79), .A2(\REGISTERS[49][1] ), .B1(n78), .B2(
        \REGISTERS[51][1] ), .C1(n75), .C2(\REGISTERS[50][1] ), .ZN(n6215) );
  AOI222_X1 U2732 ( .A1(n12), .A2(\REGISTERS[82][1] ), .B1(n10), .B2(
        \REGISTERS[84][1] ), .C1(n6), .C2(\REGISTERS[83][1] ), .ZN(n6224) );
  AOI222_X1 U2733 ( .A1(n1143), .A2(\REGISTERS[49][1] ), .B1(n1142), .B2(
        \REGISTERS[51][1] ), .C1(n1139), .C2(\REGISTERS[50][1] ), .ZN(n4772)
         );
  AOI222_X1 U2734 ( .A1(n725), .A2(\REGISTERS[82][1] ), .B1(n724), .B2(
        \REGISTERS[84][1] ), .C1(n721), .C2(\REGISTERS[83][1] ), .ZN(n4781) );
  AOI222_X1 U2735 ( .A1(n79), .A2(\REGISTERS[49][2] ), .B1(n78), .B2(
        \REGISTERS[51][2] ), .C1(n75), .C2(\REGISTERS[50][2] ), .ZN(n6174) );
  AOI222_X1 U2736 ( .A1(n12), .A2(\REGISTERS[82][2] ), .B1(n10), .B2(
        \REGISTERS[84][2] ), .C1(n6), .C2(\REGISTERS[83][2] ), .ZN(n6183) );
  AOI222_X1 U2737 ( .A1(n1143), .A2(\REGISTERS[49][2] ), .B1(n1142), .B2(
        \REGISTERS[51][2] ), .C1(n1139), .C2(\REGISTERS[50][2] ), .ZN(n4731)
         );
  AOI222_X1 U2738 ( .A1(n725), .A2(\REGISTERS[82][2] ), .B1(n724), .B2(
        \REGISTERS[84][2] ), .C1(n721), .C2(\REGISTERS[83][2] ), .ZN(n4740) );
  AOI222_X1 U2739 ( .A1(n79), .A2(\REGISTERS[49][3] ), .B1(n78), .B2(
        \REGISTERS[51][3] ), .C1(n75), .C2(\REGISTERS[50][3] ), .ZN(n6133) );
  AOI222_X1 U2740 ( .A1(n12), .A2(\REGISTERS[82][3] ), .B1(n10), .B2(
        \REGISTERS[84][3] ), .C1(n6), .C2(\REGISTERS[83][3] ), .ZN(n6142) );
  AOI222_X1 U2741 ( .A1(n1143), .A2(\REGISTERS[49][3] ), .B1(n1142), .B2(
        \REGISTERS[51][3] ), .C1(n1139), .C2(\REGISTERS[50][3] ), .ZN(n4690)
         );
  AOI222_X1 U2742 ( .A1(n725), .A2(\REGISTERS[82][3] ), .B1(n724), .B2(
        \REGISTERS[84][3] ), .C1(n721), .C2(\REGISTERS[83][3] ), .ZN(n4699) );
  AOI222_X1 U2743 ( .A1(n79), .A2(\REGISTERS[49][4] ), .B1(n78), .B2(
        \REGISTERS[51][4] ), .C1(n75), .C2(\REGISTERS[50][4] ), .ZN(n6092) );
  AOI222_X1 U2744 ( .A1(n12), .A2(\REGISTERS[82][4] ), .B1(n10), .B2(
        \REGISTERS[84][4] ), .C1(n6), .C2(\REGISTERS[83][4] ), .ZN(n6101) );
  AOI222_X1 U2745 ( .A1(n1143), .A2(\REGISTERS[49][4] ), .B1(n1142), .B2(
        \REGISTERS[51][4] ), .C1(n1139), .C2(\REGISTERS[50][4] ), .ZN(n4649)
         );
  AOI222_X1 U2746 ( .A1(n725), .A2(\REGISTERS[82][4] ), .B1(n724), .B2(
        \REGISTERS[84][4] ), .C1(n721), .C2(\REGISTERS[83][4] ), .ZN(n4658) );
  AOI222_X1 U2747 ( .A1(n79), .A2(\REGISTERS[49][5] ), .B1(n78), .B2(
        \REGISTERS[51][5] ), .C1(n75), .C2(\REGISTERS[50][5] ), .ZN(n6051) );
  AOI222_X1 U2748 ( .A1(n12), .A2(\REGISTERS[82][5] ), .B1(n10), .B2(
        \REGISTERS[84][5] ), .C1(n6), .C2(\REGISTERS[83][5] ), .ZN(n6060) );
  AOI222_X1 U2749 ( .A1(n1143), .A2(\REGISTERS[49][5] ), .B1(n1142), .B2(
        \REGISTERS[51][5] ), .C1(n1139), .C2(\REGISTERS[50][5] ), .ZN(n4608)
         );
  AOI222_X1 U2750 ( .A1(n725), .A2(\REGISTERS[82][5] ), .B1(n724), .B2(
        \REGISTERS[84][5] ), .C1(n721), .C2(\REGISTERS[83][5] ), .ZN(n4617) );
  AOI222_X1 U2751 ( .A1(n79), .A2(\REGISTERS[49][6] ), .B1(n78), .B2(
        \REGISTERS[51][6] ), .C1(n75), .C2(\REGISTERS[50][6] ), .ZN(n6010) );
  AOI222_X1 U2752 ( .A1(n12), .A2(\REGISTERS[82][6] ), .B1(n10), .B2(
        \REGISTERS[84][6] ), .C1(n6), .C2(\REGISTERS[83][6] ), .ZN(n6019) );
  AOI222_X1 U2753 ( .A1(n1143), .A2(\REGISTERS[49][6] ), .B1(n1142), .B2(
        \REGISTERS[51][6] ), .C1(n1139), .C2(\REGISTERS[50][6] ), .ZN(n4567)
         );
  AOI222_X1 U2754 ( .A1(n725), .A2(\REGISTERS[82][6] ), .B1(n724), .B2(
        \REGISTERS[84][6] ), .C1(n721), .C2(\REGISTERS[83][6] ), .ZN(n4576) );
  AOI222_X1 U2755 ( .A1(n79), .A2(\REGISTERS[49][7] ), .B1(n78), .B2(
        \REGISTERS[51][7] ), .C1(n75), .C2(\REGISTERS[50][7] ), .ZN(n5969) );
  AOI222_X1 U2756 ( .A1(n12), .A2(\REGISTERS[82][7] ), .B1(n10), .B2(
        \REGISTERS[84][7] ), .C1(n6), .C2(\REGISTERS[83][7] ), .ZN(n5978) );
  AOI222_X1 U2757 ( .A1(n1143), .A2(\REGISTERS[49][7] ), .B1(n1142), .B2(
        \REGISTERS[51][7] ), .C1(n1139), .C2(\REGISTERS[50][7] ), .ZN(n4526)
         );
  AOI222_X1 U2758 ( .A1(n725), .A2(\REGISTERS[82][7] ), .B1(n724), .B2(
        \REGISTERS[84][7] ), .C1(n721), .C2(\REGISTERS[83][7] ), .ZN(n4535) );
  AOI222_X1 U2759 ( .A1(n79), .A2(\REGISTERS[49][8] ), .B1(n77), .B2(
        \REGISTERS[51][8] ), .C1(n74), .C2(\REGISTERS[50][8] ), .ZN(n5928) );
  AOI222_X1 U2760 ( .A1(n12), .A2(\REGISTERS[82][8] ), .B1(n9), .B2(
        \REGISTERS[84][8] ), .C1(n5), .C2(\REGISTERS[83][8] ), .ZN(n5937) );
  AOI222_X1 U2761 ( .A1(n1143), .A2(\REGISTERS[49][8] ), .B1(n1141), .B2(
        \REGISTERS[51][8] ), .C1(n1138), .C2(\REGISTERS[50][8] ), .ZN(n4485)
         );
  AOI222_X1 U2762 ( .A1(n725), .A2(\REGISTERS[82][8] ), .B1(n723), .B2(
        \REGISTERS[84][8] ), .C1(n720), .C2(\REGISTERS[83][8] ), .ZN(n4494) );
  AOI222_X1 U2763 ( .A1(n79), .A2(\REGISTERS[49][9] ), .B1(n77), .B2(
        \REGISTERS[51][9] ), .C1(n74), .C2(\REGISTERS[50][9] ), .ZN(n5887) );
  AOI222_X1 U2764 ( .A1(n12), .A2(\REGISTERS[82][9] ), .B1(n9), .B2(
        \REGISTERS[84][9] ), .C1(n5), .C2(\REGISTERS[83][9] ), .ZN(n5896) );
  AOI222_X1 U2765 ( .A1(n1143), .A2(\REGISTERS[49][9] ), .B1(n1141), .B2(
        \REGISTERS[51][9] ), .C1(n1138), .C2(\REGISTERS[50][9] ), .ZN(n4444)
         );
  AOI222_X1 U2766 ( .A1(n725), .A2(\REGISTERS[82][9] ), .B1(n723), .B2(
        \REGISTERS[84][9] ), .C1(n720), .C2(\REGISTERS[83][9] ), .ZN(n4453) );
  AOI222_X1 U2767 ( .A1(n79), .A2(\REGISTERS[49][10] ), .B1(n77), .B2(
        \REGISTERS[51][10] ), .C1(n74), .C2(\REGISTERS[50][10] ), .ZN(n5846)
         );
  AOI222_X1 U2768 ( .A1(n12), .A2(\REGISTERS[82][10] ), .B1(n9), .B2(
        \REGISTERS[84][10] ), .C1(n5), .C2(\REGISTERS[83][10] ), .ZN(n5855) );
  AOI222_X1 U2769 ( .A1(n1143), .A2(\REGISTERS[49][10] ), .B1(n1141), .B2(
        \REGISTERS[51][10] ), .C1(n1138), .C2(\REGISTERS[50][10] ), .ZN(n4403)
         );
  AOI222_X1 U2770 ( .A1(n725), .A2(\REGISTERS[82][10] ), .B1(n723), .B2(
        \REGISTERS[84][10] ), .C1(n720), .C2(\REGISTERS[83][10] ), .ZN(n4412)
         );
  AOI222_X1 U2771 ( .A1(n79), .A2(\REGISTERS[49][11] ), .B1(n77), .B2(
        \REGISTERS[51][11] ), .C1(n74), .C2(\REGISTERS[50][11] ), .ZN(n5805)
         );
  AOI222_X1 U2772 ( .A1(n12), .A2(\REGISTERS[82][11] ), .B1(n9), .B2(
        \REGISTERS[84][11] ), .C1(n5), .C2(\REGISTERS[83][11] ), .ZN(n5814) );
  AOI222_X1 U2773 ( .A1(n1143), .A2(\REGISTERS[49][11] ), .B1(n1141), .B2(
        \REGISTERS[51][11] ), .C1(n1138), .C2(\REGISTERS[50][11] ), .ZN(n4362)
         );
  AOI222_X1 U2774 ( .A1(n725), .A2(\REGISTERS[82][11] ), .B1(n723), .B2(
        \REGISTERS[84][11] ), .C1(n720), .C2(\REGISTERS[83][11] ), .ZN(n4371)
         );
  AOI222_X1 U2775 ( .A1(n432), .A2(\REGISTERS[49][12] ), .B1(n77), .B2(
        \REGISTERS[51][12] ), .C1(n74), .C2(\REGISTERS[50][12] ), .ZN(n5764)
         );
  AOI222_X1 U2776 ( .A1(n13), .A2(\REGISTERS[82][12] ), .B1(n9), .B2(
        \REGISTERS[84][12] ), .C1(n5), .C2(\REGISTERS[83][12] ), .ZN(n5773) );
  AOI222_X1 U2777 ( .A1(n1144), .A2(\REGISTERS[49][12] ), .B1(n1141), .B2(
        \REGISTERS[51][12] ), .C1(n1138), .C2(\REGISTERS[50][12] ), .ZN(n4321)
         );
  AOI222_X1 U2778 ( .A1(n726), .A2(\REGISTERS[82][12] ), .B1(n723), .B2(
        \REGISTERS[84][12] ), .C1(n720), .C2(\REGISTERS[83][12] ), .ZN(n4330)
         );
  AOI222_X1 U2779 ( .A1(n432), .A2(\REGISTERS[49][13] ), .B1(n77), .B2(
        \REGISTERS[51][13] ), .C1(n74), .C2(\REGISTERS[50][13] ), .ZN(n5723)
         );
  AOI222_X1 U2780 ( .A1(n13), .A2(\REGISTERS[82][13] ), .B1(n9), .B2(
        \REGISTERS[84][13] ), .C1(n5), .C2(\REGISTERS[83][13] ), .ZN(n5732) );
  AOI222_X1 U2781 ( .A1(n1144), .A2(\REGISTERS[49][13] ), .B1(n1141), .B2(
        \REGISTERS[51][13] ), .C1(n1138), .C2(\REGISTERS[50][13] ), .ZN(n4280)
         );
  AOI222_X1 U2782 ( .A1(n726), .A2(\REGISTERS[82][13] ), .B1(n723), .B2(
        \REGISTERS[84][13] ), .C1(n720), .C2(\REGISTERS[83][13] ), .ZN(n4289)
         );
  AOI222_X1 U2783 ( .A1(n432), .A2(\REGISTERS[49][14] ), .B1(n77), .B2(
        \REGISTERS[51][14] ), .C1(n74), .C2(\REGISTERS[50][14] ), .ZN(n5682)
         );
  AOI222_X1 U2784 ( .A1(n13), .A2(\REGISTERS[82][14] ), .B1(n9), .B2(
        \REGISTERS[84][14] ), .C1(n5), .C2(\REGISTERS[83][14] ), .ZN(n5691) );
  AOI222_X1 U2785 ( .A1(n1144), .A2(\REGISTERS[49][14] ), .B1(n1141), .B2(
        \REGISTERS[51][14] ), .C1(n1138), .C2(\REGISTERS[50][14] ), .ZN(n4239)
         );
  AOI222_X1 U2786 ( .A1(n726), .A2(\REGISTERS[82][14] ), .B1(n723), .B2(
        \REGISTERS[84][14] ), .C1(n720), .C2(\REGISTERS[83][14] ), .ZN(n4248)
         );
  AOI222_X1 U2787 ( .A1(n432), .A2(\REGISTERS[49][15] ), .B1(n77), .B2(
        \REGISTERS[51][15] ), .C1(n74), .C2(\REGISTERS[50][15] ), .ZN(n5641)
         );
  AOI222_X1 U2788 ( .A1(n13), .A2(\REGISTERS[82][15] ), .B1(n9), .B2(
        \REGISTERS[84][15] ), .C1(n5), .C2(\REGISTERS[83][15] ), .ZN(n5650) );
  AOI222_X1 U2789 ( .A1(n1144), .A2(\REGISTERS[49][15] ), .B1(n1141), .B2(
        \REGISTERS[51][15] ), .C1(n1138), .C2(\REGISTERS[50][15] ), .ZN(n4198)
         );
  AOI222_X1 U2790 ( .A1(n726), .A2(\REGISTERS[82][15] ), .B1(n723), .B2(
        \REGISTERS[84][15] ), .C1(n720), .C2(\REGISTERS[83][15] ), .ZN(n4207)
         );
  AOI222_X1 U2791 ( .A1(n432), .A2(\REGISTERS[49][16] ), .B1(n77), .B2(
        \REGISTERS[51][16] ), .C1(n74), .C2(\REGISTERS[50][16] ), .ZN(n5600)
         );
  AOI222_X1 U2792 ( .A1(n13), .A2(\REGISTERS[82][16] ), .B1(n9), .B2(
        \REGISTERS[84][16] ), .C1(n5), .C2(\REGISTERS[83][16] ), .ZN(n5609) );
  AOI222_X1 U2793 ( .A1(n1144), .A2(\REGISTERS[49][16] ), .B1(n1141), .B2(
        \REGISTERS[51][16] ), .C1(n1138), .C2(\REGISTERS[50][16] ), .ZN(n4157)
         );
  AOI222_X1 U2794 ( .A1(n726), .A2(\REGISTERS[82][16] ), .B1(n723), .B2(
        \REGISTERS[84][16] ), .C1(n720), .C2(\REGISTERS[83][16] ), .ZN(n4166)
         );
  AOI222_X1 U2795 ( .A1(n432), .A2(\REGISTERS[49][17] ), .B1(n77), .B2(
        \REGISTERS[51][17] ), .C1(n74), .C2(\REGISTERS[50][17] ), .ZN(n5559)
         );
  AOI222_X1 U2796 ( .A1(n13), .A2(\REGISTERS[82][17] ), .B1(n9), .B2(
        \REGISTERS[84][17] ), .C1(n5), .C2(\REGISTERS[83][17] ), .ZN(n5568) );
  AOI222_X1 U2797 ( .A1(n1144), .A2(\REGISTERS[49][17] ), .B1(n1141), .B2(
        \REGISTERS[51][17] ), .C1(n1138), .C2(\REGISTERS[50][17] ), .ZN(n4116)
         );
  AOI222_X1 U2798 ( .A1(n726), .A2(\REGISTERS[82][17] ), .B1(n723), .B2(
        \REGISTERS[84][17] ), .C1(n720), .C2(\REGISTERS[83][17] ), .ZN(n4125)
         );
  AOI222_X1 U2799 ( .A1(n432), .A2(\REGISTERS[49][18] ), .B1(n77), .B2(
        \REGISTERS[51][18] ), .C1(n74), .C2(\REGISTERS[50][18] ), .ZN(n5518)
         );
  AOI222_X1 U2800 ( .A1(n13), .A2(\REGISTERS[82][18] ), .B1(n9), .B2(
        \REGISTERS[84][18] ), .C1(n5), .C2(\REGISTERS[83][18] ), .ZN(n5527) );
  AOI222_X1 U2801 ( .A1(n1144), .A2(\REGISTERS[49][18] ), .B1(n1141), .B2(
        \REGISTERS[51][18] ), .C1(n1138), .C2(\REGISTERS[50][18] ), .ZN(n4075)
         );
  AOI222_X1 U2802 ( .A1(n726), .A2(\REGISTERS[82][18] ), .B1(n723), .B2(
        \REGISTERS[84][18] ), .C1(n720), .C2(\REGISTERS[83][18] ), .ZN(n4084)
         );
  AOI222_X1 U2803 ( .A1(n432), .A2(\REGISTERS[49][19] ), .B1(n77), .B2(
        \REGISTERS[51][19] ), .C1(n74), .C2(\REGISTERS[50][19] ), .ZN(n5477)
         );
  AOI222_X1 U2804 ( .A1(n13), .A2(\REGISTERS[82][19] ), .B1(n9), .B2(
        \REGISTERS[84][19] ), .C1(n5), .C2(\REGISTERS[83][19] ), .ZN(n5486) );
  AOI222_X1 U2805 ( .A1(n1144), .A2(\REGISTERS[49][19] ), .B1(n1141), .B2(
        \REGISTERS[51][19] ), .C1(n1138), .C2(\REGISTERS[50][19] ), .ZN(n4034)
         );
  AOI222_X1 U2806 ( .A1(n726), .A2(\REGISTERS[82][19] ), .B1(n723), .B2(
        \REGISTERS[84][19] ), .C1(n720), .C2(\REGISTERS[83][19] ), .ZN(n4043)
         );
  AOI222_X1 U2807 ( .A1(n432), .A2(\REGISTERS[49][20] ), .B1(n76), .B2(
        \REGISTERS[51][20] ), .C1(n73), .C2(\REGISTERS[50][20] ), .ZN(n5436)
         );
  AOI222_X1 U2808 ( .A1(n13), .A2(\REGISTERS[82][20] ), .B1(n8), .B2(
        \REGISTERS[84][20] ), .C1(n4), .C2(\REGISTERS[83][20] ), .ZN(n5445) );
  AOI222_X1 U2809 ( .A1(n1144), .A2(\REGISTERS[49][20] ), .B1(n1140), .B2(
        \REGISTERS[51][20] ), .C1(n1137), .C2(\REGISTERS[50][20] ), .ZN(n3993)
         );
  AOI222_X1 U2810 ( .A1(n726), .A2(\REGISTERS[82][20] ), .B1(n722), .B2(
        \REGISTERS[84][20] ), .C1(n719), .C2(\REGISTERS[83][20] ), .ZN(n4002)
         );
  AOI222_X1 U2811 ( .A1(n432), .A2(\REGISTERS[49][21] ), .B1(n76), .B2(
        \REGISTERS[51][21] ), .C1(n73), .C2(\REGISTERS[50][21] ), .ZN(n5395)
         );
  AOI222_X1 U2812 ( .A1(n13), .A2(\REGISTERS[82][21] ), .B1(n8), .B2(
        \REGISTERS[84][21] ), .C1(n4), .C2(\REGISTERS[83][21] ), .ZN(n5404) );
  AOI222_X1 U2813 ( .A1(n1144), .A2(\REGISTERS[49][21] ), .B1(n1140), .B2(
        \REGISTERS[51][21] ), .C1(n1137), .C2(\REGISTERS[50][21] ), .ZN(n3952)
         );
  AOI222_X1 U2814 ( .A1(n726), .A2(\REGISTERS[82][21] ), .B1(n722), .B2(
        \REGISTERS[84][21] ), .C1(n719), .C2(\REGISTERS[83][21] ), .ZN(n3961)
         );
  AOI222_X1 U2815 ( .A1(n432), .A2(\REGISTERS[49][22] ), .B1(n76), .B2(
        \REGISTERS[51][22] ), .C1(n73), .C2(\REGISTERS[50][22] ), .ZN(n5354)
         );
  AOI222_X1 U2816 ( .A1(n13), .A2(\REGISTERS[82][22] ), .B1(n8), .B2(
        \REGISTERS[84][22] ), .C1(n4), .C2(\REGISTERS[83][22] ), .ZN(n5363) );
  AOI222_X1 U2817 ( .A1(n1144), .A2(\REGISTERS[49][22] ), .B1(n1140), .B2(
        \REGISTERS[51][22] ), .C1(n1137), .C2(\REGISTERS[50][22] ), .ZN(n3911)
         );
  AOI222_X1 U2818 ( .A1(n726), .A2(\REGISTERS[82][22] ), .B1(n722), .B2(
        \REGISTERS[84][22] ), .C1(n719), .C2(\REGISTERS[83][22] ), .ZN(n3920)
         );
  AOI222_X1 U2819 ( .A1(n432), .A2(\REGISTERS[49][23] ), .B1(n76), .B2(
        \REGISTERS[51][23] ), .C1(n73), .C2(\REGISTERS[50][23] ), .ZN(n5313)
         );
  AOI222_X1 U2820 ( .A1(n13), .A2(\REGISTERS[82][23] ), .B1(n8), .B2(
        \REGISTERS[84][23] ), .C1(n4), .C2(\REGISTERS[83][23] ), .ZN(n5322) );
  AOI222_X1 U2821 ( .A1(n1144), .A2(\REGISTERS[49][23] ), .B1(n1140), .B2(
        \REGISTERS[51][23] ), .C1(n1137), .C2(\REGISTERS[50][23] ), .ZN(n3870)
         );
  AOI222_X1 U2822 ( .A1(n726), .A2(\REGISTERS[82][23] ), .B1(n722), .B2(
        \REGISTERS[84][23] ), .C1(n719), .C2(\REGISTERS[83][23] ), .ZN(n3879)
         );
  AOI222_X1 U2823 ( .A1(n433), .A2(\REGISTERS[49][24] ), .B1(n76), .B2(
        \REGISTERS[51][24] ), .C1(n73), .C2(\REGISTERS[50][24] ), .ZN(n5272)
         );
  AOI222_X1 U2824 ( .A1(n14), .A2(\REGISTERS[82][24] ), .B1(n8), .B2(
        \REGISTERS[84][24] ), .C1(n4), .C2(\REGISTERS[83][24] ), .ZN(n5281) );
  AOI222_X1 U2825 ( .A1(n1145), .A2(\REGISTERS[49][24] ), .B1(n1140), .B2(
        \REGISTERS[51][24] ), .C1(n1137), .C2(\REGISTERS[50][24] ), .ZN(n3829)
         );
  AOI222_X1 U2826 ( .A1(n727), .A2(\REGISTERS[82][24] ), .B1(n722), .B2(
        \REGISTERS[84][24] ), .C1(n719), .C2(\REGISTERS[83][24] ), .ZN(n3838)
         );
  AOI222_X1 U2827 ( .A1(n433), .A2(\REGISTERS[49][25] ), .B1(n76), .B2(
        \REGISTERS[51][25] ), .C1(n73), .C2(\REGISTERS[50][25] ), .ZN(n5231)
         );
  AOI222_X1 U2828 ( .A1(n14), .A2(\REGISTERS[82][25] ), .B1(n8), .B2(
        \REGISTERS[84][25] ), .C1(n4), .C2(\REGISTERS[83][25] ), .ZN(n5240) );
  AOI222_X1 U2829 ( .A1(n1145), .A2(\REGISTERS[49][25] ), .B1(n1140), .B2(
        \REGISTERS[51][25] ), .C1(n1137), .C2(\REGISTERS[50][25] ), .ZN(n3788)
         );
  AOI222_X1 U2830 ( .A1(n727), .A2(\REGISTERS[82][25] ), .B1(n722), .B2(
        \REGISTERS[84][25] ), .C1(n719), .C2(\REGISTERS[83][25] ), .ZN(n3797)
         );
  AOI222_X1 U2831 ( .A1(n433), .A2(\REGISTERS[49][26] ), .B1(n76), .B2(
        \REGISTERS[51][26] ), .C1(n73), .C2(\REGISTERS[50][26] ), .ZN(n5190)
         );
  AOI222_X1 U2832 ( .A1(n14), .A2(\REGISTERS[82][26] ), .B1(n8), .B2(
        \REGISTERS[84][26] ), .C1(n4), .C2(\REGISTERS[83][26] ), .ZN(n5199) );
  AOI222_X1 U2833 ( .A1(n1145), .A2(\REGISTERS[49][26] ), .B1(n1140), .B2(
        \REGISTERS[51][26] ), .C1(n1137), .C2(\REGISTERS[50][26] ), .ZN(n3747)
         );
  AOI222_X1 U2834 ( .A1(n727), .A2(\REGISTERS[82][26] ), .B1(n722), .B2(
        \REGISTERS[84][26] ), .C1(n719), .C2(\REGISTERS[83][26] ), .ZN(n3756)
         );
  AOI222_X1 U2835 ( .A1(n433), .A2(\REGISTERS[49][27] ), .B1(n76), .B2(
        \REGISTERS[51][27] ), .C1(n73), .C2(\REGISTERS[50][27] ), .ZN(n5149)
         );
  AOI222_X1 U2836 ( .A1(n14), .A2(\REGISTERS[82][27] ), .B1(n8), .B2(
        \REGISTERS[84][27] ), .C1(n4), .C2(\REGISTERS[83][27] ), .ZN(n5158) );
  AOI222_X1 U2837 ( .A1(n1145), .A2(\REGISTERS[49][27] ), .B1(n1140), .B2(
        \REGISTERS[51][27] ), .C1(n1137), .C2(\REGISTERS[50][27] ), .ZN(n3706)
         );
  AOI222_X1 U2838 ( .A1(n727), .A2(\REGISTERS[82][27] ), .B1(n722), .B2(
        \REGISTERS[84][27] ), .C1(n719), .C2(\REGISTERS[83][27] ), .ZN(n3715)
         );
  AOI222_X1 U2839 ( .A1(n433), .A2(\REGISTERS[49][28] ), .B1(n76), .B2(
        \REGISTERS[51][28] ), .C1(n73), .C2(\REGISTERS[50][28] ), .ZN(n5108)
         );
  AOI222_X1 U2840 ( .A1(n14), .A2(\REGISTERS[82][28] ), .B1(n8), .B2(
        \REGISTERS[84][28] ), .C1(n4), .C2(\REGISTERS[83][28] ), .ZN(n5117) );
  AOI222_X1 U2841 ( .A1(n1145), .A2(\REGISTERS[49][28] ), .B1(n1140), .B2(
        \REGISTERS[51][28] ), .C1(n1137), .C2(\REGISTERS[50][28] ), .ZN(n3665)
         );
  AOI222_X1 U2842 ( .A1(n727), .A2(\REGISTERS[82][28] ), .B1(n722), .B2(
        \REGISTERS[84][28] ), .C1(n719), .C2(\REGISTERS[83][28] ), .ZN(n3674)
         );
  AOI222_X1 U2843 ( .A1(n433), .A2(\REGISTERS[49][29] ), .B1(n76), .B2(
        \REGISTERS[51][29] ), .C1(n73), .C2(\REGISTERS[50][29] ), .ZN(n5067)
         );
  AOI222_X1 U2844 ( .A1(n14), .A2(\REGISTERS[82][29] ), .B1(n8), .B2(
        \REGISTERS[84][29] ), .C1(n4), .C2(\REGISTERS[83][29] ), .ZN(n5076) );
  AOI222_X1 U2845 ( .A1(n1145), .A2(\REGISTERS[49][29] ), .B1(n1140), .B2(
        \REGISTERS[51][29] ), .C1(n1137), .C2(\REGISTERS[50][29] ), .ZN(n3624)
         );
  AOI222_X1 U2846 ( .A1(n727), .A2(\REGISTERS[82][29] ), .B1(n722), .B2(
        \REGISTERS[84][29] ), .C1(n719), .C2(\REGISTERS[83][29] ), .ZN(n3633)
         );
  AOI222_X1 U2847 ( .A1(n433), .A2(\REGISTERS[49][30] ), .B1(n76), .B2(
        \REGISTERS[51][30] ), .C1(n73), .C2(\REGISTERS[50][30] ), .ZN(n5026)
         );
  AOI222_X1 U2848 ( .A1(n14), .A2(\REGISTERS[82][30] ), .B1(n8), .B2(
        \REGISTERS[84][30] ), .C1(n4), .C2(\REGISTERS[83][30] ), .ZN(n5035) );
  AOI222_X1 U2849 ( .A1(n1145), .A2(\REGISTERS[49][30] ), .B1(n1140), .B2(
        \REGISTERS[51][30] ), .C1(n1137), .C2(\REGISTERS[50][30] ), .ZN(n3583)
         );
  AOI222_X1 U2850 ( .A1(n727), .A2(\REGISTERS[82][30] ), .B1(n722), .B2(
        \REGISTERS[84][30] ), .C1(n719), .C2(\REGISTERS[83][30] ), .ZN(n3592)
         );
  AOI222_X1 U2851 ( .A1(n433), .A2(\REGISTERS[49][31] ), .B1(n76), .B2(
        \REGISTERS[51][31] ), .C1(n73), .C2(\REGISTERS[50][31] ), .ZN(n4941)
         );
  AOI222_X1 U2852 ( .A1(n14), .A2(\REGISTERS[82][31] ), .B1(n8), .B2(
        \REGISTERS[84][31] ), .C1(n4), .C2(\REGISTERS[83][31] ), .ZN(n4972) );
  AOI222_X1 U2853 ( .A1(n1145), .A2(\REGISTERS[49][31] ), .B1(n1140), .B2(
        \REGISTERS[51][31] ), .C1(n1137), .C2(\REGISTERS[50][31] ), .ZN(n3498)
         );
  AOI222_X1 U2854 ( .A1(n727), .A2(\REGISTERS[82][31] ), .B1(n722), .B2(
        \REGISTERS[84][31] ), .C1(n719), .C2(\REGISTERS[83][31] ), .ZN(n3529)
         );
  NOR4_X1 U2855 ( .A1(n6292), .A2(n6293), .A3(n6294), .A4(n6295), .ZN(n6291)
         );
  OAI22_X1 U2856 ( .A1(n1871), .A2(n488), .B1(n1903), .B2(n485), .ZN(n6295) );
  OAI222_X1 U2857 ( .A1(n2159), .A2(n464), .B1(n2191), .B2(n461), .C1(n2127), 
        .C2(n458), .ZN(n6292) );
  OAI222_X1 U2858 ( .A1(n2063), .A2(n473), .B1(n2095), .B2(n470), .C1(n2031), 
        .C2(n467), .ZN(n6293) );
  NOR4_X1 U2859 ( .A1(n6305), .A2(n6306), .A3(n6307), .A4(n6308), .ZN(n6304)
         );
  OAI22_X1 U2860 ( .A1(n2223), .A2(n70), .B1(n2255), .B2(n67), .ZN(n6308) );
  OAI222_X1 U2861 ( .A1(n2511), .A2(n46), .B1(n2543), .B2(n43), .C1(n2479), 
        .C2(n40), .ZN(n6305) );
  OAI222_X1 U2862 ( .A1(n2415), .A2(n55), .B1(n2447), .B2(n52), .C1(n2383), 
        .C2(n49), .ZN(n6306) );
  NOR4_X1 U2863 ( .A1(n4849), .A2(n4850), .A3(n4851), .A4(n4852), .ZN(n4848)
         );
  OAI22_X1 U2864 ( .A1(n1871), .A2(n1296), .B1(n1903), .B2(n1197), .ZN(n4852)
         );
  OAI222_X1 U2865 ( .A1(n2159), .A2(n1176), .B1(n2191), .B2(n1173), .C1(n2127), 
        .C2(n1170), .ZN(n4849) );
  OAI222_X1 U2866 ( .A1(n2063), .A2(n1185), .B1(n2095), .B2(n1182), .C1(n2031), 
        .C2(n1179), .ZN(n4850) );
  NOR4_X1 U2867 ( .A1(n4862), .A2(n4863), .A3(n4864), .A4(n4865), .ZN(n4861)
         );
  OAI22_X1 U2868 ( .A1(n2223), .A2(n782), .B1(n2255), .B2(n779), .ZN(n4865) );
  OAI222_X1 U2869 ( .A1(n2511), .A2(n758), .B1(n2543), .B2(n755), .C1(n2479), 
        .C2(n752), .ZN(n4862) );
  OAI222_X1 U2870 ( .A1(n2415), .A2(n767), .B1(n2447), .B2(n764), .C1(n2383), 
        .C2(n761), .ZN(n4863) );
  NOR4_X1 U2871 ( .A1(n6219), .A2(n6220), .A3(n6221), .A4(n6222), .ZN(n6218)
         );
  OAI22_X1 U2872 ( .A1(n1870), .A2(n488), .B1(n1902), .B2(n485), .ZN(n6222) );
  OAI222_X1 U2873 ( .A1(n2158), .A2(n464), .B1(n2190), .B2(n461), .C1(n2126), 
        .C2(n458), .ZN(n6219) );
  OAI222_X1 U2874 ( .A1(n2062), .A2(n473), .B1(n2094), .B2(n470), .C1(n2030), 
        .C2(n467), .ZN(n6220) );
  NOR4_X1 U2875 ( .A1(n6228), .A2(n6229), .A3(n6230), .A4(n6231), .ZN(n6227)
         );
  OAI22_X1 U2876 ( .A1(n2222), .A2(n70), .B1(n2254), .B2(n67), .ZN(n6231) );
  OAI222_X1 U2877 ( .A1(n2510), .A2(n46), .B1(n2542), .B2(n43), .C1(n2478), 
        .C2(n40), .ZN(n6228) );
  OAI222_X1 U2878 ( .A1(n2414), .A2(n55), .B1(n2446), .B2(n52), .C1(n2382), 
        .C2(n49), .ZN(n6229) );
  NOR4_X1 U2879 ( .A1(n4776), .A2(n4777), .A3(n4778), .A4(n4779), .ZN(n4775)
         );
  OAI22_X1 U2880 ( .A1(n1870), .A2(n1296), .B1(n1902), .B2(n1197), .ZN(n4779)
         );
  OAI222_X1 U2881 ( .A1(n2158), .A2(n1176), .B1(n2190), .B2(n1173), .C1(n2126), 
        .C2(n1170), .ZN(n4776) );
  OAI222_X1 U2882 ( .A1(n2062), .A2(n1185), .B1(n2094), .B2(n1182), .C1(n2030), 
        .C2(n1179), .ZN(n4777) );
  NOR4_X1 U2883 ( .A1(n4785), .A2(n4786), .A3(n4787), .A4(n4788), .ZN(n4784)
         );
  OAI22_X1 U2884 ( .A1(n2222), .A2(n782), .B1(n2254), .B2(n779), .ZN(n4788) );
  OAI222_X1 U2885 ( .A1(n2510), .A2(n758), .B1(n2542), .B2(n755), .C1(n2478), 
        .C2(n752), .ZN(n4785) );
  OAI222_X1 U2886 ( .A1(n2414), .A2(n767), .B1(n2446), .B2(n764), .C1(n2382), 
        .C2(n761), .ZN(n4786) );
  NOR4_X1 U2887 ( .A1(n6178), .A2(n6179), .A3(n6180), .A4(n6181), .ZN(n6177)
         );
  OAI22_X1 U2888 ( .A1(n1869), .A2(n488), .B1(n1901), .B2(n485), .ZN(n6181) );
  OAI222_X1 U2889 ( .A1(n2157), .A2(n464), .B1(n2189), .B2(n461), .C1(n2125), 
        .C2(n458), .ZN(n6178) );
  OAI222_X1 U2890 ( .A1(n2061), .A2(n473), .B1(n2093), .B2(n470), .C1(n2029), 
        .C2(n467), .ZN(n6179) );
  NOR4_X1 U2891 ( .A1(n6187), .A2(n6188), .A3(n6189), .A4(n6190), .ZN(n6186)
         );
  OAI22_X1 U2892 ( .A1(n2221), .A2(n70), .B1(n2253), .B2(n67), .ZN(n6190) );
  OAI222_X1 U2893 ( .A1(n2509), .A2(n46), .B1(n2541), .B2(n43), .C1(n2477), 
        .C2(n40), .ZN(n6187) );
  OAI222_X1 U2894 ( .A1(n2413), .A2(n55), .B1(n2445), .B2(n52), .C1(n2381), 
        .C2(n49), .ZN(n6188) );
  NOR4_X1 U2895 ( .A1(n4735), .A2(n4736), .A3(n4737), .A4(n4738), .ZN(n4734)
         );
  OAI22_X1 U2896 ( .A1(n1869), .A2(n1296), .B1(n1901), .B2(n1197), .ZN(n4738)
         );
  OAI222_X1 U2897 ( .A1(n2157), .A2(n1176), .B1(n2189), .B2(n1173), .C1(n2125), 
        .C2(n1170), .ZN(n4735) );
  OAI222_X1 U2898 ( .A1(n2061), .A2(n1185), .B1(n2093), .B2(n1182), .C1(n2029), 
        .C2(n1179), .ZN(n4736) );
  NOR4_X1 U2899 ( .A1(n4744), .A2(n4745), .A3(n4746), .A4(n4747), .ZN(n4743)
         );
  OAI22_X1 U2900 ( .A1(n2221), .A2(n782), .B1(n2253), .B2(n779), .ZN(n4747) );
  OAI222_X1 U2901 ( .A1(n2509), .A2(n758), .B1(n2541), .B2(n755), .C1(n2477), 
        .C2(n752), .ZN(n4744) );
  OAI222_X1 U2902 ( .A1(n2413), .A2(n767), .B1(n2445), .B2(n764), .C1(n2381), 
        .C2(n761), .ZN(n4745) );
  NOR4_X1 U2903 ( .A1(n6137), .A2(n6138), .A3(n6139), .A4(n6140), .ZN(n6136)
         );
  OAI22_X1 U2904 ( .A1(n1868), .A2(n488), .B1(n1900), .B2(n485), .ZN(n6140) );
  OAI222_X1 U2905 ( .A1(n2156), .A2(n464), .B1(n2188), .B2(n461), .C1(n2124), 
        .C2(n458), .ZN(n6137) );
  OAI222_X1 U2906 ( .A1(n2060), .A2(n473), .B1(n2092), .B2(n470), .C1(n2028), 
        .C2(n467), .ZN(n6138) );
  NOR4_X1 U2907 ( .A1(n6146), .A2(n6147), .A3(n6148), .A4(n6149), .ZN(n6145)
         );
  OAI22_X1 U2908 ( .A1(n2220), .A2(n70), .B1(n2252), .B2(n67), .ZN(n6149) );
  OAI222_X1 U2909 ( .A1(n2508), .A2(n46), .B1(n2540), .B2(n43), .C1(n2476), 
        .C2(n40), .ZN(n6146) );
  OAI222_X1 U2910 ( .A1(n2412), .A2(n55), .B1(n2444), .B2(n52), .C1(n2380), 
        .C2(n49), .ZN(n6147) );
  NOR4_X1 U2911 ( .A1(n4694), .A2(n4695), .A3(n4696), .A4(n4697), .ZN(n4693)
         );
  OAI22_X1 U2912 ( .A1(n1868), .A2(n1296), .B1(n1900), .B2(n1197), .ZN(n4697)
         );
  OAI222_X1 U2913 ( .A1(n2156), .A2(n1176), .B1(n2188), .B2(n1173), .C1(n2124), 
        .C2(n1170), .ZN(n4694) );
  OAI222_X1 U2914 ( .A1(n2060), .A2(n1185), .B1(n2092), .B2(n1182), .C1(n2028), 
        .C2(n1179), .ZN(n4695) );
  NOR4_X1 U2915 ( .A1(n4703), .A2(n4704), .A3(n4705), .A4(n4706), .ZN(n4702)
         );
  OAI22_X1 U2916 ( .A1(n2220), .A2(n782), .B1(n2252), .B2(n779), .ZN(n4706) );
  OAI222_X1 U2917 ( .A1(n2508), .A2(n758), .B1(n2540), .B2(n755), .C1(n2476), 
        .C2(n752), .ZN(n4703) );
  OAI222_X1 U2918 ( .A1(n2412), .A2(n767), .B1(n2444), .B2(n764), .C1(n2380), 
        .C2(n761), .ZN(n4704) );
  NOR4_X1 U2919 ( .A1(n6096), .A2(n6097), .A3(n6098), .A4(n6099), .ZN(n6095)
         );
  OAI22_X1 U2920 ( .A1(n1867), .A2(n488), .B1(n1899), .B2(n485), .ZN(n6099) );
  OAI222_X1 U2921 ( .A1(n2155), .A2(n464), .B1(n2187), .B2(n461), .C1(n2123), 
        .C2(n458), .ZN(n6096) );
  OAI222_X1 U2922 ( .A1(n2059), .A2(n473), .B1(n2091), .B2(n470), .C1(n2027), 
        .C2(n467), .ZN(n6097) );
  NOR4_X1 U2923 ( .A1(n6105), .A2(n6106), .A3(n6107), .A4(n6108), .ZN(n6104)
         );
  OAI22_X1 U2924 ( .A1(n2219), .A2(n70), .B1(n2251), .B2(n67), .ZN(n6108) );
  OAI222_X1 U2925 ( .A1(n2507), .A2(n46), .B1(n2539), .B2(n43), .C1(n2475), 
        .C2(n40), .ZN(n6105) );
  OAI222_X1 U2926 ( .A1(n2411), .A2(n55), .B1(n2443), .B2(n52), .C1(n2379), 
        .C2(n49), .ZN(n6106) );
  NOR4_X1 U2927 ( .A1(n4653), .A2(n4654), .A3(n4655), .A4(n4656), .ZN(n4652)
         );
  OAI22_X1 U2928 ( .A1(n1867), .A2(n1296), .B1(n1899), .B2(n1197), .ZN(n4656)
         );
  OAI222_X1 U2929 ( .A1(n2155), .A2(n1176), .B1(n2187), .B2(n1173), .C1(n2123), 
        .C2(n1170), .ZN(n4653) );
  OAI222_X1 U2930 ( .A1(n2059), .A2(n1185), .B1(n2091), .B2(n1182), .C1(n2027), 
        .C2(n1179), .ZN(n4654) );
  NOR4_X1 U2931 ( .A1(n4662), .A2(n4663), .A3(n4664), .A4(n4665), .ZN(n4661)
         );
  OAI22_X1 U2932 ( .A1(n2219), .A2(n782), .B1(n2251), .B2(n779), .ZN(n4665) );
  OAI222_X1 U2933 ( .A1(n2507), .A2(n758), .B1(n2539), .B2(n755), .C1(n2475), 
        .C2(n752), .ZN(n4662) );
  OAI222_X1 U2934 ( .A1(n2411), .A2(n767), .B1(n2443), .B2(n764), .C1(n2379), 
        .C2(n761), .ZN(n4663) );
  NOR4_X1 U2935 ( .A1(n6055), .A2(n6056), .A3(n6057), .A4(n6058), .ZN(n6054)
         );
  OAI22_X1 U2936 ( .A1(n1866), .A2(n488), .B1(n1898), .B2(n485), .ZN(n6058) );
  OAI222_X1 U2937 ( .A1(n2154), .A2(n464), .B1(n2186), .B2(n461), .C1(n2122), 
        .C2(n458), .ZN(n6055) );
  OAI222_X1 U2938 ( .A1(n2058), .A2(n473), .B1(n2090), .B2(n470), .C1(n2026), 
        .C2(n467), .ZN(n6056) );
  NOR4_X1 U2939 ( .A1(n6064), .A2(n6065), .A3(n6066), .A4(n6067), .ZN(n6063)
         );
  OAI22_X1 U2940 ( .A1(n2218), .A2(n70), .B1(n2250), .B2(n67), .ZN(n6067) );
  OAI222_X1 U2941 ( .A1(n2506), .A2(n46), .B1(n2538), .B2(n43), .C1(n2474), 
        .C2(n40), .ZN(n6064) );
  OAI222_X1 U2942 ( .A1(n2410), .A2(n55), .B1(n2442), .B2(n52), .C1(n2378), 
        .C2(n49), .ZN(n6065) );
  NOR4_X1 U2943 ( .A1(n4612), .A2(n4613), .A3(n4614), .A4(n4615), .ZN(n4611)
         );
  OAI22_X1 U2944 ( .A1(n1866), .A2(n1296), .B1(n1898), .B2(n1197), .ZN(n4615)
         );
  OAI222_X1 U2945 ( .A1(n2154), .A2(n1176), .B1(n2186), .B2(n1173), .C1(n2122), 
        .C2(n1170), .ZN(n4612) );
  OAI222_X1 U2946 ( .A1(n2058), .A2(n1185), .B1(n2090), .B2(n1182), .C1(n2026), 
        .C2(n1179), .ZN(n4613) );
  NOR4_X1 U2947 ( .A1(n4621), .A2(n4622), .A3(n4623), .A4(n4624), .ZN(n4620)
         );
  OAI22_X1 U2948 ( .A1(n2218), .A2(n782), .B1(n2250), .B2(n779), .ZN(n4624) );
  OAI222_X1 U2949 ( .A1(n2506), .A2(n758), .B1(n2538), .B2(n755), .C1(n2474), 
        .C2(n752), .ZN(n4621) );
  OAI222_X1 U2950 ( .A1(n2410), .A2(n767), .B1(n2442), .B2(n764), .C1(n2378), 
        .C2(n761), .ZN(n4622) );
  NOR4_X1 U2951 ( .A1(n6014), .A2(n6015), .A3(n6016), .A4(n6017), .ZN(n6013)
         );
  OAI22_X1 U2952 ( .A1(n1865), .A2(n488), .B1(n1897), .B2(n485), .ZN(n6017) );
  OAI222_X1 U2953 ( .A1(n2153), .A2(n464), .B1(n2185), .B2(n461), .C1(n2121), 
        .C2(n458), .ZN(n6014) );
  OAI222_X1 U2954 ( .A1(n2057), .A2(n473), .B1(n2089), .B2(n470), .C1(n2025), 
        .C2(n467), .ZN(n6015) );
  NOR4_X1 U2955 ( .A1(n6023), .A2(n6024), .A3(n6025), .A4(n6026), .ZN(n6022)
         );
  OAI22_X1 U2956 ( .A1(n2217), .A2(n70), .B1(n2249), .B2(n67), .ZN(n6026) );
  OAI222_X1 U2957 ( .A1(n2505), .A2(n46), .B1(n2537), .B2(n43), .C1(n2473), 
        .C2(n40), .ZN(n6023) );
  OAI222_X1 U2958 ( .A1(n2409), .A2(n55), .B1(n2441), .B2(n52), .C1(n2377), 
        .C2(n49), .ZN(n6024) );
  NOR4_X1 U2959 ( .A1(n4571), .A2(n4572), .A3(n4573), .A4(n4574), .ZN(n4570)
         );
  OAI22_X1 U2960 ( .A1(n1865), .A2(n1296), .B1(n1897), .B2(n1197), .ZN(n4574)
         );
  OAI222_X1 U2961 ( .A1(n2153), .A2(n1176), .B1(n2185), .B2(n1173), .C1(n2121), 
        .C2(n1170), .ZN(n4571) );
  OAI222_X1 U2962 ( .A1(n2057), .A2(n1185), .B1(n2089), .B2(n1182), .C1(n2025), 
        .C2(n1179), .ZN(n4572) );
  NOR4_X1 U2963 ( .A1(n4580), .A2(n4581), .A3(n4582), .A4(n4583), .ZN(n4579)
         );
  OAI22_X1 U2964 ( .A1(n2217), .A2(n782), .B1(n2249), .B2(n779), .ZN(n4583) );
  OAI222_X1 U2965 ( .A1(n2505), .A2(n758), .B1(n2537), .B2(n755), .C1(n2473), 
        .C2(n752), .ZN(n4580) );
  OAI222_X1 U2966 ( .A1(n2409), .A2(n767), .B1(n2441), .B2(n764), .C1(n2377), 
        .C2(n761), .ZN(n4581) );
  NOR4_X1 U2967 ( .A1(n5973), .A2(n5974), .A3(n5975), .A4(n5976), .ZN(n5972)
         );
  OAI22_X1 U2968 ( .A1(n1864), .A2(n488), .B1(n1896), .B2(n485), .ZN(n5976) );
  OAI222_X1 U2969 ( .A1(n2152), .A2(n464), .B1(n2184), .B2(n461), .C1(n2120), 
        .C2(n458), .ZN(n5973) );
  OAI222_X1 U2970 ( .A1(n2056), .A2(n473), .B1(n2088), .B2(n470), .C1(n2024), 
        .C2(n467), .ZN(n5974) );
  NOR4_X1 U2971 ( .A1(n5982), .A2(n5983), .A3(n5984), .A4(n5985), .ZN(n5981)
         );
  OAI22_X1 U2972 ( .A1(n2216), .A2(n70), .B1(n2248), .B2(n67), .ZN(n5985) );
  OAI222_X1 U2973 ( .A1(n2504), .A2(n46), .B1(n2536), .B2(n43), .C1(n2472), 
        .C2(n40), .ZN(n5982) );
  OAI222_X1 U2974 ( .A1(n2408), .A2(n55), .B1(n2440), .B2(n52), .C1(n2376), 
        .C2(n49), .ZN(n5983) );
  NOR4_X1 U2975 ( .A1(n4530), .A2(n4531), .A3(n4532), .A4(n4533), .ZN(n4529)
         );
  OAI22_X1 U2976 ( .A1(n1864), .A2(n1296), .B1(n1896), .B2(n1197), .ZN(n4533)
         );
  OAI222_X1 U2977 ( .A1(n2152), .A2(n1176), .B1(n2184), .B2(n1173), .C1(n2120), 
        .C2(n1170), .ZN(n4530) );
  OAI222_X1 U2978 ( .A1(n2056), .A2(n1185), .B1(n2088), .B2(n1182), .C1(n2024), 
        .C2(n1179), .ZN(n4531) );
  NOR4_X1 U2979 ( .A1(n4539), .A2(n4540), .A3(n4541), .A4(n4542), .ZN(n4538)
         );
  OAI22_X1 U2980 ( .A1(n2216), .A2(n782), .B1(n2248), .B2(n779), .ZN(n4542) );
  OAI222_X1 U2981 ( .A1(n2504), .A2(n758), .B1(n2536), .B2(n755), .C1(n2472), 
        .C2(n752), .ZN(n4539) );
  OAI222_X1 U2982 ( .A1(n2408), .A2(n767), .B1(n2440), .B2(n764), .C1(n2376), 
        .C2(n761), .ZN(n4540) );
  NOR4_X1 U2983 ( .A1(n5932), .A2(n5933), .A3(n5934), .A4(n5935), .ZN(n5931)
         );
  OAI22_X1 U2984 ( .A1(n1863), .A2(n488), .B1(n1895), .B2(n485), .ZN(n5935) );
  OAI222_X1 U2985 ( .A1(n2151), .A2(n464), .B1(n2183), .B2(n461), .C1(n2119), 
        .C2(n458), .ZN(n5932) );
  OAI222_X1 U2986 ( .A1(n2055), .A2(n473), .B1(n2087), .B2(n470), .C1(n2023), 
        .C2(n467), .ZN(n5933) );
  NOR4_X1 U2987 ( .A1(n5941), .A2(n5942), .A3(n5943), .A4(n5944), .ZN(n5940)
         );
  OAI22_X1 U2988 ( .A1(n2215), .A2(n70), .B1(n2247), .B2(n67), .ZN(n5944) );
  OAI222_X1 U2989 ( .A1(n2503), .A2(n46), .B1(n2535), .B2(n43), .C1(n2471), 
        .C2(n40), .ZN(n5941) );
  OAI222_X1 U2990 ( .A1(n2407), .A2(n55), .B1(n2439), .B2(n52), .C1(n2375), 
        .C2(n49), .ZN(n5942) );
  NOR4_X1 U2991 ( .A1(n4489), .A2(n4490), .A3(n4491), .A4(n4492), .ZN(n4488)
         );
  OAI22_X1 U2992 ( .A1(n1863), .A2(n1296), .B1(n1895), .B2(n1197), .ZN(n4492)
         );
  OAI222_X1 U2993 ( .A1(n2151), .A2(n1176), .B1(n2183), .B2(n1173), .C1(n2119), 
        .C2(n1170), .ZN(n4489) );
  OAI222_X1 U2994 ( .A1(n2055), .A2(n1185), .B1(n2087), .B2(n1182), .C1(n2023), 
        .C2(n1179), .ZN(n4490) );
  NOR4_X1 U2995 ( .A1(n4498), .A2(n4499), .A3(n4500), .A4(n4501), .ZN(n4497)
         );
  OAI22_X1 U2996 ( .A1(n2215), .A2(n782), .B1(n2247), .B2(n779), .ZN(n4501) );
  OAI222_X1 U2997 ( .A1(n2503), .A2(n758), .B1(n2535), .B2(n755), .C1(n2471), 
        .C2(n752), .ZN(n4498) );
  OAI222_X1 U2998 ( .A1(n2407), .A2(n767), .B1(n2439), .B2(n764), .C1(n2375), 
        .C2(n761), .ZN(n4499) );
  NOR4_X1 U2999 ( .A1(n5891), .A2(n5892), .A3(n5893), .A4(n5894), .ZN(n5890)
         );
  OAI22_X1 U3000 ( .A1(n1862), .A2(n488), .B1(n1894), .B2(n485), .ZN(n5894) );
  OAI222_X1 U3001 ( .A1(n2150), .A2(n464), .B1(n2182), .B2(n461), .C1(n2118), 
        .C2(n458), .ZN(n5891) );
  OAI222_X1 U3002 ( .A1(n2054), .A2(n473), .B1(n2086), .B2(n470), .C1(n2022), 
        .C2(n467), .ZN(n5892) );
  NOR4_X1 U3003 ( .A1(n5900), .A2(n5901), .A3(n5902), .A4(n5903), .ZN(n5899)
         );
  OAI22_X1 U3004 ( .A1(n2214), .A2(n70), .B1(n2246), .B2(n67), .ZN(n5903) );
  OAI222_X1 U3005 ( .A1(n2502), .A2(n46), .B1(n2534), .B2(n43), .C1(n2470), 
        .C2(n40), .ZN(n5900) );
  OAI222_X1 U3006 ( .A1(n2406), .A2(n55), .B1(n2438), .B2(n52), .C1(n2374), 
        .C2(n49), .ZN(n5901) );
  NOR4_X1 U3007 ( .A1(n4448), .A2(n4449), .A3(n4450), .A4(n4451), .ZN(n4447)
         );
  OAI22_X1 U3008 ( .A1(n1862), .A2(n1296), .B1(n1894), .B2(n1197), .ZN(n4451)
         );
  OAI222_X1 U3009 ( .A1(n2150), .A2(n1176), .B1(n2182), .B2(n1173), .C1(n2118), 
        .C2(n1170), .ZN(n4448) );
  OAI222_X1 U3010 ( .A1(n2054), .A2(n1185), .B1(n2086), .B2(n1182), .C1(n2022), 
        .C2(n1179), .ZN(n4449) );
  NOR4_X1 U3011 ( .A1(n4457), .A2(n4458), .A3(n4459), .A4(n4460), .ZN(n4456)
         );
  OAI22_X1 U3012 ( .A1(n2214), .A2(n782), .B1(n2246), .B2(n779), .ZN(n4460) );
  OAI222_X1 U3013 ( .A1(n2502), .A2(n758), .B1(n2534), .B2(n755), .C1(n2470), 
        .C2(n752), .ZN(n4457) );
  OAI222_X1 U3014 ( .A1(n2406), .A2(n767), .B1(n2438), .B2(n764), .C1(n2374), 
        .C2(n761), .ZN(n4458) );
  NOR4_X1 U3015 ( .A1(n5850), .A2(n5851), .A3(n5852), .A4(n5853), .ZN(n5849)
         );
  OAI22_X1 U3016 ( .A1(n1861), .A2(n488), .B1(n1893), .B2(n485), .ZN(n5853) );
  OAI222_X1 U3017 ( .A1(n2149), .A2(n464), .B1(n2181), .B2(n461), .C1(n2117), 
        .C2(n458), .ZN(n5850) );
  OAI222_X1 U3018 ( .A1(n2053), .A2(n473), .B1(n2085), .B2(n470), .C1(n2021), 
        .C2(n467), .ZN(n5851) );
  NOR4_X1 U3019 ( .A1(n5859), .A2(n5860), .A3(n5861), .A4(n5862), .ZN(n5858)
         );
  OAI22_X1 U3020 ( .A1(n2213), .A2(n70), .B1(n2245), .B2(n67), .ZN(n5862) );
  OAI222_X1 U3021 ( .A1(n2501), .A2(n46), .B1(n2533), .B2(n43), .C1(n2469), 
        .C2(n40), .ZN(n5859) );
  OAI222_X1 U3022 ( .A1(n2405), .A2(n55), .B1(n2437), .B2(n52), .C1(n2373), 
        .C2(n49), .ZN(n5860) );
  NOR4_X1 U3023 ( .A1(n4407), .A2(n4408), .A3(n4409), .A4(n4410), .ZN(n4406)
         );
  OAI22_X1 U3024 ( .A1(n1861), .A2(n1296), .B1(n1893), .B2(n1197), .ZN(n4410)
         );
  OAI222_X1 U3025 ( .A1(n2149), .A2(n1176), .B1(n2181), .B2(n1173), .C1(n2117), 
        .C2(n1170), .ZN(n4407) );
  OAI222_X1 U3026 ( .A1(n2053), .A2(n1185), .B1(n2085), .B2(n1182), .C1(n2021), 
        .C2(n1179), .ZN(n4408) );
  NOR4_X1 U3027 ( .A1(n4416), .A2(n4417), .A3(n4418), .A4(n4419), .ZN(n4415)
         );
  OAI22_X1 U3028 ( .A1(n2213), .A2(n782), .B1(n2245), .B2(n779), .ZN(n4419) );
  OAI222_X1 U3029 ( .A1(n2501), .A2(n758), .B1(n2533), .B2(n755), .C1(n2469), 
        .C2(n752), .ZN(n4416) );
  OAI222_X1 U3030 ( .A1(n2405), .A2(n767), .B1(n2437), .B2(n764), .C1(n2373), 
        .C2(n761), .ZN(n4417) );
  NOR4_X1 U3031 ( .A1(n5809), .A2(n5810), .A3(n5811), .A4(n5812), .ZN(n5808)
         );
  OAI22_X1 U3032 ( .A1(n1860), .A2(n488), .B1(n1892), .B2(n485), .ZN(n5812) );
  OAI222_X1 U3033 ( .A1(n2148), .A2(n464), .B1(n2180), .B2(n461), .C1(n2116), 
        .C2(n458), .ZN(n5809) );
  OAI222_X1 U3034 ( .A1(n2052), .A2(n473), .B1(n2084), .B2(n470), .C1(n2020), 
        .C2(n467), .ZN(n5810) );
  NOR4_X1 U3035 ( .A1(n5818), .A2(n5819), .A3(n5820), .A4(n5821), .ZN(n5817)
         );
  OAI22_X1 U3036 ( .A1(n2212), .A2(n70), .B1(n2244), .B2(n67), .ZN(n5821) );
  OAI222_X1 U3037 ( .A1(n2500), .A2(n46), .B1(n2532), .B2(n43), .C1(n2468), 
        .C2(n40), .ZN(n5818) );
  OAI222_X1 U3038 ( .A1(n2404), .A2(n55), .B1(n2436), .B2(n52), .C1(n2372), 
        .C2(n49), .ZN(n5819) );
  NOR4_X1 U3039 ( .A1(n4366), .A2(n4367), .A3(n4368), .A4(n4369), .ZN(n4365)
         );
  OAI22_X1 U3040 ( .A1(n1860), .A2(n1296), .B1(n1892), .B2(n1197), .ZN(n4369)
         );
  OAI222_X1 U3041 ( .A1(n2148), .A2(n1176), .B1(n2180), .B2(n1173), .C1(n2116), 
        .C2(n1170), .ZN(n4366) );
  OAI222_X1 U3042 ( .A1(n2052), .A2(n1185), .B1(n2084), .B2(n1182), .C1(n2020), 
        .C2(n1179), .ZN(n4367) );
  NOR4_X1 U3043 ( .A1(n4375), .A2(n4376), .A3(n4377), .A4(n4378), .ZN(n4374)
         );
  OAI22_X1 U3044 ( .A1(n2212), .A2(n782), .B1(n2244), .B2(n779), .ZN(n4378) );
  OAI222_X1 U3045 ( .A1(n2500), .A2(n758), .B1(n2532), .B2(n755), .C1(n2468), 
        .C2(n752), .ZN(n4375) );
  OAI222_X1 U3046 ( .A1(n2404), .A2(n767), .B1(n2436), .B2(n764), .C1(n2372), 
        .C2(n761), .ZN(n4376) );
  NOR4_X1 U3047 ( .A1(n5768), .A2(n5769), .A3(n5770), .A4(n5771), .ZN(n5767)
         );
  OAI22_X1 U3048 ( .A1(n1859), .A2(n489), .B1(n1891), .B2(n486), .ZN(n5771) );
  OAI222_X1 U3049 ( .A1(n2147), .A2(n465), .B1(n2179), .B2(n462), .C1(n2115), 
        .C2(n459), .ZN(n5768) );
  OAI222_X1 U3050 ( .A1(n2051), .A2(n474), .B1(n2083), .B2(n471), .C1(n2019), 
        .C2(n468), .ZN(n5769) );
  NOR4_X1 U3051 ( .A1(n5777), .A2(n5778), .A3(n5779), .A4(n5780), .ZN(n5776)
         );
  OAI22_X1 U3052 ( .A1(n2211), .A2(n71), .B1(n2243), .B2(n68), .ZN(n5780) );
  OAI222_X1 U3053 ( .A1(n2499), .A2(n47), .B1(n2531), .B2(n44), .C1(n2467), 
        .C2(n41), .ZN(n5777) );
  OAI222_X1 U3054 ( .A1(n2403), .A2(n56), .B1(n2435), .B2(n53), .C1(n2371), 
        .C2(n50), .ZN(n5778) );
  NOR4_X1 U3055 ( .A1(n4325), .A2(n4326), .A3(n4327), .A4(n4328), .ZN(n4324)
         );
  OAI22_X1 U3056 ( .A1(n1859), .A2(n1297), .B1(n1891), .B2(n1198), .ZN(n4328)
         );
  OAI222_X1 U3057 ( .A1(n2147), .A2(n1177), .B1(n2179), .B2(n1174), .C1(n2115), 
        .C2(n1171), .ZN(n4325) );
  OAI222_X1 U3058 ( .A1(n2051), .A2(n1186), .B1(n2083), .B2(n1183), .C1(n2019), 
        .C2(n1180), .ZN(n4326) );
  NOR4_X1 U3059 ( .A1(n4334), .A2(n4335), .A3(n4336), .A4(n4337), .ZN(n4333)
         );
  OAI22_X1 U3060 ( .A1(n2211), .A2(n783), .B1(n2243), .B2(n780), .ZN(n4337) );
  OAI222_X1 U3061 ( .A1(n2499), .A2(n759), .B1(n2531), .B2(n756), .C1(n2467), 
        .C2(n753), .ZN(n4334) );
  OAI222_X1 U3062 ( .A1(n2403), .A2(n768), .B1(n2435), .B2(n765), .C1(n2371), 
        .C2(n762), .ZN(n4335) );
  NOR4_X1 U3063 ( .A1(n5727), .A2(n5728), .A3(n5729), .A4(n5730), .ZN(n5726)
         );
  OAI22_X1 U3064 ( .A1(n1858), .A2(n489), .B1(n1890), .B2(n486), .ZN(n5730) );
  OAI222_X1 U3065 ( .A1(n2146), .A2(n465), .B1(n2178), .B2(n462), .C1(n2114), 
        .C2(n459), .ZN(n5727) );
  OAI222_X1 U3066 ( .A1(n2050), .A2(n474), .B1(n2082), .B2(n471), .C1(n2018), 
        .C2(n468), .ZN(n5728) );
  NOR4_X1 U3067 ( .A1(n5736), .A2(n5737), .A3(n5738), .A4(n5739), .ZN(n5735)
         );
  OAI22_X1 U3068 ( .A1(n2210), .A2(n71), .B1(n2242), .B2(n68), .ZN(n5739) );
  OAI222_X1 U3069 ( .A1(n2498), .A2(n47), .B1(n2530), .B2(n44), .C1(n2466), 
        .C2(n41), .ZN(n5736) );
  OAI222_X1 U3070 ( .A1(n2402), .A2(n56), .B1(n2434), .B2(n53), .C1(n2370), 
        .C2(n50), .ZN(n5737) );
  NOR4_X1 U3071 ( .A1(n4284), .A2(n4285), .A3(n4286), .A4(n4287), .ZN(n4283)
         );
  OAI22_X1 U3072 ( .A1(n1858), .A2(n1297), .B1(n1890), .B2(n1198), .ZN(n4287)
         );
  OAI222_X1 U3073 ( .A1(n2146), .A2(n1177), .B1(n2178), .B2(n1174), .C1(n2114), 
        .C2(n1171), .ZN(n4284) );
  OAI222_X1 U3074 ( .A1(n2050), .A2(n1186), .B1(n2082), .B2(n1183), .C1(n2018), 
        .C2(n1180), .ZN(n4285) );
  NOR4_X1 U3075 ( .A1(n4293), .A2(n4294), .A3(n4295), .A4(n4296), .ZN(n4292)
         );
  OAI22_X1 U3076 ( .A1(n2210), .A2(n783), .B1(n2242), .B2(n780), .ZN(n4296) );
  OAI222_X1 U3077 ( .A1(n2498), .A2(n759), .B1(n2530), .B2(n756), .C1(n2466), 
        .C2(n753), .ZN(n4293) );
  OAI222_X1 U3078 ( .A1(n2402), .A2(n768), .B1(n2434), .B2(n765), .C1(n2370), 
        .C2(n762), .ZN(n4294) );
  NOR4_X1 U3079 ( .A1(n5686), .A2(n5687), .A3(n5688), .A4(n5689), .ZN(n5685)
         );
  OAI22_X1 U3080 ( .A1(n1857), .A2(n489), .B1(n1889), .B2(n486), .ZN(n5689) );
  OAI222_X1 U3081 ( .A1(n2145), .A2(n465), .B1(n2177), .B2(n462), .C1(n2113), 
        .C2(n459), .ZN(n5686) );
  OAI222_X1 U3082 ( .A1(n2049), .A2(n474), .B1(n2081), .B2(n471), .C1(n2017), 
        .C2(n468), .ZN(n5687) );
  NOR4_X1 U3083 ( .A1(n5695), .A2(n5696), .A3(n5697), .A4(n5698), .ZN(n5694)
         );
  OAI22_X1 U3084 ( .A1(n2209), .A2(n71), .B1(n2241), .B2(n68), .ZN(n5698) );
  OAI222_X1 U3085 ( .A1(n2497), .A2(n47), .B1(n2529), .B2(n44), .C1(n2465), 
        .C2(n41), .ZN(n5695) );
  OAI222_X1 U3086 ( .A1(n2401), .A2(n56), .B1(n2433), .B2(n53), .C1(n2369), 
        .C2(n50), .ZN(n5696) );
  NOR4_X1 U3087 ( .A1(n4243), .A2(n4244), .A3(n4245), .A4(n4246), .ZN(n4242)
         );
  OAI22_X1 U3088 ( .A1(n1857), .A2(n1297), .B1(n1889), .B2(n1198), .ZN(n4246)
         );
  OAI222_X1 U3089 ( .A1(n2145), .A2(n1177), .B1(n2177), .B2(n1174), .C1(n2113), 
        .C2(n1171), .ZN(n4243) );
  OAI222_X1 U3090 ( .A1(n2049), .A2(n1186), .B1(n2081), .B2(n1183), .C1(n2017), 
        .C2(n1180), .ZN(n4244) );
  NOR4_X1 U3091 ( .A1(n4252), .A2(n4253), .A3(n4254), .A4(n4255), .ZN(n4251)
         );
  OAI22_X1 U3092 ( .A1(n2209), .A2(n783), .B1(n2241), .B2(n780), .ZN(n4255) );
  OAI222_X1 U3093 ( .A1(n2497), .A2(n759), .B1(n2529), .B2(n756), .C1(n2465), 
        .C2(n753), .ZN(n4252) );
  OAI222_X1 U3094 ( .A1(n2401), .A2(n768), .B1(n2433), .B2(n765), .C1(n2369), 
        .C2(n762), .ZN(n4253) );
  NOR4_X1 U3095 ( .A1(n5645), .A2(n5646), .A3(n5647), .A4(n5648), .ZN(n5644)
         );
  OAI22_X1 U3096 ( .A1(n1856), .A2(n489), .B1(n1888), .B2(n486), .ZN(n5648) );
  OAI222_X1 U3097 ( .A1(n2144), .A2(n465), .B1(n2176), .B2(n462), .C1(n2112), 
        .C2(n459), .ZN(n5645) );
  OAI222_X1 U3098 ( .A1(n2048), .A2(n474), .B1(n2080), .B2(n471), .C1(n2016), 
        .C2(n468), .ZN(n5646) );
  NOR4_X1 U3099 ( .A1(n5654), .A2(n5655), .A3(n5656), .A4(n5657), .ZN(n5653)
         );
  OAI22_X1 U3100 ( .A1(n2208), .A2(n71), .B1(n2240), .B2(n68), .ZN(n5657) );
  OAI222_X1 U3101 ( .A1(n2496), .A2(n47), .B1(n2528), .B2(n44), .C1(n2464), 
        .C2(n41), .ZN(n5654) );
  OAI222_X1 U3102 ( .A1(n2400), .A2(n56), .B1(n2432), .B2(n53), .C1(n2368), 
        .C2(n50), .ZN(n5655) );
  NOR4_X1 U3103 ( .A1(n4202), .A2(n4203), .A3(n4204), .A4(n4205), .ZN(n4201)
         );
  OAI22_X1 U3104 ( .A1(n1856), .A2(n1297), .B1(n1888), .B2(n1198), .ZN(n4205)
         );
  OAI222_X1 U3105 ( .A1(n2144), .A2(n1177), .B1(n2176), .B2(n1174), .C1(n2112), 
        .C2(n1171), .ZN(n4202) );
  OAI222_X1 U3106 ( .A1(n2048), .A2(n1186), .B1(n2080), .B2(n1183), .C1(n2016), 
        .C2(n1180), .ZN(n4203) );
  NOR4_X1 U3107 ( .A1(n4211), .A2(n4212), .A3(n4213), .A4(n4214), .ZN(n4210)
         );
  OAI22_X1 U3108 ( .A1(n2208), .A2(n783), .B1(n2240), .B2(n780), .ZN(n4214) );
  OAI222_X1 U3109 ( .A1(n2496), .A2(n759), .B1(n2528), .B2(n756), .C1(n2464), 
        .C2(n753), .ZN(n4211) );
  OAI222_X1 U3110 ( .A1(n2400), .A2(n768), .B1(n2432), .B2(n765), .C1(n2368), 
        .C2(n762), .ZN(n4212) );
  NOR4_X1 U3111 ( .A1(n5604), .A2(n5605), .A3(n5606), .A4(n5607), .ZN(n5603)
         );
  OAI22_X1 U3112 ( .A1(n1855), .A2(n489), .B1(n1887), .B2(n486), .ZN(n5607) );
  OAI222_X1 U3113 ( .A1(n2143), .A2(n465), .B1(n2175), .B2(n462), .C1(n2111), 
        .C2(n459), .ZN(n5604) );
  OAI222_X1 U3114 ( .A1(n2047), .A2(n474), .B1(n2079), .B2(n471), .C1(n2015), 
        .C2(n468), .ZN(n5605) );
  NOR4_X1 U3115 ( .A1(n5613), .A2(n5614), .A3(n5615), .A4(n5616), .ZN(n5612)
         );
  OAI22_X1 U3116 ( .A1(n2207), .A2(n71), .B1(n2239), .B2(n68), .ZN(n5616) );
  OAI222_X1 U3117 ( .A1(n2495), .A2(n47), .B1(n2527), .B2(n44), .C1(n2463), 
        .C2(n41), .ZN(n5613) );
  OAI222_X1 U3118 ( .A1(n2399), .A2(n56), .B1(n2431), .B2(n53), .C1(n2367), 
        .C2(n50), .ZN(n5614) );
  NOR4_X1 U3119 ( .A1(n4161), .A2(n4162), .A3(n4163), .A4(n4164), .ZN(n4160)
         );
  OAI22_X1 U3120 ( .A1(n1855), .A2(n1297), .B1(n1887), .B2(n1198), .ZN(n4164)
         );
  OAI222_X1 U3121 ( .A1(n2143), .A2(n1177), .B1(n2175), .B2(n1174), .C1(n2111), 
        .C2(n1171), .ZN(n4161) );
  OAI222_X1 U3122 ( .A1(n2047), .A2(n1186), .B1(n2079), .B2(n1183), .C1(n2015), 
        .C2(n1180), .ZN(n4162) );
  NOR4_X1 U3123 ( .A1(n4170), .A2(n4171), .A3(n4172), .A4(n4173), .ZN(n4169)
         );
  OAI22_X1 U3124 ( .A1(n2207), .A2(n783), .B1(n2239), .B2(n780), .ZN(n4173) );
  OAI222_X1 U3125 ( .A1(n2495), .A2(n759), .B1(n2527), .B2(n756), .C1(n2463), 
        .C2(n753), .ZN(n4170) );
  OAI222_X1 U3126 ( .A1(n2399), .A2(n768), .B1(n2431), .B2(n765), .C1(n2367), 
        .C2(n762), .ZN(n4171) );
  NOR4_X1 U3127 ( .A1(n5563), .A2(n5564), .A3(n5565), .A4(n5566), .ZN(n5562)
         );
  OAI22_X1 U3128 ( .A1(n1854), .A2(n489), .B1(n1886), .B2(n486), .ZN(n5566) );
  OAI222_X1 U3129 ( .A1(n2142), .A2(n465), .B1(n2174), .B2(n462), .C1(n2110), 
        .C2(n459), .ZN(n5563) );
  OAI222_X1 U3130 ( .A1(n2046), .A2(n474), .B1(n2078), .B2(n471), .C1(n2014), 
        .C2(n468), .ZN(n5564) );
  NOR4_X1 U3131 ( .A1(n5572), .A2(n5573), .A3(n5574), .A4(n5575), .ZN(n5571)
         );
  OAI22_X1 U3132 ( .A1(n2206), .A2(n71), .B1(n2238), .B2(n68), .ZN(n5575) );
  OAI222_X1 U3133 ( .A1(n2494), .A2(n47), .B1(n2526), .B2(n44), .C1(n2462), 
        .C2(n41), .ZN(n5572) );
  OAI222_X1 U3134 ( .A1(n2398), .A2(n56), .B1(n2430), .B2(n53), .C1(n2366), 
        .C2(n50), .ZN(n5573) );
  NOR4_X1 U3135 ( .A1(n4120), .A2(n4121), .A3(n4122), .A4(n4123), .ZN(n4119)
         );
  OAI22_X1 U3136 ( .A1(n1854), .A2(n1297), .B1(n1886), .B2(n1198), .ZN(n4123)
         );
  OAI222_X1 U3137 ( .A1(n2142), .A2(n1177), .B1(n2174), .B2(n1174), .C1(n2110), 
        .C2(n1171), .ZN(n4120) );
  OAI222_X1 U3138 ( .A1(n2046), .A2(n1186), .B1(n2078), .B2(n1183), .C1(n2014), 
        .C2(n1180), .ZN(n4121) );
  NOR4_X1 U3139 ( .A1(n4129), .A2(n4130), .A3(n4131), .A4(n4132), .ZN(n4128)
         );
  OAI22_X1 U3140 ( .A1(n2206), .A2(n783), .B1(n2238), .B2(n780), .ZN(n4132) );
  OAI222_X1 U3141 ( .A1(n2494), .A2(n759), .B1(n2526), .B2(n756), .C1(n2462), 
        .C2(n753), .ZN(n4129) );
  OAI222_X1 U3142 ( .A1(n2398), .A2(n768), .B1(n2430), .B2(n765), .C1(n2366), 
        .C2(n762), .ZN(n4130) );
  NOR4_X1 U3143 ( .A1(n5522), .A2(n5523), .A3(n5524), .A4(n5525), .ZN(n5521)
         );
  OAI22_X1 U3144 ( .A1(n1853), .A2(n489), .B1(n1885), .B2(n486), .ZN(n5525) );
  OAI222_X1 U3145 ( .A1(n2141), .A2(n465), .B1(n2173), .B2(n462), .C1(n2109), 
        .C2(n459), .ZN(n5522) );
  OAI222_X1 U3146 ( .A1(n2045), .A2(n474), .B1(n2077), .B2(n471), .C1(n2013), 
        .C2(n468), .ZN(n5523) );
  NOR4_X1 U3147 ( .A1(n5531), .A2(n5532), .A3(n5533), .A4(n5534), .ZN(n5530)
         );
  OAI22_X1 U3148 ( .A1(n2205), .A2(n71), .B1(n2237), .B2(n68), .ZN(n5534) );
  OAI222_X1 U3149 ( .A1(n2493), .A2(n47), .B1(n2525), .B2(n44), .C1(n2461), 
        .C2(n41), .ZN(n5531) );
  OAI222_X1 U3150 ( .A1(n2397), .A2(n56), .B1(n2429), .B2(n53), .C1(n2365), 
        .C2(n50), .ZN(n5532) );
  NOR4_X1 U3151 ( .A1(n4079), .A2(n4080), .A3(n4081), .A4(n4082), .ZN(n4078)
         );
  OAI22_X1 U3152 ( .A1(n1853), .A2(n1297), .B1(n1885), .B2(n1198), .ZN(n4082)
         );
  OAI222_X1 U3153 ( .A1(n2141), .A2(n1177), .B1(n2173), .B2(n1174), .C1(n2109), 
        .C2(n1171), .ZN(n4079) );
  OAI222_X1 U3154 ( .A1(n2045), .A2(n1186), .B1(n2077), .B2(n1183), .C1(n2013), 
        .C2(n1180), .ZN(n4080) );
  NOR4_X1 U3155 ( .A1(n4088), .A2(n4089), .A3(n4090), .A4(n4091), .ZN(n4087)
         );
  OAI22_X1 U3156 ( .A1(n2205), .A2(n783), .B1(n2237), .B2(n780), .ZN(n4091) );
  OAI222_X1 U3157 ( .A1(n2493), .A2(n759), .B1(n2525), .B2(n756), .C1(n2461), 
        .C2(n753), .ZN(n4088) );
  OAI222_X1 U3158 ( .A1(n2397), .A2(n768), .B1(n2429), .B2(n765), .C1(n2365), 
        .C2(n762), .ZN(n4089) );
  NOR4_X1 U3159 ( .A1(n5481), .A2(n5482), .A3(n5483), .A4(n5484), .ZN(n5480)
         );
  OAI22_X1 U3160 ( .A1(n1852), .A2(n489), .B1(n1884), .B2(n486), .ZN(n5484) );
  OAI222_X1 U3161 ( .A1(n2140), .A2(n465), .B1(n2172), .B2(n462), .C1(n2108), 
        .C2(n459), .ZN(n5481) );
  OAI222_X1 U3162 ( .A1(n2044), .A2(n474), .B1(n2076), .B2(n471), .C1(n2012), 
        .C2(n468), .ZN(n5482) );
  NOR4_X1 U3163 ( .A1(n5490), .A2(n5491), .A3(n5492), .A4(n5493), .ZN(n5489)
         );
  OAI22_X1 U3164 ( .A1(n2204), .A2(n71), .B1(n2236), .B2(n68), .ZN(n5493) );
  OAI222_X1 U3165 ( .A1(n2492), .A2(n47), .B1(n2524), .B2(n44), .C1(n2460), 
        .C2(n41), .ZN(n5490) );
  OAI222_X1 U3166 ( .A1(n2396), .A2(n56), .B1(n2428), .B2(n53), .C1(n2364), 
        .C2(n50), .ZN(n5491) );
  NOR4_X1 U3167 ( .A1(n4038), .A2(n4039), .A3(n4040), .A4(n4041), .ZN(n4037)
         );
  OAI22_X1 U3168 ( .A1(n1852), .A2(n1297), .B1(n1884), .B2(n1198), .ZN(n4041)
         );
  OAI222_X1 U3169 ( .A1(n2140), .A2(n1177), .B1(n2172), .B2(n1174), .C1(n2108), 
        .C2(n1171), .ZN(n4038) );
  OAI222_X1 U3170 ( .A1(n2044), .A2(n1186), .B1(n2076), .B2(n1183), .C1(n2012), 
        .C2(n1180), .ZN(n4039) );
  NOR4_X1 U3171 ( .A1(n4047), .A2(n4048), .A3(n4049), .A4(n4050), .ZN(n4046)
         );
  OAI22_X1 U3172 ( .A1(n2204), .A2(n783), .B1(n2236), .B2(n780), .ZN(n4050) );
  OAI222_X1 U3173 ( .A1(n2492), .A2(n759), .B1(n2524), .B2(n756), .C1(n2460), 
        .C2(n753), .ZN(n4047) );
  OAI222_X1 U3174 ( .A1(n2396), .A2(n768), .B1(n2428), .B2(n765), .C1(n2364), 
        .C2(n762), .ZN(n4048) );
  NOR4_X1 U3175 ( .A1(n5440), .A2(n5441), .A3(n5442), .A4(n5443), .ZN(n5439)
         );
  OAI22_X1 U3176 ( .A1(n1851), .A2(n489), .B1(n1883), .B2(n486), .ZN(n5443) );
  OAI222_X1 U3177 ( .A1(n2139), .A2(n465), .B1(n2171), .B2(n462), .C1(n2107), 
        .C2(n459), .ZN(n5440) );
  OAI222_X1 U3178 ( .A1(n2043), .A2(n474), .B1(n2075), .B2(n471), .C1(n2011), 
        .C2(n468), .ZN(n5441) );
  NOR4_X1 U3179 ( .A1(n5449), .A2(n5450), .A3(n5451), .A4(n5452), .ZN(n5448)
         );
  OAI22_X1 U3180 ( .A1(n2203), .A2(n71), .B1(n2235), .B2(n68), .ZN(n5452) );
  OAI222_X1 U3181 ( .A1(n2491), .A2(n47), .B1(n2523), .B2(n44), .C1(n2459), 
        .C2(n41), .ZN(n5449) );
  OAI222_X1 U3182 ( .A1(n2395), .A2(n56), .B1(n2427), .B2(n53), .C1(n2363), 
        .C2(n50), .ZN(n5450) );
  NOR4_X1 U3183 ( .A1(n3997), .A2(n3998), .A3(n3999), .A4(n4000), .ZN(n3996)
         );
  OAI22_X1 U3184 ( .A1(n1851), .A2(n1297), .B1(n1883), .B2(n1198), .ZN(n4000)
         );
  OAI222_X1 U3185 ( .A1(n2139), .A2(n1177), .B1(n2171), .B2(n1174), .C1(n2107), 
        .C2(n1171), .ZN(n3997) );
  OAI222_X1 U3186 ( .A1(n2043), .A2(n1186), .B1(n2075), .B2(n1183), .C1(n2011), 
        .C2(n1180), .ZN(n3998) );
  NOR4_X1 U3187 ( .A1(n4006), .A2(n4007), .A3(n4008), .A4(n4009), .ZN(n4005)
         );
  OAI22_X1 U3188 ( .A1(n2203), .A2(n783), .B1(n2235), .B2(n780), .ZN(n4009) );
  OAI222_X1 U3189 ( .A1(n2491), .A2(n759), .B1(n2523), .B2(n756), .C1(n2459), 
        .C2(n753), .ZN(n4006) );
  OAI222_X1 U3190 ( .A1(n2395), .A2(n768), .B1(n2427), .B2(n765), .C1(n2363), 
        .C2(n762), .ZN(n4007) );
  NOR4_X1 U3191 ( .A1(n5399), .A2(n5400), .A3(n5401), .A4(n5402), .ZN(n5398)
         );
  OAI22_X1 U3192 ( .A1(n1850), .A2(n489), .B1(n1882), .B2(n486), .ZN(n5402) );
  OAI222_X1 U3193 ( .A1(n2138), .A2(n465), .B1(n2170), .B2(n462), .C1(n2106), 
        .C2(n459), .ZN(n5399) );
  OAI222_X1 U3194 ( .A1(n2042), .A2(n474), .B1(n2074), .B2(n471), .C1(n2010), 
        .C2(n468), .ZN(n5400) );
  NOR4_X1 U3195 ( .A1(n5408), .A2(n5409), .A3(n5410), .A4(n5411), .ZN(n5407)
         );
  OAI22_X1 U3196 ( .A1(n2202), .A2(n71), .B1(n2234), .B2(n68), .ZN(n5411) );
  OAI222_X1 U3197 ( .A1(n2490), .A2(n47), .B1(n2522), .B2(n44), .C1(n2458), 
        .C2(n41), .ZN(n5408) );
  OAI222_X1 U3198 ( .A1(n2394), .A2(n56), .B1(n2426), .B2(n53), .C1(n2362), 
        .C2(n50), .ZN(n5409) );
  NOR4_X1 U3199 ( .A1(n3956), .A2(n3957), .A3(n3958), .A4(n3959), .ZN(n3955)
         );
  OAI22_X1 U3200 ( .A1(n1850), .A2(n1297), .B1(n1882), .B2(n1198), .ZN(n3959)
         );
  OAI222_X1 U3201 ( .A1(n2138), .A2(n1177), .B1(n2170), .B2(n1174), .C1(n2106), 
        .C2(n1171), .ZN(n3956) );
  OAI222_X1 U3202 ( .A1(n2042), .A2(n1186), .B1(n2074), .B2(n1183), .C1(n2010), 
        .C2(n1180), .ZN(n3957) );
  NOR4_X1 U3203 ( .A1(n3965), .A2(n3966), .A3(n3967), .A4(n3968), .ZN(n3964)
         );
  OAI22_X1 U3204 ( .A1(n2202), .A2(n783), .B1(n2234), .B2(n780), .ZN(n3968) );
  OAI222_X1 U3205 ( .A1(n2490), .A2(n759), .B1(n2522), .B2(n756), .C1(n2458), 
        .C2(n753), .ZN(n3965) );
  OAI222_X1 U3206 ( .A1(n2394), .A2(n768), .B1(n2426), .B2(n765), .C1(n2362), 
        .C2(n762), .ZN(n3966) );
  NOR4_X1 U3207 ( .A1(n5358), .A2(n5359), .A3(n5360), .A4(n5361), .ZN(n5357)
         );
  OAI22_X1 U3208 ( .A1(n1849), .A2(n489), .B1(n1881), .B2(n486), .ZN(n5361) );
  OAI222_X1 U3209 ( .A1(n2137), .A2(n465), .B1(n2169), .B2(n462), .C1(n2105), 
        .C2(n459), .ZN(n5358) );
  OAI222_X1 U3210 ( .A1(n2041), .A2(n474), .B1(n2073), .B2(n471), .C1(n2009), 
        .C2(n468), .ZN(n5359) );
  NOR4_X1 U3211 ( .A1(n5367), .A2(n5368), .A3(n5369), .A4(n5370), .ZN(n5366)
         );
  OAI22_X1 U3212 ( .A1(n2201), .A2(n71), .B1(n2233), .B2(n68), .ZN(n5370) );
  OAI222_X1 U3213 ( .A1(n2489), .A2(n47), .B1(n2521), .B2(n44), .C1(n2457), 
        .C2(n41), .ZN(n5367) );
  OAI222_X1 U3214 ( .A1(n2393), .A2(n56), .B1(n2425), .B2(n53), .C1(n2361), 
        .C2(n50), .ZN(n5368) );
  NOR4_X1 U3215 ( .A1(n3915), .A2(n3916), .A3(n3917), .A4(n3918), .ZN(n3914)
         );
  OAI22_X1 U3216 ( .A1(n1849), .A2(n1297), .B1(n1881), .B2(n1198), .ZN(n3918)
         );
  OAI222_X1 U3217 ( .A1(n2137), .A2(n1177), .B1(n2169), .B2(n1174), .C1(n2105), 
        .C2(n1171), .ZN(n3915) );
  OAI222_X1 U3218 ( .A1(n2041), .A2(n1186), .B1(n2073), .B2(n1183), .C1(n2009), 
        .C2(n1180), .ZN(n3916) );
  NOR4_X1 U3219 ( .A1(n3924), .A2(n3925), .A3(n3926), .A4(n3927), .ZN(n3923)
         );
  OAI22_X1 U3220 ( .A1(n2201), .A2(n783), .B1(n2233), .B2(n780), .ZN(n3927) );
  OAI222_X1 U3221 ( .A1(n2489), .A2(n759), .B1(n2521), .B2(n756), .C1(n2457), 
        .C2(n753), .ZN(n3924) );
  OAI222_X1 U3222 ( .A1(n2393), .A2(n768), .B1(n2425), .B2(n765), .C1(n2361), 
        .C2(n762), .ZN(n3925) );
  NOR4_X1 U3223 ( .A1(n5317), .A2(n5318), .A3(n5319), .A4(n5320), .ZN(n5316)
         );
  OAI22_X1 U3224 ( .A1(n1848), .A2(n489), .B1(n1880), .B2(n486), .ZN(n5320) );
  OAI222_X1 U3225 ( .A1(n2136), .A2(n465), .B1(n2168), .B2(n462), .C1(n2104), 
        .C2(n459), .ZN(n5317) );
  OAI222_X1 U3226 ( .A1(n2040), .A2(n474), .B1(n2072), .B2(n471), .C1(n2008), 
        .C2(n468), .ZN(n5318) );
  NOR4_X1 U3227 ( .A1(n5326), .A2(n5327), .A3(n5328), .A4(n5329), .ZN(n5325)
         );
  OAI22_X1 U3228 ( .A1(n2200), .A2(n71), .B1(n2232), .B2(n68), .ZN(n5329) );
  OAI222_X1 U3229 ( .A1(n2488), .A2(n47), .B1(n2520), .B2(n44), .C1(n2456), 
        .C2(n41), .ZN(n5326) );
  OAI222_X1 U3230 ( .A1(n2392), .A2(n56), .B1(n2424), .B2(n53), .C1(n2360), 
        .C2(n50), .ZN(n5327) );
  NOR4_X1 U3231 ( .A1(n3874), .A2(n3875), .A3(n3876), .A4(n3877), .ZN(n3873)
         );
  OAI22_X1 U3232 ( .A1(n1848), .A2(n1297), .B1(n1880), .B2(n1198), .ZN(n3877)
         );
  OAI222_X1 U3233 ( .A1(n2136), .A2(n1177), .B1(n2168), .B2(n1174), .C1(n2104), 
        .C2(n1171), .ZN(n3874) );
  OAI222_X1 U3234 ( .A1(n2040), .A2(n1186), .B1(n2072), .B2(n1183), .C1(n2008), 
        .C2(n1180), .ZN(n3875) );
  NOR4_X1 U3235 ( .A1(n3883), .A2(n3884), .A3(n3885), .A4(n3886), .ZN(n3882)
         );
  OAI22_X1 U3236 ( .A1(n2200), .A2(n783), .B1(n2232), .B2(n780), .ZN(n3886) );
  OAI222_X1 U3237 ( .A1(n2488), .A2(n759), .B1(n2520), .B2(n756), .C1(n2456), 
        .C2(n753), .ZN(n3883) );
  OAI222_X1 U3238 ( .A1(n2392), .A2(n768), .B1(n2424), .B2(n765), .C1(n2360), 
        .C2(n762), .ZN(n3884) );
  NOR4_X1 U3239 ( .A1(n5276), .A2(n5277), .A3(n5278), .A4(n5279), .ZN(n5275)
         );
  OAI22_X1 U3240 ( .A1(n1847), .A2(n490), .B1(n1879), .B2(n487), .ZN(n5279) );
  OAI222_X1 U3241 ( .A1(n2135), .A2(n466), .B1(n2167), .B2(n463), .C1(n2103), 
        .C2(n460), .ZN(n5276) );
  OAI222_X1 U3242 ( .A1(n2039), .A2(n475), .B1(n2071), .B2(n472), .C1(n2007), 
        .C2(n469), .ZN(n5277) );
  NOR4_X1 U3243 ( .A1(n5285), .A2(n5286), .A3(n5287), .A4(n5288), .ZN(n5284)
         );
  OAI22_X1 U3244 ( .A1(n2199), .A2(n72), .B1(n2231), .B2(n69), .ZN(n5288) );
  OAI222_X1 U3245 ( .A1(n2487), .A2(n48), .B1(n2519), .B2(n45), .C1(n2455), 
        .C2(n42), .ZN(n5285) );
  OAI222_X1 U3246 ( .A1(n2391), .A2(n57), .B1(n2423), .B2(n54), .C1(n2359), 
        .C2(n51), .ZN(n5286) );
  NOR4_X1 U3247 ( .A1(n3833), .A2(n3834), .A3(n3835), .A4(n3836), .ZN(n3832)
         );
  OAI22_X1 U3248 ( .A1(n1847), .A2(n1298), .B1(n1879), .B2(n1199), .ZN(n3836)
         );
  OAI222_X1 U3249 ( .A1(n2135), .A2(n1178), .B1(n2167), .B2(n1175), .C1(n2103), 
        .C2(n1172), .ZN(n3833) );
  OAI222_X1 U3250 ( .A1(n2039), .A2(n1187), .B1(n2071), .B2(n1184), .C1(n2007), 
        .C2(n1181), .ZN(n3834) );
  NOR4_X1 U3251 ( .A1(n3842), .A2(n3843), .A3(n3844), .A4(n3845), .ZN(n3841)
         );
  OAI22_X1 U3252 ( .A1(n2199), .A2(n1136), .B1(n2231), .B2(n781), .ZN(n3845)
         );
  OAI222_X1 U3253 ( .A1(n2487), .A2(n760), .B1(n2519), .B2(n757), .C1(n2455), 
        .C2(n754), .ZN(n3842) );
  OAI222_X1 U3254 ( .A1(n2391), .A2(n769), .B1(n2423), .B2(n766), .C1(n2359), 
        .C2(n763), .ZN(n3843) );
  NOR4_X1 U3255 ( .A1(n5235), .A2(n5236), .A3(n5237), .A4(n5238), .ZN(n5234)
         );
  OAI22_X1 U3256 ( .A1(n1846), .A2(n490), .B1(n1878), .B2(n487), .ZN(n5238) );
  OAI222_X1 U3257 ( .A1(n2134), .A2(n466), .B1(n2166), .B2(n463), .C1(n2102), 
        .C2(n460), .ZN(n5235) );
  OAI222_X1 U3258 ( .A1(n2038), .A2(n475), .B1(n2070), .B2(n472), .C1(n2006), 
        .C2(n469), .ZN(n5236) );
  NOR4_X1 U3259 ( .A1(n5244), .A2(n5245), .A3(n5246), .A4(n5247), .ZN(n5243)
         );
  OAI22_X1 U3260 ( .A1(n2198), .A2(n72), .B1(n2230), .B2(n69), .ZN(n5247) );
  OAI222_X1 U3261 ( .A1(n2486), .A2(n48), .B1(n2518), .B2(n45), .C1(n2454), 
        .C2(n42), .ZN(n5244) );
  OAI222_X1 U3262 ( .A1(n2390), .A2(n57), .B1(n2422), .B2(n54), .C1(n2358), 
        .C2(n51), .ZN(n5245) );
  NOR4_X1 U3263 ( .A1(n3792), .A2(n3793), .A3(n3794), .A4(n3795), .ZN(n3791)
         );
  OAI22_X1 U3264 ( .A1(n1846), .A2(n1298), .B1(n1878), .B2(n1199), .ZN(n3795)
         );
  OAI222_X1 U3265 ( .A1(n2134), .A2(n1178), .B1(n2166), .B2(n1175), .C1(n2102), 
        .C2(n1172), .ZN(n3792) );
  OAI222_X1 U3266 ( .A1(n2038), .A2(n1187), .B1(n2070), .B2(n1184), .C1(n2006), 
        .C2(n1181), .ZN(n3793) );
  NOR4_X1 U3267 ( .A1(n3801), .A2(n3802), .A3(n3803), .A4(n3804), .ZN(n3800)
         );
  OAI22_X1 U3268 ( .A1(n2198), .A2(n1136), .B1(n2230), .B2(n781), .ZN(n3804)
         );
  OAI222_X1 U3269 ( .A1(n2486), .A2(n760), .B1(n2518), .B2(n757), .C1(n2454), 
        .C2(n754), .ZN(n3801) );
  OAI222_X1 U3270 ( .A1(n2390), .A2(n769), .B1(n2422), .B2(n766), .C1(n2358), 
        .C2(n763), .ZN(n3802) );
  NOR4_X1 U3271 ( .A1(n5194), .A2(n5195), .A3(n5196), .A4(n5197), .ZN(n5193)
         );
  OAI22_X1 U3272 ( .A1(n1845), .A2(n490), .B1(n1877), .B2(n487), .ZN(n5197) );
  OAI222_X1 U3273 ( .A1(n2133), .A2(n466), .B1(n2165), .B2(n463), .C1(n2101), 
        .C2(n460), .ZN(n5194) );
  OAI222_X1 U3274 ( .A1(n2037), .A2(n475), .B1(n2069), .B2(n472), .C1(n2005), 
        .C2(n469), .ZN(n5195) );
  NOR4_X1 U3275 ( .A1(n5203), .A2(n5204), .A3(n5205), .A4(n5206), .ZN(n5202)
         );
  OAI22_X1 U3276 ( .A1(n2197), .A2(n72), .B1(n2229), .B2(n69), .ZN(n5206) );
  OAI222_X1 U3277 ( .A1(n2485), .A2(n48), .B1(n2517), .B2(n45), .C1(n2453), 
        .C2(n42), .ZN(n5203) );
  OAI222_X1 U3278 ( .A1(n2389), .A2(n57), .B1(n2421), .B2(n54), .C1(n2357), 
        .C2(n51), .ZN(n5204) );
  NOR4_X1 U3279 ( .A1(n3751), .A2(n3752), .A3(n3753), .A4(n3754), .ZN(n3750)
         );
  OAI22_X1 U3280 ( .A1(n1845), .A2(n1298), .B1(n1877), .B2(n1199), .ZN(n3754)
         );
  OAI222_X1 U3281 ( .A1(n2133), .A2(n1178), .B1(n2165), .B2(n1175), .C1(n2101), 
        .C2(n1172), .ZN(n3751) );
  OAI222_X1 U3282 ( .A1(n2037), .A2(n1187), .B1(n2069), .B2(n1184), .C1(n2005), 
        .C2(n1181), .ZN(n3752) );
  NOR4_X1 U3283 ( .A1(n3760), .A2(n3761), .A3(n3762), .A4(n3763), .ZN(n3759)
         );
  OAI22_X1 U3284 ( .A1(n2197), .A2(n1136), .B1(n2229), .B2(n781), .ZN(n3763)
         );
  OAI222_X1 U3285 ( .A1(n2485), .A2(n760), .B1(n2517), .B2(n757), .C1(n2453), 
        .C2(n754), .ZN(n3760) );
  OAI222_X1 U3286 ( .A1(n2389), .A2(n769), .B1(n2421), .B2(n766), .C1(n2357), 
        .C2(n763), .ZN(n3761) );
  NOR4_X1 U3287 ( .A1(n5153), .A2(n5154), .A3(n5155), .A4(n5156), .ZN(n5152)
         );
  OAI22_X1 U3288 ( .A1(n1844), .A2(n490), .B1(n1876), .B2(n487), .ZN(n5156) );
  OAI222_X1 U3289 ( .A1(n2132), .A2(n466), .B1(n2164), .B2(n463), .C1(n2100), 
        .C2(n460), .ZN(n5153) );
  OAI222_X1 U3290 ( .A1(n2036), .A2(n475), .B1(n2068), .B2(n472), .C1(n2004), 
        .C2(n469), .ZN(n5154) );
  NOR4_X1 U3291 ( .A1(n5162), .A2(n5163), .A3(n5164), .A4(n5165), .ZN(n5161)
         );
  OAI22_X1 U3292 ( .A1(n2196), .A2(n72), .B1(n2228), .B2(n69), .ZN(n5165) );
  OAI222_X1 U3293 ( .A1(n2484), .A2(n48), .B1(n2516), .B2(n45), .C1(n2452), 
        .C2(n42), .ZN(n5162) );
  OAI222_X1 U3294 ( .A1(n2388), .A2(n57), .B1(n2420), .B2(n54), .C1(n2356), 
        .C2(n51), .ZN(n5163) );
  NOR4_X1 U3295 ( .A1(n3710), .A2(n3711), .A3(n3712), .A4(n3713), .ZN(n3709)
         );
  OAI22_X1 U3296 ( .A1(n1844), .A2(n1298), .B1(n1876), .B2(n1199), .ZN(n3713)
         );
  OAI222_X1 U3297 ( .A1(n2132), .A2(n1178), .B1(n2164), .B2(n1175), .C1(n2100), 
        .C2(n1172), .ZN(n3710) );
  OAI222_X1 U3298 ( .A1(n2036), .A2(n1187), .B1(n2068), .B2(n1184), .C1(n2004), 
        .C2(n1181), .ZN(n3711) );
  NOR4_X1 U3299 ( .A1(n3719), .A2(n3720), .A3(n3721), .A4(n3722), .ZN(n3718)
         );
  OAI22_X1 U3300 ( .A1(n2196), .A2(n1136), .B1(n2228), .B2(n781), .ZN(n3722)
         );
  OAI222_X1 U3301 ( .A1(n2484), .A2(n760), .B1(n2516), .B2(n757), .C1(n2452), 
        .C2(n754), .ZN(n3719) );
  OAI222_X1 U3302 ( .A1(n2388), .A2(n769), .B1(n2420), .B2(n766), .C1(n2356), 
        .C2(n763), .ZN(n3720) );
  NOR4_X1 U3303 ( .A1(n5112), .A2(n5113), .A3(n5114), .A4(n5115), .ZN(n5111)
         );
  OAI22_X1 U3304 ( .A1(n1843), .A2(n490), .B1(n1875), .B2(n487), .ZN(n5115) );
  OAI222_X1 U3305 ( .A1(n2131), .A2(n466), .B1(n2163), .B2(n463), .C1(n2099), 
        .C2(n460), .ZN(n5112) );
  OAI222_X1 U3306 ( .A1(n2035), .A2(n475), .B1(n2067), .B2(n472), .C1(n2003), 
        .C2(n469), .ZN(n5113) );
  NOR4_X1 U3307 ( .A1(n5121), .A2(n5122), .A3(n5123), .A4(n5124), .ZN(n5120)
         );
  OAI22_X1 U3308 ( .A1(n2195), .A2(n72), .B1(n2227), .B2(n69), .ZN(n5124) );
  OAI222_X1 U3309 ( .A1(n2483), .A2(n48), .B1(n2515), .B2(n45), .C1(n2451), 
        .C2(n42), .ZN(n5121) );
  OAI222_X1 U3310 ( .A1(n2387), .A2(n57), .B1(n2419), .B2(n54), .C1(n2355), 
        .C2(n51), .ZN(n5122) );
  NOR4_X1 U3311 ( .A1(n3669), .A2(n3670), .A3(n3671), .A4(n3672), .ZN(n3668)
         );
  OAI22_X1 U3312 ( .A1(n1843), .A2(n1298), .B1(n1875), .B2(n1199), .ZN(n3672)
         );
  OAI222_X1 U3313 ( .A1(n2131), .A2(n1178), .B1(n2163), .B2(n1175), .C1(n2099), 
        .C2(n1172), .ZN(n3669) );
  OAI222_X1 U3314 ( .A1(n2035), .A2(n1187), .B1(n2067), .B2(n1184), .C1(n2003), 
        .C2(n1181), .ZN(n3670) );
  NOR4_X1 U3315 ( .A1(n3678), .A2(n3679), .A3(n3680), .A4(n3681), .ZN(n3677)
         );
  OAI22_X1 U3316 ( .A1(n2195), .A2(n1136), .B1(n2227), .B2(n781), .ZN(n3681)
         );
  OAI222_X1 U3317 ( .A1(n2483), .A2(n760), .B1(n2515), .B2(n757), .C1(n2451), 
        .C2(n754), .ZN(n3678) );
  OAI222_X1 U3318 ( .A1(n2387), .A2(n769), .B1(n2419), .B2(n766), .C1(n2355), 
        .C2(n763), .ZN(n3679) );
  NOR4_X1 U3319 ( .A1(n5071), .A2(n5072), .A3(n5073), .A4(n5074), .ZN(n5070)
         );
  OAI22_X1 U3320 ( .A1(n1842), .A2(n490), .B1(n1874), .B2(n487), .ZN(n5074) );
  OAI222_X1 U3321 ( .A1(n2130), .A2(n466), .B1(n2162), .B2(n463), .C1(n2098), 
        .C2(n460), .ZN(n5071) );
  OAI222_X1 U3322 ( .A1(n2034), .A2(n475), .B1(n2066), .B2(n472), .C1(n2002), 
        .C2(n469), .ZN(n5072) );
  NOR4_X1 U3323 ( .A1(n5080), .A2(n5081), .A3(n5082), .A4(n5083), .ZN(n5079)
         );
  OAI22_X1 U3324 ( .A1(n2194), .A2(n72), .B1(n2226), .B2(n69), .ZN(n5083) );
  OAI222_X1 U3325 ( .A1(n2482), .A2(n48), .B1(n2514), .B2(n45), .C1(n2450), 
        .C2(n42), .ZN(n5080) );
  OAI222_X1 U3326 ( .A1(n2386), .A2(n57), .B1(n2418), .B2(n54), .C1(n2354), 
        .C2(n51), .ZN(n5081) );
  NOR4_X1 U3327 ( .A1(n3628), .A2(n3629), .A3(n3630), .A4(n3631), .ZN(n3627)
         );
  OAI22_X1 U3328 ( .A1(n1842), .A2(n1298), .B1(n1874), .B2(n1199), .ZN(n3631)
         );
  OAI222_X1 U3329 ( .A1(n2130), .A2(n1178), .B1(n2162), .B2(n1175), .C1(n2098), 
        .C2(n1172), .ZN(n3628) );
  OAI222_X1 U3330 ( .A1(n2034), .A2(n1187), .B1(n2066), .B2(n1184), .C1(n2002), 
        .C2(n1181), .ZN(n3629) );
  NOR4_X1 U3331 ( .A1(n3637), .A2(n3638), .A3(n3639), .A4(n3640), .ZN(n3636)
         );
  OAI22_X1 U3332 ( .A1(n2194), .A2(n1136), .B1(n2226), .B2(n781), .ZN(n3640)
         );
  OAI222_X1 U3333 ( .A1(n2482), .A2(n760), .B1(n2514), .B2(n757), .C1(n2450), 
        .C2(n754), .ZN(n3637) );
  OAI222_X1 U3334 ( .A1(n2386), .A2(n769), .B1(n2418), .B2(n766), .C1(n2354), 
        .C2(n763), .ZN(n3638) );
  NOR4_X1 U3335 ( .A1(n5030), .A2(n5031), .A3(n5032), .A4(n5033), .ZN(n5029)
         );
  OAI22_X1 U3336 ( .A1(n1841), .A2(n490), .B1(n1873), .B2(n487), .ZN(n5033) );
  OAI222_X1 U3337 ( .A1(n2129), .A2(n466), .B1(n2161), .B2(n463), .C1(n2097), 
        .C2(n460), .ZN(n5030) );
  OAI222_X1 U3338 ( .A1(n2033), .A2(n475), .B1(n2065), .B2(n472), .C1(n2001), 
        .C2(n469), .ZN(n5031) );
  NOR4_X1 U3339 ( .A1(n5039), .A2(n5040), .A3(n5041), .A4(n5042), .ZN(n5038)
         );
  OAI22_X1 U3340 ( .A1(n2193), .A2(n72), .B1(n2225), .B2(n69), .ZN(n5042) );
  OAI222_X1 U3341 ( .A1(n2481), .A2(n48), .B1(n2513), .B2(n45), .C1(n2449), 
        .C2(n42), .ZN(n5039) );
  OAI222_X1 U3342 ( .A1(n2385), .A2(n57), .B1(n2417), .B2(n54), .C1(n2353), 
        .C2(n51), .ZN(n5040) );
  NOR4_X1 U3343 ( .A1(n3587), .A2(n3588), .A3(n3589), .A4(n3590), .ZN(n3586)
         );
  OAI22_X1 U3344 ( .A1(n1841), .A2(n1298), .B1(n1873), .B2(n1199), .ZN(n3590)
         );
  OAI222_X1 U3345 ( .A1(n2129), .A2(n1178), .B1(n2161), .B2(n1175), .C1(n2097), 
        .C2(n1172), .ZN(n3587) );
  OAI222_X1 U3346 ( .A1(n2033), .A2(n1187), .B1(n2065), .B2(n1184), .C1(n2001), 
        .C2(n1181), .ZN(n3588) );
  NOR4_X1 U3347 ( .A1(n3596), .A2(n3597), .A3(n3598), .A4(n3599), .ZN(n3595)
         );
  OAI22_X1 U3348 ( .A1(n2193), .A2(n1136), .B1(n2225), .B2(n781), .ZN(n3599)
         );
  OAI222_X1 U3349 ( .A1(n2481), .A2(n760), .B1(n2513), .B2(n757), .C1(n2449), 
        .C2(n754), .ZN(n3596) );
  OAI222_X1 U3350 ( .A1(n2385), .A2(n769), .B1(n2417), .B2(n766), .C1(n2353), 
        .C2(n763), .ZN(n3597) );
  NOR4_X1 U3351 ( .A1(n4945), .A2(n4946), .A3(n4947), .A4(n4948), .ZN(n4944)
         );
  OAI22_X1 U3352 ( .A1(n1840), .A2(n490), .B1(n1872), .B2(n487), .ZN(n4948) );
  OAI222_X1 U3353 ( .A1(n2128), .A2(n466), .B1(n2160), .B2(n463), .C1(n2096), 
        .C2(n460), .ZN(n4945) );
  OAI222_X1 U3354 ( .A1(n2032), .A2(n475), .B1(n2064), .B2(n472), .C1(n2000), 
        .C2(n469), .ZN(n4946) );
  NOR4_X1 U3355 ( .A1(n4976), .A2(n4977), .A3(n4978), .A4(n4979), .ZN(n4975)
         );
  OAI22_X1 U3356 ( .A1(n2192), .A2(n72), .B1(n2224), .B2(n69), .ZN(n4979) );
  OAI222_X1 U3357 ( .A1(n2480), .A2(n48), .B1(n2512), .B2(n45), .C1(n2448), 
        .C2(n42), .ZN(n4976) );
  OAI222_X1 U3358 ( .A1(n2384), .A2(n57), .B1(n2416), .B2(n54), .C1(n2352), 
        .C2(n51), .ZN(n4977) );
  NOR4_X1 U3359 ( .A1(n3502), .A2(n3503), .A3(n3504), .A4(n3505), .ZN(n3501)
         );
  OAI22_X1 U3360 ( .A1(n1840), .A2(n1298), .B1(n1872), .B2(n1199), .ZN(n3505)
         );
  OAI222_X1 U3361 ( .A1(n2128), .A2(n1178), .B1(n2160), .B2(n1175), .C1(n2096), 
        .C2(n1172), .ZN(n3502) );
  OAI222_X1 U3362 ( .A1(n2032), .A2(n1187), .B1(n2064), .B2(n1184), .C1(n2000), 
        .C2(n1181), .ZN(n3503) );
  NOR4_X1 U3363 ( .A1(n3533), .A2(n3534), .A3(n3535), .A4(n3536), .ZN(n3532)
         );
  OAI22_X1 U3364 ( .A1(n2192), .A2(n1136), .B1(n2224), .B2(n781), .ZN(n3536)
         );
  OAI222_X1 U3365 ( .A1(n2480), .A2(n760), .B1(n2512), .B2(n757), .C1(n2448), 
        .C2(n754), .ZN(n3533) );
  OAI222_X1 U3366 ( .A1(n2384), .A2(n769), .B1(n2416), .B2(n766), .C1(n2352), 
        .C2(n763), .ZN(n3534) );
  AOI22_X1 U3367 ( .A1(N2161), .A2(n3391), .B1(N2154), .B2(N2151), .ZN(n3406)
         );
  AOI22_X1 U3368 ( .A1(N2163), .A2(n3391), .B1(N2156), .B2(N2151), .ZN(n3359)
         );
  INV_X1 U3369 ( .A(ADD_WR[3]), .ZN(N2163) );
  AOI22_X1 U3370 ( .A1(N2160), .A2(n3391), .B1(N2153), .B2(N2151), .ZN(n3405)
         );
  AOI22_X1 U3371 ( .A1(N2162), .A2(n3391), .B1(N2155), .B2(N2151), .ZN(n3377)
         );
  AOI221_X1 U3372 ( .B1(n455), .B2(\REGISTERS[45][0] ), .C1(n452), .C2(
        \REGISTERS[44][0] ), .A(n6299), .ZN(n6290) );
  OAI222_X1 U3373 ( .A1(n1615), .A2(n449), .B1(n1647), .B2(n446), .C1(n1583), 
        .C2(n443), .ZN(n6299) );
  AOI221_X1 U3374 ( .B1(n37), .B2(\REGISTERS[78][0] ), .C1(n34), .C2(
        \REGISTERS[77][0] ), .A(n6311), .ZN(n6303) );
  OAI222_X1 U3375 ( .A1(n2671), .A2(n31), .B1(n2703), .B2(n28), .C1(n2639), 
        .C2(n25), .ZN(n6311) );
  AOI221_X1 U3376 ( .B1(n1167), .B2(\REGISTERS[45][0] ), .C1(n1164), .C2(
        \REGISTERS[44][0] ), .A(n4856), .ZN(n4847) );
  OAI222_X1 U3377 ( .A1(n1615), .A2(n1161), .B1(n1647), .B2(n1158), .C1(n1583), 
        .C2(n1155), .ZN(n4856) );
  AOI221_X1 U3378 ( .B1(n749), .B2(\REGISTERS[78][0] ), .C1(n746), .C2(
        \REGISTERS[77][0] ), .A(n4868), .ZN(n4860) );
  OAI222_X1 U3379 ( .A1(n2671), .A2(n743), .B1(n2703), .B2(n740), .C1(n2639), 
        .C2(n737), .ZN(n4868) );
  AOI221_X1 U3380 ( .B1(n455), .B2(\REGISTERS[45][1] ), .C1(n452), .C2(
        \REGISTERS[44][1] ), .A(n6223), .ZN(n6217) );
  OAI222_X1 U3381 ( .A1(n1614), .A2(n449), .B1(n1646), .B2(n446), .C1(n1582), 
        .C2(n443), .ZN(n6223) );
  AOI221_X1 U3382 ( .B1(n37), .B2(\REGISTERS[78][1] ), .C1(n34), .C2(
        \REGISTERS[77][1] ), .A(n6232), .ZN(n6226) );
  OAI222_X1 U3383 ( .A1(n2670), .A2(n31), .B1(n2702), .B2(n28), .C1(n2638), 
        .C2(n25), .ZN(n6232) );
  AOI221_X1 U3384 ( .B1(n1167), .B2(\REGISTERS[45][1] ), .C1(n1164), .C2(
        \REGISTERS[44][1] ), .A(n4780), .ZN(n4774) );
  OAI222_X1 U3385 ( .A1(n1614), .A2(n1161), .B1(n1646), .B2(n1158), .C1(n1582), 
        .C2(n1155), .ZN(n4780) );
  AOI221_X1 U3386 ( .B1(n749), .B2(\REGISTERS[78][1] ), .C1(n746), .C2(
        \REGISTERS[77][1] ), .A(n4789), .ZN(n4783) );
  OAI222_X1 U3387 ( .A1(n2670), .A2(n743), .B1(n2702), .B2(n740), .C1(n2638), 
        .C2(n737), .ZN(n4789) );
  AOI221_X1 U3388 ( .B1(n455), .B2(\REGISTERS[45][2] ), .C1(n452), .C2(
        \REGISTERS[44][2] ), .A(n6182), .ZN(n6176) );
  OAI222_X1 U3389 ( .A1(n1613), .A2(n449), .B1(n1645), .B2(n446), .C1(n1581), 
        .C2(n443), .ZN(n6182) );
  AOI221_X1 U3390 ( .B1(n37), .B2(\REGISTERS[78][2] ), .C1(n34), .C2(
        \REGISTERS[77][2] ), .A(n6191), .ZN(n6185) );
  OAI222_X1 U3391 ( .A1(n2669), .A2(n31), .B1(n2701), .B2(n28), .C1(n2637), 
        .C2(n25), .ZN(n6191) );
  AOI221_X1 U3392 ( .B1(n1167), .B2(\REGISTERS[45][2] ), .C1(n1164), .C2(
        \REGISTERS[44][2] ), .A(n4739), .ZN(n4733) );
  OAI222_X1 U3393 ( .A1(n1613), .A2(n1161), .B1(n1645), .B2(n1158), .C1(n1581), 
        .C2(n1155), .ZN(n4739) );
  AOI221_X1 U3394 ( .B1(n749), .B2(\REGISTERS[78][2] ), .C1(n746), .C2(
        \REGISTERS[77][2] ), .A(n4748), .ZN(n4742) );
  OAI222_X1 U3395 ( .A1(n2669), .A2(n743), .B1(n2701), .B2(n740), .C1(n2637), 
        .C2(n737), .ZN(n4748) );
  AOI221_X1 U3396 ( .B1(n455), .B2(\REGISTERS[45][3] ), .C1(n452), .C2(
        \REGISTERS[44][3] ), .A(n6141), .ZN(n6135) );
  OAI222_X1 U3397 ( .A1(n1612), .A2(n449), .B1(n1644), .B2(n446), .C1(n1580), 
        .C2(n443), .ZN(n6141) );
  AOI221_X1 U3398 ( .B1(n37), .B2(\REGISTERS[78][3] ), .C1(n34), .C2(
        \REGISTERS[77][3] ), .A(n6150), .ZN(n6144) );
  OAI222_X1 U3399 ( .A1(n2668), .A2(n31), .B1(n2700), .B2(n28), .C1(n2636), 
        .C2(n25), .ZN(n6150) );
  AOI221_X1 U3400 ( .B1(n1167), .B2(\REGISTERS[45][3] ), .C1(n1164), .C2(
        \REGISTERS[44][3] ), .A(n4698), .ZN(n4692) );
  OAI222_X1 U3401 ( .A1(n1612), .A2(n1161), .B1(n1644), .B2(n1158), .C1(n1580), 
        .C2(n1155), .ZN(n4698) );
  AOI221_X1 U3402 ( .B1(n749), .B2(\REGISTERS[78][3] ), .C1(n746), .C2(
        \REGISTERS[77][3] ), .A(n4707), .ZN(n4701) );
  OAI222_X1 U3403 ( .A1(n2668), .A2(n743), .B1(n2700), .B2(n740), .C1(n2636), 
        .C2(n737), .ZN(n4707) );
  AOI221_X1 U3404 ( .B1(n455), .B2(\REGISTERS[45][4] ), .C1(n452), .C2(
        \REGISTERS[44][4] ), .A(n6100), .ZN(n6094) );
  OAI222_X1 U3405 ( .A1(n1611), .A2(n449), .B1(n1643), .B2(n446), .C1(n1579), 
        .C2(n443), .ZN(n6100) );
  AOI221_X1 U3406 ( .B1(n37), .B2(\REGISTERS[78][4] ), .C1(n34), .C2(
        \REGISTERS[77][4] ), .A(n6109), .ZN(n6103) );
  OAI222_X1 U3407 ( .A1(n2667), .A2(n31), .B1(n2699), .B2(n28), .C1(n2635), 
        .C2(n25), .ZN(n6109) );
  AOI221_X1 U3408 ( .B1(n1167), .B2(\REGISTERS[45][4] ), .C1(n1164), .C2(
        \REGISTERS[44][4] ), .A(n4657), .ZN(n4651) );
  OAI222_X1 U3409 ( .A1(n1611), .A2(n1161), .B1(n1643), .B2(n1158), .C1(n1579), 
        .C2(n1155), .ZN(n4657) );
  AOI221_X1 U3410 ( .B1(n749), .B2(\REGISTERS[78][4] ), .C1(n746), .C2(
        \REGISTERS[77][4] ), .A(n4666), .ZN(n4660) );
  OAI222_X1 U3411 ( .A1(n2667), .A2(n743), .B1(n2699), .B2(n740), .C1(n2635), 
        .C2(n737), .ZN(n4666) );
  AOI221_X1 U3412 ( .B1(n455), .B2(\REGISTERS[45][5] ), .C1(n452), .C2(
        \REGISTERS[44][5] ), .A(n6059), .ZN(n6053) );
  OAI222_X1 U3413 ( .A1(n1610), .A2(n449), .B1(n1642), .B2(n446), .C1(n1578), 
        .C2(n443), .ZN(n6059) );
  AOI221_X1 U3414 ( .B1(n37), .B2(\REGISTERS[78][5] ), .C1(n34), .C2(
        \REGISTERS[77][5] ), .A(n6068), .ZN(n6062) );
  OAI222_X1 U3415 ( .A1(n2666), .A2(n31), .B1(n2698), .B2(n28), .C1(n2634), 
        .C2(n25), .ZN(n6068) );
  AOI221_X1 U3416 ( .B1(n1167), .B2(\REGISTERS[45][5] ), .C1(n1164), .C2(
        \REGISTERS[44][5] ), .A(n4616), .ZN(n4610) );
  OAI222_X1 U3417 ( .A1(n1610), .A2(n1161), .B1(n1642), .B2(n1158), .C1(n1578), 
        .C2(n1155), .ZN(n4616) );
  AOI221_X1 U3418 ( .B1(n749), .B2(\REGISTERS[78][5] ), .C1(n746), .C2(
        \REGISTERS[77][5] ), .A(n4625), .ZN(n4619) );
  OAI222_X1 U3419 ( .A1(n2666), .A2(n743), .B1(n2698), .B2(n740), .C1(n2634), 
        .C2(n737), .ZN(n4625) );
  AOI221_X1 U3420 ( .B1(n455), .B2(\REGISTERS[45][6] ), .C1(n452), .C2(
        \REGISTERS[44][6] ), .A(n6018), .ZN(n6012) );
  OAI222_X1 U3421 ( .A1(n1609), .A2(n449), .B1(n1641), .B2(n446), .C1(n1577), 
        .C2(n443), .ZN(n6018) );
  AOI221_X1 U3422 ( .B1(n37), .B2(\REGISTERS[78][6] ), .C1(n34), .C2(
        \REGISTERS[77][6] ), .A(n6027), .ZN(n6021) );
  OAI222_X1 U3423 ( .A1(n2665), .A2(n31), .B1(n2697), .B2(n28), .C1(n2633), 
        .C2(n25), .ZN(n6027) );
  AOI221_X1 U3424 ( .B1(n1167), .B2(\REGISTERS[45][6] ), .C1(n1164), .C2(
        \REGISTERS[44][6] ), .A(n4575), .ZN(n4569) );
  OAI222_X1 U3425 ( .A1(n1609), .A2(n1161), .B1(n1641), .B2(n1158), .C1(n1577), 
        .C2(n1155), .ZN(n4575) );
  AOI221_X1 U3426 ( .B1(n749), .B2(\REGISTERS[78][6] ), .C1(n746), .C2(
        \REGISTERS[77][6] ), .A(n4584), .ZN(n4578) );
  OAI222_X1 U3427 ( .A1(n2665), .A2(n743), .B1(n2697), .B2(n740), .C1(n2633), 
        .C2(n737), .ZN(n4584) );
  AOI221_X1 U3428 ( .B1(n455), .B2(\REGISTERS[45][7] ), .C1(n452), .C2(
        \REGISTERS[44][7] ), .A(n5977), .ZN(n5971) );
  OAI222_X1 U3429 ( .A1(n1608), .A2(n449), .B1(n1640), .B2(n446), .C1(n1576), 
        .C2(n443), .ZN(n5977) );
  AOI221_X1 U3430 ( .B1(n37), .B2(\REGISTERS[78][7] ), .C1(n34), .C2(
        \REGISTERS[77][7] ), .A(n5986), .ZN(n5980) );
  OAI222_X1 U3431 ( .A1(n2664), .A2(n31), .B1(n2696), .B2(n28), .C1(n2632), 
        .C2(n25), .ZN(n5986) );
  AOI221_X1 U3432 ( .B1(n1167), .B2(\REGISTERS[45][7] ), .C1(n1164), .C2(
        \REGISTERS[44][7] ), .A(n4534), .ZN(n4528) );
  OAI222_X1 U3433 ( .A1(n1608), .A2(n1161), .B1(n1640), .B2(n1158), .C1(n1576), 
        .C2(n1155), .ZN(n4534) );
  AOI221_X1 U3434 ( .B1(n749), .B2(\REGISTERS[78][7] ), .C1(n746), .C2(
        \REGISTERS[77][7] ), .A(n4543), .ZN(n4537) );
  OAI222_X1 U3435 ( .A1(n2664), .A2(n743), .B1(n2696), .B2(n740), .C1(n2632), 
        .C2(n737), .ZN(n4543) );
  AOI221_X1 U3436 ( .B1(n455), .B2(\REGISTERS[45][8] ), .C1(n452), .C2(
        \REGISTERS[44][8] ), .A(n5936), .ZN(n5930) );
  OAI222_X1 U3437 ( .A1(n1607), .A2(n449), .B1(n1639), .B2(n446), .C1(n1575), 
        .C2(n443), .ZN(n5936) );
  AOI221_X1 U3438 ( .B1(n37), .B2(\REGISTERS[78][8] ), .C1(n34), .C2(
        \REGISTERS[77][8] ), .A(n5945), .ZN(n5939) );
  OAI222_X1 U3439 ( .A1(n2663), .A2(n31), .B1(n2695), .B2(n28), .C1(n2631), 
        .C2(n25), .ZN(n5945) );
  AOI221_X1 U3440 ( .B1(n1167), .B2(\REGISTERS[45][8] ), .C1(n1164), .C2(
        \REGISTERS[44][8] ), .A(n4493), .ZN(n4487) );
  OAI222_X1 U3441 ( .A1(n1607), .A2(n1161), .B1(n1639), .B2(n1158), .C1(n1575), 
        .C2(n1155), .ZN(n4493) );
  AOI221_X1 U3442 ( .B1(n749), .B2(\REGISTERS[78][8] ), .C1(n746), .C2(
        \REGISTERS[77][8] ), .A(n4502), .ZN(n4496) );
  OAI222_X1 U3443 ( .A1(n2663), .A2(n743), .B1(n2695), .B2(n740), .C1(n2631), 
        .C2(n737), .ZN(n4502) );
  AOI221_X1 U3444 ( .B1(n455), .B2(\REGISTERS[45][9] ), .C1(n452), .C2(
        \REGISTERS[44][9] ), .A(n5895), .ZN(n5889) );
  OAI222_X1 U3445 ( .A1(n1606), .A2(n449), .B1(n1638), .B2(n446), .C1(n1574), 
        .C2(n443), .ZN(n5895) );
  AOI221_X1 U3446 ( .B1(n37), .B2(\REGISTERS[78][9] ), .C1(n34), .C2(
        \REGISTERS[77][9] ), .A(n5904), .ZN(n5898) );
  OAI222_X1 U3447 ( .A1(n2662), .A2(n31), .B1(n2694), .B2(n28), .C1(n2630), 
        .C2(n25), .ZN(n5904) );
  AOI221_X1 U3448 ( .B1(n1167), .B2(\REGISTERS[45][9] ), .C1(n1164), .C2(
        \REGISTERS[44][9] ), .A(n4452), .ZN(n4446) );
  OAI222_X1 U3449 ( .A1(n1606), .A2(n1161), .B1(n1638), .B2(n1158), .C1(n1574), 
        .C2(n1155), .ZN(n4452) );
  AOI221_X1 U3450 ( .B1(n749), .B2(\REGISTERS[78][9] ), .C1(n746), .C2(
        \REGISTERS[77][9] ), .A(n4461), .ZN(n4455) );
  OAI222_X1 U3451 ( .A1(n2662), .A2(n743), .B1(n2694), .B2(n740), .C1(n2630), 
        .C2(n737), .ZN(n4461) );
  AOI221_X1 U3452 ( .B1(n455), .B2(\REGISTERS[45][10] ), .C1(n452), .C2(
        \REGISTERS[44][10] ), .A(n5854), .ZN(n5848) );
  OAI222_X1 U3453 ( .A1(n1605), .A2(n449), .B1(n1637), .B2(n446), .C1(n1573), 
        .C2(n443), .ZN(n5854) );
  AOI221_X1 U3454 ( .B1(n37), .B2(\REGISTERS[78][10] ), .C1(n34), .C2(
        \REGISTERS[77][10] ), .A(n5863), .ZN(n5857) );
  OAI222_X1 U3455 ( .A1(n2661), .A2(n31), .B1(n2693), .B2(n28), .C1(n2629), 
        .C2(n25), .ZN(n5863) );
  AOI221_X1 U3456 ( .B1(n1167), .B2(\REGISTERS[45][10] ), .C1(n1164), .C2(
        \REGISTERS[44][10] ), .A(n4411), .ZN(n4405) );
  OAI222_X1 U3457 ( .A1(n1605), .A2(n1161), .B1(n1637), .B2(n1158), .C1(n1573), 
        .C2(n1155), .ZN(n4411) );
  AOI221_X1 U3458 ( .B1(n749), .B2(\REGISTERS[78][10] ), .C1(n746), .C2(
        \REGISTERS[77][10] ), .A(n4420), .ZN(n4414) );
  OAI222_X1 U3459 ( .A1(n2661), .A2(n743), .B1(n2693), .B2(n740), .C1(n2629), 
        .C2(n737), .ZN(n4420) );
  AOI221_X1 U3460 ( .B1(n455), .B2(\REGISTERS[45][11] ), .C1(n452), .C2(
        \REGISTERS[44][11] ), .A(n5813), .ZN(n5807) );
  OAI222_X1 U3461 ( .A1(n1604), .A2(n449), .B1(n1636), .B2(n446), .C1(n1572), 
        .C2(n443), .ZN(n5813) );
  AOI221_X1 U3462 ( .B1(n37), .B2(\REGISTERS[78][11] ), .C1(n34), .C2(
        \REGISTERS[77][11] ), .A(n5822), .ZN(n5816) );
  OAI222_X1 U3463 ( .A1(n2660), .A2(n31), .B1(n2692), .B2(n28), .C1(n2628), 
        .C2(n25), .ZN(n5822) );
  AOI221_X1 U3464 ( .B1(n1167), .B2(\REGISTERS[45][11] ), .C1(n1164), .C2(
        \REGISTERS[44][11] ), .A(n4370), .ZN(n4364) );
  OAI222_X1 U3465 ( .A1(n1604), .A2(n1161), .B1(n1636), .B2(n1158), .C1(n1572), 
        .C2(n1155), .ZN(n4370) );
  AOI221_X1 U3466 ( .B1(n749), .B2(\REGISTERS[78][11] ), .C1(n746), .C2(
        \REGISTERS[77][11] ), .A(n4379), .ZN(n4373) );
  OAI222_X1 U3467 ( .A1(n2660), .A2(n743), .B1(n2692), .B2(n740), .C1(n2628), 
        .C2(n737), .ZN(n4379) );
  AOI221_X1 U3468 ( .B1(n456), .B2(\REGISTERS[45][12] ), .C1(n453), .C2(
        \REGISTERS[44][12] ), .A(n5772), .ZN(n5766) );
  OAI222_X1 U3469 ( .A1(n1603), .A2(n450), .B1(n1635), .B2(n447), .C1(n1571), 
        .C2(n444), .ZN(n5772) );
  AOI221_X1 U3470 ( .B1(n38), .B2(\REGISTERS[78][12] ), .C1(n35), .C2(
        \REGISTERS[77][12] ), .A(n5781), .ZN(n5775) );
  OAI222_X1 U3471 ( .A1(n2659), .A2(n32), .B1(n2691), .B2(n29), .C1(n2627), 
        .C2(n26), .ZN(n5781) );
  AOI221_X1 U3472 ( .B1(n1168), .B2(\REGISTERS[45][12] ), .C1(n1165), .C2(
        \REGISTERS[44][12] ), .A(n4329), .ZN(n4323) );
  OAI222_X1 U3473 ( .A1(n1603), .A2(n1162), .B1(n1635), .B2(n1159), .C1(n1571), 
        .C2(n1156), .ZN(n4329) );
  AOI221_X1 U3474 ( .B1(n750), .B2(\REGISTERS[78][12] ), .C1(n747), .C2(
        \REGISTERS[77][12] ), .A(n4338), .ZN(n4332) );
  OAI222_X1 U3475 ( .A1(n2659), .A2(n744), .B1(n2691), .B2(n741), .C1(n2627), 
        .C2(n738), .ZN(n4338) );
  AOI221_X1 U3476 ( .B1(n456), .B2(\REGISTERS[45][13] ), .C1(n453), .C2(
        \REGISTERS[44][13] ), .A(n5731), .ZN(n5725) );
  OAI222_X1 U3477 ( .A1(n1602), .A2(n450), .B1(n1634), .B2(n447), .C1(n1570), 
        .C2(n444), .ZN(n5731) );
  AOI221_X1 U3478 ( .B1(n38), .B2(\REGISTERS[78][13] ), .C1(n35), .C2(
        \REGISTERS[77][13] ), .A(n5740), .ZN(n5734) );
  OAI222_X1 U3479 ( .A1(n2658), .A2(n32), .B1(n2690), .B2(n29), .C1(n2626), 
        .C2(n26), .ZN(n5740) );
  AOI221_X1 U3480 ( .B1(n1168), .B2(\REGISTERS[45][13] ), .C1(n1165), .C2(
        \REGISTERS[44][13] ), .A(n4288), .ZN(n4282) );
  OAI222_X1 U3481 ( .A1(n1602), .A2(n1162), .B1(n1634), .B2(n1159), .C1(n1570), 
        .C2(n1156), .ZN(n4288) );
  AOI221_X1 U3482 ( .B1(n750), .B2(\REGISTERS[78][13] ), .C1(n747), .C2(
        \REGISTERS[77][13] ), .A(n4297), .ZN(n4291) );
  OAI222_X1 U3483 ( .A1(n2658), .A2(n744), .B1(n2690), .B2(n741), .C1(n2626), 
        .C2(n738), .ZN(n4297) );
  AOI221_X1 U3484 ( .B1(n456), .B2(\REGISTERS[45][14] ), .C1(n453), .C2(
        \REGISTERS[44][14] ), .A(n5690), .ZN(n5684) );
  OAI222_X1 U3485 ( .A1(n1601), .A2(n450), .B1(n1633), .B2(n447), .C1(n1569), 
        .C2(n444), .ZN(n5690) );
  AOI221_X1 U3486 ( .B1(n38), .B2(\REGISTERS[78][14] ), .C1(n35), .C2(
        \REGISTERS[77][14] ), .A(n5699), .ZN(n5693) );
  OAI222_X1 U3487 ( .A1(n2657), .A2(n32), .B1(n2689), .B2(n29), .C1(n2625), 
        .C2(n26), .ZN(n5699) );
  AOI221_X1 U3488 ( .B1(n1168), .B2(\REGISTERS[45][14] ), .C1(n1165), .C2(
        \REGISTERS[44][14] ), .A(n4247), .ZN(n4241) );
  OAI222_X1 U3489 ( .A1(n1601), .A2(n1162), .B1(n1633), .B2(n1159), .C1(n1569), 
        .C2(n1156), .ZN(n4247) );
  AOI221_X1 U3490 ( .B1(n750), .B2(\REGISTERS[78][14] ), .C1(n747), .C2(
        \REGISTERS[77][14] ), .A(n4256), .ZN(n4250) );
  OAI222_X1 U3491 ( .A1(n2657), .A2(n744), .B1(n2689), .B2(n741), .C1(n2625), 
        .C2(n738), .ZN(n4256) );
  AOI221_X1 U3492 ( .B1(n456), .B2(\REGISTERS[45][15] ), .C1(n453), .C2(
        \REGISTERS[44][15] ), .A(n5649), .ZN(n5643) );
  OAI222_X1 U3493 ( .A1(n1600), .A2(n450), .B1(n1632), .B2(n447), .C1(n1568), 
        .C2(n444), .ZN(n5649) );
  AOI221_X1 U3494 ( .B1(n38), .B2(\REGISTERS[78][15] ), .C1(n35), .C2(
        \REGISTERS[77][15] ), .A(n5658), .ZN(n5652) );
  OAI222_X1 U3495 ( .A1(n2656), .A2(n32), .B1(n2688), .B2(n29), .C1(n2624), 
        .C2(n26), .ZN(n5658) );
  AOI221_X1 U3496 ( .B1(n1168), .B2(\REGISTERS[45][15] ), .C1(n1165), .C2(
        \REGISTERS[44][15] ), .A(n4206), .ZN(n4200) );
  OAI222_X1 U3497 ( .A1(n1600), .A2(n1162), .B1(n1632), .B2(n1159), .C1(n1568), 
        .C2(n1156), .ZN(n4206) );
  AOI221_X1 U3498 ( .B1(n750), .B2(\REGISTERS[78][15] ), .C1(n747), .C2(
        \REGISTERS[77][15] ), .A(n4215), .ZN(n4209) );
  OAI222_X1 U3499 ( .A1(n2656), .A2(n744), .B1(n2688), .B2(n741), .C1(n2624), 
        .C2(n738), .ZN(n4215) );
  AOI221_X1 U3500 ( .B1(n456), .B2(\REGISTERS[45][16] ), .C1(n453), .C2(
        \REGISTERS[44][16] ), .A(n5608), .ZN(n5602) );
  OAI222_X1 U3501 ( .A1(n1599), .A2(n450), .B1(n1631), .B2(n447), .C1(n1567), 
        .C2(n444), .ZN(n5608) );
  AOI221_X1 U3502 ( .B1(n38), .B2(\REGISTERS[78][16] ), .C1(n35), .C2(
        \REGISTERS[77][16] ), .A(n5617), .ZN(n5611) );
  OAI222_X1 U3503 ( .A1(n2655), .A2(n32), .B1(n2687), .B2(n29), .C1(n2623), 
        .C2(n26), .ZN(n5617) );
  AOI221_X1 U3504 ( .B1(n1168), .B2(\REGISTERS[45][16] ), .C1(n1165), .C2(
        \REGISTERS[44][16] ), .A(n4165), .ZN(n4159) );
  OAI222_X1 U3505 ( .A1(n1599), .A2(n1162), .B1(n1631), .B2(n1159), .C1(n1567), 
        .C2(n1156), .ZN(n4165) );
  AOI221_X1 U3506 ( .B1(n750), .B2(\REGISTERS[78][16] ), .C1(n747), .C2(
        \REGISTERS[77][16] ), .A(n4174), .ZN(n4168) );
  OAI222_X1 U3507 ( .A1(n2655), .A2(n744), .B1(n2687), .B2(n741), .C1(n2623), 
        .C2(n738), .ZN(n4174) );
  AOI221_X1 U3508 ( .B1(n456), .B2(\REGISTERS[45][17] ), .C1(n453), .C2(
        \REGISTERS[44][17] ), .A(n5567), .ZN(n5561) );
  OAI222_X1 U3509 ( .A1(n1598), .A2(n450), .B1(n1630), .B2(n447), .C1(n1566), 
        .C2(n444), .ZN(n5567) );
  AOI221_X1 U3510 ( .B1(n38), .B2(\REGISTERS[78][17] ), .C1(n35), .C2(
        \REGISTERS[77][17] ), .A(n5576), .ZN(n5570) );
  OAI222_X1 U3511 ( .A1(n2654), .A2(n32), .B1(n2686), .B2(n29), .C1(n2622), 
        .C2(n26), .ZN(n5576) );
  AOI221_X1 U3512 ( .B1(n1168), .B2(\REGISTERS[45][17] ), .C1(n1165), .C2(
        \REGISTERS[44][17] ), .A(n4124), .ZN(n4118) );
  OAI222_X1 U3513 ( .A1(n1598), .A2(n1162), .B1(n1630), .B2(n1159), .C1(n1566), 
        .C2(n1156), .ZN(n4124) );
  AOI221_X1 U3514 ( .B1(n750), .B2(\REGISTERS[78][17] ), .C1(n747), .C2(
        \REGISTERS[77][17] ), .A(n4133), .ZN(n4127) );
  OAI222_X1 U3515 ( .A1(n2654), .A2(n744), .B1(n2686), .B2(n741), .C1(n2622), 
        .C2(n738), .ZN(n4133) );
  AOI221_X1 U3516 ( .B1(n456), .B2(\REGISTERS[45][18] ), .C1(n453), .C2(
        \REGISTERS[44][18] ), .A(n5526), .ZN(n5520) );
  OAI222_X1 U3517 ( .A1(n1597), .A2(n450), .B1(n1629), .B2(n447), .C1(n1565), 
        .C2(n444), .ZN(n5526) );
  AOI221_X1 U3518 ( .B1(n38), .B2(\REGISTERS[78][18] ), .C1(n35), .C2(
        \REGISTERS[77][18] ), .A(n5535), .ZN(n5529) );
  OAI222_X1 U3519 ( .A1(n2653), .A2(n32), .B1(n2685), .B2(n29), .C1(n2621), 
        .C2(n26), .ZN(n5535) );
  AOI221_X1 U3520 ( .B1(n1168), .B2(\REGISTERS[45][18] ), .C1(n1165), .C2(
        \REGISTERS[44][18] ), .A(n4083), .ZN(n4077) );
  OAI222_X1 U3521 ( .A1(n1597), .A2(n1162), .B1(n1629), .B2(n1159), .C1(n1565), 
        .C2(n1156), .ZN(n4083) );
  AOI221_X1 U3522 ( .B1(n750), .B2(\REGISTERS[78][18] ), .C1(n747), .C2(
        \REGISTERS[77][18] ), .A(n4092), .ZN(n4086) );
  OAI222_X1 U3523 ( .A1(n2653), .A2(n744), .B1(n2685), .B2(n741), .C1(n2621), 
        .C2(n738), .ZN(n4092) );
  AOI221_X1 U3524 ( .B1(n456), .B2(\REGISTERS[45][19] ), .C1(n453), .C2(
        \REGISTERS[44][19] ), .A(n5485), .ZN(n5479) );
  OAI222_X1 U3525 ( .A1(n1596), .A2(n450), .B1(n1628), .B2(n447), .C1(n1564), 
        .C2(n444), .ZN(n5485) );
  AOI221_X1 U3526 ( .B1(n38), .B2(\REGISTERS[78][19] ), .C1(n35), .C2(
        \REGISTERS[77][19] ), .A(n5494), .ZN(n5488) );
  OAI222_X1 U3527 ( .A1(n2652), .A2(n32), .B1(n2684), .B2(n29), .C1(n2620), 
        .C2(n26), .ZN(n5494) );
  AOI221_X1 U3528 ( .B1(n1168), .B2(\REGISTERS[45][19] ), .C1(n1165), .C2(
        \REGISTERS[44][19] ), .A(n4042), .ZN(n4036) );
  OAI222_X1 U3529 ( .A1(n1596), .A2(n1162), .B1(n1628), .B2(n1159), .C1(n1564), 
        .C2(n1156), .ZN(n4042) );
  AOI221_X1 U3530 ( .B1(n750), .B2(\REGISTERS[78][19] ), .C1(n747), .C2(
        \REGISTERS[77][19] ), .A(n4051), .ZN(n4045) );
  OAI222_X1 U3531 ( .A1(n2652), .A2(n744), .B1(n2684), .B2(n741), .C1(n2620), 
        .C2(n738), .ZN(n4051) );
  AOI221_X1 U3532 ( .B1(n456), .B2(\REGISTERS[45][20] ), .C1(n453), .C2(
        \REGISTERS[44][20] ), .A(n5444), .ZN(n5438) );
  OAI222_X1 U3533 ( .A1(n1595), .A2(n450), .B1(n1627), .B2(n447), .C1(n1563), 
        .C2(n444), .ZN(n5444) );
  AOI221_X1 U3534 ( .B1(n38), .B2(\REGISTERS[78][20] ), .C1(n35), .C2(
        \REGISTERS[77][20] ), .A(n5453), .ZN(n5447) );
  OAI222_X1 U3535 ( .A1(n2651), .A2(n32), .B1(n2683), .B2(n29), .C1(n2619), 
        .C2(n26), .ZN(n5453) );
  AOI221_X1 U3536 ( .B1(n1168), .B2(\REGISTERS[45][20] ), .C1(n1165), .C2(
        \REGISTERS[44][20] ), .A(n4001), .ZN(n3995) );
  OAI222_X1 U3537 ( .A1(n1595), .A2(n1162), .B1(n1627), .B2(n1159), .C1(n1563), 
        .C2(n1156), .ZN(n4001) );
  AOI221_X1 U3538 ( .B1(n750), .B2(\REGISTERS[78][20] ), .C1(n747), .C2(
        \REGISTERS[77][20] ), .A(n4010), .ZN(n4004) );
  OAI222_X1 U3539 ( .A1(n2651), .A2(n744), .B1(n2683), .B2(n741), .C1(n2619), 
        .C2(n738), .ZN(n4010) );
  AOI221_X1 U3540 ( .B1(n456), .B2(\REGISTERS[45][21] ), .C1(n453), .C2(
        \REGISTERS[44][21] ), .A(n5403), .ZN(n5397) );
  OAI222_X1 U3541 ( .A1(n1594), .A2(n450), .B1(n1626), .B2(n447), .C1(n1562), 
        .C2(n444), .ZN(n5403) );
  AOI221_X1 U3542 ( .B1(n38), .B2(\REGISTERS[78][21] ), .C1(n35), .C2(
        \REGISTERS[77][21] ), .A(n5412), .ZN(n5406) );
  OAI222_X1 U3543 ( .A1(n2650), .A2(n32), .B1(n2682), .B2(n29), .C1(n2618), 
        .C2(n26), .ZN(n5412) );
  AOI221_X1 U3544 ( .B1(n1168), .B2(\REGISTERS[45][21] ), .C1(n1165), .C2(
        \REGISTERS[44][21] ), .A(n3960), .ZN(n3954) );
  OAI222_X1 U3545 ( .A1(n1594), .A2(n1162), .B1(n1626), .B2(n1159), .C1(n1562), 
        .C2(n1156), .ZN(n3960) );
  AOI221_X1 U3546 ( .B1(n750), .B2(\REGISTERS[78][21] ), .C1(n747), .C2(
        \REGISTERS[77][21] ), .A(n3969), .ZN(n3963) );
  OAI222_X1 U3547 ( .A1(n2650), .A2(n744), .B1(n2682), .B2(n741), .C1(n2618), 
        .C2(n738), .ZN(n3969) );
  AOI221_X1 U3548 ( .B1(n456), .B2(\REGISTERS[45][22] ), .C1(n453), .C2(
        \REGISTERS[44][22] ), .A(n5362), .ZN(n5356) );
  OAI222_X1 U3549 ( .A1(n1593), .A2(n450), .B1(n1625), .B2(n447), .C1(n1561), 
        .C2(n444), .ZN(n5362) );
  AOI221_X1 U3550 ( .B1(n38), .B2(\REGISTERS[78][22] ), .C1(n35), .C2(
        \REGISTERS[77][22] ), .A(n5371), .ZN(n5365) );
  OAI222_X1 U3551 ( .A1(n2649), .A2(n32), .B1(n2681), .B2(n29), .C1(n2617), 
        .C2(n26), .ZN(n5371) );
  AOI221_X1 U3552 ( .B1(n1168), .B2(\REGISTERS[45][22] ), .C1(n1165), .C2(
        \REGISTERS[44][22] ), .A(n3919), .ZN(n3913) );
  OAI222_X1 U3553 ( .A1(n1593), .A2(n1162), .B1(n1625), .B2(n1159), .C1(n1561), 
        .C2(n1156), .ZN(n3919) );
  AOI221_X1 U3554 ( .B1(n750), .B2(\REGISTERS[78][22] ), .C1(n747), .C2(
        \REGISTERS[77][22] ), .A(n3928), .ZN(n3922) );
  OAI222_X1 U3555 ( .A1(n2649), .A2(n744), .B1(n2681), .B2(n741), .C1(n2617), 
        .C2(n738), .ZN(n3928) );
  AOI221_X1 U3556 ( .B1(n456), .B2(\REGISTERS[45][23] ), .C1(n453), .C2(
        \REGISTERS[44][23] ), .A(n5321), .ZN(n5315) );
  OAI222_X1 U3557 ( .A1(n1592), .A2(n450), .B1(n1624), .B2(n447), .C1(n1560), 
        .C2(n444), .ZN(n5321) );
  AOI221_X1 U3558 ( .B1(n38), .B2(\REGISTERS[78][23] ), .C1(n35), .C2(
        \REGISTERS[77][23] ), .A(n5330), .ZN(n5324) );
  OAI222_X1 U3559 ( .A1(n2648), .A2(n32), .B1(n2680), .B2(n29), .C1(n2616), 
        .C2(n26), .ZN(n5330) );
  AOI221_X1 U3560 ( .B1(n1168), .B2(\REGISTERS[45][23] ), .C1(n1165), .C2(
        \REGISTERS[44][23] ), .A(n3878), .ZN(n3872) );
  OAI222_X1 U3561 ( .A1(n1592), .A2(n1162), .B1(n1624), .B2(n1159), .C1(n1560), 
        .C2(n1156), .ZN(n3878) );
  AOI221_X1 U3562 ( .B1(n750), .B2(\REGISTERS[78][23] ), .C1(n747), .C2(
        \REGISTERS[77][23] ), .A(n3887), .ZN(n3881) );
  OAI222_X1 U3563 ( .A1(n2648), .A2(n744), .B1(n2680), .B2(n741), .C1(n2616), 
        .C2(n738), .ZN(n3887) );
  AOI221_X1 U3564 ( .B1(n457), .B2(\REGISTERS[45][24] ), .C1(n454), .C2(
        \REGISTERS[44][24] ), .A(n5280), .ZN(n5274) );
  OAI222_X1 U3565 ( .A1(n1591), .A2(n451), .B1(n1623), .B2(n448), .C1(n1559), 
        .C2(n445), .ZN(n5280) );
  AOI221_X1 U3566 ( .B1(n39), .B2(\REGISTERS[78][24] ), .C1(n36), .C2(
        \REGISTERS[77][24] ), .A(n5289), .ZN(n5283) );
  OAI222_X1 U3567 ( .A1(n2647), .A2(n33), .B1(n2679), .B2(n30), .C1(n2615), 
        .C2(n27), .ZN(n5289) );
  AOI221_X1 U3568 ( .B1(n1169), .B2(\REGISTERS[45][24] ), .C1(n1166), .C2(
        \REGISTERS[44][24] ), .A(n3837), .ZN(n3831) );
  OAI222_X1 U3569 ( .A1(n1591), .A2(n1163), .B1(n1623), .B2(n1160), .C1(n1559), 
        .C2(n1157), .ZN(n3837) );
  AOI221_X1 U3570 ( .B1(n751), .B2(\REGISTERS[78][24] ), .C1(n748), .C2(
        \REGISTERS[77][24] ), .A(n3846), .ZN(n3840) );
  OAI222_X1 U3571 ( .A1(n2647), .A2(n745), .B1(n2679), .B2(n742), .C1(n2615), 
        .C2(n739), .ZN(n3846) );
  AOI221_X1 U3572 ( .B1(n457), .B2(\REGISTERS[45][25] ), .C1(n454), .C2(
        \REGISTERS[44][25] ), .A(n5239), .ZN(n5233) );
  OAI222_X1 U3573 ( .A1(n1590), .A2(n451), .B1(n1622), .B2(n448), .C1(n1558), 
        .C2(n445), .ZN(n5239) );
  AOI221_X1 U3574 ( .B1(n39), .B2(\REGISTERS[78][25] ), .C1(n36), .C2(
        \REGISTERS[77][25] ), .A(n5248), .ZN(n5242) );
  OAI222_X1 U3575 ( .A1(n2646), .A2(n33), .B1(n2678), .B2(n30), .C1(n2614), 
        .C2(n27), .ZN(n5248) );
  AOI221_X1 U3576 ( .B1(n1169), .B2(\REGISTERS[45][25] ), .C1(n1166), .C2(
        \REGISTERS[44][25] ), .A(n3796), .ZN(n3790) );
  OAI222_X1 U3577 ( .A1(n1590), .A2(n1163), .B1(n1622), .B2(n1160), .C1(n1558), 
        .C2(n1157), .ZN(n3796) );
  AOI221_X1 U3578 ( .B1(n751), .B2(\REGISTERS[78][25] ), .C1(n748), .C2(
        \REGISTERS[77][25] ), .A(n3805), .ZN(n3799) );
  OAI222_X1 U3579 ( .A1(n2646), .A2(n745), .B1(n2678), .B2(n742), .C1(n2614), 
        .C2(n739), .ZN(n3805) );
  AOI221_X1 U3580 ( .B1(n457), .B2(\REGISTERS[45][26] ), .C1(n454), .C2(
        \REGISTERS[44][26] ), .A(n5198), .ZN(n5192) );
  OAI222_X1 U3581 ( .A1(n1589), .A2(n451), .B1(n1621), .B2(n448), .C1(n1557), 
        .C2(n445), .ZN(n5198) );
  AOI221_X1 U3582 ( .B1(n39), .B2(\REGISTERS[78][26] ), .C1(n36), .C2(
        \REGISTERS[77][26] ), .A(n5207), .ZN(n5201) );
  OAI222_X1 U3583 ( .A1(n2645), .A2(n33), .B1(n2677), .B2(n30), .C1(n2613), 
        .C2(n27), .ZN(n5207) );
  AOI221_X1 U3584 ( .B1(n1169), .B2(\REGISTERS[45][26] ), .C1(n1166), .C2(
        \REGISTERS[44][26] ), .A(n3755), .ZN(n3749) );
  OAI222_X1 U3585 ( .A1(n1589), .A2(n1163), .B1(n1621), .B2(n1160), .C1(n1557), 
        .C2(n1157), .ZN(n3755) );
  AOI221_X1 U3586 ( .B1(n751), .B2(\REGISTERS[78][26] ), .C1(n748), .C2(
        \REGISTERS[77][26] ), .A(n3764), .ZN(n3758) );
  OAI222_X1 U3587 ( .A1(n2645), .A2(n745), .B1(n2677), .B2(n742), .C1(n2613), 
        .C2(n739), .ZN(n3764) );
  AOI221_X1 U3588 ( .B1(n457), .B2(\REGISTERS[45][27] ), .C1(n454), .C2(
        \REGISTERS[44][27] ), .A(n5157), .ZN(n5151) );
  OAI222_X1 U3589 ( .A1(n1588), .A2(n451), .B1(n1620), .B2(n448), .C1(n1556), 
        .C2(n445), .ZN(n5157) );
  AOI221_X1 U3590 ( .B1(n39), .B2(\REGISTERS[78][27] ), .C1(n36), .C2(
        \REGISTERS[77][27] ), .A(n5166), .ZN(n5160) );
  OAI222_X1 U3591 ( .A1(n2644), .A2(n33), .B1(n2676), .B2(n30), .C1(n2612), 
        .C2(n27), .ZN(n5166) );
  AOI221_X1 U3592 ( .B1(n1169), .B2(\REGISTERS[45][27] ), .C1(n1166), .C2(
        \REGISTERS[44][27] ), .A(n3714), .ZN(n3708) );
  OAI222_X1 U3593 ( .A1(n1588), .A2(n1163), .B1(n1620), .B2(n1160), .C1(n1556), 
        .C2(n1157), .ZN(n3714) );
  AOI221_X1 U3594 ( .B1(n751), .B2(\REGISTERS[78][27] ), .C1(n748), .C2(
        \REGISTERS[77][27] ), .A(n3723), .ZN(n3717) );
  OAI222_X1 U3595 ( .A1(n2644), .A2(n745), .B1(n2676), .B2(n742), .C1(n2612), 
        .C2(n739), .ZN(n3723) );
  AOI221_X1 U3596 ( .B1(n457), .B2(\REGISTERS[45][28] ), .C1(n454), .C2(
        \REGISTERS[44][28] ), .A(n5116), .ZN(n5110) );
  OAI222_X1 U3597 ( .A1(n1587), .A2(n451), .B1(n1619), .B2(n448), .C1(n1555), 
        .C2(n445), .ZN(n5116) );
  AOI221_X1 U3598 ( .B1(n39), .B2(\REGISTERS[78][28] ), .C1(n36), .C2(
        \REGISTERS[77][28] ), .A(n5125), .ZN(n5119) );
  OAI222_X1 U3599 ( .A1(n2643), .A2(n33), .B1(n2675), .B2(n30), .C1(n2611), 
        .C2(n27), .ZN(n5125) );
  AOI221_X1 U3600 ( .B1(n1169), .B2(\REGISTERS[45][28] ), .C1(n1166), .C2(
        \REGISTERS[44][28] ), .A(n3673), .ZN(n3667) );
  OAI222_X1 U3601 ( .A1(n1587), .A2(n1163), .B1(n1619), .B2(n1160), .C1(n1555), 
        .C2(n1157), .ZN(n3673) );
  AOI221_X1 U3602 ( .B1(n751), .B2(\REGISTERS[78][28] ), .C1(n748), .C2(
        \REGISTERS[77][28] ), .A(n3682), .ZN(n3676) );
  OAI222_X1 U3603 ( .A1(n2643), .A2(n745), .B1(n2675), .B2(n742), .C1(n2611), 
        .C2(n739), .ZN(n3682) );
  AOI221_X1 U3604 ( .B1(n457), .B2(\REGISTERS[45][29] ), .C1(n454), .C2(
        \REGISTERS[44][29] ), .A(n5075), .ZN(n5069) );
  OAI222_X1 U3605 ( .A1(n1586), .A2(n451), .B1(n1618), .B2(n448), .C1(n1554), 
        .C2(n445), .ZN(n5075) );
  AOI221_X1 U3606 ( .B1(n39), .B2(\REGISTERS[78][29] ), .C1(n36), .C2(
        \REGISTERS[77][29] ), .A(n5084), .ZN(n5078) );
  OAI222_X1 U3607 ( .A1(n2642), .A2(n33), .B1(n2674), .B2(n30), .C1(n2610), 
        .C2(n27), .ZN(n5084) );
  AOI221_X1 U3608 ( .B1(n1169), .B2(\REGISTERS[45][29] ), .C1(n1166), .C2(
        \REGISTERS[44][29] ), .A(n3632), .ZN(n3626) );
  OAI222_X1 U3609 ( .A1(n1586), .A2(n1163), .B1(n1618), .B2(n1160), .C1(n1554), 
        .C2(n1157), .ZN(n3632) );
  AOI221_X1 U3610 ( .B1(n751), .B2(\REGISTERS[78][29] ), .C1(n748), .C2(
        \REGISTERS[77][29] ), .A(n3641), .ZN(n3635) );
  OAI222_X1 U3611 ( .A1(n2642), .A2(n745), .B1(n2674), .B2(n742), .C1(n2610), 
        .C2(n739), .ZN(n3641) );
  AOI221_X1 U3612 ( .B1(n457), .B2(\REGISTERS[45][30] ), .C1(n454), .C2(
        \REGISTERS[44][30] ), .A(n5034), .ZN(n5028) );
  OAI222_X1 U3613 ( .A1(n1585), .A2(n451), .B1(n1617), .B2(n448), .C1(n1553), 
        .C2(n445), .ZN(n5034) );
  AOI221_X1 U3614 ( .B1(n39), .B2(\REGISTERS[78][30] ), .C1(n36), .C2(
        \REGISTERS[77][30] ), .A(n5043), .ZN(n5037) );
  OAI222_X1 U3615 ( .A1(n2641), .A2(n33), .B1(n2673), .B2(n30), .C1(n2609), 
        .C2(n27), .ZN(n5043) );
  AOI221_X1 U3616 ( .B1(n1169), .B2(\REGISTERS[45][30] ), .C1(n1166), .C2(
        \REGISTERS[44][30] ), .A(n3591), .ZN(n3585) );
  OAI222_X1 U3617 ( .A1(n1585), .A2(n1163), .B1(n1617), .B2(n1160), .C1(n1553), 
        .C2(n1157), .ZN(n3591) );
  AOI221_X1 U3618 ( .B1(n751), .B2(\REGISTERS[78][30] ), .C1(n748), .C2(
        \REGISTERS[77][30] ), .A(n3600), .ZN(n3594) );
  OAI222_X1 U3619 ( .A1(n2641), .A2(n745), .B1(n2673), .B2(n742), .C1(n2609), 
        .C2(n739), .ZN(n3600) );
  AOI221_X1 U3620 ( .B1(n457), .B2(\REGISTERS[45][31] ), .C1(n454), .C2(
        \REGISTERS[44][31] ), .A(n4962), .ZN(n4943) );
  OAI222_X1 U3621 ( .A1(n1584), .A2(n451), .B1(n1616), .B2(n448), .C1(n1552), 
        .C2(n445), .ZN(n4962) );
  AOI221_X1 U3622 ( .B1(n39), .B2(\REGISTERS[78][31] ), .C1(n36), .C2(
        \REGISTERS[77][31] ), .A(n4993), .ZN(n4974) );
  OAI222_X1 U3623 ( .A1(n2640), .A2(n33), .B1(n2672), .B2(n30), .C1(n2608), 
        .C2(n27), .ZN(n4993) );
  AOI221_X1 U3624 ( .B1(n1169), .B2(\REGISTERS[45][31] ), .C1(n1166), .C2(
        \REGISTERS[44][31] ), .A(n3519), .ZN(n3500) );
  OAI222_X1 U3625 ( .A1(n1584), .A2(n1163), .B1(n1616), .B2(n1160), .C1(n1552), 
        .C2(n1157), .ZN(n3519) );
  AOI221_X1 U3626 ( .B1(n751), .B2(\REGISTERS[78][31] ), .C1(n748), .C2(
        \REGISTERS[77][31] ), .A(n3550), .ZN(n3531) );
  OAI222_X1 U3627 ( .A1(n2640), .A2(n745), .B1(n2672), .B2(n742), .C1(n2608), 
        .C2(n739), .ZN(n3550) );
  AND3_X1 U3628 ( .A1(WR), .A2(ENABLE), .A3(wr_signal), .ZN(n3106) );
  OAI22_X1 U3629 ( .A1(n87), .A2(n718), .B1(n119), .B2(n715), .ZN(n5261) );
  OAI22_X1 U3630 ( .A1(n791), .A2(n652), .B1(n823), .B2(n649), .ZN(n5270) );
  OAI22_X1 U3631 ( .A1(n87), .A2(n1430), .B1(n119), .B2(n1427), .ZN(n3818) );
  OAI22_X1 U3632 ( .A1(n791), .A2(n1364), .B1(n823), .B2(n1361), .ZN(n3827) );
  OAI22_X1 U3633 ( .A1(n86), .A2(n718), .B1(n118), .B2(n715), .ZN(n5220) );
  OAI22_X1 U3634 ( .A1(n790), .A2(n652), .B1(n822), .B2(n649), .ZN(n5229) );
  OAI22_X1 U3635 ( .A1(n86), .A2(n1430), .B1(n118), .B2(n1427), .ZN(n3777) );
  OAI22_X1 U3636 ( .A1(n790), .A2(n1364), .B1(n822), .B2(n1361), .ZN(n3786) );
  OAI22_X1 U3637 ( .A1(n85), .A2(n718), .B1(n117), .B2(n715), .ZN(n5179) );
  OAI22_X1 U3638 ( .A1(n789), .A2(n652), .B1(n821), .B2(n649), .ZN(n5188) );
  OAI22_X1 U3639 ( .A1(n85), .A2(n1430), .B1(n117), .B2(n1427), .ZN(n3736) );
  OAI22_X1 U3640 ( .A1(n789), .A2(n1364), .B1(n821), .B2(n1361), .ZN(n3745) );
  OAI22_X1 U3641 ( .A1(n84), .A2(n718), .B1(n116), .B2(n715), .ZN(n5138) );
  OAI22_X1 U3642 ( .A1(n788), .A2(n652), .B1(n820), .B2(n649), .ZN(n5147) );
  OAI22_X1 U3643 ( .A1(n84), .A2(n1430), .B1(n116), .B2(n1427), .ZN(n3695) );
  OAI22_X1 U3644 ( .A1(n788), .A2(n1364), .B1(n820), .B2(n1361), .ZN(n3704) );
  OAI22_X1 U3645 ( .A1(n83), .A2(n718), .B1(n115), .B2(n715), .ZN(n5097) );
  OAI22_X1 U3646 ( .A1(n787), .A2(n652), .B1(n819), .B2(n649), .ZN(n5106) );
  OAI22_X1 U3647 ( .A1(n83), .A2(n1430), .B1(n115), .B2(n1427), .ZN(n3654) );
  OAI22_X1 U3648 ( .A1(n787), .A2(n1364), .B1(n819), .B2(n1361), .ZN(n3663) );
  OAI22_X1 U3649 ( .A1(n82), .A2(n718), .B1(n114), .B2(n715), .ZN(n5056) );
  OAI22_X1 U3650 ( .A1(n786), .A2(n652), .B1(n818), .B2(n649), .ZN(n5065) );
  OAI22_X1 U3651 ( .A1(n82), .A2(n1430), .B1(n114), .B2(n1427), .ZN(n3613) );
  OAI22_X1 U3652 ( .A1(n786), .A2(n1364), .B1(n818), .B2(n1361), .ZN(n3622) );
  OAI22_X1 U3653 ( .A1(n81), .A2(n718), .B1(n113), .B2(n715), .ZN(n5015) );
  OAI22_X1 U3654 ( .A1(n785), .A2(n652), .B1(n817), .B2(n649), .ZN(n5024) );
  OAI22_X1 U3655 ( .A1(n81), .A2(n1430), .B1(n113), .B2(n1427), .ZN(n3572) );
  OAI22_X1 U3656 ( .A1(n785), .A2(n1364), .B1(n817), .B2(n1361), .ZN(n3581) );
  OAI22_X1 U3657 ( .A1(n80), .A2(n718), .B1(n112), .B2(n715), .ZN(n4886) );
  OAI22_X1 U3658 ( .A1(n784), .A2(n652), .B1(n816), .B2(n649), .ZN(n4917) );
  OAI22_X1 U3659 ( .A1(n80), .A2(n1430), .B1(n112), .B2(n1427), .ZN(n3443) );
  OAI22_X1 U3660 ( .A1(n784), .A2(n1364), .B1(n816), .B2(n1361), .ZN(n3474) );
  OAI22_X1 U3661 ( .A1(n111), .A2(n716), .B1(n143), .B2(n713), .ZN(n6245) );
  OAI22_X1 U3662 ( .A1(n815), .A2(n650), .B1(n847), .B2(n647), .ZN(n6276) );
  OAI22_X1 U3663 ( .A1(n111), .A2(n1428), .B1(n143), .B2(n1425), .ZN(n4802) );
  OAI22_X1 U3664 ( .A1(n815), .A2(n1362), .B1(n847), .B2(n1359), .ZN(n4833) );
  OAI22_X1 U3665 ( .A1(n110), .A2(n716), .B1(n142), .B2(n713), .ZN(n6204) );
  OAI22_X1 U3666 ( .A1(n814), .A2(n650), .B1(n846), .B2(n647), .ZN(n6213) );
  OAI22_X1 U3667 ( .A1(n110), .A2(n1428), .B1(n142), .B2(n1425), .ZN(n4761) );
  OAI22_X1 U3668 ( .A1(n814), .A2(n1362), .B1(n846), .B2(n1359), .ZN(n4770) );
  OAI22_X1 U3669 ( .A1(n109), .A2(n716), .B1(n141), .B2(n713), .ZN(n6163) );
  OAI22_X1 U3670 ( .A1(n813), .A2(n650), .B1(n845), .B2(n647), .ZN(n6172) );
  OAI22_X1 U3671 ( .A1(n109), .A2(n1428), .B1(n141), .B2(n1425), .ZN(n4720) );
  OAI22_X1 U3672 ( .A1(n813), .A2(n1362), .B1(n845), .B2(n1359), .ZN(n4729) );
  OAI22_X1 U3673 ( .A1(n108), .A2(n716), .B1(n140), .B2(n713), .ZN(n6122) );
  OAI22_X1 U3674 ( .A1(n812), .A2(n650), .B1(n844), .B2(n647), .ZN(n6131) );
  OAI22_X1 U3675 ( .A1(n108), .A2(n1428), .B1(n140), .B2(n1425), .ZN(n4679) );
  OAI22_X1 U3676 ( .A1(n812), .A2(n1362), .B1(n844), .B2(n1359), .ZN(n4688) );
  OAI22_X1 U3677 ( .A1(n107), .A2(n716), .B1(n139), .B2(n713), .ZN(n6081) );
  OAI22_X1 U3678 ( .A1(n811), .A2(n650), .B1(n843), .B2(n647), .ZN(n6090) );
  OAI22_X1 U3679 ( .A1(n107), .A2(n1428), .B1(n139), .B2(n1425), .ZN(n4638) );
  OAI22_X1 U3680 ( .A1(n811), .A2(n1362), .B1(n843), .B2(n1359), .ZN(n4647) );
  OAI22_X1 U3681 ( .A1(n106), .A2(n716), .B1(n138), .B2(n713), .ZN(n6040) );
  OAI22_X1 U3682 ( .A1(n810), .A2(n650), .B1(n842), .B2(n647), .ZN(n6049) );
  OAI22_X1 U3683 ( .A1(n106), .A2(n1428), .B1(n138), .B2(n1425), .ZN(n4597) );
  OAI22_X1 U3684 ( .A1(n810), .A2(n1362), .B1(n842), .B2(n1359), .ZN(n4606) );
  OAI22_X1 U3685 ( .A1(n105), .A2(n716), .B1(n137), .B2(n713), .ZN(n5999) );
  OAI22_X1 U3686 ( .A1(n809), .A2(n650), .B1(n841), .B2(n647), .ZN(n6008) );
  OAI22_X1 U3687 ( .A1(n105), .A2(n1428), .B1(n137), .B2(n1425), .ZN(n4556) );
  OAI22_X1 U3688 ( .A1(n809), .A2(n1362), .B1(n841), .B2(n1359), .ZN(n4565) );
  OAI22_X1 U3689 ( .A1(n104), .A2(n716), .B1(n136), .B2(n713), .ZN(n5958) );
  OAI22_X1 U3690 ( .A1(n808), .A2(n650), .B1(n840), .B2(n647), .ZN(n5967) );
  OAI22_X1 U3691 ( .A1(n104), .A2(n1428), .B1(n136), .B2(n1425), .ZN(n4515) );
  OAI22_X1 U3692 ( .A1(n808), .A2(n1362), .B1(n840), .B2(n1359), .ZN(n4524) );
  OAI22_X1 U3693 ( .A1(n103), .A2(n716), .B1(n135), .B2(n713), .ZN(n5917) );
  OAI22_X1 U3694 ( .A1(n807), .A2(n650), .B1(n839), .B2(n647), .ZN(n5926) );
  OAI22_X1 U3695 ( .A1(n103), .A2(n1428), .B1(n135), .B2(n1425), .ZN(n4474) );
  OAI22_X1 U3696 ( .A1(n807), .A2(n1362), .B1(n839), .B2(n1359), .ZN(n4483) );
  OAI22_X1 U3697 ( .A1(n102), .A2(n716), .B1(n134), .B2(n713), .ZN(n5876) );
  OAI22_X1 U3698 ( .A1(n806), .A2(n650), .B1(n838), .B2(n647), .ZN(n5885) );
  OAI22_X1 U3699 ( .A1(n102), .A2(n1428), .B1(n134), .B2(n1425), .ZN(n4433) );
  OAI22_X1 U3700 ( .A1(n806), .A2(n1362), .B1(n838), .B2(n1359), .ZN(n4442) );
  OAI22_X1 U3701 ( .A1(n101), .A2(n716), .B1(n133), .B2(n713), .ZN(n5835) );
  OAI22_X1 U3702 ( .A1(n805), .A2(n650), .B1(n837), .B2(n647), .ZN(n5844) );
  OAI22_X1 U3703 ( .A1(n101), .A2(n1428), .B1(n133), .B2(n1425), .ZN(n4392) );
  OAI22_X1 U3704 ( .A1(n805), .A2(n1362), .B1(n837), .B2(n1359), .ZN(n4401) );
  OAI22_X1 U3705 ( .A1(n100), .A2(n716), .B1(n132), .B2(n713), .ZN(n5794) );
  OAI22_X1 U3706 ( .A1(n804), .A2(n650), .B1(n836), .B2(n647), .ZN(n5803) );
  OAI22_X1 U3707 ( .A1(n100), .A2(n1428), .B1(n132), .B2(n1425), .ZN(n4351) );
  OAI22_X1 U3708 ( .A1(n804), .A2(n1362), .B1(n836), .B2(n1359), .ZN(n4360) );
  OAI22_X1 U3709 ( .A1(n99), .A2(n717), .B1(n131), .B2(n714), .ZN(n5753) );
  OAI22_X1 U3710 ( .A1(n803), .A2(n651), .B1(n835), .B2(n648), .ZN(n5762) );
  OAI22_X1 U3711 ( .A1(n99), .A2(n1429), .B1(n131), .B2(n1426), .ZN(n4310) );
  OAI22_X1 U3712 ( .A1(n803), .A2(n1363), .B1(n835), .B2(n1360), .ZN(n4319) );
  OAI22_X1 U3713 ( .A1(n98), .A2(n717), .B1(n130), .B2(n714), .ZN(n5712) );
  OAI22_X1 U3714 ( .A1(n802), .A2(n651), .B1(n834), .B2(n648), .ZN(n5721) );
  OAI22_X1 U3715 ( .A1(n98), .A2(n1429), .B1(n130), .B2(n1426), .ZN(n4269) );
  OAI22_X1 U3716 ( .A1(n802), .A2(n1363), .B1(n834), .B2(n1360), .ZN(n4278) );
  OAI22_X1 U3717 ( .A1(n97), .A2(n717), .B1(n129), .B2(n714), .ZN(n5671) );
  OAI22_X1 U3718 ( .A1(n801), .A2(n651), .B1(n833), .B2(n648), .ZN(n5680) );
  OAI22_X1 U3719 ( .A1(n97), .A2(n1429), .B1(n129), .B2(n1426), .ZN(n4228) );
  OAI22_X1 U3720 ( .A1(n801), .A2(n1363), .B1(n833), .B2(n1360), .ZN(n4237) );
  OAI22_X1 U3721 ( .A1(n96), .A2(n717), .B1(n128), .B2(n714), .ZN(n5630) );
  OAI22_X1 U3722 ( .A1(n800), .A2(n651), .B1(n832), .B2(n648), .ZN(n5639) );
  OAI22_X1 U3723 ( .A1(n96), .A2(n1429), .B1(n128), .B2(n1426), .ZN(n4187) );
  OAI22_X1 U3724 ( .A1(n800), .A2(n1363), .B1(n832), .B2(n1360), .ZN(n4196) );
  OAI22_X1 U3725 ( .A1(n95), .A2(n717), .B1(n127), .B2(n714), .ZN(n5589) );
  OAI22_X1 U3726 ( .A1(n799), .A2(n651), .B1(n831), .B2(n648), .ZN(n5598) );
  OAI22_X1 U3727 ( .A1(n95), .A2(n1429), .B1(n127), .B2(n1426), .ZN(n4146) );
  OAI22_X1 U3728 ( .A1(n799), .A2(n1363), .B1(n831), .B2(n1360), .ZN(n4155) );
  OAI22_X1 U3729 ( .A1(n94), .A2(n717), .B1(n126), .B2(n714), .ZN(n5548) );
  OAI22_X1 U3730 ( .A1(n798), .A2(n651), .B1(n830), .B2(n648), .ZN(n5557) );
  OAI22_X1 U3731 ( .A1(n94), .A2(n1429), .B1(n126), .B2(n1426), .ZN(n4105) );
  OAI22_X1 U3732 ( .A1(n798), .A2(n1363), .B1(n830), .B2(n1360), .ZN(n4114) );
  OAI22_X1 U3733 ( .A1(n93), .A2(n717), .B1(n125), .B2(n714), .ZN(n5507) );
  OAI22_X1 U3734 ( .A1(n797), .A2(n651), .B1(n829), .B2(n648), .ZN(n5516) );
  OAI22_X1 U3735 ( .A1(n93), .A2(n1429), .B1(n125), .B2(n1426), .ZN(n4064) );
  OAI22_X1 U3736 ( .A1(n797), .A2(n1363), .B1(n829), .B2(n1360), .ZN(n4073) );
  OAI22_X1 U3737 ( .A1(n92), .A2(n717), .B1(n124), .B2(n714), .ZN(n5466) );
  OAI22_X1 U3738 ( .A1(n796), .A2(n651), .B1(n828), .B2(n648), .ZN(n5475) );
  OAI22_X1 U3739 ( .A1(n92), .A2(n1429), .B1(n124), .B2(n1426), .ZN(n4023) );
  OAI22_X1 U3740 ( .A1(n796), .A2(n1363), .B1(n828), .B2(n1360), .ZN(n4032) );
  OAI22_X1 U3741 ( .A1(n91), .A2(n717), .B1(n123), .B2(n714), .ZN(n5425) );
  OAI22_X1 U3742 ( .A1(n795), .A2(n651), .B1(n827), .B2(n648), .ZN(n5434) );
  OAI22_X1 U3743 ( .A1(n91), .A2(n1429), .B1(n123), .B2(n1426), .ZN(n3982) );
  OAI22_X1 U3744 ( .A1(n795), .A2(n1363), .B1(n827), .B2(n1360), .ZN(n3991) );
  OAI22_X1 U3745 ( .A1(n90), .A2(n717), .B1(n122), .B2(n714), .ZN(n5384) );
  OAI22_X1 U3746 ( .A1(n794), .A2(n651), .B1(n826), .B2(n648), .ZN(n5393) );
  OAI22_X1 U3747 ( .A1(n90), .A2(n1429), .B1(n122), .B2(n1426), .ZN(n3941) );
  OAI22_X1 U3748 ( .A1(n794), .A2(n1363), .B1(n826), .B2(n1360), .ZN(n3950) );
  OAI22_X1 U3749 ( .A1(n89), .A2(n717), .B1(n121), .B2(n714), .ZN(n5343) );
  OAI22_X1 U3750 ( .A1(n793), .A2(n651), .B1(n825), .B2(n648), .ZN(n5352) );
  OAI22_X1 U3751 ( .A1(n89), .A2(n1429), .B1(n121), .B2(n1426), .ZN(n3900) );
  OAI22_X1 U3752 ( .A1(n793), .A2(n1363), .B1(n825), .B2(n1360), .ZN(n3909) );
  OAI22_X1 U3753 ( .A1(n88), .A2(n717), .B1(n120), .B2(n714), .ZN(n5302) );
  OAI22_X1 U3754 ( .A1(n792), .A2(n651), .B1(n824), .B2(n648), .ZN(n5311) );
  OAI22_X1 U3755 ( .A1(n88), .A2(n1429), .B1(n120), .B2(n1426), .ZN(n3859) );
  OAI22_X1 U3756 ( .A1(n792), .A2(n1363), .B1(n824), .B2(n1360), .ZN(n3868) );
  NAND4_X1 U3757 ( .A1(n6238), .A2(n6239), .A3(n6240), .A4(n6241), .ZN(n6237)
         );
  AOI221_X1 U3758 ( .B1(n683), .B2(\REGISTERS[12][0] ), .C1(n680), .C2(
        \REGISTERS[11][0] ), .A(n6258), .ZN(n6240) );
  NOR4_X1 U3759 ( .A1(n6242), .A2(n6243), .A3(n6244), .A4(n6245), .ZN(n6241)
         );
  AOI222_X1 U3760 ( .A1(n659), .A2(\REGISTERS[16][0] ), .B1(n658), .B2(
        \REGISTERS[18][0] ), .C1(n655), .C2(\REGISTERS[17][0] ), .ZN(n6238) );
  NAND4_X1 U3761 ( .A1(n4795), .A2(n4796), .A3(n4797), .A4(n4798), .ZN(n4794)
         );
  AOI221_X1 U3762 ( .B1(n1395), .B2(\REGISTERS[12][0] ), .C1(n1392), .C2(
        \REGISTERS[11][0] ), .A(n4815), .ZN(n4797) );
  NOR4_X1 U3763 ( .A1(n4799), .A2(n4800), .A3(n4801), .A4(n4802), .ZN(n4798)
         );
  AOI222_X1 U3764 ( .A1(n1371), .A2(\REGISTERS[16][0] ), .B1(n1370), .B2(
        \REGISTERS[18][0] ), .C1(n1367), .C2(\REGISTERS[17][0] ), .ZN(n4795)
         );
  NAND4_X1 U3765 ( .A1(n6197), .A2(n6198), .A3(n6199), .A4(n6200), .ZN(n6196)
         );
  AOI221_X1 U3766 ( .B1(n683), .B2(\REGISTERS[12][1] ), .C1(n680), .C2(
        \REGISTERS[11][1] ), .A(n6205), .ZN(n6199) );
  NOR4_X1 U3767 ( .A1(n6201), .A2(n6202), .A3(n6203), .A4(n6204), .ZN(n6200)
         );
  AOI222_X1 U3768 ( .A1(n659), .A2(\REGISTERS[16][1] ), .B1(n658), .B2(
        \REGISTERS[18][1] ), .C1(n655), .C2(\REGISTERS[17][1] ), .ZN(n6197) );
  NAND4_X1 U3769 ( .A1(n4754), .A2(n4755), .A3(n4756), .A4(n4757), .ZN(n4753)
         );
  AOI221_X1 U3770 ( .B1(n1395), .B2(\REGISTERS[12][1] ), .C1(n1392), .C2(
        \REGISTERS[11][1] ), .A(n4762), .ZN(n4756) );
  NOR4_X1 U3771 ( .A1(n4758), .A2(n4759), .A3(n4760), .A4(n4761), .ZN(n4757)
         );
  AOI222_X1 U3772 ( .A1(n1371), .A2(\REGISTERS[16][1] ), .B1(n1370), .B2(
        \REGISTERS[18][1] ), .C1(n1367), .C2(\REGISTERS[17][1] ), .ZN(n4754)
         );
  NAND4_X1 U3773 ( .A1(n6156), .A2(n6157), .A3(n6158), .A4(n6159), .ZN(n6155)
         );
  AOI221_X1 U3774 ( .B1(n683), .B2(\REGISTERS[12][2] ), .C1(n680), .C2(
        \REGISTERS[11][2] ), .A(n6164), .ZN(n6158) );
  NOR4_X1 U3775 ( .A1(n6160), .A2(n6161), .A3(n6162), .A4(n6163), .ZN(n6159)
         );
  AOI222_X1 U3776 ( .A1(n659), .A2(\REGISTERS[16][2] ), .B1(n658), .B2(
        \REGISTERS[18][2] ), .C1(n655), .C2(\REGISTERS[17][2] ), .ZN(n6156) );
  NAND4_X1 U3777 ( .A1(n4713), .A2(n4714), .A3(n4715), .A4(n4716), .ZN(n4712)
         );
  AOI221_X1 U3778 ( .B1(n1395), .B2(\REGISTERS[12][2] ), .C1(n1392), .C2(
        \REGISTERS[11][2] ), .A(n4721), .ZN(n4715) );
  NOR4_X1 U3779 ( .A1(n4717), .A2(n4718), .A3(n4719), .A4(n4720), .ZN(n4716)
         );
  AOI222_X1 U3780 ( .A1(n1371), .A2(\REGISTERS[16][2] ), .B1(n1370), .B2(
        \REGISTERS[18][2] ), .C1(n1367), .C2(\REGISTERS[17][2] ), .ZN(n4713)
         );
  NAND4_X1 U3781 ( .A1(n6115), .A2(n6116), .A3(n6117), .A4(n6118), .ZN(n6114)
         );
  AOI221_X1 U3782 ( .B1(n683), .B2(\REGISTERS[12][3] ), .C1(n680), .C2(
        \REGISTERS[11][3] ), .A(n6123), .ZN(n6117) );
  NOR4_X1 U3783 ( .A1(n6119), .A2(n6120), .A3(n6121), .A4(n6122), .ZN(n6118)
         );
  AOI222_X1 U3784 ( .A1(n659), .A2(\REGISTERS[16][3] ), .B1(n658), .B2(
        \REGISTERS[18][3] ), .C1(n655), .C2(\REGISTERS[17][3] ), .ZN(n6115) );
  NAND4_X1 U3785 ( .A1(n4672), .A2(n4673), .A3(n4674), .A4(n4675), .ZN(n4671)
         );
  AOI221_X1 U3786 ( .B1(n1395), .B2(\REGISTERS[12][3] ), .C1(n1392), .C2(
        \REGISTERS[11][3] ), .A(n4680), .ZN(n4674) );
  NOR4_X1 U3787 ( .A1(n4676), .A2(n4677), .A3(n4678), .A4(n4679), .ZN(n4675)
         );
  AOI222_X1 U3788 ( .A1(n1371), .A2(\REGISTERS[16][3] ), .B1(n1370), .B2(
        \REGISTERS[18][3] ), .C1(n1367), .C2(\REGISTERS[17][3] ), .ZN(n4672)
         );
  NAND4_X1 U3789 ( .A1(n6074), .A2(n6075), .A3(n6076), .A4(n6077), .ZN(n6073)
         );
  AOI221_X1 U3790 ( .B1(n683), .B2(\REGISTERS[12][4] ), .C1(n680), .C2(
        \REGISTERS[11][4] ), .A(n6082), .ZN(n6076) );
  NOR4_X1 U3791 ( .A1(n6078), .A2(n6079), .A3(n6080), .A4(n6081), .ZN(n6077)
         );
  AOI222_X1 U3792 ( .A1(n659), .A2(\REGISTERS[16][4] ), .B1(n658), .B2(
        \REGISTERS[18][4] ), .C1(n655), .C2(\REGISTERS[17][4] ), .ZN(n6074) );
  NAND4_X1 U3793 ( .A1(n4631), .A2(n4632), .A3(n4633), .A4(n4634), .ZN(n4630)
         );
  AOI221_X1 U3794 ( .B1(n1395), .B2(\REGISTERS[12][4] ), .C1(n1392), .C2(
        \REGISTERS[11][4] ), .A(n4639), .ZN(n4633) );
  NOR4_X1 U3795 ( .A1(n4635), .A2(n4636), .A3(n4637), .A4(n4638), .ZN(n4634)
         );
  AOI222_X1 U3796 ( .A1(n1371), .A2(\REGISTERS[16][4] ), .B1(n1370), .B2(
        \REGISTERS[18][4] ), .C1(n1367), .C2(\REGISTERS[17][4] ), .ZN(n4631)
         );
  NAND4_X1 U3797 ( .A1(n6033), .A2(n6034), .A3(n6035), .A4(n6036), .ZN(n6032)
         );
  AOI221_X1 U3798 ( .B1(n683), .B2(\REGISTERS[12][5] ), .C1(n680), .C2(
        \REGISTERS[11][5] ), .A(n6041), .ZN(n6035) );
  NOR4_X1 U3799 ( .A1(n6037), .A2(n6038), .A3(n6039), .A4(n6040), .ZN(n6036)
         );
  AOI222_X1 U3800 ( .A1(n659), .A2(\REGISTERS[16][5] ), .B1(n658), .B2(
        \REGISTERS[18][5] ), .C1(n655), .C2(\REGISTERS[17][5] ), .ZN(n6033) );
  NAND4_X1 U3801 ( .A1(n4590), .A2(n4591), .A3(n4592), .A4(n4593), .ZN(n4589)
         );
  AOI221_X1 U3802 ( .B1(n1395), .B2(\REGISTERS[12][5] ), .C1(n1392), .C2(
        \REGISTERS[11][5] ), .A(n4598), .ZN(n4592) );
  NOR4_X1 U3803 ( .A1(n4594), .A2(n4595), .A3(n4596), .A4(n4597), .ZN(n4593)
         );
  AOI222_X1 U3804 ( .A1(n1371), .A2(\REGISTERS[16][5] ), .B1(n1370), .B2(
        \REGISTERS[18][5] ), .C1(n1367), .C2(\REGISTERS[17][5] ), .ZN(n4590)
         );
  NAND4_X1 U3805 ( .A1(n5992), .A2(n5993), .A3(n5994), .A4(n5995), .ZN(n5991)
         );
  AOI221_X1 U3806 ( .B1(n683), .B2(\REGISTERS[12][6] ), .C1(n680), .C2(
        \REGISTERS[11][6] ), .A(n6000), .ZN(n5994) );
  NOR4_X1 U3807 ( .A1(n5996), .A2(n5997), .A3(n5998), .A4(n5999), .ZN(n5995)
         );
  AOI222_X1 U3808 ( .A1(n659), .A2(\REGISTERS[16][6] ), .B1(n658), .B2(
        \REGISTERS[18][6] ), .C1(n655), .C2(\REGISTERS[17][6] ), .ZN(n5992) );
  NAND4_X1 U3809 ( .A1(n4549), .A2(n4550), .A3(n4551), .A4(n4552), .ZN(n4548)
         );
  AOI221_X1 U3810 ( .B1(n1395), .B2(\REGISTERS[12][6] ), .C1(n1392), .C2(
        \REGISTERS[11][6] ), .A(n4557), .ZN(n4551) );
  NOR4_X1 U3811 ( .A1(n4553), .A2(n4554), .A3(n4555), .A4(n4556), .ZN(n4552)
         );
  AOI222_X1 U3812 ( .A1(n1371), .A2(\REGISTERS[16][6] ), .B1(n1370), .B2(
        \REGISTERS[18][6] ), .C1(n1367), .C2(\REGISTERS[17][6] ), .ZN(n4549)
         );
  NAND4_X1 U3813 ( .A1(n5951), .A2(n5952), .A3(n5953), .A4(n5954), .ZN(n5950)
         );
  AOI221_X1 U3814 ( .B1(n683), .B2(\REGISTERS[12][7] ), .C1(n680), .C2(
        \REGISTERS[11][7] ), .A(n5959), .ZN(n5953) );
  NOR4_X1 U3815 ( .A1(n5955), .A2(n5956), .A3(n5957), .A4(n5958), .ZN(n5954)
         );
  AOI222_X1 U3816 ( .A1(n659), .A2(\REGISTERS[16][7] ), .B1(n658), .B2(
        \REGISTERS[18][7] ), .C1(n655), .C2(\REGISTERS[17][7] ), .ZN(n5951) );
  NAND4_X1 U3817 ( .A1(n4508), .A2(n4509), .A3(n4510), .A4(n4511), .ZN(n4507)
         );
  AOI221_X1 U3818 ( .B1(n1395), .B2(\REGISTERS[12][7] ), .C1(n1392), .C2(
        \REGISTERS[11][7] ), .A(n4516), .ZN(n4510) );
  NOR4_X1 U3819 ( .A1(n4512), .A2(n4513), .A3(n4514), .A4(n4515), .ZN(n4511)
         );
  AOI222_X1 U3820 ( .A1(n1371), .A2(\REGISTERS[16][7] ), .B1(n1370), .B2(
        \REGISTERS[18][7] ), .C1(n1367), .C2(\REGISTERS[17][7] ), .ZN(n4508)
         );
  NAND4_X1 U3821 ( .A1(n5910), .A2(n5911), .A3(n5912), .A4(n5913), .ZN(n5909)
         );
  AOI221_X1 U3822 ( .B1(n683), .B2(\REGISTERS[12][8] ), .C1(n680), .C2(
        \REGISTERS[11][8] ), .A(n5918), .ZN(n5912) );
  NOR4_X1 U3823 ( .A1(n5914), .A2(n5915), .A3(n5916), .A4(n5917), .ZN(n5913)
         );
  AOI222_X1 U3824 ( .A1(n659), .A2(\REGISTERS[16][8] ), .B1(n657), .B2(
        \REGISTERS[18][8] ), .C1(n654), .C2(\REGISTERS[17][8] ), .ZN(n5910) );
  NAND4_X1 U3825 ( .A1(n4467), .A2(n4468), .A3(n4469), .A4(n4470), .ZN(n4466)
         );
  AOI221_X1 U3826 ( .B1(n1395), .B2(\REGISTERS[12][8] ), .C1(n1392), .C2(
        \REGISTERS[11][8] ), .A(n4475), .ZN(n4469) );
  NOR4_X1 U3827 ( .A1(n4471), .A2(n4472), .A3(n4473), .A4(n4474), .ZN(n4470)
         );
  AOI222_X1 U3828 ( .A1(n1371), .A2(\REGISTERS[16][8] ), .B1(n1369), .B2(
        \REGISTERS[18][8] ), .C1(n1366), .C2(\REGISTERS[17][8] ), .ZN(n4467)
         );
  NAND4_X1 U3829 ( .A1(n5869), .A2(n5870), .A3(n5871), .A4(n5872), .ZN(n5868)
         );
  AOI221_X1 U3830 ( .B1(n683), .B2(\REGISTERS[12][9] ), .C1(n680), .C2(
        \REGISTERS[11][9] ), .A(n5877), .ZN(n5871) );
  NOR4_X1 U3831 ( .A1(n5873), .A2(n5874), .A3(n5875), .A4(n5876), .ZN(n5872)
         );
  AOI222_X1 U3832 ( .A1(n659), .A2(\REGISTERS[16][9] ), .B1(n657), .B2(
        \REGISTERS[18][9] ), .C1(n654), .C2(\REGISTERS[17][9] ), .ZN(n5869) );
  NAND4_X1 U3833 ( .A1(n4426), .A2(n4427), .A3(n4428), .A4(n4429), .ZN(n4425)
         );
  AOI221_X1 U3834 ( .B1(n1395), .B2(\REGISTERS[12][9] ), .C1(n1392), .C2(
        \REGISTERS[11][9] ), .A(n4434), .ZN(n4428) );
  NOR4_X1 U3835 ( .A1(n4430), .A2(n4431), .A3(n4432), .A4(n4433), .ZN(n4429)
         );
  AOI222_X1 U3836 ( .A1(n1371), .A2(\REGISTERS[16][9] ), .B1(n1369), .B2(
        \REGISTERS[18][9] ), .C1(n1366), .C2(\REGISTERS[17][9] ), .ZN(n4426)
         );
  NAND4_X1 U3837 ( .A1(n5828), .A2(n5829), .A3(n5830), .A4(n5831), .ZN(n5827)
         );
  AOI221_X1 U3838 ( .B1(n683), .B2(\REGISTERS[12][10] ), .C1(n680), .C2(
        \REGISTERS[11][10] ), .A(n5836), .ZN(n5830) );
  NOR4_X1 U3839 ( .A1(n5832), .A2(n5833), .A3(n5834), .A4(n5835), .ZN(n5831)
         );
  AOI222_X1 U3840 ( .A1(n659), .A2(\REGISTERS[16][10] ), .B1(n657), .B2(
        \REGISTERS[18][10] ), .C1(n654), .C2(\REGISTERS[17][10] ), .ZN(n5828)
         );
  NAND4_X1 U3841 ( .A1(n4385), .A2(n4386), .A3(n4387), .A4(n4388), .ZN(n4384)
         );
  AOI221_X1 U3842 ( .B1(n1395), .B2(\REGISTERS[12][10] ), .C1(n1392), .C2(
        \REGISTERS[11][10] ), .A(n4393), .ZN(n4387) );
  NOR4_X1 U3843 ( .A1(n4389), .A2(n4390), .A3(n4391), .A4(n4392), .ZN(n4388)
         );
  AOI222_X1 U3844 ( .A1(n1371), .A2(\REGISTERS[16][10] ), .B1(n1369), .B2(
        \REGISTERS[18][10] ), .C1(n1366), .C2(\REGISTERS[17][10] ), .ZN(n4385)
         );
  NAND4_X1 U3845 ( .A1(n5787), .A2(n5788), .A3(n5789), .A4(n5790), .ZN(n5786)
         );
  AOI221_X1 U3846 ( .B1(n683), .B2(\REGISTERS[12][11] ), .C1(n680), .C2(
        \REGISTERS[11][11] ), .A(n5795), .ZN(n5789) );
  NOR4_X1 U3847 ( .A1(n5791), .A2(n5792), .A3(n5793), .A4(n5794), .ZN(n5790)
         );
  AOI222_X1 U3848 ( .A1(n659), .A2(\REGISTERS[16][11] ), .B1(n657), .B2(
        \REGISTERS[18][11] ), .C1(n654), .C2(\REGISTERS[17][11] ), .ZN(n5787)
         );
  NAND4_X1 U3849 ( .A1(n4344), .A2(n4345), .A3(n4346), .A4(n4347), .ZN(n4343)
         );
  AOI221_X1 U3850 ( .B1(n1395), .B2(\REGISTERS[12][11] ), .C1(n1392), .C2(
        \REGISTERS[11][11] ), .A(n4352), .ZN(n4346) );
  NOR4_X1 U3851 ( .A1(n4348), .A2(n4349), .A3(n4350), .A4(n4351), .ZN(n4347)
         );
  AOI222_X1 U3852 ( .A1(n1371), .A2(\REGISTERS[16][11] ), .B1(n1369), .B2(
        \REGISTERS[18][11] ), .C1(n1366), .C2(\REGISTERS[17][11] ), .ZN(n4344)
         );
  NAND4_X1 U3853 ( .A1(n5746), .A2(n5747), .A3(n5748), .A4(n5749), .ZN(n5745)
         );
  AOI221_X1 U3854 ( .B1(n684), .B2(\REGISTERS[12][12] ), .C1(n681), .C2(
        \REGISTERS[11][12] ), .A(n5754), .ZN(n5748) );
  NOR4_X1 U3855 ( .A1(n5750), .A2(n5751), .A3(n5752), .A4(n5753), .ZN(n5749)
         );
  AOI222_X1 U3856 ( .A1(n660), .A2(\REGISTERS[16][12] ), .B1(n657), .B2(
        \REGISTERS[18][12] ), .C1(n654), .C2(\REGISTERS[17][12] ), .ZN(n5746)
         );
  NAND4_X1 U3857 ( .A1(n4303), .A2(n4304), .A3(n4305), .A4(n4306), .ZN(n4302)
         );
  AOI221_X1 U3858 ( .B1(n1396), .B2(\REGISTERS[12][12] ), .C1(n1393), .C2(
        \REGISTERS[11][12] ), .A(n4311), .ZN(n4305) );
  NOR4_X1 U3859 ( .A1(n4307), .A2(n4308), .A3(n4309), .A4(n4310), .ZN(n4306)
         );
  AOI222_X1 U3860 ( .A1(n1372), .A2(\REGISTERS[16][12] ), .B1(n1369), .B2(
        \REGISTERS[18][12] ), .C1(n1366), .C2(\REGISTERS[17][12] ), .ZN(n4303)
         );
  NAND4_X1 U3861 ( .A1(n5705), .A2(n5706), .A3(n5707), .A4(n5708), .ZN(n5704)
         );
  AOI221_X1 U3862 ( .B1(n684), .B2(\REGISTERS[12][13] ), .C1(n681), .C2(
        \REGISTERS[11][13] ), .A(n5713), .ZN(n5707) );
  NOR4_X1 U3863 ( .A1(n5709), .A2(n5710), .A3(n5711), .A4(n5712), .ZN(n5708)
         );
  AOI222_X1 U3864 ( .A1(n660), .A2(\REGISTERS[16][13] ), .B1(n657), .B2(
        \REGISTERS[18][13] ), .C1(n654), .C2(\REGISTERS[17][13] ), .ZN(n5705)
         );
  NAND4_X1 U3865 ( .A1(n4262), .A2(n4263), .A3(n4264), .A4(n4265), .ZN(n4261)
         );
  AOI221_X1 U3866 ( .B1(n1396), .B2(\REGISTERS[12][13] ), .C1(n1393), .C2(
        \REGISTERS[11][13] ), .A(n4270), .ZN(n4264) );
  NOR4_X1 U3867 ( .A1(n4266), .A2(n4267), .A3(n4268), .A4(n4269), .ZN(n4265)
         );
  AOI222_X1 U3868 ( .A1(n1372), .A2(\REGISTERS[16][13] ), .B1(n1369), .B2(
        \REGISTERS[18][13] ), .C1(n1366), .C2(\REGISTERS[17][13] ), .ZN(n4262)
         );
  NAND4_X1 U3869 ( .A1(n5664), .A2(n5665), .A3(n5666), .A4(n5667), .ZN(n5663)
         );
  AOI221_X1 U3870 ( .B1(n684), .B2(\REGISTERS[12][14] ), .C1(n681), .C2(
        \REGISTERS[11][14] ), .A(n5672), .ZN(n5666) );
  NOR4_X1 U3871 ( .A1(n5668), .A2(n5669), .A3(n5670), .A4(n5671), .ZN(n5667)
         );
  AOI222_X1 U3872 ( .A1(n660), .A2(\REGISTERS[16][14] ), .B1(n657), .B2(
        \REGISTERS[18][14] ), .C1(n654), .C2(\REGISTERS[17][14] ), .ZN(n5664)
         );
  NAND4_X1 U3873 ( .A1(n4221), .A2(n4222), .A3(n4223), .A4(n4224), .ZN(n4220)
         );
  AOI221_X1 U3874 ( .B1(n1396), .B2(\REGISTERS[12][14] ), .C1(n1393), .C2(
        \REGISTERS[11][14] ), .A(n4229), .ZN(n4223) );
  NOR4_X1 U3875 ( .A1(n4225), .A2(n4226), .A3(n4227), .A4(n4228), .ZN(n4224)
         );
  AOI222_X1 U3876 ( .A1(n1372), .A2(\REGISTERS[16][14] ), .B1(n1369), .B2(
        \REGISTERS[18][14] ), .C1(n1366), .C2(\REGISTERS[17][14] ), .ZN(n4221)
         );
  NAND4_X1 U3877 ( .A1(n5623), .A2(n5624), .A3(n5625), .A4(n5626), .ZN(n5622)
         );
  AOI221_X1 U3878 ( .B1(n684), .B2(\REGISTERS[12][15] ), .C1(n681), .C2(
        \REGISTERS[11][15] ), .A(n5631), .ZN(n5625) );
  NOR4_X1 U3879 ( .A1(n5627), .A2(n5628), .A3(n5629), .A4(n5630), .ZN(n5626)
         );
  AOI222_X1 U3880 ( .A1(n660), .A2(\REGISTERS[16][15] ), .B1(n657), .B2(
        \REGISTERS[18][15] ), .C1(n654), .C2(\REGISTERS[17][15] ), .ZN(n5623)
         );
  NAND4_X1 U3881 ( .A1(n4180), .A2(n4181), .A3(n4182), .A4(n4183), .ZN(n4179)
         );
  AOI221_X1 U3882 ( .B1(n1396), .B2(\REGISTERS[12][15] ), .C1(n1393), .C2(
        \REGISTERS[11][15] ), .A(n4188), .ZN(n4182) );
  NOR4_X1 U3883 ( .A1(n4184), .A2(n4185), .A3(n4186), .A4(n4187), .ZN(n4183)
         );
  AOI222_X1 U3884 ( .A1(n1372), .A2(\REGISTERS[16][15] ), .B1(n1369), .B2(
        \REGISTERS[18][15] ), .C1(n1366), .C2(\REGISTERS[17][15] ), .ZN(n4180)
         );
  NAND4_X1 U3885 ( .A1(n5582), .A2(n5583), .A3(n5584), .A4(n5585), .ZN(n5581)
         );
  AOI221_X1 U3886 ( .B1(n684), .B2(\REGISTERS[12][16] ), .C1(n681), .C2(
        \REGISTERS[11][16] ), .A(n5590), .ZN(n5584) );
  NOR4_X1 U3887 ( .A1(n5586), .A2(n5587), .A3(n5588), .A4(n5589), .ZN(n5585)
         );
  AOI222_X1 U3888 ( .A1(n660), .A2(\REGISTERS[16][16] ), .B1(n657), .B2(
        \REGISTERS[18][16] ), .C1(n654), .C2(\REGISTERS[17][16] ), .ZN(n5582)
         );
  NAND4_X1 U3889 ( .A1(n4139), .A2(n4140), .A3(n4141), .A4(n4142), .ZN(n4138)
         );
  AOI221_X1 U3890 ( .B1(n1396), .B2(\REGISTERS[12][16] ), .C1(n1393), .C2(
        \REGISTERS[11][16] ), .A(n4147), .ZN(n4141) );
  NOR4_X1 U3891 ( .A1(n4143), .A2(n4144), .A3(n4145), .A4(n4146), .ZN(n4142)
         );
  AOI222_X1 U3892 ( .A1(n1372), .A2(\REGISTERS[16][16] ), .B1(n1369), .B2(
        \REGISTERS[18][16] ), .C1(n1366), .C2(\REGISTERS[17][16] ), .ZN(n4139)
         );
  NAND4_X1 U3893 ( .A1(n5541), .A2(n5542), .A3(n5543), .A4(n5544), .ZN(n5540)
         );
  AOI221_X1 U3894 ( .B1(n684), .B2(\REGISTERS[12][17] ), .C1(n681), .C2(
        \REGISTERS[11][17] ), .A(n5549), .ZN(n5543) );
  NOR4_X1 U3895 ( .A1(n5545), .A2(n5546), .A3(n5547), .A4(n5548), .ZN(n5544)
         );
  AOI222_X1 U3896 ( .A1(n660), .A2(\REGISTERS[16][17] ), .B1(n657), .B2(
        \REGISTERS[18][17] ), .C1(n654), .C2(\REGISTERS[17][17] ), .ZN(n5541)
         );
  NAND4_X1 U3897 ( .A1(n4098), .A2(n4099), .A3(n4100), .A4(n4101), .ZN(n4097)
         );
  AOI221_X1 U3898 ( .B1(n1396), .B2(\REGISTERS[12][17] ), .C1(n1393), .C2(
        \REGISTERS[11][17] ), .A(n4106), .ZN(n4100) );
  NOR4_X1 U3899 ( .A1(n4102), .A2(n4103), .A3(n4104), .A4(n4105), .ZN(n4101)
         );
  AOI222_X1 U3900 ( .A1(n1372), .A2(\REGISTERS[16][17] ), .B1(n1369), .B2(
        \REGISTERS[18][17] ), .C1(n1366), .C2(\REGISTERS[17][17] ), .ZN(n4098)
         );
  NAND4_X1 U3901 ( .A1(n5500), .A2(n5501), .A3(n5502), .A4(n5503), .ZN(n5499)
         );
  AOI221_X1 U3902 ( .B1(n684), .B2(\REGISTERS[12][18] ), .C1(n681), .C2(
        \REGISTERS[11][18] ), .A(n5508), .ZN(n5502) );
  NOR4_X1 U3903 ( .A1(n5504), .A2(n5505), .A3(n5506), .A4(n5507), .ZN(n5503)
         );
  AOI222_X1 U3904 ( .A1(n660), .A2(\REGISTERS[16][18] ), .B1(n657), .B2(
        \REGISTERS[18][18] ), .C1(n654), .C2(\REGISTERS[17][18] ), .ZN(n5500)
         );
  NAND4_X1 U3905 ( .A1(n4057), .A2(n4058), .A3(n4059), .A4(n4060), .ZN(n4056)
         );
  AOI221_X1 U3906 ( .B1(n1396), .B2(\REGISTERS[12][18] ), .C1(n1393), .C2(
        \REGISTERS[11][18] ), .A(n4065), .ZN(n4059) );
  NOR4_X1 U3907 ( .A1(n4061), .A2(n4062), .A3(n4063), .A4(n4064), .ZN(n4060)
         );
  AOI222_X1 U3908 ( .A1(n1372), .A2(\REGISTERS[16][18] ), .B1(n1369), .B2(
        \REGISTERS[18][18] ), .C1(n1366), .C2(\REGISTERS[17][18] ), .ZN(n4057)
         );
  NAND4_X1 U3909 ( .A1(n5459), .A2(n5460), .A3(n5461), .A4(n5462), .ZN(n5458)
         );
  AOI221_X1 U3910 ( .B1(n684), .B2(\REGISTERS[12][19] ), .C1(n681), .C2(
        \REGISTERS[11][19] ), .A(n5467), .ZN(n5461) );
  NOR4_X1 U3911 ( .A1(n5463), .A2(n5464), .A3(n5465), .A4(n5466), .ZN(n5462)
         );
  AOI222_X1 U3912 ( .A1(n660), .A2(\REGISTERS[16][19] ), .B1(n657), .B2(
        \REGISTERS[18][19] ), .C1(n654), .C2(\REGISTERS[17][19] ), .ZN(n5459)
         );
  NAND4_X1 U3913 ( .A1(n4016), .A2(n4017), .A3(n4018), .A4(n4019), .ZN(n4015)
         );
  AOI221_X1 U3914 ( .B1(n1396), .B2(\REGISTERS[12][19] ), .C1(n1393), .C2(
        \REGISTERS[11][19] ), .A(n4024), .ZN(n4018) );
  NOR4_X1 U3915 ( .A1(n4020), .A2(n4021), .A3(n4022), .A4(n4023), .ZN(n4019)
         );
  AOI222_X1 U3916 ( .A1(n1372), .A2(\REGISTERS[16][19] ), .B1(n1369), .B2(
        \REGISTERS[18][19] ), .C1(n1366), .C2(\REGISTERS[17][19] ), .ZN(n4016)
         );
  NAND4_X1 U3917 ( .A1(n5418), .A2(n5419), .A3(n5420), .A4(n5421), .ZN(n5417)
         );
  AOI221_X1 U3918 ( .B1(n684), .B2(\REGISTERS[12][20] ), .C1(n681), .C2(
        \REGISTERS[11][20] ), .A(n5426), .ZN(n5420) );
  NOR4_X1 U3919 ( .A1(n5422), .A2(n5423), .A3(n5424), .A4(n5425), .ZN(n5421)
         );
  AOI222_X1 U3920 ( .A1(n660), .A2(\REGISTERS[16][20] ), .B1(n656), .B2(
        \REGISTERS[18][20] ), .C1(n653), .C2(\REGISTERS[17][20] ), .ZN(n5418)
         );
  NAND4_X1 U3921 ( .A1(n3975), .A2(n3976), .A3(n3977), .A4(n3978), .ZN(n3974)
         );
  AOI221_X1 U3922 ( .B1(n1396), .B2(\REGISTERS[12][20] ), .C1(n1393), .C2(
        \REGISTERS[11][20] ), .A(n3983), .ZN(n3977) );
  NOR4_X1 U3923 ( .A1(n3979), .A2(n3980), .A3(n3981), .A4(n3982), .ZN(n3978)
         );
  AOI222_X1 U3924 ( .A1(n1372), .A2(\REGISTERS[16][20] ), .B1(n1368), .B2(
        \REGISTERS[18][20] ), .C1(n1365), .C2(\REGISTERS[17][20] ), .ZN(n3975)
         );
  NAND4_X1 U3925 ( .A1(n5377), .A2(n5378), .A3(n5379), .A4(n5380), .ZN(n5376)
         );
  AOI221_X1 U3926 ( .B1(n684), .B2(\REGISTERS[12][21] ), .C1(n681), .C2(
        \REGISTERS[11][21] ), .A(n5385), .ZN(n5379) );
  NOR4_X1 U3927 ( .A1(n5381), .A2(n5382), .A3(n5383), .A4(n5384), .ZN(n5380)
         );
  AOI222_X1 U3928 ( .A1(n660), .A2(\REGISTERS[16][21] ), .B1(n656), .B2(
        \REGISTERS[18][21] ), .C1(n653), .C2(\REGISTERS[17][21] ), .ZN(n5377)
         );
  NAND4_X1 U3929 ( .A1(n3934), .A2(n3935), .A3(n3936), .A4(n3937), .ZN(n3933)
         );
  AOI221_X1 U3930 ( .B1(n1396), .B2(\REGISTERS[12][21] ), .C1(n1393), .C2(
        \REGISTERS[11][21] ), .A(n3942), .ZN(n3936) );
  NOR4_X1 U3931 ( .A1(n3938), .A2(n3939), .A3(n3940), .A4(n3941), .ZN(n3937)
         );
  AOI222_X1 U3932 ( .A1(n1372), .A2(\REGISTERS[16][21] ), .B1(n1368), .B2(
        \REGISTERS[18][21] ), .C1(n1365), .C2(\REGISTERS[17][21] ), .ZN(n3934)
         );
  NAND4_X1 U3933 ( .A1(n5336), .A2(n5337), .A3(n5338), .A4(n5339), .ZN(n5335)
         );
  AOI221_X1 U3934 ( .B1(n684), .B2(\REGISTERS[12][22] ), .C1(n681), .C2(
        \REGISTERS[11][22] ), .A(n5344), .ZN(n5338) );
  NOR4_X1 U3935 ( .A1(n5340), .A2(n5341), .A3(n5342), .A4(n5343), .ZN(n5339)
         );
  AOI222_X1 U3936 ( .A1(n660), .A2(\REGISTERS[16][22] ), .B1(n656), .B2(
        \REGISTERS[18][22] ), .C1(n653), .C2(\REGISTERS[17][22] ), .ZN(n5336)
         );
  NAND4_X1 U3937 ( .A1(n3893), .A2(n3894), .A3(n3895), .A4(n3896), .ZN(n3892)
         );
  AOI221_X1 U3938 ( .B1(n1396), .B2(\REGISTERS[12][22] ), .C1(n1393), .C2(
        \REGISTERS[11][22] ), .A(n3901), .ZN(n3895) );
  NOR4_X1 U3939 ( .A1(n3897), .A2(n3898), .A3(n3899), .A4(n3900), .ZN(n3896)
         );
  AOI222_X1 U3940 ( .A1(n1372), .A2(\REGISTERS[16][22] ), .B1(n1368), .B2(
        \REGISTERS[18][22] ), .C1(n1365), .C2(\REGISTERS[17][22] ), .ZN(n3893)
         );
  NAND4_X1 U3941 ( .A1(n5295), .A2(n5296), .A3(n5297), .A4(n5298), .ZN(n5294)
         );
  AOI221_X1 U3942 ( .B1(n684), .B2(\REGISTERS[12][23] ), .C1(n681), .C2(
        \REGISTERS[11][23] ), .A(n5303), .ZN(n5297) );
  NOR4_X1 U3943 ( .A1(n5299), .A2(n5300), .A3(n5301), .A4(n5302), .ZN(n5298)
         );
  AOI222_X1 U3944 ( .A1(n660), .A2(\REGISTERS[16][23] ), .B1(n656), .B2(
        \REGISTERS[18][23] ), .C1(n653), .C2(\REGISTERS[17][23] ), .ZN(n5295)
         );
  NAND4_X1 U3945 ( .A1(n3852), .A2(n3853), .A3(n3854), .A4(n3855), .ZN(n3851)
         );
  AOI221_X1 U3946 ( .B1(n1396), .B2(\REGISTERS[12][23] ), .C1(n1393), .C2(
        \REGISTERS[11][23] ), .A(n3860), .ZN(n3854) );
  NOR4_X1 U3947 ( .A1(n3856), .A2(n3857), .A3(n3858), .A4(n3859), .ZN(n3855)
         );
  AOI222_X1 U3948 ( .A1(n1372), .A2(\REGISTERS[16][23] ), .B1(n1368), .B2(
        \REGISTERS[18][23] ), .C1(n1365), .C2(\REGISTERS[17][23] ), .ZN(n3852)
         );
  NAND4_X1 U3949 ( .A1(n5254), .A2(n5255), .A3(n5256), .A4(n5257), .ZN(n5253)
         );
  AOI221_X1 U3950 ( .B1(n685), .B2(\REGISTERS[12][24] ), .C1(n682), .C2(
        \REGISTERS[11][24] ), .A(n5262), .ZN(n5256) );
  NOR4_X1 U3951 ( .A1(n5258), .A2(n5259), .A3(n5260), .A4(n5261), .ZN(n5257)
         );
  AOI222_X1 U3952 ( .A1(n661), .A2(\REGISTERS[16][24] ), .B1(n656), .B2(
        \REGISTERS[18][24] ), .C1(n653), .C2(\REGISTERS[17][24] ), .ZN(n5254)
         );
  NAND4_X1 U3953 ( .A1(n3811), .A2(n3812), .A3(n3813), .A4(n3814), .ZN(n3810)
         );
  AOI221_X1 U3954 ( .B1(n1397), .B2(\REGISTERS[12][24] ), .C1(n1394), .C2(
        \REGISTERS[11][24] ), .A(n3819), .ZN(n3813) );
  NOR4_X1 U3955 ( .A1(n3815), .A2(n3816), .A3(n3817), .A4(n3818), .ZN(n3814)
         );
  AOI222_X1 U3956 ( .A1(n1373), .A2(\REGISTERS[16][24] ), .B1(n1368), .B2(
        \REGISTERS[18][24] ), .C1(n1365), .C2(\REGISTERS[17][24] ), .ZN(n3811)
         );
  NAND4_X1 U3957 ( .A1(n5213), .A2(n5214), .A3(n5215), .A4(n5216), .ZN(n5212)
         );
  AOI221_X1 U3958 ( .B1(n685), .B2(\REGISTERS[12][25] ), .C1(n682), .C2(
        \REGISTERS[11][25] ), .A(n5221), .ZN(n5215) );
  NOR4_X1 U3959 ( .A1(n5217), .A2(n5218), .A3(n5219), .A4(n5220), .ZN(n5216)
         );
  AOI222_X1 U3960 ( .A1(n661), .A2(\REGISTERS[16][25] ), .B1(n656), .B2(
        \REGISTERS[18][25] ), .C1(n653), .C2(\REGISTERS[17][25] ), .ZN(n5213)
         );
  NAND4_X1 U3961 ( .A1(n3770), .A2(n3771), .A3(n3772), .A4(n3773), .ZN(n3769)
         );
  AOI221_X1 U3962 ( .B1(n1397), .B2(\REGISTERS[12][25] ), .C1(n1394), .C2(
        \REGISTERS[11][25] ), .A(n3778), .ZN(n3772) );
  NOR4_X1 U3963 ( .A1(n3774), .A2(n3775), .A3(n3776), .A4(n3777), .ZN(n3773)
         );
  AOI222_X1 U3964 ( .A1(n1373), .A2(\REGISTERS[16][25] ), .B1(n1368), .B2(
        \REGISTERS[18][25] ), .C1(n1365), .C2(\REGISTERS[17][25] ), .ZN(n3770)
         );
  NAND4_X1 U3965 ( .A1(n5172), .A2(n5173), .A3(n5174), .A4(n5175), .ZN(n5171)
         );
  AOI221_X1 U3966 ( .B1(n685), .B2(\REGISTERS[12][26] ), .C1(n682), .C2(
        \REGISTERS[11][26] ), .A(n5180), .ZN(n5174) );
  NOR4_X1 U3967 ( .A1(n5176), .A2(n5177), .A3(n5178), .A4(n5179), .ZN(n5175)
         );
  AOI222_X1 U3968 ( .A1(n661), .A2(\REGISTERS[16][26] ), .B1(n656), .B2(
        \REGISTERS[18][26] ), .C1(n653), .C2(\REGISTERS[17][26] ), .ZN(n5172)
         );
  NAND4_X1 U3969 ( .A1(n3729), .A2(n3730), .A3(n3731), .A4(n3732), .ZN(n3728)
         );
  AOI221_X1 U3970 ( .B1(n1397), .B2(\REGISTERS[12][26] ), .C1(n1394), .C2(
        \REGISTERS[11][26] ), .A(n3737), .ZN(n3731) );
  NOR4_X1 U3971 ( .A1(n3733), .A2(n3734), .A3(n3735), .A4(n3736), .ZN(n3732)
         );
  AOI222_X1 U3972 ( .A1(n1373), .A2(\REGISTERS[16][26] ), .B1(n1368), .B2(
        \REGISTERS[18][26] ), .C1(n1365), .C2(\REGISTERS[17][26] ), .ZN(n3729)
         );
  NAND4_X1 U3973 ( .A1(n5131), .A2(n5132), .A3(n5133), .A4(n5134), .ZN(n5130)
         );
  AOI221_X1 U3974 ( .B1(n685), .B2(\REGISTERS[12][27] ), .C1(n682), .C2(
        \REGISTERS[11][27] ), .A(n5139), .ZN(n5133) );
  NOR4_X1 U3975 ( .A1(n5135), .A2(n5136), .A3(n5137), .A4(n5138), .ZN(n5134)
         );
  AOI222_X1 U3976 ( .A1(n661), .A2(\REGISTERS[16][27] ), .B1(n656), .B2(
        \REGISTERS[18][27] ), .C1(n653), .C2(\REGISTERS[17][27] ), .ZN(n5131)
         );
  NAND4_X1 U3977 ( .A1(n3688), .A2(n3689), .A3(n3690), .A4(n3691), .ZN(n3687)
         );
  AOI221_X1 U3978 ( .B1(n1397), .B2(\REGISTERS[12][27] ), .C1(n1394), .C2(
        \REGISTERS[11][27] ), .A(n3696), .ZN(n3690) );
  NOR4_X1 U3979 ( .A1(n3692), .A2(n3693), .A3(n3694), .A4(n3695), .ZN(n3691)
         );
  AOI222_X1 U3980 ( .A1(n1373), .A2(\REGISTERS[16][27] ), .B1(n1368), .B2(
        \REGISTERS[18][27] ), .C1(n1365), .C2(\REGISTERS[17][27] ), .ZN(n3688)
         );
  NAND4_X1 U3981 ( .A1(n5090), .A2(n5091), .A3(n5092), .A4(n5093), .ZN(n5089)
         );
  AOI221_X1 U3982 ( .B1(n685), .B2(\REGISTERS[12][28] ), .C1(n682), .C2(
        \REGISTERS[11][28] ), .A(n5098), .ZN(n5092) );
  NOR4_X1 U3983 ( .A1(n5094), .A2(n5095), .A3(n5096), .A4(n5097), .ZN(n5093)
         );
  AOI222_X1 U3984 ( .A1(n661), .A2(\REGISTERS[16][28] ), .B1(n656), .B2(
        \REGISTERS[18][28] ), .C1(n653), .C2(\REGISTERS[17][28] ), .ZN(n5090)
         );
  NAND4_X1 U3985 ( .A1(n3647), .A2(n3648), .A3(n3649), .A4(n3650), .ZN(n3646)
         );
  AOI221_X1 U3986 ( .B1(n1397), .B2(\REGISTERS[12][28] ), .C1(n1394), .C2(
        \REGISTERS[11][28] ), .A(n3655), .ZN(n3649) );
  NOR4_X1 U3987 ( .A1(n3651), .A2(n3652), .A3(n3653), .A4(n3654), .ZN(n3650)
         );
  AOI222_X1 U3988 ( .A1(n1373), .A2(\REGISTERS[16][28] ), .B1(n1368), .B2(
        \REGISTERS[18][28] ), .C1(n1365), .C2(\REGISTERS[17][28] ), .ZN(n3647)
         );
  NAND4_X1 U3989 ( .A1(n5049), .A2(n5050), .A3(n5051), .A4(n5052), .ZN(n5048)
         );
  AOI221_X1 U3990 ( .B1(n685), .B2(\REGISTERS[12][29] ), .C1(n682), .C2(
        \REGISTERS[11][29] ), .A(n5057), .ZN(n5051) );
  NOR4_X1 U3991 ( .A1(n5053), .A2(n5054), .A3(n5055), .A4(n5056), .ZN(n5052)
         );
  AOI222_X1 U3992 ( .A1(n661), .A2(\REGISTERS[16][29] ), .B1(n656), .B2(
        \REGISTERS[18][29] ), .C1(n653), .C2(\REGISTERS[17][29] ), .ZN(n5049)
         );
  NAND4_X1 U3993 ( .A1(n3606), .A2(n3607), .A3(n3608), .A4(n3609), .ZN(n3605)
         );
  AOI221_X1 U3994 ( .B1(n1397), .B2(\REGISTERS[12][29] ), .C1(n1394), .C2(
        \REGISTERS[11][29] ), .A(n3614), .ZN(n3608) );
  NOR4_X1 U3995 ( .A1(n3610), .A2(n3611), .A3(n3612), .A4(n3613), .ZN(n3609)
         );
  AOI222_X1 U3996 ( .A1(n1373), .A2(\REGISTERS[16][29] ), .B1(n1368), .B2(
        \REGISTERS[18][29] ), .C1(n1365), .C2(\REGISTERS[17][29] ), .ZN(n3606)
         );
  NAND4_X1 U3997 ( .A1(n5008), .A2(n5009), .A3(n5010), .A4(n5011), .ZN(n5007)
         );
  AOI221_X1 U3998 ( .B1(n685), .B2(\REGISTERS[12][30] ), .C1(n682), .C2(
        \REGISTERS[11][30] ), .A(n5016), .ZN(n5010) );
  NOR4_X1 U3999 ( .A1(n5012), .A2(n5013), .A3(n5014), .A4(n5015), .ZN(n5011)
         );
  AOI222_X1 U4000 ( .A1(n661), .A2(\REGISTERS[16][30] ), .B1(n656), .B2(
        \REGISTERS[18][30] ), .C1(n653), .C2(\REGISTERS[17][30] ), .ZN(n5008)
         );
  NAND4_X1 U4001 ( .A1(n3565), .A2(n3566), .A3(n3567), .A4(n3568), .ZN(n3564)
         );
  AOI221_X1 U4002 ( .B1(n1397), .B2(\REGISTERS[12][30] ), .C1(n1394), .C2(
        \REGISTERS[11][30] ), .A(n3573), .ZN(n3567) );
  NOR4_X1 U4003 ( .A1(n3569), .A2(n3570), .A3(n3571), .A4(n3572), .ZN(n3568)
         );
  AOI222_X1 U4004 ( .A1(n1373), .A2(\REGISTERS[16][30] ), .B1(n1368), .B2(
        \REGISTERS[18][30] ), .C1(n1365), .C2(\REGISTERS[17][30] ), .ZN(n3565)
         );
  NAND4_X1 U4005 ( .A1(n4879), .A2(n4880), .A3(n4881), .A4(n4882), .ZN(n4878)
         );
  AOI221_X1 U4006 ( .B1(n685), .B2(\REGISTERS[12][31] ), .C1(n682), .C2(
        \REGISTERS[11][31] ), .A(n4900), .ZN(n4881) );
  NOR4_X1 U4007 ( .A1(n4883), .A2(n4884), .A3(n4885), .A4(n4886), .ZN(n4882)
         );
  AOI222_X1 U4008 ( .A1(n661), .A2(\REGISTERS[16][31] ), .B1(n656), .B2(
        \REGISTERS[18][31] ), .C1(n653), .C2(\REGISTERS[17][31] ), .ZN(n4879)
         );
  NAND4_X1 U4009 ( .A1(n3436), .A2(n3437), .A3(n3438), .A4(n3439), .ZN(n3435)
         );
  AOI221_X1 U4010 ( .B1(n1397), .B2(\REGISTERS[12][31] ), .C1(n1394), .C2(
        \REGISTERS[11][31] ), .A(n3457), .ZN(n3438) );
  NOR4_X1 U4011 ( .A1(n3440), .A2(n3441), .A3(n3442), .A4(n3443), .ZN(n3439)
         );
  AOI222_X1 U4012 ( .A1(n1373), .A2(\REGISTERS[16][31] ), .B1(n1368), .B2(
        \REGISTERS[18][31] ), .C1(n1365), .C2(\REGISTERS[17][31] ), .ZN(n3436)
         );
  NAND4_X1 U4013 ( .A1(n6269), .A2(n6270), .A3(n6271), .A4(n6272), .ZN(n6236)
         );
  AOI221_X1 U4014 ( .B1(n617), .B2(\REGISTERS[34][0] ), .C1(n614), .C2(
        \REGISTERS[33][0] ), .A(n6282), .ZN(n6271) );
  NOR4_X1 U4015 ( .A1(n6273), .A2(n6274), .A3(n6275), .A4(n6276), .ZN(n6272)
         );
  AOI222_X1 U4016 ( .A1(n593), .A2(\REGISTERS[38][0] ), .B1(n592), .B2(
        \REGISTERS[40][0] ), .C1(n493), .C2(\REGISTERS[39][0] ), .ZN(n6269) );
  NAND4_X1 U4017 ( .A1(n4826), .A2(n4827), .A3(n4828), .A4(n4829), .ZN(n4793)
         );
  AOI221_X1 U4018 ( .B1(n1329), .B2(\REGISTERS[34][0] ), .C1(n1326), .C2(
        \REGISTERS[33][0] ), .A(n4839), .ZN(n4828) );
  NOR4_X1 U4019 ( .A1(n4830), .A2(n4831), .A3(n4832), .A4(n4833), .ZN(n4829)
         );
  AOI222_X1 U4020 ( .A1(n1305), .A2(\REGISTERS[38][0] ), .B1(n1304), .B2(
        \REGISTERS[40][0] ), .C1(n1301), .C2(\REGISTERS[39][0] ), .ZN(n4826)
         );
  NAND4_X1 U4021 ( .A1(n6206), .A2(n6207), .A3(n6208), .A4(n6209), .ZN(n6195)
         );
  AOI221_X1 U4022 ( .B1(n617), .B2(\REGISTERS[34][1] ), .C1(n614), .C2(
        \REGISTERS[33][1] ), .A(n6214), .ZN(n6208) );
  NOR4_X1 U4023 ( .A1(n6210), .A2(n6211), .A3(n6212), .A4(n6213), .ZN(n6209)
         );
  AOI222_X1 U4024 ( .A1(n593), .A2(\REGISTERS[38][1] ), .B1(n592), .B2(
        \REGISTERS[40][1] ), .C1(n493), .C2(\REGISTERS[39][1] ), .ZN(n6206) );
  NAND4_X1 U4025 ( .A1(n4763), .A2(n4764), .A3(n4765), .A4(n4766), .ZN(n4752)
         );
  AOI221_X1 U4026 ( .B1(n1329), .B2(\REGISTERS[34][1] ), .C1(n1326), .C2(
        \REGISTERS[33][1] ), .A(n4771), .ZN(n4765) );
  NOR4_X1 U4027 ( .A1(n4767), .A2(n4768), .A3(n4769), .A4(n4770), .ZN(n4766)
         );
  AOI222_X1 U4028 ( .A1(n1305), .A2(\REGISTERS[38][1] ), .B1(n1304), .B2(
        \REGISTERS[40][1] ), .C1(n1301), .C2(\REGISTERS[39][1] ), .ZN(n4763)
         );
  NAND4_X1 U4029 ( .A1(n6165), .A2(n6166), .A3(n6167), .A4(n6168), .ZN(n6154)
         );
  AOI221_X1 U4030 ( .B1(n617), .B2(\REGISTERS[34][2] ), .C1(n614), .C2(
        \REGISTERS[33][2] ), .A(n6173), .ZN(n6167) );
  NOR4_X1 U4031 ( .A1(n6169), .A2(n6170), .A3(n6171), .A4(n6172), .ZN(n6168)
         );
  AOI222_X1 U4032 ( .A1(n593), .A2(\REGISTERS[38][2] ), .B1(n592), .B2(
        \REGISTERS[40][2] ), .C1(n493), .C2(\REGISTERS[39][2] ), .ZN(n6165) );
  NAND4_X1 U4033 ( .A1(n4722), .A2(n4723), .A3(n4724), .A4(n4725), .ZN(n4711)
         );
  AOI221_X1 U4034 ( .B1(n1329), .B2(\REGISTERS[34][2] ), .C1(n1326), .C2(
        \REGISTERS[33][2] ), .A(n4730), .ZN(n4724) );
  NOR4_X1 U4035 ( .A1(n4726), .A2(n4727), .A3(n4728), .A4(n4729), .ZN(n4725)
         );
  AOI222_X1 U4036 ( .A1(n1305), .A2(\REGISTERS[38][2] ), .B1(n1304), .B2(
        \REGISTERS[40][2] ), .C1(n1301), .C2(\REGISTERS[39][2] ), .ZN(n4722)
         );
  NAND4_X1 U4037 ( .A1(n6124), .A2(n6125), .A3(n6126), .A4(n6127), .ZN(n6113)
         );
  AOI221_X1 U4038 ( .B1(n617), .B2(\REGISTERS[34][3] ), .C1(n614), .C2(
        \REGISTERS[33][3] ), .A(n6132), .ZN(n6126) );
  NOR4_X1 U4039 ( .A1(n6128), .A2(n6129), .A3(n6130), .A4(n6131), .ZN(n6127)
         );
  AOI222_X1 U4040 ( .A1(n593), .A2(\REGISTERS[38][3] ), .B1(n592), .B2(
        \REGISTERS[40][3] ), .C1(n493), .C2(\REGISTERS[39][3] ), .ZN(n6124) );
  NAND4_X1 U4041 ( .A1(n4681), .A2(n4682), .A3(n4683), .A4(n4684), .ZN(n4670)
         );
  AOI221_X1 U4042 ( .B1(n1329), .B2(\REGISTERS[34][3] ), .C1(n1326), .C2(
        \REGISTERS[33][3] ), .A(n4689), .ZN(n4683) );
  NOR4_X1 U4043 ( .A1(n4685), .A2(n4686), .A3(n4687), .A4(n4688), .ZN(n4684)
         );
  AOI222_X1 U4044 ( .A1(n1305), .A2(\REGISTERS[38][3] ), .B1(n1304), .B2(
        \REGISTERS[40][3] ), .C1(n1301), .C2(\REGISTERS[39][3] ), .ZN(n4681)
         );
  NAND4_X1 U4045 ( .A1(n6083), .A2(n6084), .A3(n6085), .A4(n6086), .ZN(n6072)
         );
  AOI221_X1 U4046 ( .B1(n617), .B2(\REGISTERS[34][4] ), .C1(n614), .C2(
        \REGISTERS[33][4] ), .A(n6091), .ZN(n6085) );
  NOR4_X1 U4047 ( .A1(n6087), .A2(n6088), .A3(n6089), .A4(n6090), .ZN(n6086)
         );
  AOI222_X1 U4048 ( .A1(n593), .A2(\REGISTERS[38][4] ), .B1(n592), .B2(
        \REGISTERS[40][4] ), .C1(n493), .C2(\REGISTERS[39][4] ), .ZN(n6083) );
  NAND4_X1 U4049 ( .A1(n4640), .A2(n4641), .A3(n4642), .A4(n4643), .ZN(n4629)
         );
  AOI221_X1 U4050 ( .B1(n1329), .B2(\REGISTERS[34][4] ), .C1(n1326), .C2(
        \REGISTERS[33][4] ), .A(n4648), .ZN(n4642) );
  NOR4_X1 U4051 ( .A1(n4644), .A2(n4645), .A3(n4646), .A4(n4647), .ZN(n4643)
         );
  AOI222_X1 U4052 ( .A1(n1305), .A2(\REGISTERS[38][4] ), .B1(n1304), .B2(
        \REGISTERS[40][4] ), .C1(n1301), .C2(\REGISTERS[39][4] ), .ZN(n4640)
         );
  NAND4_X1 U4053 ( .A1(n6042), .A2(n6043), .A3(n6044), .A4(n6045), .ZN(n6031)
         );
  AOI221_X1 U4054 ( .B1(n617), .B2(\REGISTERS[34][5] ), .C1(n614), .C2(
        \REGISTERS[33][5] ), .A(n6050), .ZN(n6044) );
  NOR4_X1 U4055 ( .A1(n6046), .A2(n6047), .A3(n6048), .A4(n6049), .ZN(n6045)
         );
  AOI222_X1 U4056 ( .A1(n593), .A2(\REGISTERS[38][5] ), .B1(n592), .B2(
        \REGISTERS[40][5] ), .C1(n493), .C2(\REGISTERS[39][5] ), .ZN(n6042) );
  NAND4_X1 U4057 ( .A1(n4599), .A2(n4600), .A3(n4601), .A4(n4602), .ZN(n4588)
         );
  AOI221_X1 U4058 ( .B1(n1329), .B2(\REGISTERS[34][5] ), .C1(n1326), .C2(
        \REGISTERS[33][5] ), .A(n4607), .ZN(n4601) );
  NOR4_X1 U4059 ( .A1(n4603), .A2(n4604), .A3(n4605), .A4(n4606), .ZN(n4602)
         );
  AOI222_X1 U4060 ( .A1(n1305), .A2(\REGISTERS[38][5] ), .B1(n1304), .B2(
        \REGISTERS[40][5] ), .C1(n1301), .C2(\REGISTERS[39][5] ), .ZN(n4599)
         );
  NAND4_X1 U4061 ( .A1(n6001), .A2(n6002), .A3(n6003), .A4(n6004), .ZN(n5990)
         );
  AOI221_X1 U4062 ( .B1(n617), .B2(\REGISTERS[34][6] ), .C1(n614), .C2(
        \REGISTERS[33][6] ), .A(n6009), .ZN(n6003) );
  NOR4_X1 U4063 ( .A1(n6005), .A2(n6006), .A3(n6007), .A4(n6008), .ZN(n6004)
         );
  AOI222_X1 U4064 ( .A1(n593), .A2(\REGISTERS[38][6] ), .B1(n592), .B2(
        \REGISTERS[40][6] ), .C1(n493), .C2(\REGISTERS[39][6] ), .ZN(n6001) );
  NAND4_X1 U4065 ( .A1(n4558), .A2(n4559), .A3(n4560), .A4(n4561), .ZN(n4547)
         );
  AOI221_X1 U4066 ( .B1(n1329), .B2(\REGISTERS[34][6] ), .C1(n1326), .C2(
        \REGISTERS[33][6] ), .A(n4566), .ZN(n4560) );
  NOR4_X1 U4067 ( .A1(n4562), .A2(n4563), .A3(n4564), .A4(n4565), .ZN(n4561)
         );
  AOI222_X1 U4068 ( .A1(n1305), .A2(\REGISTERS[38][6] ), .B1(n1304), .B2(
        \REGISTERS[40][6] ), .C1(n1301), .C2(\REGISTERS[39][6] ), .ZN(n4558)
         );
  NAND4_X1 U4069 ( .A1(n5960), .A2(n5961), .A3(n5962), .A4(n5963), .ZN(n5949)
         );
  AOI221_X1 U4070 ( .B1(n617), .B2(\REGISTERS[34][7] ), .C1(n614), .C2(
        \REGISTERS[33][7] ), .A(n5968), .ZN(n5962) );
  NOR4_X1 U4071 ( .A1(n5964), .A2(n5965), .A3(n5966), .A4(n5967), .ZN(n5963)
         );
  AOI222_X1 U4072 ( .A1(n593), .A2(\REGISTERS[38][7] ), .B1(n592), .B2(
        \REGISTERS[40][7] ), .C1(n493), .C2(\REGISTERS[39][7] ), .ZN(n5960) );
  NAND4_X1 U4073 ( .A1(n4517), .A2(n4518), .A3(n4519), .A4(n4520), .ZN(n4506)
         );
  AOI221_X1 U4074 ( .B1(n1329), .B2(\REGISTERS[34][7] ), .C1(n1326), .C2(
        \REGISTERS[33][7] ), .A(n4525), .ZN(n4519) );
  NOR4_X1 U4075 ( .A1(n4521), .A2(n4522), .A3(n4523), .A4(n4524), .ZN(n4520)
         );
  AOI222_X1 U4076 ( .A1(n1305), .A2(\REGISTERS[38][7] ), .B1(n1304), .B2(
        \REGISTERS[40][7] ), .C1(n1301), .C2(\REGISTERS[39][7] ), .ZN(n4517)
         );
  NAND4_X1 U4077 ( .A1(n5919), .A2(n5920), .A3(n5921), .A4(n5922), .ZN(n5908)
         );
  AOI221_X1 U4078 ( .B1(n617), .B2(\REGISTERS[34][8] ), .C1(n614), .C2(
        \REGISTERS[33][8] ), .A(n5927), .ZN(n5921) );
  NOR4_X1 U4079 ( .A1(n5923), .A2(n5924), .A3(n5925), .A4(n5926), .ZN(n5922)
         );
  AOI222_X1 U4080 ( .A1(n593), .A2(\REGISTERS[38][8] ), .B1(n495), .B2(
        \REGISTERS[40][8] ), .C1(n492), .C2(\REGISTERS[39][8] ), .ZN(n5919) );
  NAND4_X1 U4081 ( .A1(n4476), .A2(n4477), .A3(n4478), .A4(n4479), .ZN(n4465)
         );
  AOI221_X1 U4082 ( .B1(n1329), .B2(\REGISTERS[34][8] ), .C1(n1326), .C2(
        \REGISTERS[33][8] ), .A(n4484), .ZN(n4478) );
  NOR4_X1 U4083 ( .A1(n4480), .A2(n4481), .A3(n4482), .A4(n4483), .ZN(n4479)
         );
  AOI222_X1 U4084 ( .A1(n1305), .A2(\REGISTERS[38][8] ), .B1(n1303), .B2(
        \REGISTERS[40][8] ), .C1(n1300), .C2(\REGISTERS[39][8] ), .ZN(n4476)
         );
  NAND4_X1 U4085 ( .A1(n5878), .A2(n5879), .A3(n5880), .A4(n5881), .ZN(n5867)
         );
  AOI221_X1 U4086 ( .B1(n617), .B2(\REGISTERS[34][9] ), .C1(n614), .C2(
        \REGISTERS[33][9] ), .A(n5886), .ZN(n5880) );
  NOR4_X1 U4087 ( .A1(n5882), .A2(n5883), .A3(n5884), .A4(n5885), .ZN(n5881)
         );
  AOI222_X1 U4088 ( .A1(n593), .A2(\REGISTERS[38][9] ), .B1(n495), .B2(
        \REGISTERS[40][9] ), .C1(n492), .C2(\REGISTERS[39][9] ), .ZN(n5878) );
  NAND4_X1 U4089 ( .A1(n4435), .A2(n4436), .A3(n4437), .A4(n4438), .ZN(n4424)
         );
  AOI221_X1 U4090 ( .B1(n1329), .B2(\REGISTERS[34][9] ), .C1(n1326), .C2(
        \REGISTERS[33][9] ), .A(n4443), .ZN(n4437) );
  NOR4_X1 U4091 ( .A1(n4439), .A2(n4440), .A3(n4441), .A4(n4442), .ZN(n4438)
         );
  AOI222_X1 U4092 ( .A1(n1305), .A2(\REGISTERS[38][9] ), .B1(n1303), .B2(
        \REGISTERS[40][9] ), .C1(n1300), .C2(\REGISTERS[39][9] ), .ZN(n4435)
         );
  NAND4_X1 U4093 ( .A1(n5837), .A2(n5838), .A3(n5839), .A4(n5840), .ZN(n5826)
         );
  AOI221_X1 U4094 ( .B1(n617), .B2(\REGISTERS[34][10] ), .C1(n614), .C2(
        \REGISTERS[33][10] ), .A(n5845), .ZN(n5839) );
  NOR4_X1 U4095 ( .A1(n5841), .A2(n5842), .A3(n5843), .A4(n5844), .ZN(n5840)
         );
  AOI222_X1 U4096 ( .A1(n593), .A2(\REGISTERS[38][10] ), .B1(n495), .B2(
        \REGISTERS[40][10] ), .C1(n492), .C2(\REGISTERS[39][10] ), .ZN(n5837)
         );
  NAND4_X1 U4097 ( .A1(n4394), .A2(n4395), .A3(n4396), .A4(n4397), .ZN(n4383)
         );
  AOI221_X1 U4098 ( .B1(n1329), .B2(\REGISTERS[34][10] ), .C1(n1326), .C2(
        \REGISTERS[33][10] ), .A(n4402), .ZN(n4396) );
  NOR4_X1 U4099 ( .A1(n4398), .A2(n4399), .A3(n4400), .A4(n4401), .ZN(n4397)
         );
  AOI222_X1 U4100 ( .A1(n1305), .A2(\REGISTERS[38][10] ), .B1(n1303), .B2(
        \REGISTERS[40][10] ), .C1(n1300), .C2(\REGISTERS[39][10] ), .ZN(n4394)
         );
  NAND4_X1 U4101 ( .A1(n5796), .A2(n5797), .A3(n5798), .A4(n5799), .ZN(n5785)
         );
  AOI221_X1 U4102 ( .B1(n617), .B2(\REGISTERS[34][11] ), .C1(n614), .C2(
        \REGISTERS[33][11] ), .A(n5804), .ZN(n5798) );
  NOR4_X1 U4103 ( .A1(n5800), .A2(n5801), .A3(n5802), .A4(n5803), .ZN(n5799)
         );
  AOI222_X1 U4104 ( .A1(n593), .A2(\REGISTERS[38][11] ), .B1(n495), .B2(
        \REGISTERS[40][11] ), .C1(n492), .C2(\REGISTERS[39][11] ), .ZN(n5796)
         );
  NAND4_X1 U4105 ( .A1(n4353), .A2(n4354), .A3(n4355), .A4(n4356), .ZN(n4342)
         );
  AOI221_X1 U4106 ( .B1(n1329), .B2(\REGISTERS[34][11] ), .C1(n1326), .C2(
        \REGISTERS[33][11] ), .A(n4361), .ZN(n4355) );
  NOR4_X1 U4107 ( .A1(n4357), .A2(n4358), .A3(n4359), .A4(n4360), .ZN(n4356)
         );
  AOI222_X1 U4108 ( .A1(n1305), .A2(\REGISTERS[38][11] ), .B1(n1303), .B2(
        \REGISTERS[40][11] ), .C1(n1300), .C2(\REGISTERS[39][11] ), .ZN(n4353)
         );
  NAND4_X1 U4109 ( .A1(n5755), .A2(n5756), .A3(n5757), .A4(n5758), .ZN(n5744)
         );
  AOI221_X1 U4110 ( .B1(n618), .B2(\REGISTERS[34][12] ), .C1(n615), .C2(
        \REGISTERS[33][12] ), .A(n5763), .ZN(n5757) );
  NOR4_X1 U4111 ( .A1(n5759), .A2(n5760), .A3(n5761), .A4(n5762), .ZN(n5758)
         );
  AOI222_X1 U4112 ( .A1(n594), .A2(\REGISTERS[38][12] ), .B1(n495), .B2(
        \REGISTERS[40][12] ), .C1(n492), .C2(\REGISTERS[39][12] ), .ZN(n5755)
         );
  NAND4_X1 U4113 ( .A1(n4312), .A2(n4313), .A3(n4314), .A4(n4315), .ZN(n4301)
         );
  AOI221_X1 U4114 ( .B1(n1330), .B2(\REGISTERS[34][12] ), .C1(n1327), .C2(
        \REGISTERS[33][12] ), .A(n4320), .ZN(n4314) );
  NOR4_X1 U4115 ( .A1(n4316), .A2(n4317), .A3(n4318), .A4(n4319), .ZN(n4315)
         );
  AOI222_X1 U4116 ( .A1(n1306), .A2(\REGISTERS[38][12] ), .B1(n1303), .B2(
        \REGISTERS[40][12] ), .C1(n1300), .C2(\REGISTERS[39][12] ), .ZN(n4312)
         );
  NAND4_X1 U4117 ( .A1(n5714), .A2(n5715), .A3(n5716), .A4(n5717), .ZN(n5703)
         );
  AOI221_X1 U4118 ( .B1(n618), .B2(\REGISTERS[34][13] ), .C1(n615), .C2(
        \REGISTERS[33][13] ), .A(n5722), .ZN(n5716) );
  NOR4_X1 U4119 ( .A1(n5718), .A2(n5719), .A3(n5720), .A4(n5721), .ZN(n5717)
         );
  AOI222_X1 U4120 ( .A1(n594), .A2(\REGISTERS[38][13] ), .B1(n495), .B2(
        \REGISTERS[40][13] ), .C1(n492), .C2(\REGISTERS[39][13] ), .ZN(n5714)
         );
  NAND4_X1 U4121 ( .A1(n4271), .A2(n4272), .A3(n4273), .A4(n4274), .ZN(n4260)
         );
  AOI221_X1 U4122 ( .B1(n1330), .B2(\REGISTERS[34][13] ), .C1(n1327), .C2(
        \REGISTERS[33][13] ), .A(n4279), .ZN(n4273) );
  NOR4_X1 U4123 ( .A1(n4275), .A2(n4276), .A3(n4277), .A4(n4278), .ZN(n4274)
         );
  AOI222_X1 U4124 ( .A1(n1306), .A2(\REGISTERS[38][13] ), .B1(n1303), .B2(
        \REGISTERS[40][13] ), .C1(n1300), .C2(\REGISTERS[39][13] ), .ZN(n4271)
         );
  NAND4_X1 U4125 ( .A1(n5673), .A2(n5674), .A3(n5675), .A4(n5676), .ZN(n5662)
         );
  AOI221_X1 U4126 ( .B1(n618), .B2(\REGISTERS[34][14] ), .C1(n615), .C2(
        \REGISTERS[33][14] ), .A(n5681), .ZN(n5675) );
  NOR4_X1 U4127 ( .A1(n5677), .A2(n5678), .A3(n5679), .A4(n5680), .ZN(n5676)
         );
  AOI222_X1 U4128 ( .A1(n594), .A2(\REGISTERS[38][14] ), .B1(n495), .B2(
        \REGISTERS[40][14] ), .C1(n492), .C2(\REGISTERS[39][14] ), .ZN(n5673)
         );
  NAND4_X1 U4129 ( .A1(n4230), .A2(n4231), .A3(n4232), .A4(n4233), .ZN(n4219)
         );
  AOI221_X1 U4130 ( .B1(n1330), .B2(\REGISTERS[34][14] ), .C1(n1327), .C2(
        \REGISTERS[33][14] ), .A(n4238), .ZN(n4232) );
  NOR4_X1 U4131 ( .A1(n4234), .A2(n4235), .A3(n4236), .A4(n4237), .ZN(n4233)
         );
  AOI222_X1 U4132 ( .A1(n1306), .A2(\REGISTERS[38][14] ), .B1(n1303), .B2(
        \REGISTERS[40][14] ), .C1(n1300), .C2(\REGISTERS[39][14] ), .ZN(n4230)
         );
  NAND4_X1 U4133 ( .A1(n5632), .A2(n5633), .A3(n5634), .A4(n5635), .ZN(n5621)
         );
  AOI221_X1 U4134 ( .B1(n618), .B2(\REGISTERS[34][15] ), .C1(n615), .C2(
        \REGISTERS[33][15] ), .A(n5640), .ZN(n5634) );
  NOR4_X1 U4135 ( .A1(n5636), .A2(n5637), .A3(n5638), .A4(n5639), .ZN(n5635)
         );
  AOI222_X1 U4136 ( .A1(n594), .A2(\REGISTERS[38][15] ), .B1(n495), .B2(
        \REGISTERS[40][15] ), .C1(n492), .C2(\REGISTERS[39][15] ), .ZN(n5632)
         );
  NAND4_X1 U4137 ( .A1(n4189), .A2(n4190), .A3(n4191), .A4(n4192), .ZN(n4178)
         );
  AOI221_X1 U4138 ( .B1(n1330), .B2(\REGISTERS[34][15] ), .C1(n1327), .C2(
        \REGISTERS[33][15] ), .A(n4197), .ZN(n4191) );
  NOR4_X1 U4139 ( .A1(n4193), .A2(n4194), .A3(n4195), .A4(n4196), .ZN(n4192)
         );
  AOI222_X1 U4140 ( .A1(n1306), .A2(\REGISTERS[38][15] ), .B1(n1303), .B2(
        \REGISTERS[40][15] ), .C1(n1300), .C2(\REGISTERS[39][15] ), .ZN(n4189)
         );
  NAND4_X1 U4141 ( .A1(n5591), .A2(n5592), .A3(n5593), .A4(n5594), .ZN(n5580)
         );
  AOI221_X1 U4142 ( .B1(n618), .B2(\REGISTERS[34][16] ), .C1(n615), .C2(
        \REGISTERS[33][16] ), .A(n5599), .ZN(n5593) );
  NOR4_X1 U4143 ( .A1(n5595), .A2(n5596), .A3(n5597), .A4(n5598), .ZN(n5594)
         );
  AOI222_X1 U4144 ( .A1(n594), .A2(\REGISTERS[38][16] ), .B1(n495), .B2(
        \REGISTERS[40][16] ), .C1(n492), .C2(\REGISTERS[39][16] ), .ZN(n5591)
         );
  NAND4_X1 U4145 ( .A1(n4148), .A2(n4149), .A3(n4150), .A4(n4151), .ZN(n4137)
         );
  AOI221_X1 U4146 ( .B1(n1330), .B2(\REGISTERS[34][16] ), .C1(n1327), .C2(
        \REGISTERS[33][16] ), .A(n4156), .ZN(n4150) );
  NOR4_X1 U4147 ( .A1(n4152), .A2(n4153), .A3(n4154), .A4(n4155), .ZN(n4151)
         );
  AOI222_X1 U4148 ( .A1(n1306), .A2(\REGISTERS[38][16] ), .B1(n1303), .B2(
        \REGISTERS[40][16] ), .C1(n1300), .C2(\REGISTERS[39][16] ), .ZN(n4148)
         );
  NAND4_X1 U4149 ( .A1(n5550), .A2(n5551), .A3(n5552), .A4(n5553), .ZN(n5539)
         );
  AOI221_X1 U4150 ( .B1(n618), .B2(\REGISTERS[34][17] ), .C1(n615), .C2(
        \REGISTERS[33][17] ), .A(n5558), .ZN(n5552) );
  NOR4_X1 U4151 ( .A1(n5554), .A2(n5555), .A3(n5556), .A4(n5557), .ZN(n5553)
         );
  AOI222_X1 U4152 ( .A1(n594), .A2(\REGISTERS[38][17] ), .B1(n495), .B2(
        \REGISTERS[40][17] ), .C1(n492), .C2(\REGISTERS[39][17] ), .ZN(n5550)
         );
  NAND4_X1 U4153 ( .A1(n4107), .A2(n4108), .A3(n4109), .A4(n4110), .ZN(n4096)
         );
  AOI221_X1 U4154 ( .B1(n1330), .B2(\REGISTERS[34][17] ), .C1(n1327), .C2(
        \REGISTERS[33][17] ), .A(n4115), .ZN(n4109) );
  NOR4_X1 U4155 ( .A1(n4111), .A2(n4112), .A3(n4113), .A4(n4114), .ZN(n4110)
         );
  AOI222_X1 U4156 ( .A1(n1306), .A2(\REGISTERS[38][17] ), .B1(n1303), .B2(
        \REGISTERS[40][17] ), .C1(n1300), .C2(\REGISTERS[39][17] ), .ZN(n4107)
         );
  NAND4_X1 U4157 ( .A1(n5509), .A2(n5510), .A3(n5511), .A4(n5512), .ZN(n5498)
         );
  AOI221_X1 U4158 ( .B1(n618), .B2(\REGISTERS[34][18] ), .C1(n615), .C2(
        \REGISTERS[33][18] ), .A(n5517), .ZN(n5511) );
  NOR4_X1 U4159 ( .A1(n5513), .A2(n5514), .A3(n5515), .A4(n5516), .ZN(n5512)
         );
  AOI222_X1 U4160 ( .A1(n594), .A2(\REGISTERS[38][18] ), .B1(n495), .B2(
        \REGISTERS[40][18] ), .C1(n492), .C2(\REGISTERS[39][18] ), .ZN(n5509)
         );
  NAND4_X1 U4161 ( .A1(n4066), .A2(n4067), .A3(n4068), .A4(n4069), .ZN(n4055)
         );
  AOI221_X1 U4162 ( .B1(n1330), .B2(\REGISTERS[34][18] ), .C1(n1327), .C2(
        \REGISTERS[33][18] ), .A(n4074), .ZN(n4068) );
  NOR4_X1 U4163 ( .A1(n4070), .A2(n4071), .A3(n4072), .A4(n4073), .ZN(n4069)
         );
  AOI222_X1 U4164 ( .A1(n1306), .A2(\REGISTERS[38][18] ), .B1(n1303), .B2(
        \REGISTERS[40][18] ), .C1(n1300), .C2(\REGISTERS[39][18] ), .ZN(n4066)
         );
  NAND4_X1 U4165 ( .A1(n5468), .A2(n5469), .A3(n5470), .A4(n5471), .ZN(n5457)
         );
  AOI221_X1 U4166 ( .B1(n618), .B2(\REGISTERS[34][19] ), .C1(n615), .C2(
        \REGISTERS[33][19] ), .A(n5476), .ZN(n5470) );
  NOR4_X1 U4167 ( .A1(n5472), .A2(n5473), .A3(n5474), .A4(n5475), .ZN(n5471)
         );
  AOI222_X1 U4168 ( .A1(n594), .A2(\REGISTERS[38][19] ), .B1(n495), .B2(
        \REGISTERS[40][19] ), .C1(n492), .C2(\REGISTERS[39][19] ), .ZN(n5468)
         );
  NAND4_X1 U4169 ( .A1(n4025), .A2(n4026), .A3(n4027), .A4(n4028), .ZN(n4014)
         );
  AOI221_X1 U4170 ( .B1(n1330), .B2(\REGISTERS[34][19] ), .C1(n1327), .C2(
        \REGISTERS[33][19] ), .A(n4033), .ZN(n4027) );
  NOR4_X1 U4171 ( .A1(n4029), .A2(n4030), .A3(n4031), .A4(n4032), .ZN(n4028)
         );
  AOI222_X1 U4172 ( .A1(n1306), .A2(\REGISTERS[38][19] ), .B1(n1303), .B2(
        \REGISTERS[40][19] ), .C1(n1300), .C2(\REGISTERS[39][19] ), .ZN(n4025)
         );
  NAND4_X1 U4173 ( .A1(n5427), .A2(n5428), .A3(n5429), .A4(n5430), .ZN(n5416)
         );
  AOI221_X1 U4174 ( .B1(n618), .B2(\REGISTERS[34][20] ), .C1(n615), .C2(
        \REGISTERS[33][20] ), .A(n5435), .ZN(n5429) );
  NOR4_X1 U4175 ( .A1(n5431), .A2(n5432), .A3(n5433), .A4(n5434), .ZN(n5430)
         );
  AOI222_X1 U4176 ( .A1(n594), .A2(\REGISTERS[38][20] ), .B1(n494), .B2(
        \REGISTERS[40][20] ), .C1(n491), .C2(\REGISTERS[39][20] ), .ZN(n5427)
         );
  NAND4_X1 U4177 ( .A1(n3984), .A2(n3985), .A3(n3986), .A4(n3987), .ZN(n3973)
         );
  AOI221_X1 U4178 ( .B1(n1330), .B2(\REGISTERS[34][20] ), .C1(n1327), .C2(
        \REGISTERS[33][20] ), .A(n3992), .ZN(n3986) );
  NOR4_X1 U4179 ( .A1(n3988), .A2(n3989), .A3(n3990), .A4(n3991), .ZN(n3987)
         );
  AOI222_X1 U4180 ( .A1(n1306), .A2(\REGISTERS[38][20] ), .B1(n1302), .B2(
        \REGISTERS[40][20] ), .C1(n1299), .C2(\REGISTERS[39][20] ), .ZN(n3984)
         );
  NAND4_X1 U4181 ( .A1(n5386), .A2(n5387), .A3(n5388), .A4(n5389), .ZN(n5375)
         );
  AOI221_X1 U4182 ( .B1(n618), .B2(\REGISTERS[34][21] ), .C1(n615), .C2(
        \REGISTERS[33][21] ), .A(n5394), .ZN(n5388) );
  NOR4_X1 U4183 ( .A1(n5390), .A2(n5391), .A3(n5392), .A4(n5393), .ZN(n5389)
         );
  AOI222_X1 U4184 ( .A1(n594), .A2(\REGISTERS[38][21] ), .B1(n494), .B2(
        \REGISTERS[40][21] ), .C1(n491), .C2(\REGISTERS[39][21] ), .ZN(n5386)
         );
  NAND4_X1 U4185 ( .A1(n3943), .A2(n3944), .A3(n3945), .A4(n3946), .ZN(n3932)
         );
  AOI221_X1 U4186 ( .B1(n1330), .B2(\REGISTERS[34][21] ), .C1(n1327), .C2(
        \REGISTERS[33][21] ), .A(n3951), .ZN(n3945) );
  NOR4_X1 U4187 ( .A1(n3947), .A2(n3948), .A3(n3949), .A4(n3950), .ZN(n3946)
         );
  AOI222_X1 U4188 ( .A1(n1306), .A2(\REGISTERS[38][21] ), .B1(n1302), .B2(
        \REGISTERS[40][21] ), .C1(n1299), .C2(\REGISTERS[39][21] ), .ZN(n3943)
         );
  NAND4_X1 U4189 ( .A1(n5345), .A2(n5346), .A3(n5347), .A4(n5348), .ZN(n5334)
         );
  AOI221_X1 U4190 ( .B1(n618), .B2(\REGISTERS[34][22] ), .C1(n615), .C2(
        \REGISTERS[33][22] ), .A(n5353), .ZN(n5347) );
  NOR4_X1 U4191 ( .A1(n5349), .A2(n5350), .A3(n5351), .A4(n5352), .ZN(n5348)
         );
  AOI222_X1 U4192 ( .A1(n594), .A2(\REGISTERS[38][22] ), .B1(n494), .B2(
        \REGISTERS[40][22] ), .C1(n491), .C2(\REGISTERS[39][22] ), .ZN(n5345)
         );
  NAND4_X1 U4193 ( .A1(n3902), .A2(n3903), .A3(n3904), .A4(n3905), .ZN(n3891)
         );
  AOI221_X1 U4194 ( .B1(n1330), .B2(\REGISTERS[34][22] ), .C1(n1327), .C2(
        \REGISTERS[33][22] ), .A(n3910), .ZN(n3904) );
  NOR4_X1 U4195 ( .A1(n3906), .A2(n3907), .A3(n3908), .A4(n3909), .ZN(n3905)
         );
  AOI222_X1 U4196 ( .A1(n1306), .A2(\REGISTERS[38][22] ), .B1(n1302), .B2(
        \REGISTERS[40][22] ), .C1(n1299), .C2(\REGISTERS[39][22] ), .ZN(n3902)
         );
  NAND4_X1 U4197 ( .A1(n5304), .A2(n5305), .A3(n5306), .A4(n5307), .ZN(n5293)
         );
  AOI221_X1 U4198 ( .B1(n618), .B2(\REGISTERS[34][23] ), .C1(n615), .C2(
        \REGISTERS[33][23] ), .A(n5312), .ZN(n5306) );
  NOR4_X1 U4199 ( .A1(n5308), .A2(n5309), .A3(n5310), .A4(n5311), .ZN(n5307)
         );
  AOI222_X1 U4200 ( .A1(n594), .A2(\REGISTERS[38][23] ), .B1(n494), .B2(
        \REGISTERS[40][23] ), .C1(n491), .C2(\REGISTERS[39][23] ), .ZN(n5304)
         );
  NAND4_X1 U4201 ( .A1(n3861), .A2(n3862), .A3(n3863), .A4(n3864), .ZN(n3850)
         );
  AOI221_X1 U4202 ( .B1(n1330), .B2(\REGISTERS[34][23] ), .C1(n1327), .C2(
        \REGISTERS[33][23] ), .A(n3869), .ZN(n3863) );
  NOR4_X1 U4203 ( .A1(n3865), .A2(n3866), .A3(n3867), .A4(n3868), .ZN(n3864)
         );
  AOI222_X1 U4204 ( .A1(n1306), .A2(\REGISTERS[38][23] ), .B1(n1302), .B2(
        \REGISTERS[40][23] ), .C1(n1299), .C2(\REGISTERS[39][23] ), .ZN(n3861)
         );
  NAND4_X1 U4205 ( .A1(n5263), .A2(n5264), .A3(n5265), .A4(n5266), .ZN(n5252)
         );
  AOI221_X1 U4206 ( .B1(n619), .B2(\REGISTERS[34][24] ), .C1(n616), .C2(
        \REGISTERS[33][24] ), .A(n5271), .ZN(n5265) );
  NOR4_X1 U4207 ( .A1(n5267), .A2(n5268), .A3(n5269), .A4(n5270), .ZN(n5266)
         );
  AOI222_X1 U4208 ( .A1(n595), .A2(\REGISTERS[38][24] ), .B1(n494), .B2(
        \REGISTERS[40][24] ), .C1(n491), .C2(\REGISTERS[39][24] ), .ZN(n5263)
         );
  NAND4_X1 U4209 ( .A1(n3820), .A2(n3821), .A3(n3822), .A4(n3823), .ZN(n3809)
         );
  AOI221_X1 U4210 ( .B1(n1331), .B2(\REGISTERS[34][24] ), .C1(n1328), .C2(
        \REGISTERS[33][24] ), .A(n3828), .ZN(n3822) );
  NOR4_X1 U4211 ( .A1(n3824), .A2(n3825), .A3(n3826), .A4(n3827), .ZN(n3823)
         );
  AOI222_X1 U4212 ( .A1(n1307), .A2(\REGISTERS[38][24] ), .B1(n1302), .B2(
        \REGISTERS[40][24] ), .C1(n1299), .C2(\REGISTERS[39][24] ), .ZN(n3820)
         );
  NAND4_X1 U4213 ( .A1(n5222), .A2(n5223), .A3(n5224), .A4(n5225), .ZN(n5211)
         );
  AOI221_X1 U4214 ( .B1(n619), .B2(\REGISTERS[34][25] ), .C1(n616), .C2(
        \REGISTERS[33][25] ), .A(n5230), .ZN(n5224) );
  NOR4_X1 U4215 ( .A1(n5226), .A2(n5227), .A3(n5228), .A4(n5229), .ZN(n5225)
         );
  AOI222_X1 U4216 ( .A1(n595), .A2(\REGISTERS[38][25] ), .B1(n494), .B2(
        \REGISTERS[40][25] ), .C1(n491), .C2(\REGISTERS[39][25] ), .ZN(n5222)
         );
  NAND4_X1 U4217 ( .A1(n3779), .A2(n3780), .A3(n3781), .A4(n3782), .ZN(n3768)
         );
  AOI221_X1 U4218 ( .B1(n1331), .B2(\REGISTERS[34][25] ), .C1(n1328), .C2(
        \REGISTERS[33][25] ), .A(n3787), .ZN(n3781) );
  NOR4_X1 U4219 ( .A1(n3783), .A2(n3784), .A3(n3785), .A4(n3786), .ZN(n3782)
         );
  AOI222_X1 U4220 ( .A1(n1307), .A2(\REGISTERS[38][25] ), .B1(n1302), .B2(
        \REGISTERS[40][25] ), .C1(n1299), .C2(\REGISTERS[39][25] ), .ZN(n3779)
         );
  NAND4_X1 U4221 ( .A1(n5181), .A2(n5182), .A3(n5183), .A4(n5184), .ZN(n5170)
         );
  AOI221_X1 U4222 ( .B1(n619), .B2(\REGISTERS[34][26] ), .C1(n616), .C2(
        \REGISTERS[33][26] ), .A(n5189), .ZN(n5183) );
  NOR4_X1 U4223 ( .A1(n5185), .A2(n5186), .A3(n5187), .A4(n5188), .ZN(n5184)
         );
  AOI222_X1 U4224 ( .A1(n595), .A2(\REGISTERS[38][26] ), .B1(n494), .B2(
        \REGISTERS[40][26] ), .C1(n491), .C2(\REGISTERS[39][26] ), .ZN(n5181)
         );
  NAND4_X1 U4225 ( .A1(n3738), .A2(n3739), .A3(n3740), .A4(n3741), .ZN(n3727)
         );
  AOI221_X1 U4226 ( .B1(n1331), .B2(\REGISTERS[34][26] ), .C1(n1328), .C2(
        \REGISTERS[33][26] ), .A(n3746), .ZN(n3740) );
  NOR4_X1 U4227 ( .A1(n3742), .A2(n3743), .A3(n3744), .A4(n3745), .ZN(n3741)
         );
  AOI222_X1 U4228 ( .A1(n1307), .A2(\REGISTERS[38][26] ), .B1(n1302), .B2(
        \REGISTERS[40][26] ), .C1(n1299), .C2(\REGISTERS[39][26] ), .ZN(n3738)
         );
  NAND4_X1 U4229 ( .A1(n5140), .A2(n5141), .A3(n5142), .A4(n5143), .ZN(n5129)
         );
  AOI221_X1 U4230 ( .B1(n619), .B2(\REGISTERS[34][27] ), .C1(n616), .C2(
        \REGISTERS[33][27] ), .A(n5148), .ZN(n5142) );
  NOR4_X1 U4231 ( .A1(n5144), .A2(n5145), .A3(n5146), .A4(n5147), .ZN(n5143)
         );
  AOI222_X1 U4232 ( .A1(n595), .A2(\REGISTERS[38][27] ), .B1(n494), .B2(
        \REGISTERS[40][27] ), .C1(n491), .C2(\REGISTERS[39][27] ), .ZN(n5140)
         );
  NAND4_X1 U4233 ( .A1(n3697), .A2(n3698), .A3(n3699), .A4(n3700), .ZN(n3686)
         );
  AOI221_X1 U4234 ( .B1(n1331), .B2(\REGISTERS[34][27] ), .C1(n1328), .C2(
        \REGISTERS[33][27] ), .A(n3705), .ZN(n3699) );
  NOR4_X1 U4235 ( .A1(n3701), .A2(n3702), .A3(n3703), .A4(n3704), .ZN(n3700)
         );
  AOI222_X1 U4236 ( .A1(n1307), .A2(\REGISTERS[38][27] ), .B1(n1302), .B2(
        \REGISTERS[40][27] ), .C1(n1299), .C2(\REGISTERS[39][27] ), .ZN(n3697)
         );
  NAND4_X1 U4237 ( .A1(n5099), .A2(n5100), .A3(n5101), .A4(n5102), .ZN(n5088)
         );
  AOI221_X1 U4238 ( .B1(n619), .B2(\REGISTERS[34][28] ), .C1(n616), .C2(
        \REGISTERS[33][28] ), .A(n5107), .ZN(n5101) );
  NOR4_X1 U4239 ( .A1(n5103), .A2(n5104), .A3(n5105), .A4(n5106), .ZN(n5102)
         );
  AOI222_X1 U4240 ( .A1(n595), .A2(\REGISTERS[38][28] ), .B1(n494), .B2(
        \REGISTERS[40][28] ), .C1(n491), .C2(\REGISTERS[39][28] ), .ZN(n5099)
         );
  NAND4_X1 U4241 ( .A1(n3656), .A2(n3657), .A3(n3658), .A4(n3659), .ZN(n3645)
         );
  AOI221_X1 U4242 ( .B1(n1331), .B2(\REGISTERS[34][28] ), .C1(n1328), .C2(
        \REGISTERS[33][28] ), .A(n3664), .ZN(n3658) );
  NOR4_X1 U4243 ( .A1(n3660), .A2(n3661), .A3(n3662), .A4(n3663), .ZN(n3659)
         );
  AOI222_X1 U4244 ( .A1(n1307), .A2(\REGISTERS[38][28] ), .B1(n1302), .B2(
        \REGISTERS[40][28] ), .C1(n1299), .C2(\REGISTERS[39][28] ), .ZN(n3656)
         );
  NAND4_X1 U4245 ( .A1(n5058), .A2(n5059), .A3(n5060), .A4(n5061), .ZN(n5047)
         );
  AOI221_X1 U4246 ( .B1(n619), .B2(\REGISTERS[34][29] ), .C1(n616), .C2(
        \REGISTERS[33][29] ), .A(n5066), .ZN(n5060) );
  NOR4_X1 U4247 ( .A1(n5062), .A2(n5063), .A3(n5064), .A4(n5065), .ZN(n5061)
         );
  AOI222_X1 U4248 ( .A1(n595), .A2(\REGISTERS[38][29] ), .B1(n494), .B2(
        \REGISTERS[40][29] ), .C1(n491), .C2(\REGISTERS[39][29] ), .ZN(n5058)
         );
  NAND4_X1 U4249 ( .A1(n3615), .A2(n3616), .A3(n3617), .A4(n3618), .ZN(n3604)
         );
  AOI221_X1 U4250 ( .B1(n1331), .B2(\REGISTERS[34][29] ), .C1(n1328), .C2(
        \REGISTERS[33][29] ), .A(n3623), .ZN(n3617) );
  NOR4_X1 U4251 ( .A1(n3619), .A2(n3620), .A3(n3621), .A4(n3622), .ZN(n3618)
         );
  AOI222_X1 U4252 ( .A1(n1307), .A2(\REGISTERS[38][29] ), .B1(n1302), .B2(
        \REGISTERS[40][29] ), .C1(n1299), .C2(\REGISTERS[39][29] ), .ZN(n3615)
         );
  NAND4_X1 U4253 ( .A1(n5017), .A2(n5018), .A3(n5019), .A4(n5020), .ZN(n5006)
         );
  AOI221_X1 U4254 ( .B1(n619), .B2(\REGISTERS[34][30] ), .C1(n616), .C2(
        \REGISTERS[33][30] ), .A(n5025), .ZN(n5019) );
  NOR4_X1 U4255 ( .A1(n5021), .A2(n5022), .A3(n5023), .A4(n5024), .ZN(n5020)
         );
  AOI222_X1 U4256 ( .A1(n595), .A2(\REGISTERS[38][30] ), .B1(n494), .B2(
        \REGISTERS[40][30] ), .C1(n491), .C2(\REGISTERS[39][30] ), .ZN(n5017)
         );
  NAND4_X1 U4257 ( .A1(n3574), .A2(n3575), .A3(n3576), .A4(n3577), .ZN(n3563)
         );
  AOI221_X1 U4258 ( .B1(n1331), .B2(\REGISTERS[34][30] ), .C1(n1328), .C2(
        \REGISTERS[33][30] ), .A(n3582), .ZN(n3576) );
  NOR4_X1 U4259 ( .A1(n3578), .A2(n3579), .A3(n3580), .A4(n3581), .ZN(n3577)
         );
  AOI222_X1 U4260 ( .A1(n1307), .A2(\REGISTERS[38][30] ), .B1(n1302), .B2(
        \REGISTERS[40][30] ), .C1(n1299), .C2(\REGISTERS[39][30] ), .ZN(n3574)
         );
  NAND4_X1 U4261 ( .A1(n4910), .A2(n4911), .A3(n4912), .A4(n4913), .ZN(n4877)
         );
  AOI221_X1 U4262 ( .B1(n619), .B2(\REGISTERS[34][31] ), .C1(n616), .C2(
        \REGISTERS[33][31] ), .A(n4931), .ZN(n4912) );
  NOR4_X1 U4263 ( .A1(n4914), .A2(n4915), .A3(n4916), .A4(n4917), .ZN(n4913)
         );
  AOI222_X1 U4264 ( .A1(n595), .A2(\REGISTERS[38][31] ), .B1(n494), .B2(
        \REGISTERS[40][31] ), .C1(n491), .C2(\REGISTERS[39][31] ), .ZN(n4910)
         );
  NAND4_X1 U4265 ( .A1(n3467), .A2(n3468), .A3(n3469), .A4(n3470), .ZN(n3434)
         );
  AOI221_X1 U4266 ( .B1(n1331), .B2(\REGISTERS[34][31] ), .C1(n1328), .C2(
        \REGISTERS[33][31] ), .A(n3488), .ZN(n3469) );
  NOR4_X1 U4267 ( .A1(n3471), .A2(n3472), .A3(n3473), .A4(n3474), .ZN(n3470)
         );
  AOI222_X1 U4268 ( .A1(n1307), .A2(\REGISTERS[38][31] ), .B1(n1302), .B2(
        \REGISTERS[40][31] ), .C1(n1299), .C2(\REGISTERS[39][31] ), .ZN(n3467)
         );
  OR2_X1 U4269 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(N8430) );
  OR2_X1 U4270 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(N8574) );
  OR2_X1 U4271 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .ZN(N2166) );
  OR2_X1 U4272 ( .A1(RD1), .A2(n3333), .ZN(N8702) );
  OR2_X1 U4273 ( .A1(RD2), .A2(n3333), .ZN(N8735) );
  CLKBUF_X1 U4306 ( .A(DATAIN[0]), .Z(n1797) );
  CLKBUF_X1 U4307 ( .A(DATAIN[0]), .Z(n1798) );
  CLKBUF_X1 U4308 ( .A(DATAIN[0]), .Z(n1799) );
  CLKBUF_X1 U4309 ( .A(DATAIN[1]), .Z(n1808) );
  CLKBUF_X1 U4310 ( .A(DATAIN[1]), .Z(n1809) );
  CLKBUF_X1 U4311 ( .A(DATAIN[1]), .Z(n1810) );
  CLKBUF_X1 U4312 ( .A(DATAIN[2]), .Z(n1819) );
  CLKBUF_X1 U4313 ( .A(DATAIN[2]), .Z(n1820) );
  CLKBUF_X1 U4314 ( .A(DATAIN[2]), .Z(n1821) );
  CLKBUF_X1 U4315 ( .A(DATAIN[3]), .Z(n1830) );
  CLKBUF_X1 U4316 ( .A(DATAIN[3]), .Z(n1831) );
  CLKBUF_X1 U4317 ( .A(DATAIN[3]), .Z(n1832) );
  CLKBUF_X1 U4318 ( .A(DATAIN[4]), .Z(n2545) );
  CLKBUF_X1 U4319 ( .A(DATAIN[4]), .Z(n2546) );
  CLKBUF_X1 U4320 ( .A(DATAIN[4]), .Z(n2547) );
  CLKBUF_X1 U4321 ( .A(DATAIN[5]), .Z(n2556) );
  CLKBUF_X1 U4322 ( .A(DATAIN[5]), .Z(n2557) );
  CLKBUF_X1 U4323 ( .A(DATAIN[5]), .Z(n2558) );
  CLKBUF_X1 U4324 ( .A(DATAIN[6]), .Z(n2567) );
  CLKBUF_X1 U4325 ( .A(DATAIN[6]), .Z(n2568) );
  CLKBUF_X1 U4326 ( .A(DATAIN[6]), .Z(n2569) );
  CLKBUF_X1 U4327 ( .A(DATAIN[7]), .Z(n2578) );
  CLKBUF_X1 U4328 ( .A(DATAIN[7]), .Z(n2579) );
  CLKBUF_X1 U4329 ( .A(DATAIN[7]), .Z(n2580) );
  CLKBUF_X1 U4330 ( .A(DATAIN[8]), .Z(n2589) );
  CLKBUF_X1 U4331 ( .A(DATAIN[8]), .Z(n2590) );
  CLKBUF_X1 U4332 ( .A(DATAIN[8]), .Z(n2591) );
  CLKBUF_X1 U4333 ( .A(DATAIN[9]), .Z(n2600) );
  CLKBUF_X1 U4334 ( .A(DATAIN[9]), .Z(n2601) );
  CLKBUF_X1 U4335 ( .A(DATAIN[9]), .Z(n2602) );
  CLKBUF_X1 U4336 ( .A(DATAIN[10]), .Z(n2707) );
  CLKBUF_X1 U4337 ( .A(DATAIN[10]), .Z(n2708) );
  CLKBUF_X1 U4338 ( .A(DATAIN[10]), .Z(n2709) );
  CLKBUF_X1 U4339 ( .A(DATAIN[11]), .Z(n2718) );
  CLKBUF_X1 U4340 ( .A(DATAIN[11]), .Z(n2719) );
  CLKBUF_X1 U4341 ( .A(DATAIN[11]), .Z(n2720) );
  CLKBUF_X1 U4342 ( .A(DATAIN[12]), .Z(n2729) );
  CLKBUF_X1 U4343 ( .A(DATAIN[12]), .Z(n2730) );
  CLKBUF_X1 U4344 ( .A(DATAIN[12]), .Z(n2731) );
  CLKBUF_X1 U4345 ( .A(DATAIN[13]), .Z(n2740) );
  CLKBUF_X1 U4346 ( .A(DATAIN[13]), .Z(n2741) );
  CLKBUF_X1 U4347 ( .A(DATAIN[13]), .Z(n2742) );
  CLKBUF_X1 U4348 ( .A(DATAIN[14]), .Z(n2751) );
  CLKBUF_X1 U4349 ( .A(DATAIN[14]), .Z(n2752) );
  CLKBUF_X1 U4350 ( .A(DATAIN[14]), .Z(n2753) );
  CLKBUF_X1 U4351 ( .A(DATAIN[15]), .Z(n2762) );
  CLKBUF_X1 U4352 ( .A(DATAIN[15]), .Z(n2763) );
  CLKBUF_X1 U4353 ( .A(DATAIN[15]), .Z(n2764) );
  CLKBUF_X1 U4354 ( .A(DATAIN[16]), .Z(n2773) );
  CLKBUF_X1 U4355 ( .A(DATAIN[16]), .Z(n2774) );
  CLKBUF_X1 U4356 ( .A(DATAIN[16]), .Z(n2775) );
  CLKBUF_X1 U4357 ( .A(DATAIN[17]), .Z(n2784) );
  CLKBUF_X1 U4358 ( .A(DATAIN[17]), .Z(n2785) );
  CLKBUF_X1 U4359 ( .A(DATAIN[17]), .Z(n2786) );
  CLKBUF_X1 U4360 ( .A(DATAIN[18]), .Z(n2795) );
  CLKBUF_X1 U4361 ( .A(DATAIN[18]), .Z(n2796) );
  CLKBUF_X1 U4362 ( .A(DATAIN[18]), .Z(n2797) );
  CLKBUF_X1 U4363 ( .A(DATAIN[19]), .Z(n2806) );
  CLKBUF_X1 U4364 ( .A(DATAIN[19]), .Z(n2807) );
  CLKBUF_X1 U4365 ( .A(DATAIN[19]), .Z(n2808) );
  CLKBUF_X1 U4366 ( .A(DATAIN[20]), .Z(n2817) );
  CLKBUF_X1 U4367 ( .A(DATAIN[20]), .Z(n2818) );
  CLKBUF_X1 U4368 ( .A(DATAIN[20]), .Z(n2819) );
  CLKBUF_X1 U4369 ( .A(DATAIN[21]), .Z(n2828) );
  CLKBUF_X1 U4370 ( .A(DATAIN[21]), .Z(n2829) );
  CLKBUF_X1 U4371 ( .A(DATAIN[21]), .Z(n2830) );
  CLKBUF_X1 U4372 ( .A(DATAIN[22]), .Z(n2839) );
  CLKBUF_X1 U4373 ( .A(DATAIN[22]), .Z(n2840) );
  CLKBUF_X1 U4374 ( .A(DATAIN[22]), .Z(n2841) );
  CLKBUF_X1 U4375 ( .A(DATAIN[23]), .Z(n2850) );
  CLKBUF_X1 U4376 ( .A(DATAIN[23]), .Z(n2851) );
  CLKBUF_X1 U4377 ( .A(DATAIN[23]), .Z(n2852) );
  CLKBUF_X1 U4378 ( .A(DATAIN[24]), .Z(n2861) );
  CLKBUF_X1 U4379 ( .A(DATAIN[24]), .Z(n2862) );
  CLKBUF_X1 U4380 ( .A(DATAIN[24]), .Z(n2863) );
  CLKBUF_X1 U4381 ( .A(DATAIN[25]), .Z(n2872) );
  CLKBUF_X1 U4382 ( .A(DATAIN[25]), .Z(n2873) );
  CLKBUF_X1 U4383 ( .A(DATAIN[25]), .Z(n2874) );
  CLKBUF_X1 U4384 ( .A(DATAIN[26]), .Z(n2883) );
  CLKBUF_X1 U4385 ( .A(DATAIN[26]), .Z(n2884) );
  CLKBUF_X1 U4386 ( .A(DATAIN[26]), .Z(n2885) );
  CLKBUF_X1 U4387 ( .A(DATAIN[27]), .Z(n2894) );
  CLKBUF_X1 U4388 ( .A(DATAIN[27]), .Z(n2895) );
  CLKBUF_X1 U4389 ( .A(DATAIN[27]), .Z(n2896) );
  CLKBUF_X1 U4390 ( .A(DATAIN[28]), .Z(n2906) );
  CLKBUF_X1 U4391 ( .A(DATAIN[28]), .Z(n2907) );
  CLKBUF_X1 U4392 ( .A(DATAIN[28]), .Z(n2908) );
  CLKBUF_X1 U4393 ( .A(DATAIN[29]), .Z(n2922) );
  CLKBUF_X1 U4394 ( .A(DATAIN[29]), .Z(n2923) );
  CLKBUF_X1 U4395 ( .A(DATAIN[29]), .Z(n2924) );
  CLKBUF_X1 U4396 ( .A(DATAIN[30]), .Z(n2933) );
  CLKBUF_X1 U4397 ( .A(DATAIN[30]), .Z(n2934) );
  CLKBUF_X1 U4398 ( .A(DATAIN[30]), .Z(n2935) );
  CLKBUF_X1 U4399 ( .A(DATAIN[31]), .Z(n2944) );
  CLKBUF_X1 U4400 ( .A(DATAIN[31]), .Z(n2945) );
  CLKBUF_X1 U4401 ( .A(DATAIN[31]), .Z(n2946) );
  INV_X1 U4402 ( .A(n3302), .ZN(n2956) );
  INV_X1 U4403 ( .A(n3301), .ZN(n2957) );
  INV_X1 U4404 ( .A(n3301), .ZN(n2958) );
  INV_X1 U4405 ( .A(n3301), .ZN(n2959) );
  INV_X1 U4406 ( .A(n3301), .ZN(n2960) );
  INV_X1 U4407 ( .A(n3301), .ZN(n2961) );
  INV_X1 U4408 ( .A(n3301), .ZN(n2962) );
  INV_X1 U4409 ( .A(n3301), .ZN(n2963) );
  INV_X1 U4410 ( .A(n3300), .ZN(n2964) );
  INV_X1 U4411 ( .A(n3300), .ZN(n2965) );
  INV_X1 U4412 ( .A(n3300), .ZN(n2966) );
  INV_X1 U4413 ( .A(n3300), .ZN(n2967) );
  INV_X1 U4414 ( .A(n3300), .ZN(n2968) );
  INV_X1 U4415 ( .A(n3300), .ZN(n2969) );
  INV_X1 U4416 ( .A(n3300), .ZN(n2970) );
  INV_X1 U4417 ( .A(n3298), .ZN(n2971) );
  INV_X1 U4418 ( .A(n3298), .ZN(n2972) );
  INV_X1 U4419 ( .A(n3298), .ZN(n2973) );
  INV_X1 U4420 ( .A(n3298), .ZN(n2974) );
  INV_X1 U4421 ( .A(n3298), .ZN(n2975) );
  INV_X1 U4422 ( .A(n3298), .ZN(n2976) );
  INV_X1 U4423 ( .A(n3298), .ZN(n2977) );
  INV_X1 U4424 ( .A(n3297), .ZN(n2978) );
  INV_X1 U4425 ( .A(n3297), .ZN(n2979) );
  INV_X1 U4426 ( .A(n3297), .ZN(n2980) );
  INV_X1 U4427 ( .A(n3297), .ZN(n2981) );
  INV_X1 U4428 ( .A(n3297), .ZN(n2982) );
  INV_X1 U4429 ( .A(n3297), .ZN(n2983) );
  INV_X1 U4430 ( .A(n3297), .ZN(n2984) );
  INV_X1 U4431 ( .A(n3296), .ZN(n2985) );
  INV_X1 U4432 ( .A(n3296), .ZN(n2986) );
  INV_X1 U4433 ( .A(n3296), .ZN(n2987) );
  INV_X1 U4434 ( .A(n3296), .ZN(n2988) );
  INV_X1 U4435 ( .A(n3296), .ZN(n2989) );
  INV_X1 U4436 ( .A(n3296), .ZN(n2990) );
  INV_X1 U4437 ( .A(n3296), .ZN(n2991) );
  INV_X1 U4438 ( .A(n3294), .ZN(n2992) );
  INV_X1 U4439 ( .A(n3294), .ZN(n2993) );
  INV_X1 U4440 ( .A(n3294), .ZN(n2994) );
  INV_X1 U4441 ( .A(n3294), .ZN(n2995) );
  INV_X1 U4442 ( .A(n3294), .ZN(n2997) );
  INV_X1 U4443 ( .A(n3294), .ZN(n2998) );
  INV_X1 U4444 ( .A(n3293), .ZN(n2999) );
  INV_X1 U4445 ( .A(n3293), .ZN(n3000) );
  INV_X1 U4446 ( .A(n3293), .ZN(n3001) );
  INV_X1 U4447 ( .A(n3293), .ZN(n3002) );
  INV_X1 U4448 ( .A(n3293), .ZN(n3003) );
  INV_X1 U4449 ( .A(n3293), .ZN(n3004) );
  INV_X1 U4450 ( .A(n3293), .ZN(n3005) );
  INV_X1 U4451 ( .A(n3292), .ZN(n3006) );
  INV_X1 U4452 ( .A(n3292), .ZN(n3007) );
  INV_X1 U4453 ( .A(n3292), .ZN(n3008) );
  INV_X1 U4454 ( .A(n3292), .ZN(n3009) );
  INV_X1 U4455 ( .A(n3292), .ZN(n3010) );
  INV_X1 U4456 ( .A(n3292), .ZN(n3011) );
  INV_X1 U4457 ( .A(n3292), .ZN(n3012) );
  INV_X1 U4458 ( .A(n3290), .ZN(n3013) );
  INV_X1 U4459 ( .A(n3290), .ZN(n3014) );
  INV_X1 U4460 ( .A(n3290), .ZN(n3015) );
  INV_X1 U4461 ( .A(n3290), .ZN(n3016) );
  INV_X1 U4462 ( .A(n3290), .ZN(n3017) );
  INV_X1 U4463 ( .A(n3290), .ZN(n3018) );
  INV_X1 U4464 ( .A(n3290), .ZN(n3019) );
  INV_X1 U4465 ( .A(n3289), .ZN(n3020) );
  INV_X1 U4466 ( .A(n3289), .ZN(n3021) );
  INV_X1 U4467 ( .A(n3289), .ZN(n3022) );
  INV_X1 U4468 ( .A(n3289), .ZN(n3023) );
  INV_X1 U4469 ( .A(n3289), .ZN(n3024) );
  INV_X1 U4470 ( .A(n3289), .ZN(n3025) );
  INV_X1 U4471 ( .A(n3288), .ZN(n3026) );
  INV_X1 U4472 ( .A(n3288), .ZN(n3027) );
  INV_X1 U4473 ( .A(n3288), .ZN(n3028) );
  INV_X1 U4474 ( .A(n3288), .ZN(n3031) );
  INV_X1 U4475 ( .A(n3288), .ZN(n3032) );
  INV_X1 U4476 ( .A(n3288), .ZN(n3034) );
  INV_X1 U4477 ( .A(n3288), .ZN(n3036) );
  INV_X1 U4478 ( .A(n3286), .ZN(n3037) );
  INV_X1 U4479 ( .A(n3286), .ZN(n3039) );
  INV_X1 U4480 ( .A(n3286), .ZN(n3041) );
  INV_X1 U4481 ( .A(n3286), .ZN(n3042) );
  INV_X1 U4482 ( .A(n3286), .ZN(n3044) );
  INV_X1 U4483 ( .A(n3286), .ZN(n3046) );
  INV_X1 U4484 ( .A(n3294), .ZN(n3047) );
  INV_X1 U4485 ( .A(n3331), .ZN(n3049) );
  INV_X1 U4486 ( .A(n3331), .ZN(n3051) );
  INV_X1 U4487 ( .A(n3331), .ZN(n3052) );
  INV_X1 U4488 ( .A(n3331), .ZN(n3054) );
  INV_X1 U4489 ( .A(n3331), .ZN(n3056) );
  INV_X1 U4490 ( .A(n3331), .ZN(n3057) );
  INV_X1 U4491 ( .A(n3330), .ZN(n3059) );
  INV_X1 U4492 ( .A(n3331), .ZN(n3061) );
  INV_X1 U4493 ( .A(n3330), .ZN(n3062) );
  INV_X1 U4494 ( .A(n3330), .ZN(n3064) );
  INV_X1 U4495 ( .A(n3330), .ZN(n3066) );
  INV_X1 U4496 ( .A(n3330), .ZN(n3067) );
  INV_X1 U4497 ( .A(n3330), .ZN(n3069) );
  INV_X1 U4498 ( .A(n3330), .ZN(n3071) );
  INV_X1 U4499 ( .A(n3329), .ZN(n3072) );
  INV_X1 U4500 ( .A(n3329), .ZN(n3074) );
  INV_X1 U4501 ( .A(n3329), .ZN(n3076) );
  INV_X1 U4502 ( .A(n3329), .ZN(n3077) );
  INV_X1 U4503 ( .A(n3329), .ZN(n3079) );
  INV_X1 U4504 ( .A(n3329), .ZN(n3081) );
  INV_X1 U4505 ( .A(n3327), .ZN(n3082) );
  INV_X1 U4506 ( .A(n3329), .ZN(n3084) );
  INV_X1 U4507 ( .A(n3327), .ZN(n3086) );
  INV_X1 U4508 ( .A(n3327), .ZN(n3087) );
  INV_X1 U4509 ( .A(n3327), .ZN(n3089) );
  INV_X1 U4510 ( .A(n3327), .ZN(n3091) );
  INV_X1 U4511 ( .A(n3327), .ZN(n3092) );
  INV_X1 U4512 ( .A(n3327), .ZN(n3094) );
  INV_X1 U4513 ( .A(n3326), .ZN(n3096) );
  INV_X1 U4514 ( .A(n3326), .ZN(n3097) );
  INV_X1 U4515 ( .A(n3326), .ZN(n3099) );
  INV_X1 U4516 ( .A(n3326), .ZN(n3101) );
  INV_X1 U4517 ( .A(n3326), .ZN(n3102) );
  INV_X1 U4518 ( .A(n3326), .ZN(n3104) );
  INV_X1 U4519 ( .A(n3326), .ZN(n3110) );
  INV_X1 U4520 ( .A(n3325), .ZN(n3111) );
  INV_X1 U4521 ( .A(n3325), .ZN(n3113) );
  INV_X1 U4522 ( .A(n3325), .ZN(n3115) );
  INV_X1 U4523 ( .A(n3325), .ZN(n3116) );
  INV_X1 U4524 ( .A(n3325), .ZN(n3118) );
  INV_X1 U4525 ( .A(n3325), .ZN(n3119) );
  INV_X1 U4526 ( .A(n3325), .ZN(n3120) );
  INV_X1 U4527 ( .A(n3323), .ZN(n3122) );
  INV_X1 U4528 ( .A(n3323), .ZN(n3123) );
  INV_X1 U4529 ( .A(n3323), .ZN(n3124) );
  INV_X1 U4530 ( .A(n3323), .ZN(n3126) );
  INV_X1 U4531 ( .A(n3323), .ZN(n3127) );
  INV_X1 U4532 ( .A(n3323), .ZN(n3128) );
  INV_X1 U4533 ( .A(n3323), .ZN(n3130) );
  INV_X1 U4534 ( .A(n3322), .ZN(n3131) );
  INV_X1 U4535 ( .A(n3322), .ZN(n3132) );
  INV_X1 U4536 ( .A(n3322), .ZN(n3134) );
  INV_X1 U4537 ( .A(n3322), .ZN(n3135) );
  INV_X1 U4538 ( .A(n3322), .ZN(n3136) );
  INV_X1 U4539 ( .A(n3322), .ZN(n3138) );
  INV_X1 U4540 ( .A(n3322), .ZN(n3139) );
  INV_X1 U4541 ( .A(n3321), .ZN(n3140) );
  INV_X1 U4542 ( .A(n3321), .ZN(n3142) );
  INV_X1 U4543 ( .A(n3321), .ZN(n3143) );
  INV_X1 U4544 ( .A(n3321), .ZN(n3144) );
  INV_X1 U4545 ( .A(n3321), .ZN(n3146) );
  INV_X1 U4546 ( .A(n3321), .ZN(n3147) );
  INV_X1 U4547 ( .A(n3321), .ZN(n3148) );
  INV_X1 U4548 ( .A(n3319), .ZN(n3150) );
  INV_X1 U4549 ( .A(n3319), .ZN(n3151) );
  INV_X1 U4550 ( .A(n3319), .ZN(n3152) );
  INV_X1 U4551 ( .A(n3319), .ZN(n3154) );
  INV_X1 U4552 ( .A(n3319), .ZN(n3155) );
  INV_X1 U4553 ( .A(n3319), .ZN(n3156) );
  INV_X1 U4554 ( .A(n3319), .ZN(n3158) );
  INV_X1 U4555 ( .A(n3318), .ZN(n3159) );
  INV_X1 U4556 ( .A(n3318), .ZN(n3160) );
  INV_X1 U4557 ( .A(n3318), .ZN(n3162) );
  INV_X1 U4558 ( .A(n3318), .ZN(n3163) );
  INV_X1 U4559 ( .A(n3318), .ZN(n3164) );
  INV_X1 U4560 ( .A(n3318), .ZN(n3166) );
  INV_X1 U4561 ( .A(n3317), .ZN(n3167) );
  INV_X1 U4562 ( .A(n3317), .ZN(n3168) );
  INV_X1 U4563 ( .A(n3317), .ZN(n3170) );
  INV_X1 U4564 ( .A(n3317), .ZN(n3171) );
  INV_X1 U4565 ( .A(n3317), .ZN(n3172) );
  INV_X1 U4566 ( .A(n3317), .ZN(n3174) );
  INV_X1 U4567 ( .A(n3317), .ZN(n3175) );
  INV_X1 U4568 ( .A(n3315), .ZN(n3176) );
  INV_X1 U4569 ( .A(n3315), .ZN(n3178) );
  INV_X1 U4570 ( .A(n3315), .ZN(n3180) );
  INV_X1 U4571 ( .A(n3315), .ZN(n3181) );
  INV_X1 U4572 ( .A(n3315), .ZN(n3183) );
  INV_X1 U4573 ( .A(n3315), .ZN(n3184) );
  INV_X1 U4574 ( .A(n3315), .ZN(n3185) );
  INV_X1 U4575 ( .A(n3314), .ZN(n3187) );
  INV_X1 U4576 ( .A(n3314), .ZN(n3188) );
  INV_X1 U4577 ( .A(n3314), .ZN(n3189) );
  INV_X1 U4578 ( .A(n3314), .ZN(n3191) );
  INV_X1 U4579 ( .A(n3314), .ZN(n3192) );
  INV_X1 U4580 ( .A(n3314), .ZN(n3193) );
  INV_X1 U4581 ( .A(n3314), .ZN(n3195) );
  INV_X1 U4582 ( .A(n3313), .ZN(n3196) );
  INV_X1 U4583 ( .A(n3313), .ZN(n3197) );
  INV_X1 U4584 ( .A(n3313), .ZN(n3199) );
  INV_X1 U4585 ( .A(n3313), .ZN(n3200) );
  INV_X1 U4586 ( .A(n3313), .ZN(n3201) );
  INV_X1 U4587 ( .A(n3313), .ZN(n3203) );
  INV_X1 U4588 ( .A(n3313), .ZN(n3204) );
  INV_X1 U4589 ( .A(n3311), .ZN(n3205) );
  INV_X1 U4590 ( .A(n3311), .ZN(n3207) );
  INV_X1 U4591 ( .A(n3311), .ZN(n3208) );
  INV_X1 U4592 ( .A(n3311), .ZN(n3209) );
  INV_X1 U4593 ( .A(n3311), .ZN(n3211) );
  INV_X1 U4594 ( .A(n3311), .ZN(n3212) );
  INV_X1 U4595 ( .A(n3311), .ZN(n3213) );
  INV_X1 U4596 ( .A(n3310), .ZN(n3215) );
  INV_X1 U4597 ( .A(n3310), .ZN(n3216) );
  INV_X1 U4598 ( .A(n3310), .ZN(n3217) );
  INV_X1 U4599 ( .A(n3310), .ZN(n3219) );
  INV_X1 U4600 ( .A(n3310), .ZN(n3220) );
  INV_X1 U4601 ( .A(n3310), .ZN(n3221) );
  INV_X1 U4602 ( .A(n3310), .ZN(n3223) );
  INV_X1 U4603 ( .A(n3308), .ZN(n3224) );
  INV_X1 U4604 ( .A(n3308), .ZN(n3225) );
  INV_X1 U4605 ( .A(n3308), .ZN(n3227) );
  INV_X1 U4606 ( .A(n3308), .ZN(n3228) );
  INV_X1 U4607 ( .A(n3308), .ZN(n3229) );
  INV_X1 U4608 ( .A(n3308), .ZN(n3231) );
  INV_X1 U4609 ( .A(n3308), .ZN(n3232) );
  INV_X1 U4610 ( .A(n3306), .ZN(n3233) );
  INV_X1 U4611 ( .A(n3306), .ZN(n3235) );
  INV_X1 U4612 ( .A(n3306), .ZN(n3236) );
  INV_X1 U4613 ( .A(n3306), .ZN(n3237) );
  INV_X1 U4614 ( .A(n3306), .ZN(n3239) );
  INV_X1 U4615 ( .A(n3306), .ZN(n3240) );
  INV_X1 U4616 ( .A(n3306), .ZN(n3241) );
  INV_X1 U4617 ( .A(n3305), .ZN(n3243) );
  INV_X1 U4618 ( .A(n3305), .ZN(n3245) );
  INV_X1 U4619 ( .A(n3305), .ZN(n3246) );
  INV_X1 U4620 ( .A(n3305), .ZN(n3248) );
  INV_X1 U4621 ( .A(n3305), .ZN(n3249) );
  INV_X1 U4622 ( .A(n3305), .ZN(n3250) );
  INV_X1 U4623 ( .A(n3305), .ZN(n3252) );
  INV_X1 U4624 ( .A(n3304), .ZN(n3253) );
  INV_X1 U4625 ( .A(n3304), .ZN(n3254) );
  INV_X1 U4626 ( .A(n3304), .ZN(n3256) );
  INV_X1 U4627 ( .A(n3304), .ZN(n3257) );
  INV_X1 U4628 ( .A(n3304), .ZN(n3258) );
  INV_X1 U4629 ( .A(n3304), .ZN(n3260) );
  INV_X1 U4630 ( .A(n3304), .ZN(n3261) );
  INV_X1 U4631 ( .A(n3318), .ZN(n3262) );
  INV_X1 U4632 ( .A(n3286), .ZN(n3264) );
  NAND2_X1 U4633 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .ZN(N2151) );
  NAND2_X1 U4634 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(N8415) );
  NAND2_X1 U4635 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(N8559) );
  MUX2_X1 U4636 ( .A(\REGISTERS[87][31] ), .B(n2947), .S(n1431), .Z(n9101) );
  MUX2_X1 U4637 ( .A(\REGISTERS[87][30] ), .B(n2936), .S(n1431), .Z(n9102) );
  MUX2_X1 U4638 ( .A(\REGISTERS[87][29] ), .B(n2925), .S(n1431), .Z(n9103) );
  MUX2_X1 U4639 ( .A(\REGISTERS[87][28] ), .B(n2909), .S(n1431), .Z(n9104) );
  MUX2_X1 U4640 ( .A(\REGISTERS[87][27] ), .B(n2897), .S(n1431), .Z(n9105) );
  MUX2_X1 U4641 ( .A(\REGISTERS[87][26] ), .B(n2886), .S(n1431), .Z(n9106) );
  MUX2_X1 U4642 ( .A(\REGISTERS[87][25] ), .B(n2875), .S(n1431), .Z(n9107) );
  MUX2_X1 U4643 ( .A(\REGISTERS[87][24] ), .B(n2864), .S(n1431), .Z(n9108) );
  MUX2_X1 U4644 ( .A(\REGISTERS[87][23] ), .B(n2853), .S(n1431), .Z(n9109) );
  MUX2_X1 U4645 ( .A(\REGISTERS[87][22] ), .B(n2842), .S(n1431), .Z(n9110) );
  MUX2_X1 U4646 ( .A(\REGISTERS[87][21] ), .B(n2831), .S(n1431), .Z(n9111) );
  MUX2_X1 U4647 ( .A(\REGISTERS[87][20] ), .B(n2820), .S(n1431), .Z(n9112) );
  MUX2_X1 U4648 ( .A(\REGISTERS[87][19] ), .B(n2809), .S(n1432), .Z(n9113) );
  MUX2_X1 U4649 ( .A(\REGISTERS[87][18] ), .B(n2798), .S(n1432), .Z(n9114) );
  MUX2_X1 U4650 ( .A(\REGISTERS[87][17] ), .B(n2787), .S(n1432), .Z(n9115) );
  MUX2_X1 U4651 ( .A(\REGISTERS[87][16] ), .B(n2776), .S(n1432), .Z(n9116) );
  MUX2_X1 U4652 ( .A(\REGISTERS[87][15] ), .B(n2765), .S(n1432), .Z(n9117) );
  MUX2_X1 U4653 ( .A(\REGISTERS[87][14] ), .B(n2754), .S(n1432), .Z(n9118) );
  MUX2_X1 U4654 ( .A(\REGISTERS[87][13] ), .B(n2743), .S(n1432), .Z(n9119) );
  MUX2_X1 U4655 ( .A(\REGISTERS[87][12] ), .B(n2732), .S(n1432), .Z(n9120) );
  MUX2_X1 U4656 ( .A(\REGISTERS[87][11] ), .B(n2721), .S(n1432), .Z(n9121) );
  MUX2_X1 U4657 ( .A(\REGISTERS[87][10] ), .B(n2710), .S(n1432), .Z(n9122) );
  MUX2_X1 U4658 ( .A(\REGISTERS[87][9] ), .B(n2603), .S(n1432), .Z(n9123) );
  MUX2_X1 U4659 ( .A(\REGISTERS[87][8] ), .B(n2592), .S(n1432), .Z(n9124) );
  MUX2_X1 U4660 ( .A(\REGISTERS[87][7] ), .B(n2581), .S(n1433), .Z(n9125) );
  MUX2_X1 U4661 ( .A(\REGISTERS[87][6] ), .B(n2570), .S(n1433), .Z(n9126) );
  MUX2_X1 U4662 ( .A(\REGISTERS[87][5] ), .B(n2559), .S(n1433), .Z(n9127) );
  MUX2_X1 U4663 ( .A(\REGISTERS[87][4] ), .B(n2548), .S(n1433), .Z(n9128) );
  MUX2_X1 U4664 ( .A(\REGISTERS[87][3] ), .B(n1833), .S(n1433), .Z(n9129) );
  MUX2_X1 U4665 ( .A(\REGISTERS[87][2] ), .B(n1822), .S(n1433), .Z(n9130) );
  MUX2_X1 U4666 ( .A(\REGISTERS[87][1] ), .B(n1811), .S(n1433), .Z(n9131) );
  MUX2_X1 U4667 ( .A(\REGISTERS[87][0] ), .B(n1800), .S(n1433), .Z(n9132) );
  MUX2_X1 U4668 ( .A(\REGISTERS[86][31] ), .B(n2947), .S(n1434), .Z(n9069) );
  MUX2_X1 U4669 ( .A(\REGISTERS[86][30] ), .B(n2936), .S(n1434), .Z(n9070) );
  MUX2_X1 U4670 ( .A(\REGISTERS[86][29] ), .B(n2925), .S(n1434), .Z(n9071) );
  MUX2_X1 U4671 ( .A(\REGISTERS[86][28] ), .B(n2909), .S(n1434), .Z(n9072) );
  MUX2_X1 U4672 ( .A(\REGISTERS[86][27] ), .B(n2897), .S(n1434), .Z(n9073) );
  MUX2_X1 U4673 ( .A(\REGISTERS[86][26] ), .B(n2886), .S(n1434), .Z(n9074) );
  MUX2_X1 U4674 ( .A(\REGISTERS[86][25] ), .B(n2875), .S(n1434), .Z(n9075) );
  MUX2_X1 U4675 ( .A(\REGISTERS[86][24] ), .B(n2864), .S(n1434), .Z(n9076) );
  MUX2_X1 U4676 ( .A(\REGISTERS[86][23] ), .B(n2853), .S(n1434), .Z(n9077) );
  MUX2_X1 U4677 ( .A(\REGISTERS[86][22] ), .B(n2842), .S(n1434), .Z(n9078) );
  MUX2_X1 U4678 ( .A(\REGISTERS[86][21] ), .B(n2831), .S(n1434), .Z(n9079) );
  MUX2_X1 U4679 ( .A(\REGISTERS[86][20] ), .B(n2820), .S(n1434), .Z(n9080) );
  MUX2_X1 U4680 ( .A(\REGISTERS[86][19] ), .B(n2809), .S(n1435), .Z(n9081) );
  MUX2_X1 U4681 ( .A(\REGISTERS[86][18] ), .B(n2798), .S(n1435), .Z(n9082) );
  MUX2_X1 U4682 ( .A(\REGISTERS[86][17] ), .B(n2787), .S(n1435), .Z(n9083) );
  MUX2_X1 U4683 ( .A(\REGISTERS[86][16] ), .B(n2776), .S(n1435), .Z(n9084) );
  MUX2_X1 U4684 ( .A(\REGISTERS[86][15] ), .B(n2765), .S(n1435), .Z(n9085) );
  MUX2_X1 U4685 ( .A(\REGISTERS[86][14] ), .B(n2754), .S(n1435), .Z(n9086) );
  MUX2_X1 U4686 ( .A(\REGISTERS[86][13] ), .B(n2743), .S(n1435), .Z(n9087) );
  MUX2_X1 U4687 ( .A(\REGISTERS[86][12] ), .B(n2732), .S(n1435), .Z(n9088) );
  MUX2_X1 U4688 ( .A(\REGISTERS[86][11] ), .B(n2721), .S(n1435), .Z(n9089) );
  MUX2_X1 U4689 ( .A(\REGISTERS[86][10] ), .B(n2710), .S(n1435), .Z(n9090) );
  MUX2_X1 U4690 ( .A(\REGISTERS[86][9] ), .B(n2603), .S(n1435), .Z(n9091) );
  MUX2_X1 U4691 ( .A(\REGISTERS[86][8] ), .B(n2592), .S(n1435), .Z(n9092) );
  MUX2_X1 U4692 ( .A(\REGISTERS[86][7] ), .B(n2581), .S(n1436), .Z(n9093) );
  MUX2_X1 U4693 ( .A(\REGISTERS[86][6] ), .B(n2570), .S(n1436), .Z(n9094) );
  MUX2_X1 U4694 ( .A(\REGISTERS[86][5] ), .B(n2559), .S(n1436), .Z(n9095) );
  MUX2_X1 U4695 ( .A(\REGISTERS[86][4] ), .B(n2548), .S(n1436), .Z(n9096) );
  MUX2_X1 U4696 ( .A(\REGISTERS[86][3] ), .B(n1833), .S(n1436), .Z(n9097) );
  MUX2_X1 U4697 ( .A(\REGISTERS[86][2] ), .B(n1822), .S(n1436), .Z(n9098) );
  MUX2_X1 U4698 ( .A(\REGISTERS[86][1] ), .B(n1811), .S(n1436), .Z(n9099) );
  MUX2_X1 U4699 ( .A(\REGISTERS[86][0] ), .B(n1800), .S(n1436), .Z(n9100) );
  MUX2_X1 U4700 ( .A(\REGISTERS[85][31] ), .B(n2947), .S(n1437), .Z(n9037) );
  MUX2_X1 U4701 ( .A(\REGISTERS[85][30] ), .B(n2936), .S(n1437), .Z(n9038) );
  MUX2_X1 U4702 ( .A(\REGISTERS[85][29] ), .B(n2925), .S(n1437), .Z(n9039) );
  MUX2_X1 U4703 ( .A(\REGISTERS[85][28] ), .B(n2909), .S(n1437), .Z(n9040) );
  MUX2_X1 U4704 ( .A(\REGISTERS[85][27] ), .B(n2897), .S(n1437), .Z(n9041) );
  MUX2_X1 U4705 ( .A(\REGISTERS[85][26] ), .B(n2886), .S(n1437), .Z(n9042) );
  MUX2_X1 U4706 ( .A(\REGISTERS[85][25] ), .B(n2875), .S(n1437), .Z(n9043) );
  MUX2_X1 U4707 ( .A(\REGISTERS[85][24] ), .B(n2864), .S(n1437), .Z(n9044) );
  MUX2_X1 U4708 ( .A(\REGISTERS[85][23] ), .B(n2853), .S(n1437), .Z(n9045) );
  MUX2_X1 U4709 ( .A(\REGISTERS[85][22] ), .B(n2842), .S(n1437), .Z(n9046) );
  MUX2_X1 U4710 ( .A(\REGISTERS[85][21] ), .B(n2831), .S(n1437), .Z(n9047) );
  MUX2_X1 U4711 ( .A(\REGISTERS[85][20] ), .B(n2820), .S(n1437), .Z(n9048) );
  MUX2_X1 U4712 ( .A(\REGISTERS[85][19] ), .B(n2809), .S(n1438), .Z(n9049) );
  MUX2_X1 U4713 ( .A(\REGISTERS[85][18] ), .B(n2798), .S(n1438), .Z(n9050) );
  MUX2_X1 U4714 ( .A(\REGISTERS[85][17] ), .B(n2787), .S(n1438), .Z(n9051) );
  MUX2_X1 U4715 ( .A(\REGISTERS[85][16] ), .B(n2776), .S(n1438), .Z(n9052) );
  MUX2_X1 U4716 ( .A(\REGISTERS[85][15] ), .B(n2765), .S(n1438), .Z(n9053) );
  MUX2_X1 U4717 ( .A(\REGISTERS[85][14] ), .B(n2754), .S(n1438), .Z(n9054) );
  MUX2_X1 U4718 ( .A(\REGISTERS[85][13] ), .B(n2743), .S(n1438), .Z(n9055) );
  MUX2_X1 U4719 ( .A(\REGISTERS[85][12] ), .B(n2732), .S(n1438), .Z(n9056) );
  MUX2_X1 U4720 ( .A(\REGISTERS[85][11] ), .B(n2721), .S(n1438), .Z(n9057) );
  MUX2_X1 U4721 ( .A(\REGISTERS[85][10] ), .B(n2710), .S(n1438), .Z(n9058) );
  MUX2_X1 U4722 ( .A(\REGISTERS[85][9] ), .B(n2603), .S(n1438), .Z(n9059) );
  MUX2_X1 U4723 ( .A(\REGISTERS[85][8] ), .B(n2592), .S(n1438), .Z(n9060) );
  MUX2_X1 U4724 ( .A(\REGISTERS[85][7] ), .B(n2581), .S(n1439), .Z(n9061) );
  MUX2_X1 U4725 ( .A(\REGISTERS[85][6] ), .B(n2570), .S(n1439), .Z(n9062) );
  MUX2_X1 U4726 ( .A(\REGISTERS[85][5] ), .B(n2559), .S(n1439), .Z(n9063) );
  MUX2_X1 U4727 ( .A(\REGISTERS[85][4] ), .B(n2548), .S(n1439), .Z(n9064) );
  MUX2_X1 U4728 ( .A(\REGISTERS[85][3] ), .B(n1833), .S(n1439), .Z(n9065) );
  MUX2_X1 U4729 ( .A(\REGISTERS[85][2] ), .B(n1822), .S(n1439), .Z(n9066) );
  MUX2_X1 U4730 ( .A(\REGISTERS[85][1] ), .B(n1811), .S(n1439), .Z(n9067) );
  MUX2_X1 U4731 ( .A(\REGISTERS[85][0] ), .B(n1800), .S(n1439), .Z(n9068) );
  MUX2_X1 U4732 ( .A(\REGISTERS[84][31] ), .B(n2947), .S(n1440), .Z(n9005) );
  MUX2_X1 U4733 ( .A(\REGISTERS[84][30] ), .B(n2936), .S(n1440), .Z(n9006) );
  MUX2_X1 U4734 ( .A(\REGISTERS[84][29] ), .B(n2925), .S(n1440), .Z(n9007) );
  MUX2_X1 U4735 ( .A(\REGISTERS[84][28] ), .B(n2909), .S(n1440), .Z(n9008) );
  MUX2_X1 U4736 ( .A(\REGISTERS[84][27] ), .B(n2897), .S(n1440), .Z(n9009) );
  MUX2_X1 U4737 ( .A(\REGISTERS[84][26] ), .B(n2886), .S(n1440), .Z(n9010) );
  MUX2_X1 U4738 ( .A(\REGISTERS[84][25] ), .B(n2875), .S(n1440), .Z(n9011) );
  MUX2_X1 U4739 ( .A(\REGISTERS[84][24] ), .B(n2864), .S(n1440), .Z(n9012) );
  MUX2_X1 U4740 ( .A(\REGISTERS[84][23] ), .B(n2853), .S(n1440), .Z(n9013) );
  MUX2_X1 U4741 ( .A(\REGISTERS[84][22] ), .B(n2842), .S(n1440), .Z(n9014) );
  MUX2_X1 U4742 ( .A(\REGISTERS[84][21] ), .B(n2831), .S(n1440), .Z(n9015) );
  MUX2_X1 U4743 ( .A(\REGISTERS[84][20] ), .B(n2820), .S(n1440), .Z(n9016) );
  MUX2_X1 U4744 ( .A(\REGISTERS[84][19] ), .B(n2809), .S(n1441), .Z(n9017) );
  MUX2_X1 U4745 ( .A(\REGISTERS[84][18] ), .B(n2798), .S(n1441), .Z(n9018) );
  MUX2_X1 U4746 ( .A(\REGISTERS[84][17] ), .B(n2787), .S(n1441), .Z(n9019) );
  MUX2_X1 U4747 ( .A(\REGISTERS[84][16] ), .B(n2776), .S(n1441), .Z(n9020) );
  MUX2_X1 U4748 ( .A(\REGISTERS[84][15] ), .B(n2765), .S(n1441), .Z(n9021) );
  MUX2_X1 U4749 ( .A(\REGISTERS[84][14] ), .B(n2754), .S(n1441), .Z(n9022) );
  MUX2_X1 U4750 ( .A(\REGISTERS[84][13] ), .B(n2743), .S(n1441), .Z(n9023) );
  MUX2_X1 U4751 ( .A(\REGISTERS[84][12] ), .B(n2732), .S(n1441), .Z(n9024) );
  MUX2_X1 U4752 ( .A(\REGISTERS[84][11] ), .B(n2721), .S(n1441), .Z(n9025) );
  MUX2_X1 U4753 ( .A(\REGISTERS[84][10] ), .B(n2710), .S(n1441), .Z(n9026) );
  MUX2_X1 U4754 ( .A(\REGISTERS[84][9] ), .B(n2603), .S(n1441), .Z(n9027) );
  MUX2_X1 U4755 ( .A(\REGISTERS[84][8] ), .B(n2592), .S(n1441), .Z(n9028) );
  MUX2_X1 U4756 ( .A(\REGISTERS[84][7] ), .B(n2581), .S(n1442), .Z(n9029) );
  MUX2_X1 U4757 ( .A(\REGISTERS[84][6] ), .B(n2570), .S(n1442), .Z(n9030) );
  MUX2_X1 U4758 ( .A(\REGISTERS[84][5] ), .B(n2559), .S(n1442), .Z(n9031) );
  MUX2_X1 U4759 ( .A(\REGISTERS[84][4] ), .B(n2548), .S(n1442), .Z(n9032) );
  MUX2_X1 U4760 ( .A(\REGISTERS[84][3] ), .B(n1833), .S(n1442), .Z(n9033) );
  MUX2_X1 U4761 ( .A(\REGISTERS[84][2] ), .B(n1822), .S(n1442), .Z(n9034) );
  MUX2_X1 U4762 ( .A(\REGISTERS[84][1] ), .B(n1811), .S(n1442), .Z(n9035) );
  MUX2_X1 U4763 ( .A(\REGISTERS[84][0] ), .B(n1800), .S(n1442), .Z(n9036) );
  MUX2_X1 U4764 ( .A(\REGISTERS[83][31] ), .B(n2947), .S(n1443), .Z(n8973) );
  MUX2_X1 U4765 ( .A(\REGISTERS[83][30] ), .B(n2936), .S(n1443), .Z(n8974) );
  MUX2_X1 U4766 ( .A(\REGISTERS[83][29] ), .B(n2925), .S(n1443), .Z(n8975) );
  MUX2_X1 U4767 ( .A(\REGISTERS[83][28] ), .B(n2909), .S(n1443), .Z(n8976) );
  MUX2_X1 U4768 ( .A(\REGISTERS[83][27] ), .B(n2897), .S(n1443), .Z(n8977) );
  MUX2_X1 U4769 ( .A(\REGISTERS[83][26] ), .B(n2886), .S(n1443), .Z(n8978) );
  MUX2_X1 U4770 ( .A(\REGISTERS[83][25] ), .B(n2875), .S(n1443), .Z(n8979) );
  MUX2_X1 U4771 ( .A(\REGISTERS[83][24] ), .B(n2864), .S(n1443), .Z(n8980) );
  MUX2_X1 U4772 ( .A(\REGISTERS[83][23] ), .B(n2853), .S(n1443), .Z(n8981) );
  MUX2_X1 U4773 ( .A(\REGISTERS[83][22] ), .B(n2842), .S(n1443), .Z(n8982) );
  MUX2_X1 U4774 ( .A(\REGISTERS[83][21] ), .B(n2831), .S(n1443), .Z(n8983) );
  MUX2_X1 U4775 ( .A(\REGISTERS[83][20] ), .B(n2820), .S(n1443), .Z(n8984) );
  MUX2_X1 U4776 ( .A(\REGISTERS[83][19] ), .B(n2809), .S(n1444), .Z(n8985) );
  MUX2_X1 U4777 ( .A(\REGISTERS[83][18] ), .B(n2798), .S(n1444), .Z(n8986) );
  MUX2_X1 U4778 ( .A(\REGISTERS[83][17] ), .B(n2787), .S(n1444), .Z(n8987) );
  MUX2_X1 U4779 ( .A(\REGISTERS[83][16] ), .B(n2776), .S(n1444), .Z(n8988) );
  MUX2_X1 U4780 ( .A(\REGISTERS[83][15] ), .B(n2765), .S(n1444), .Z(n8989) );
  MUX2_X1 U4781 ( .A(\REGISTERS[83][14] ), .B(n2754), .S(n1444), .Z(n8990) );
  MUX2_X1 U4782 ( .A(\REGISTERS[83][13] ), .B(n2743), .S(n1444), .Z(n8991) );
  MUX2_X1 U4783 ( .A(\REGISTERS[83][12] ), .B(n2732), .S(n1444), .Z(n8992) );
  MUX2_X1 U4784 ( .A(\REGISTERS[83][11] ), .B(n2721), .S(n1444), .Z(n8993) );
  MUX2_X1 U4785 ( .A(\REGISTERS[83][10] ), .B(n2710), .S(n1444), .Z(n8994) );
  MUX2_X1 U4786 ( .A(\REGISTERS[83][9] ), .B(n2603), .S(n1444), .Z(n8995) );
  MUX2_X1 U4787 ( .A(\REGISTERS[83][8] ), .B(n2592), .S(n1444), .Z(n8996) );
  MUX2_X1 U4788 ( .A(\REGISTERS[83][7] ), .B(n2581), .S(n1445), .Z(n8997) );
  MUX2_X1 U4789 ( .A(\REGISTERS[83][6] ), .B(n2570), .S(n1445), .Z(n8998) );
  MUX2_X1 U4790 ( .A(\REGISTERS[83][5] ), .B(n2559), .S(n1445), .Z(n8999) );
  MUX2_X1 U4791 ( .A(\REGISTERS[83][4] ), .B(n2548), .S(n1445), .Z(n9000) );
  MUX2_X1 U4792 ( .A(\REGISTERS[83][3] ), .B(n1833), .S(n1445), .Z(n9001) );
  MUX2_X1 U4793 ( .A(\REGISTERS[83][2] ), .B(n1822), .S(n1445), .Z(n9002) );
  MUX2_X1 U4794 ( .A(\REGISTERS[83][1] ), .B(n1811), .S(n1445), .Z(n9003) );
  MUX2_X1 U4795 ( .A(\REGISTERS[83][0] ), .B(n1800), .S(n1445), .Z(n9004) );
  MUX2_X1 U4796 ( .A(\REGISTERS[82][31] ), .B(n2947), .S(n1446), .Z(n8941) );
  MUX2_X1 U4797 ( .A(\REGISTERS[82][30] ), .B(n2936), .S(n1446), .Z(n8942) );
  MUX2_X1 U4798 ( .A(\REGISTERS[82][29] ), .B(n2925), .S(n1446), .Z(n8943) );
  MUX2_X1 U4799 ( .A(\REGISTERS[82][28] ), .B(n2909), .S(n1446), .Z(n8944) );
  MUX2_X1 U4800 ( .A(\REGISTERS[82][27] ), .B(n2897), .S(n1446), .Z(n8945) );
  MUX2_X1 U4801 ( .A(\REGISTERS[82][26] ), .B(n2886), .S(n1446), .Z(n8946) );
  MUX2_X1 U4802 ( .A(\REGISTERS[82][25] ), .B(n2875), .S(n1446), .Z(n8947) );
  MUX2_X1 U4803 ( .A(\REGISTERS[82][24] ), .B(n2864), .S(n1446), .Z(n8948) );
  MUX2_X1 U4804 ( .A(\REGISTERS[82][23] ), .B(n2853), .S(n1446), .Z(n8949) );
  MUX2_X1 U4805 ( .A(\REGISTERS[82][22] ), .B(n2842), .S(n1446), .Z(n8950) );
  MUX2_X1 U4806 ( .A(\REGISTERS[82][21] ), .B(n2831), .S(n1446), .Z(n8951) );
  MUX2_X1 U4807 ( .A(\REGISTERS[82][20] ), .B(n2820), .S(n1446), .Z(n8952) );
  MUX2_X1 U4808 ( .A(\REGISTERS[82][19] ), .B(n2809), .S(n1447), .Z(n8953) );
  MUX2_X1 U4809 ( .A(\REGISTERS[82][18] ), .B(n2798), .S(n1447), .Z(n8954) );
  MUX2_X1 U4810 ( .A(\REGISTERS[82][17] ), .B(n2787), .S(n1447), .Z(n8955) );
  MUX2_X1 U4811 ( .A(\REGISTERS[82][16] ), .B(n2776), .S(n1447), .Z(n8956) );
  MUX2_X1 U4812 ( .A(\REGISTERS[82][15] ), .B(n2765), .S(n1447), .Z(n8957) );
  MUX2_X1 U4813 ( .A(\REGISTERS[82][14] ), .B(n2754), .S(n1447), .Z(n8958) );
  MUX2_X1 U4814 ( .A(\REGISTERS[82][13] ), .B(n2743), .S(n1447), .Z(n8959) );
  MUX2_X1 U4815 ( .A(\REGISTERS[82][12] ), .B(n2732), .S(n1447), .Z(n8960) );
  MUX2_X1 U4816 ( .A(\REGISTERS[82][11] ), .B(n2721), .S(n1447), .Z(n8961) );
  MUX2_X1 U4817 ( .A(\REGISTERS[82][10] ), .B(n2710), .S(n1447), .Z(n8962) );
  MUX2_X1 U4818 ( .A(\REGISTERS[82][9] ), .B(n2603), .S(n1447), .Z(n8963) );
  MUX2_X1 U4819 ( .A(\REGISTERS[82][8] ), .B(n2592), .S(n1447), .Z(n8964) );
  MUX2_X1 U4820 ( .A(\REGISTERS[82][7] ), .B(n2581), .S(n1448), .Z(n8965) );
  MUX2_X1 U4821 ( .A(\REGISTERS[82][6] ), .B(n2570), .S(n1448), .Z(n8966) );
  MUX2_X1 U4822 ( .A(\REGISTERS[82][5] ), .B(n2559), .S(n1448), .Z(n8967) );
  MUX2_X1 U4823 ( .A(\REGISTERS[82][4] ), .B(n2548), .S(n1448), .Z(n8968) );
  MUX2_X1 U4824 ( .A(\REGISTERS[82][3] ), .B(n1833), .S(n1448), .Z(n8969) );
  MUX2_X1 U4825 ( .A(\REGISTERS[82][2] ), .B(n1822), .S(n1448), .Z(n8970) );
  MUX2_X1 U4826 ( .A(\REGISTERS[82][1] ), .B(n1811), .S(n1448), .Z(n8971) );
  MUX2_X1 U4827 ( .A(\REGISTERS[82][0] ), .B(n1800), .S(n1448), .Z(n8972) );
  MUX2_X1 U4828 ( .A(n10886), .B(n2947), .S(n1449), .Z(n8909) );
  MUX2_X1 U4829 ( .A(n10887), .B(n2936), .S(n1449), .Z(n8910) );
  MUX2_X1 U4830 ( .A(n10888), .B(n2925), .S(n1449), .Z(n8911) );
  MUX2_X1 U4831 ( .A(n10889), .B(n2909), .S(n1449), .Z(n8912) );
  MUX2_X1 U4832 ( .A(n10890), .B(n2897), .S(n1449), .Z(n8913) );
  MUX2_X1 U4833 ( .A(n10891), .B(n2886), .S(n1449), .Z(n8914) );
  MUX2_X1 U4834 ( .A(n10892), .B(n2875), .S(n1449), .Z(n8915) );
  MUX2_X1 U4835 ( .A(n10893), .B(n2864), .S(n1449), .Z(n8916) );
  MUX2_X1 U4836 ( .A(n10894), .B(n2853), .S(n1449), .Z(n8917) );
  MUX2_X1 U4837 ( .A(n10895), .B(n2842), .S(n1449), .Z(n8918) );
  MUX2_X1 U4838 ( .A(n10896), .B(n2831), .S(n1449), .Z(n8919) );
  MUX2_X1 U4839 ( .A(n10897), .B(n2820), .S(n1449), .Z(n8920) );
  MUX2_X1 U4840 ( .A(n10898), .B(n2809), .S(n1450), .Z(n8921) );
  MUX2_X1 U4841 ( .A(n10899), .B(n2798), .S(n1450), .Z(n8922) );
  MUX2_X1 U4842 ( .A(n10900), .B(n2787), .S(n1450), .Z(n8923) );
  MUX2_X1 U4843 ( .A(n10901), .B(n2776), .S(n1450), .Z(n8924) );
  MUX2_X1 U4844 ( .A(n10902), .B(n2765), .S(n1450), .Z(n8925) );
  MUX2_X1 U4845 ( .A(n10903), .B(n2754), .S(n1450), .Z(n8926) );
  MUX2_X1 U4846 ( .A(n10904), .B(n2743), .S(n1450), .Z(n8927) );
  MUX2_X1 U4847 ( .A(n10905), .B(n2732), .S(n1450), .Z(n8928) );
  MUX2_X1 U4848 ( .A(n10906), .B(n2721), .S(n1450), .Z(n8929) );
  MUX2_X1 U4849 ( .A(n10907), .B(n2710), .S(n1450), .Z(n8930) );
  MUX2_X1 U4850 ( .A(n10908), .B(n2603), .S(n1450), .Z(n8931) );
  MUX2_X1 U4851 ( .A(n10909), .B(n2592), .S(n1450), .Z(n8932) );
  MUX2_X1 U4852 ( .A(n10910), .B(n2581), .S(n1451), .Z(n8933) );
  MUX2_X1 U4853 ( .A(n10911), .B(n2570), .S(n1451), .Z(n8934) );
  MUX2_X1 U4854 ( .A(n10912), .B(n2559), .S(n1451), .Z(n8935) );
  MUX2_X1 U4855 ( .A(n10913), .B(n2548), .S(n1451), .Z(n8936) );
  MUX2_X1 U4856 ( .A(n10914), .B(n1833), .S(n1451), .Z(n8937) );
  MUX2_X1 U4857 ( .A(n10915), .B(n1822), .S(n1451), .Z(n8938) );
  MUX2_X1 U4858 ( .A(n10916), .B(n1811), .S(n1451), .Z(n8939) );
  MUX2_X1 U4859 ( .A(n10917), .B(n1800), .S(n1451), .Z(n8940) );
  MUX2_X1 U4860 ( .A(n10854), .B(n2947), .S(n1452), .Z(n8877) );
  MUX2_X1 U4861 ( .A(n10855), .B(n2936), .S(n1452), .Z(n8878) );
  MUX2_X1 U4862 ( .A(n10856), .B(n2925), .S(n1452), .Z(n8879) );
  MUX2_X1 U4863 ( .A(n10857), .B(n2909), .S(n1452), .Z(n8880) );
  MUX2_X1 U4864 ( .A(n10858), .B(n2897), .S(n1452), .Z(n8881) );
  MUX2_X1 U4865 ( .A(n10859), .B(n2886), .S(n1452), .Z(n8882) );
  MUX2_X1 U4866 ( .A(n10860), .B(n2875), .S(n1452), .Z(n8883) );
  MUX2_X1 U4867 ( .A(n10861), .B(n2864), .S(n1452), .Z(n8884) );
  MUX2_X1 U4868 ( .A(n10862), .B(n2853), .S(n1452), .Z(n8885) );
  MUX2_X1 U4869 ( .A(n10863), .B(n2842), .S(n1452), .Z(n8886) );
  MUX2_X1 U4870 ( .A(n10864), .B(n2831), .S(n1452), .Z(n8887) );
  MUX2_X1 U4871 ( .A(n10865), .B(n2820), .S(n1452), .Z(n8888) );
  MUX2_X1 U4872 ( .A(n10866), .B(n2809), .S(n1453), .Z(n8889) );
  MUX2_X1 U4873 ( .A(n10867), .B(n2798), .S(n1453), .Z(n8890) );
  MUX2_X1 U4874 ( .A(n10868), .B(n2787), .S(n1453), .Z(n8891) );
  MUX2_X1 U4875 ( .A(n10869), .B(n2776), .S(n1453), .Z(n8892) );
  MUX2_X1 U4876 ( .A(n10870), .B(n2765), .S(n1453), .Z(n8893) );
  MUX2_X1 U4877 ( .A(n10871), .B(n2754), .S(n1453), .Z(n8894) );
  MUX2_X1 U4878 ( .A(n10872), .B(n2743), .S(n1453), .Z(n8895) );
  MUX2_X1 U4879 ( .A(n10873), .B(n2732), .S(n1453), .Z(n8896) );
  MUX2_X1 U4880 ( .A(n10874), .B(n2721), .S(n1453), .Z(n8897) );
  MUX2_X1 U4881 ( .A(n10875), .B(n2710), .S(n1453), .Z(n8898) );
  MUX2_X1 U4882 ( .A(n10876), .B(n2603), .S(n1453), .Z(n8899) );
  MUX2_X1 U4883 ( .A(n10877), .B(n2592), .S(n1453), .Z(n8900) );
  MUX2_X1 U4884 ( .A(n10878), .B(n2581), .S(n1454), .Z(n8901) );
  MUX2_X1 U4885 ( .A(n10879), .B(n2570), .S(n1454), .Z(n8902) );
  MUX2_X1 U4886 ( .A(n10880), .B(n2559), .S(n1454), .Z(n8903) );
  MUX2_X1 U4887 ( .A(n10881), .B(n2548), .S(n1454), .Z(n8904) );
  MUX2_X1 U4888 ( .A(n10882), .B(n1833), .S(n1454), .Z(n8905) );
  MUX2_X1 U4889 ( .A(n10883), .B(n1822), .S(n1454), .Z(n8906) );
  MUX2_X1 U4890 ( .A(n10884), .B(n1811), .S(n1454), .Z(n8907) );
  MUX2_X1 U4891 ( .A(n10885), .B(n1800), .S(n1454), .Z(n8908) );
  MUX2_X1 U4892 ( .A(n10822), .B(n2947), .S(n1455), .Z(n8845) );
  MUX2_X1 U4893 ( .A(n10823), .B(n2936), .S(n1455), .Z(n8846) );
  MUX2_X1 U4894 ( .A(n10824), .B(n2925), .S(n1455), .Z(n8847) );
  MUX2_X1 U4895 ( .A(n10825), .B(n2909), .S(n1455), .Z(n8848) );
  MUX2_X1 U4896 ( .A(n10826), .B(n2897), .S(n1455), .Z(n8849) );
  MUX2_X1 U4897 ( .A(n10827), .B(n2886), .S(n1455), .Z(n8850) );
  MUX2_X1 U4898 ( .A(n10828), .B(n2875), .S(n1455), .Z(n8851) );
  MUX2_X1 U4899 ( .A(n10829), .B(n2864), .S(n1455), .Z(n8852) );
  MUX2_X1 U4900 ( .A(n10830), .B(n2853), .S(n1455), .Z(n8853) );
  MUX2_X1 U4901 ( .A(n10831), .B(n2842), .S(n1455), .Z(n8854) );
  MUX2_X1 U4902 ( .A(n10832), .B(n2831), .S(n1455), .Z(n8855) );
  MUX2_X1 U4903 ( .A(n10833), .B(n2820), .S(n1455), .Z(n8856) );
  MUX2_X1 U4904 ( .A(n10834), .B(n2809), .S(n1456), .Z(n8857) );
  MUX2_X1 U4905 ( .A(n10835), .B(n2798), .S(n1456), .Z(n8858) );
  MUX2_X1 U4906 ( .A(n10836), .B(n2787), .S(n1456), .Z(n8859) );
  MUX2_X1 U4907 ( .A(n10837), .B(n2776), .S(n1456), .Z(n8860) );
  MUX2_X1 U4908 ( .A(n10838), .B(n2765), .S(n1456), .Z(n8861) );
  MUX2_X1 U4909 ( .A(n10839), .B(n2754), .S(n1456), .Z(n8862) );
  MUX2_X1 U4910 ( .A(n10840), .B(n2743), .S(n1456), .Z(n8863) );
  MUX2_X1 U4911 ( .A(n10841), .B(n2732), .S(n1456), .Z(n8864) );
  MUX2_X1 U4912 ( .A(n10842), .B(n2721), .S(n1456), .Z(n8865) );
  MUX2_X1 U4913 ( .A(n10843), .B(n2710), .S(n1456), .Z(n8866) );
  MUX2_X1 U4914 ( .A(n10844), .B(n2603), .S(n1456), .Z(n8867) );
  MUX2_X1 U4915 ( .A(n10845), .B(n2592), .S(n1456), .Z(n8868) );
  MUX2_X1 U4916 ( .A(n10846), .B(n2581), .S(n1457), .Z(n8869) );
  MUX2_X1 U4917 ( .A(n10847), .B(n2570), .S(n1457), .Z(n8870) );
  MUX2_X1 U4918 ( .A(n10848), .B(n2559), .S(n1457), .Z(n8871) );
  MUX2_X1 U4919 ( .A(n10849), .B(n2548), .S(n1457), .Z(n8872) );
  MUX2_X1 U4920 ( .A(n10850), .B(n1833), .S(n1457), .Z(n8873) );
  MUX2_X1 U4921 ( .A(n10851), .B(n1822), .S(n1457), .Z(n8874) );
  MUX2_X1 U4922 ( .A(n10852), .B(n1811), .S(n1457), .Z(n8875) );
  MUX2_X1 U4923 ( .A(n10853), .B(n1800), .S(n1457), .Z(n8876) );
  MUX2_X1 U4924 ( .A(\REGISTERS[78][31] ), .B(n2947), .S(n1458), .Z(n8813) );
  MUX2_X1 U4925 ( .A(\REGISTERS[78][30] ), .B(n2936), .S(n1458), .Z(n8814) );
  MUX2_X1 U4926 ( .A(\REGISTERS[78][29] ), .B(n2925), .S(n1458), .Z(n8815) );
  MUX2_X1 U4927 ( .A(\REGISTERS[78][28] ), .B(n2909), .S(n1458), .Z(n8816) );
  MUX2_X1 U4928 ( .A(\REGISTERS[78][27] ), .B(n2897), .S(n1458), .Z(n8817) );
  MUX2_X1 U4929 ( .A(\REGISTERS[78][26] ), .B(n2886), .S(n1458), .Z(n8818) );
  MUX2_X1 U4930 ( .A(\REGISTERS[78][25] ), .B(n2875), .S(n1458), .Z(n8819) );
  MUX2_X1 U4931 ( .A(\REGISTERS[78][24] ), .B(n2864), .S(n1458), .Z(n8820) );
  MUX2_X1 U4932 ( .A(\REGISTERS[78][23] ), .B(n2853), .S(n1458), .Z(n8821) );
  MUX2_X1 U4933 ( .A(\REGISTERS[78][22] ), .B(n2842), .S(n1458), .Z(n8822) );
  MUX2_X1 U4934 ( .A(\REGISTERS[78][21] ), .B(n2831), .S(n1458), .Z(n8823) );
  MUX2_X1 U4935 ( .A(\REGISTERS[78][20] ), .B(n2820), .S(n1458), .Z(n8824) );
  MUX2_X1 U4936 ( .A(\REGISTERS[78][19] ), .B(n2809), .S(n1459), .Z(n8825) );
  MUX2_X1 U4937 ( .A(\REGISTERS[78][18] ), .B(n2798), .S(n1459), .Z(n8826) );
  MUX2_X1 U4938 ( .A(\REGISTERS[78][17] ), .B(n2787), .S(n1459), .Z(n8827) );
  MUX2_X1 U4939 ( .A(\REGISTERS[78][16] ), .B(n2776), .S(n1459), .Z(n8828) );
  MUX2_X1 U4940 ( .A(\REGISTERS[78][15] ), .B(n2765), .S(n1459), .Z(n8829) );
  MUX2_X1 U4941 ( .A(\REGISTERS[78][14] ), .B(n2754), .S(n1459), .Z(n8830) );
  MUX2_X1 U4942 ( .A(\REGISTERS[78][13] ), .B(n2743), .S(n1459), .Z(n8831) );
  MUX2_X1 U4943 ( .A(\REGISTERS[78][12] ), .B(n2732), .S(n1459), .Z(n8832) );
  MUX2_X1 U4944 ( .A(\REGISTERS[78][11] ), .B(n2721), .S(n1459), .Z(n8833) );
  MUX2_X1 U4945 ( .A(\REGISTERS[78][10] ), .B(n2710), .S(n1459), .Z(n8834) );
  MUX2_X1 U4946 ( .A(\REGISTERS[78][9] ), .B(n2603), .S(n1459), .Z(n8835) );
  MUX2_X1 U4947 ( .A(\REGISTERS[78][8] ), .B(n2592), .S(n1459), .Z(n8836) );
  MUX2_X1 U4948 ( .A(\REGISTERS[78][7] ), .B(n2581), .S(n1460), .Z(n8837) );
  MUX2_X1 U4949 ( .A(\REGISTERS[78][6] ), .B(n2570), .S(n1460), .Z(n8838) );
  MUX2_X1 U4950 ( .A(\REGISTERS[78][5] ), .B(n2559), .S(n1460), .Z(n8839) );
  MUX2_X1 U4951 ( .A(\REGISTERS[78][4] ), .B(n2548), .S(n1460), .Z(n8840) );
  MUX2_X1 U4952 ( .A(\REGISTERS[78][3] ), .B(n1833), .S(n1460), .Z(n8841) );
  MUX2_X1 U4953 ( .A(\REGISTERS[78][2] ), .B(n1822), .S(n1460), .Z(n8842) );
  MUX2_X1 U4954 ( .A(\REGISTERS[78][1] ), .B(n1811), .S(n1460), .Z(n8843) );
  MUX2_X1 U4955 ( .A(\REGISTERS[78][0] ), .B(n1800), .S(n1460), .Z(n8844) );
  MUX2_X1 U4956 ( .A(\REGISTERS[77][31] ), .B(n2947), .S(n1461), .Z(n8781) );
  MUX2_X1 U4957 ( .A(\REGISTERS[77][30] ), .B(n2936), .S(n1461), .Z(n8782) );
  MUX2_X1 U4958 ( .A(\REGISTERS[77][29] ), .B(n2925), .S(n1461), .Z(n8783) );
  MUX2_X1 U4959 ( .A(\REGISTERS[77][28] ), .B(n2909), .S(n1461), .Z(n8784) );
  MUX2_X1 U4960 ( .A(\REGISTERS[77][27] ), .B(n2897), .S(n1461), .Z(n8785) );
  MUX2_X1 U4961 ( .A(\REGISTERS[77][26] ), .B(n2886), .S(n1461), .Z(n8786) );
  MUX2_X1 U4962 ( .A(\REGISTERS[77][25] ), .B(n2875), .S(n1461), .Z(n8787) );
  MUX2_X1 U4963 ( .A(\REGISTERS[77][24] ), .B(n2864), .S(n1461), .Z(n8788) );
  MUX2_X1 U4964 ( .A(\REGISTERS[77][23] ), .B(n2853), .S(n1461), .Z(n8789) );
  MUX2_X1 U4965 ( .A(\REGISTERS[77][22] ), .B(n2842), .S(n1461), .Z(n8790) );
  MUX2_X1 U4966 ( .A(\REGISTERS[77][21] ), .B(n2831), .S(n1461), .Z(n8791) );
  MUX2_X1 U4967 ( .A(\REGISTERS[77][20] ), .B(n2820), .S(n1461), .Z(n8792) );
  MUX2_X1 U4968 ( .A(\REGISTERS[77][19] ), .B(n2809), .S(n1462), .Z(n8793) );
  MUX2_X1 U4969 ( .A(\REGISTERS[77][18] ), .B(n2798), .S(n1462), .Z(n8794) );
  MUX2_X1 U4970 ( .A(\REGISTERS[77][17] ), .B(n2787), .S(n1462), .Z(n8795) );
  MUX2_X1 U4971 ( .A(\REGISTERS[77][16] ), .B(n2776), .S(n1462), .Z(n8796) );
  MUX2_X1 U4972 ( .A(\REGISTERS[77][15] ), .B(n2765), .S(n1462), .Z(n8797) );
  MUX2_X1 U4973 ( .A(\REGISTERS[77][14] ), .B(n2754), .S(n1462), .Z(n8798) );
  MUX2_X1 U4974 ( .A(\REGISTERS[77][13] ), .B(n2743), .S(n1462), .Z(n8799) );
  MUX2_X1 U4975 ( .A(\REGISTERS[77][12] ), .B(n2732), .S(n1462), .Z(n8800) );
  MUX2_X1 U4976 ( .A(\REGISTERS[77][11] ), .B(n2721), .S(n1462), .Z(n8801) );
  MUX2_X1 U4977 ( .A(\REGISTERS[77][10] ), .B(n2710), .S(n1462), .Z(n8802) );
  MUX2_X1 U4978 ( .A(\REGISTERS[77][9] ), .B(n2603), .S(n1462), .Z(n8803) );
  MUX2_X1 U4979 ( .A(\REGISTERS[77][8] ), .B(n2592), .S(n1462), .Z(n8804) );
  MUX2_X1 U4980 ( .A(\REGISTERS[77][7] ), .B(n2581), .S(n1463), .Z(n8805) );
  MUX2_X1 U4981 ( .A(\REGISTERS[77][6] ), .B(n2570), .S(n1463), .Z(n8806) );
  MUX2_X1 U4982 ( .A(\REGISTERS[77][5] ), .B(n2559), .S(n1463), .Z(n8807) );
  MUX2_X1 U4983 ( .A(\REGISTERS[77][4] ), .B(n2548), .S(n1463), .Z(n8808) );
  MUX2_X1 U4984 ( .A(\REGISTERS[77][3] ), .B(n1833), .S(n1463), .Z(n8809) );
  MUX2_X1 U4985 ( .A(\REGISTERS[77][2] ), .B(n1822), .S(n1463), .Z(n8810) );
  MUX2_X1 U4986 ( .A(\REGISTERS[77][1] ), .B(n1811), .S(n1463), .Z(n8811) );
  MUX2_X1 U4987 ( .A(\REGISTERS[77][0] ), .B(n1800), .S(n1463), .Z(n8812) );
  MUX2_X1 U4988 ( .A(n10790), .B(n2948), .S(n1464), .Z(n8749) );
  MUX2_X1 U4989 ( .A(n10791), .B(n2937), .S(n1464), .Z(n8750) );
  MUX2_X1 U4990 ( .A(n10792), .B(n2926), .S(n1464), .Z(n8751) );
  MUX2_X1 U4991 ( .A(n10793), .B(n2910), .S(n1464), .Z(n8752) );
  MUX2_X1 U4992 ( .A(n10794), .B(n2899), .S(n1464), .Z(n8753) );
  MUX2_X1 U4993 ( .A(n10795), .B(n2887), .S(n1464), .Z(n8754) );
  MUX2_X1 U4994 ( .A(n10796), .B(n2876), .S(n1464), .Z(n8755) );
  MUX2_X1 U4995 ( .A(n10797), .B(n2865), .S(n1464), .Z(n8756) );
  MUX2_X1 U4996 ( .A(n10798), .B(n2854), .S(n1464), .Z(n8757) );
  MUX2_X1 U4997 ( .A(n10799), .B(n2843), .S(n1464), .Z(n8758) );
  MUX2_X1 U4998 ( .A(n10800), .B(n2832), .S(n1464), .Z(n8759) );
  MUX2_X1 U4999 ( .A(n10801), .B(n2821), .S(n1464), .Z(n8760) );
  MUX2_X1 U5000 ( .A(n10802), .B(n2810), .S(n1465), .Z(n8761) );
  MUX2_X1 U5001 ( .A(n10803), .B(n2799), .S(n1465), .Z(n8762) );
  MUX2_X1 U5002 ( .A(n10804), .B(n2788), .S(n1465), .Z(n8763) );
  MUX2_X1 U5003 ( .A(n10805), .B(n2777), .S(n1465), .Z(n8764) );
  MUX2_X1 U5004 ( .A(n10806), .B(n2766), .S(n1465), .Z(n8765) );
  MUX2_X1 U5005 ( .A(n10807), .B(n2755), .S(n1465), .Z(n8766) );
  MUX2_X1 U5006 ( .A(n10808), .B(n2744), .S(n1465), .Z(n8767) );
  MUX2_X1 U5007 ( .A(n10809), .B(n2733), .S(n1465), .Z(n8768) );
  MUX2_X1 U5008 ( .A(n10810), .B(n2722), .S(n1465), .Z(n8769) );
  MUX2_X1 U5009 ( .A(n10811), .B(n2711), .S(n1465), .Z(n8770) );
  MUX2_X1 U5010 ( .A(n10812), .B(n2604), .S(n1465), .Z(n8771) );
  MUX2_X1 U5011 ( .A(n10813), .B(n2593), .S(n1465), .Z(n8772) );
  MUX2_X1 U5012 ( .A(n10814), .B(n2582), .S(n1466), .Z(n8773) );
  MUX2_X1 U5013 ( .A(n10815), .B(n2571), .S(n1466), .Z(n8774) );
  MUX2_X1 U5014 ( .A(n10816), .B(n2560), .S(n1466), .Z(n8775) );
  MUX2_X1 U5015 ( .A(n10817), .B(n2549), .S(n1466), .Z(n8776) );
  MUX2_X1 U5016 ( .A(n10818), .B(n1834), .S(n1466), .Z(n8777) );
  MUX2_X1 U5017 ( .A(n10819), .B(n1823), .S(n1466), .Z(n8778) );
  MUX2_X1 U5018 ( .A(n10820), .B(n1812), .S(n1466), .Z(n8779) );
  MUX2_X1 U5019 ( .A(n10821), .B(n1801), .S(n1466), .Z(n8780) );
  MUX2_X1 U5020 ( .A(n10758), .B(n2948), .S(n1467), .Z(n8717) );
  MUX2_X1 U5021 ( .A(n10759), .B(n2937), .S(n1467), .Z(n8718) );
  MUX2_X1 U5022 ( .A(n10760), .B(n2926), .S(n1467), .Z(n8719) );
  MUX2_X1 U5023 ( .A(n10761), .B(n2910), .S(n1467), .Z(n8720) );
  MUX2_X1 U5024 ( .A(n10762), .B(n2899), .S(n1467), .Z(n8721) );
  MUX2_X1 U5025 ( .A(n10763), .B(n2887), .S(n1467), .Z(n8722) );
  MUX2_X1 U5026 ( .A(n10764), .B(n2876), .S(n1467), .Z(n8723) );
  MUX2_X1 U5027 ( .A(n10765), .B(n2865), .S(n1467), .Z(n8724) );
  MUX2_X1 U5028 ( .A(n10766), .B(n2854), .S(n1467), .Z(n8725) );
  MUX2_X1 U5029 ( .A(n10767), .B(n2843), .S(n1467), .Z(n8726) );
  MUX2_X1 U5030 ( .A(n10768), .B(n2832), .S(n1467), .Z(n8727) );
  MUX2_X1 U5031 ( .A(n10769), .B(n2821), .S(n1467), .Z(n8728) );
  MUX2_X1 U5032 ( .A(n10770), .B(n2810), .S(n1468), .Z(n8729) );
  MUX2_X1 U5033 ( .A(n10771), .B(n2799), .S(n1468), .Z(n8730) );
  MUX2_X1 U5034 ( .A(n10772), .B(n2788), .S(n1468), .Z(n8731) );
  MUX2_X1 U5035 ( .A(n10773), .B(n2777), .S(n1468), .Z(n8732) );
  MUX2_X1 U5036 ( .A(n10774), .B(n2766), .S(n1468), .Z(n8733) );
  MUX2_X1 U5037 ( .A(n10775), .B(n2755), .S(n1468), .Z(n8734) );
  MUX2_X1 U5038 ( .A(n10776), .B(n2744), .S(n1468), .Z(n8735) );
  MUX2_X1 U5039 ( .A(n10777), .B(n2733), .S(n1468), .Z(n8736) );
  MUX2_X1 U5040 ( .A(n10778), .B(n2722), .S(n1468), .Z(n8737) );
  MUX2_X1 U5041 ( .A(n10779), .B(n2711), .S(n1468), .Z(n8738) );
  MUX2_X1 U5042 ( .A(n10780), .B(n2604), .S(n1468), .Z(n8739) );
  MUX2_X1 U5043 ( .A(n10781), .B(n2593), .S(n1468), .Z(n8740) );
  MUX2_X1 U5044 ( .A(n10782), .B(n2582), .S(n1469), .Z(n8741) );
  MUX2_X1 U5045 ( .A(n10783), .B(n2571), .S(n1469), .Z(n8742) );
  MUX2_X1 U5046 ( .A(n10784), .B(n2560), .S(n1469), .Z(n8743) );
  MUX2_X1 U5047 ( .A(n10785), .B(n2549), .S(n1469), .Z(n8744) );
  MUX2_X1 U5048 ( .A(n10786), .B(n1834), .S(n1469), .Z(n8745) );
  MUX2_X1 U5049 ( .A(n10787), .B(n1823), .S(n1469), .Z(n8746) );
  MUX2_X1 U5050 ( .A(n10788), .B(n1812), .S(n1469), .Z(n8747) );
  MUX2_X1 U5051 ( .A(n10789), .B(n1801), .S(n1469), .Z(n8748) );
  MUX2_X1 U5052 ( .A(n10726), .B(n2948), .S(n1470), .Z(n8685) );
  MUX2_X1 U5053 ( .A(n10727), .B(n2937), .S(n1470), .Z(n8686) );
  MUX2_X1 U5054 ( .A(n10728), .B(n2926), .S(n1470), .Z(n8687) );
  MUX2_X1 U5055 ( .A(n10729), .B(n2910), .S(n1470), .Z(n8688) );
  MUX2_X1 U5056 ( .A(n10730), .B(n2899), .S(n1470), .Z(n8689) );
  MUX2_X1 U5057 ( .A(n10731), .B(n2887), .S(n1470), .Z(n8690) );
  MUX2_X1 U5058 ( .A(n10732), .B(n2876), .S(n1470), .Z(n8691) );
  MUX2_X1 U5059 ( .A(n10733), .B(n2865), .S(n1470), .Z(n8692) );
  MUX2_X1 U5060 ( .A(n10734), .B(n2854), .S(n1470), .Z(n8693) );
  MUX2_X1 U5061 ( .A(n10735), .B(n2843), .S(n1470), .Z(n8694) );
  MUX2_X1 U5062 ( .A(n10736), .B(n2832), .S(n1470), .Z(n8695) );
  MUX2_X1 U5063 ( .A(n10737), .B(n2821), .S(n1470), .Z(n8696) );
  MUX2_X1 U5064 ( .A(n10738), .B(n2810), .S(n1471), .Z(n8697) );
  MUX2_X1 U5065 ( .A(n10739), .B(n2799), .S(n1471), .Z(n8698) );
  MUX2_X1 U5066 ( .A(n10740), .B(n2788), .S(n1471), .Z(n8699) );
  MUX2_X1 U5067 ( .A(n10741), .B(n2777), .S(n1471), .Z(n8700) );
  MUX2_X1 U5068 ( .A(n10742), .B(n2766), .S(n1471), .Z(n8701) );
  MUX2_X1 U5069 ( .A(n10743), .B(n2755), .S(n1471), .Z(n8702) );
  MUX2_X1 U5070 ( .A(n10744), .B(n2744), .S(n1471), .Z(n8703) );
  MUX2_X1 U5071 ( .A(n10745), .B(n2733), .S(n1471), .Z(n8704) );
  MUX2_X1 U5072 ( .A(n10746), .B(n2722), .S(n1471), .Z(n8705) );
  MUX2_X1 U5073 ( .A(n10747), .B(n2711), .S(n1471), .Z(n8706) );
  MUX2_X1 U5074 ( .A(n10748), .B(n2604), .S(n1471), .Z(n8707) );
  MUX2_X1 U5075 ( .A(n10749), .B(n2593), .S(n1471), .Z(n8708) );
  MUX2_X1 U5076 ( .A(n10750), .B(n2582), .S(n1472), .Z(n8709) );
  MUX2_X1 U5077 ( .A(n10751), .B(n2571), .S(n1472), .Z(n8710) );
  MUX2_X1 U5078 ( .A(n10752), .B(n2560), .S(n1472), .Z(n8711) );
  MUX2_X1 U5079 ( .A(n10753), .B(n2549), .S(n1472), .Z(n8712) );
  MUX2_X1 U5080 ( .A(n10754), .B(n1834), .S(n1472), .Z(n8713) );
  MUX2_X1 U5081 ( .A(n10755), .B(n1823), .S(n1472), .Z(n8714) );
  MUX2_X1 U5082 ( .A(n10756), .B(n1812), .S(n1472), .Z(n8715) );
  MUX2_X1 U5083 ( .A(n10757), .B(n1801), .S(n1472), .Z(n8716) );
  MUX2_X1 U5084 ( .A(n10694), .B(n2948), .S(n1473), .Z(n8653) );
  MUX2_X1 U5085 ( .A(n10695), .B(n2937), .S(n1473), .Z(n8654) );
  MUX2_X1 U5086 ( .A(n10696), .B(n2926), .S(n1473), .Z(n8655) );
  MUX2_X1 U5087 ( .A(n10697), .B(n2910), .S(n1473), .Z(n8656) );
  MUX2_X1 U5088 ( .A(n10698), .B(n2899), .S(n1473), .Z(n8657) );
  MUX2_X1 U5089 ( .A(n10699), .B(n2887), .S(n1473), .Z(n8658) );
  MUX2_X1 U5090 ( .A(n10700), .B(n2876), .S(n1473), .Z(n8659) );
  MUX2_X1 U5091 ( .A(n10701), .B(n2865), .S(n1473), .Z(n8660) );
  MUX2_X1 U5092 ( .A(n10702), .B(n2854), .S(n1473), .Z(n8661) );
  MUX2_X1 U5093 ( .A(n10703), .B(n2843), .S(n1473), .Z(n8662) );
  MUX2_X1 U5094 ( .A(n10704), .B(n2832), .S(n1473), .Z(n8663) );
  MUX2_X1 U5095 ( .A(n10705), .B(n2821), .S(n1473), .Z(n8664) );
  MUX2_X1 U5096 ( .A(n10706), .B(n2810), .S(n1474), .Z(n8665) );
  MUX2_X1 U5097 ( .A(n10707), .B(n2799), .S(n1474), .Z(n8666) );
  MUX2_X1 U5098 ( .A(n10708), .B(n2788), .S(n1474), .Z(n8667) );
  MUX2_X1 U5099 ( .A(n10709), .B(n2777), .S(n1474), .Z(n8668) );
  MUX2_X1 U5100 ( .A(n10710), .B(n2766), .S(n1474), .Z(n8669) );
  MUX2_X1 U5101 ( .A(n10711), .B(n2755), .S(n1474), .Z(n8670) );
  MUX2_X1 U5102 ( .A(n10712), .B(n2744), .S(n1474), .Z(n8671) );
  MUX2_X1 U5103 ( .A(n10713), .B(n2733), .S(n1474), .Z(n8672) );
  MUX2_X1 U5104 ( .A(n10714), .B(n2722), .S(n1474), .Z(n8673) );
  MUX2_X1 U5105 ( .A(n10715), .B(n2711), .S(n1474), .Z(n8674) );
  MUX2_X1 U5106 ( .A(n10716), .B(n2604), .S(n1474), .Z(n8675) );
  MUX2_X1 U5107 ( .A(n10717), .B(n2593), .S(n1474), .Z(n8676) );
  MUX2_X1 U5108 ( .A(n10718), .B(n2582), .S(n1475), .Z(n8677) );
  MUX2_X1 U5109 ( .A(n10719), .B(n2571), .S(n1475), .Z(n8678) );
  MUX2_X1 U5110 ( .A(n10720), .B(n2560), .S(n1475), .Z(n8679) );
  MUX2_X1 U5111 ( .A(n10721), .B(n2549), .S(n1475), .Z(n8680) );
  MUX2_X1 U5112 ( .A(n10722), .B(n1834), .S(n1475), .Z(n8681) );
  MUX2_X1 U5113 ( .A(n10723), .B(n1823), .S(n1475), .Z(n8682) );
  MUX2_X1 U5114 ( .A(n10724), .B(n1812), .S(n1475), .Z(n8683) );
  MUX2_X1 U5115 ( .A(n10725), .B(n1801), .S(n1475), .Z(n8684) );
  MUX2_X1 U5116 ( .A(n10662), .B(n2948), .S(n1476), .Z(n8621) );
  MUX2_X1 U5117 ( .A(n10663), .B(n2937), .S(n1476), .Z(n8622) );
  MUX2_X1 U5118 ( .A(n10664), .B(n2926), .S(n1476), .Z(n8623) );
  MUX2_X1 U5119 ( .A(n10665), .B(n2910), .S(n1476), .Z(n8624) );
  MUX2_X1 U5120 ( .A(n10666), .B(n2899), .S(n1476), .Z(n8625) );
  MUX2_X1 U5121 ( .A(n10667), .B(n2887), .S(n1476), .Z(n8626) );
  MUX2_X1 U5122 ( .A(n10668), .B(n2876), .S(n1476), .Z(n8627) );
  MUX2_X1 U5123 ( .A(n10669), .B(n2865), .S(n1476), .Z(n8628) );
  MUX2_X1 U5124 ( .A(n10670), .B(n2854), .S(n1476), .Z(n8629) );
  MUX2_X1 U5125 ( .A(n10671), .B(n2843), .S(n1476), .Z(n8630) );
  MUX2_X1 U5126 ( .A(n10672), .B(n2832), .S(n1476), .Z(n8631) );
  MUX2_X1 U5127 ( .A(n10673), .B(n2821), .S(n1476), .Z(n8632) );
  MUX2_X1 U5128 ( .A(n10674), .B(n2810), .S(n1477), .Z(n8633) );
  MUX2_X1 U5129 ( .A(n10675), .B(n2799), .S(n1477), .Z(n8634) );
  MUX2_X1 U5130 ( .A(n10676), .B(n2788), .S(n1477), .Z(n8635) );
  MUX2_X1 U5131 ( .A(n10677), .B(n2777), .S(n1477), .Z(n8636) );
  MUX2_X1 U5132 ( .A(n10678), .B(n2766), .S(n1477), .Z(n8637) );
  MUX2_X1 U5133 ( .A(n10679), .B(n2755), .S(n1477), .Z(n8638) );
  MUX2_X1 U5134 ( .A(n10680), .B(n2744), .S(n1477), .Z(n8639) );
  MUX2_X1 U5135 ( .A(n10681), .B(n2733), .S(n1477), .Z(n8640) );
  MUX2_X1 U5136 ( .A(n10682), .B(n2722), .S(n1477), .Z(n8641) );
  MUX2_X1 U5137 ( .A(n10683), .B(n2711), .S(n1477), .Z(n8642) );
  MUX2_X1 U5138 ( .A(n10684), .B(n2604), .S(n1477), .Z(n8643) );
  MUX2_X1 U5139 ( .A(n10685), .B(n2593), .S(n1477), .Z(n8644) );
  MUX2_X1 U5140 ( .A(n10686), .B(n2582), .S(n1478), .Z(n8645) );
  MUX2_X1 U5141 ( .A(n10687), .B(n2571), .S(n1478), .Z(n8646) );
  MUX2_X1 U5142 ( .A(n10688), .B(n2560), .S(n1478), .Z(n8647) );
  MUX2_X1 U5143 ( .A(n10689), .B(n2549), .S(n1478), .Z(n8648) );
  MUX2_X1 U5144 ( .A(n10690), .B(n1834), .S(n1478), .Z(n8649) );
  MUX2_X1 U5145 ( .A(n10691), .B(n1823), .S(n1478), .Z(n8650) );
  MUX2_X1 U5146 ( .A(n10692), .B(n1812), .S(n1478), .Z(n8651) );
  MUX2_X1 U5147 ( .A(n10693), .B(n1801), .S(n1478), .Z(n8652) );
  MUX2_X1 U5148 ( .A(n10630), .B(n2948), .S(n1479), .Z(n8589) );
  MUX2_X1 U5149 ( .A(n10631), .B(n2937), .S(n1479), .Z(n8590) );
  MUX2_X1 U5150 ( .A(n10632), .B(n2926), .S(n1479), .Z(n8591) );
  MUX2_X1 U5151 ( .A(n10633), .B(n2910), .S(n1479), .Z(n8592) );
  MUX2_X1 U5152 ( .A(n10634), .B(n2899), .S(n1479), .Z(n8593) );
  MUX2_X1 U5153 ( .A(n10635), .B(n2887), .S(n1479), .Z(n8594) );
  MUX2_X1 U5154 ( .A(n10636), .B(n2876), .S(n1479), .Z(n8595) );
  MUX2_X1 U5155 ( .A(n10637), .B(n2865), .S(n1479), .Z(n8596) );
  MUX2_X1 U5156 ( .A(n10638), .B(n2854), .S(n1479), .Z(n8597) );
  MUX2_X1 U5157 ( .A(n10639), .B(n2843), .S(n1479), .Z(n8598) );
  MUX2_X1 U5158 ( .A(n10640), .B(n2832), .S(n1479), .Z(n8599) );
  MUX2_X1 U5159 ( .A(n10641), .B(n2821), .S(n1479), .Z(n8600) );
  MUX2_X1 U5160 ( .A(n10642), .B(n2810), .S(n1480), .Z(n8601) );
  MUX2_X1 U5161 ( .A(n10643), .B(n2799), .S(n1480), .Z(n8602) );
  MUX2_X1 U5162 ( .A(n10644), .B(n2788), .S(n1480), .Z(n8603) );
  MUX2_X1 U5163 ( .A(n10645), .B(n2777), .S(n1480), .Z(n8604) );
  MUX2_X1 U5164 ( .A(n10646), .B(n2766), .S(n1480), .Z(n8605) );
  MUX2_X1 U5165 ( .A(n10647), .B(n2755), .S(n1480), .Z(n8606) );
  MUX2_X1 U5166 ( .A(n10648), .B(n2744), .S(n1480), .Z(n8607) );
  MUX2_X1 U5167 ( .A(n10649), .B(n2733), .S(n1480), .Z(n8608) );
  MUX2_X1 U5168 ( .A(n10650), .B(n2722), .S(n1480), .Z(n8609) );
  MUX2_X1 U5169 ( .A(n10651), .B(n2711), .S(n1480), .Z(n8610) );
  MUX2_X1 U5170 ( .A(n10652), .B(n2604), .S(n1480), .Z(n8611) );
  MUX2_X1 U5171 ( .A(n10653), .B(n2593), .S(n1480), .Z(n8612) );
  MUX2_X1 U5172 ( .A(n10654), .B(n2582), .S(n1481), .Z(n8613) );
  MUX2_X1 U5173 ( .A(n10655), .B(n2571), .S(n1481), .Z(n8614) );
  MUX2_X1 U5174 ( .A(n10656), .B(n2560), .S(n1481), .Z(n8615) );
  MUX2_X1 U5175 ( .A(n10657), .B(n2549), .S(n1481), .Z(n8616) );
  MUX2_X1 U5176 ( .A(n10658), .B(n1834), .S(n1481), .Z(n8617) );
  MUX2_X1 U5177 ( .A(n10659), .B(n1823), .S(n1481), .Z(n8618) );
  MUX2_X1 U5178 ( .A(n10660), .B(n1812), .S(n1481), .Z(n8619) );
  MUX2_X1 U5179 ( .A(n10661), .B(n1801), .S(n1481), .Z(n8620) );
  MUX2_X1 U5180 ( .A(n10598), .B(n2948), .S(n1482), .Z(n8557) );
  MUX2_X1 U5181 ( .A(n10599), .B(n2937), .S(n1482), .Z(n8558) );
  MUX2_X1 U5182 ( .A(n10600), .B(n2926), .S(n1482), .Z(n8559) );
  MUX2_X1 U5183 ( .A(n10601), .B(n2910), .S(n1482), .Z(n8560) );
  MUX2_X1 U5184 ( .A(n10602), .B(n2899), .S(n1482), .Z(n8561) );
  MUX2_X1 U5185 ( .A(n10603), .B(n2887), .S(n1482), .Z(n8562) );
  MUX2_X1 U5186 ( .A(n10604), .B(n2876), .S(n1482), .Z(n8563) );
  MUX2_X1 U5187 ( .A(n10605), .B(n2865), .S(n1482), .Z(n8564) );
  MUX2_X1 U5188 ( .A(n10606), .B(n2854), .S(n1482), .Z(n8565) );
  MUX2_X1 U5189 ( .A(n10607), .B(n2843), .S(n1482), .Z(n8566) );
  MUX2_X1 U5190 ( .A(n10608), .B(n2832), .S(n1482), .Z(n8567) );
  MUX2_X1 U5191 ( .A(n10609), .B(n2821), .S(n1482), .Z(n8568) );
  MUX2_X1 U5192 ( .A(n10610), .B(n2810), .S(n1483), .Z(n8569) );
  MUX2_X1 U5193 ( .A(n10611), .B(n2799), .S(n1483), .Z(n8570) );
  MUX2_X1 U5194 ( .A(n10612), .B(n2788), .S(n1483), .Z(n8571) );
  MUX2_X1 U5195 ( .A(n10613), .B(n2777), .S(n1483), .Z(n8572) );
  MUX2_X1 U5196 ( .A(n10614), .B(n2766), .S(n1483), .Z(n8573) );
  MUX2_X1 U5197 ( .A(n10615), .B(n2755), .S(n1483), .Z(n8574) );
  MUX2_X1 U5198 ( .A(n10616), .B(n2744), .S(n1483), .Z(n8575) );
  MUX2_X1 U5199 ( .A(n10617), .B(n2733), .S(n1483), .Z(n8576) );
  MUX2_X1 U5200 ( .A(n10618), .B(n2722), .S(n1483), .Z(n8577) );
  MUX2_X1 U5201 ( .A(n10619), .B(n2711), .S(n1483), .Z(n8578) );
  MUX2_X1 U5202 ( .A(n10620), .B(n2604), .S(n1483), .Z(n8579) );
  MUX2_X1 U5203 ( .A(n10621), .B(n2593), .S(n1483), .Z(n8580) );
  MUX2_X1 U5204 ( .A(n10622), .B(n2582), .S(n1484), .Z(n8581) );
  MUX2_X1 U5205 ( .A(n10623), .B(n2571), .S(n1484), .Z(n8582) );
  MUX2_X1 U5206 ( .A(n10624), .B(n2560), .S(n1484), .Z(n8583) );
  MUX2_X1 U5207 ( .A(n10625), .B(n2549), .S(n1484), .Z(n8584) );
  MUX2_X1 U5208 ( .A(n10626), .B(n1834), .S(n1484), .Z(n8585) );
  MUX2_X1 U5209 ( .A(n10627), .B(n1823), .S(n1484), .Z(n8586) );
  MUX2_X1 U5210 ( .A(n10628), .B(n1812), .S(n1484), .Z(n8587) );
  MUX2_X1 U5211 ( .A(n10629), .B(n1801), .S(n1484), .Z(n8588) );
  MUX2_X1 U5212 ( .A(n10566), .B(n2948), .S(n1485), .Z(n8525) );
  MUX2_X1 U5213 ( .A(n10567), .B(n2937), .S(n1485), .Z(n8526) );
  MUX2_X1 U5214 ( .A(n10568), .B(n2926), .S(n1485), .Z(n8527) );
  MUX2_X1 U5215 ( .A(n10569), .B(n2910), .S(n1485), .Z(n8528) );
  MUX2_X1 U5216 ( .A(n10570), .B(n2899), .S(n1485), .Z(n8529) );
  MUX2_X1 U5217 ( .A(n10571), .B(n2887), .S(n1485), .Z(n8530) );
  MUX2_X1 U5218 ( .A(n10572), .B(n2876), .S(n1485), .Z(n8531) );
  MUX2_X1 U5219 ( .A(n10573), .B(n2865), .S(n1485), .Z(n8532) );
  MUX2_X1 U5220 ( .A(n10574), .B(n2854), .S(n1485), .Z(n8533) );
  MUX2_X1 U5221 ( .A(n10575), .B(n2843), .S(n1485), .Z(n8534) );
  MUX2_X1 U5222 ( .A(n10576), .B(n2832), .S(n1485), .Z(n8535) );
  MUX2_X1 U5223 ( .A(n10577), .B(n2821), .S(n1485), .Z(n8536) );
  MUX2_X1 U5224 ( .A(n10578), .B(n2810), .S(n1486), .Z(n8537) );
  MUX2_X1 U5225 ( .A(n10579), .B(n2799), .S(n1486), .Z(n8538) );
  MUX2_X1 U5226 ( .A(n10580), .B(n2788), .S(n1486), .Z(n8539) );
  MUX2_X1 U5227 ( .A(n10581), .B(n2777), .S(n1486), .Z(n8540) );
  MUX2_X1 U5228 ( .A(n10582), .B(n2766), .S(n1486), .Z(n8541) );
  MUX2_X1 U5229 ( .A(n10583), .B(n2755), .S(n1486), .Z(n8542) );
  MUX2_X1 U5230 ( .A(n10584), .B(n2744), .S(n1486), .Z(n8543) );
  MUX2_X1 U5231 ( .A(n10585), .B(n2733), .S(n1486), .Z(n8544) );
  MUX2_X1 U5232 ( .A(n10586), .B(n2722), .S(n1486), .Z(n8545) );
  MUX2_X1 U5233 ( .A(n10587), .B(n2711), .S(n1486), .Z(n8546) );
  MUX2_X1 U5234 ( .A(n10588), .B(n2604), .S(n1486), .Z(n8547) );
  MUX2_X1 U5235 ( .A(n10589), .B(n2593), .S(n1486), .Z(n8548) );
  MUX2_X1 U5236 ( .A(n10590), .B(n2582), .S(n1487), .Z(n8549) );
  MUX2_X1 U5237 ( .A(n10591), .B(n2571), .S(n1487), .Z(n8550) );
  MUX2_X1 U5238 ( .A(n10592), .B(n2560), .S(n1487), .Z(n8551) );
  MUX2_X1 U5239 ( .A(n10593), .B(n2549), .S(n1487), .Z(n8552) );
  MUX2_X1 U5240 ( .A(n10594), .B(n1834), .S(n1487), .Z(n8553) );
  MUX2_X1 U5241 ( .A(n10595), .B(n1823), .S(n1487), .Z(n8554) );
  MUX2_X1 U5242 ( .A(n10596), .B(n1812), .S(n1487), .Z(n8555) );
  MUX2_X1 U5243 ( .A(n10597), .B(n1801), .S(n1487), .Z(n8556) );
  MUX2_X1 U5244 ( .A(n10534), .B(n2948), .S(n1488), .Z(n8493) );
  MUX2_X1 U5245 ( .A(n10535), .B(n2937), .S(n1488), .Z(n8494) );
  MUX2_X1 U5246 ( .A(n10536), .B(n2926), .S(n1488), .Z(n8495) );
  MUX2_X1 U5247 ( .A(n10537), .B(n2910), .S(n1488), .Z(n8496) );
  MUX2_X1 U5248 ( .A(n10538), .B(n2899), .S(n1488), .Z(n8497) );
  MUX2_X1 U5249 ( .A(n10539), .B(n2887), .S(n1488), .Z(n8498) );
  MUX2_X1 U5250 ( .A(n10540), .B(n2876), .S(n1488), .Z(n8499) );
  MUX2_X1 U5251 ( .A(n10541), .B(n2865), .S(n1488), .Z(n8500) );
  MUX2_X1 U5252 ( .A(n10542), .B(n2854), .S(n1488), .Z(n8501) );
  MUX2_X1 U5253 ( .A(n10543), .B(n2843), .S(n1488), .Z(n8502) );
  MUX2_X1 U5254 ( .A(n10544), .B(n2832), .S(n1488), .Z(n8503) );
  MUX2_X1 U5255 ( .A(n10545), .B(n2821), .S(n1488), .Z(n8504) );
  MUX2_X1 U5256 ( .A(n10546), .B(n2810), .S(n1489), .Z(n8505) );
  MUX2_X1 U5257 ( .A(n10547), .B(n2799), .S(n1489), .Z(n8506) );
  MUX2_X1 U5258 ( .A(n10548), .B(n2788), .S(n1489), .Z(n8507) );
  MUX2_X1 U5259 ( .A(n10549), .B(n2777), .S(n1489), .Z(n8508) );
  MUX2_X1 U5260 ( .A(n10550), .B(n2766), .S(n1489), .Z(n8509) );
  MUX2_X1 U5261 ( .A(n10551), .B(n2755), .S(n1489), .Z(n8510) );
  MUX2_X1 U5262 ( .A(n10552), .B(n2744), .S(n1489), .Z(n8511) );
  MUX2_X1 U5263 ( .A(n10553), .B(n2733), .S(n1489), .Z(n8512) );
  MUX2_X1 U5264 ( .A(n10554), .B(n2722), .S(n1489), .Z(n8513) );
  MUX2_X1 U5265 ( .A(n10555), .B(n2711), .S(n1489), .Z(n8514) );
  MUX2_X1 U5266 ( .A(n10556), .B(n2604), .S(n1489), .Z(n8515) );
  MUX2_X1 U5267 ( .A(n10557), .B(n2593), .S(n1489), .Z(n8516) );
  MUX2_X1 U5268 ( .A(n10558), .B(n2582), .S(n1490), .Z(n8517) );
  MUX2_X1 U5269 ( .A(n10559), .B(n2571), .S(n1490), .Z(n8518) );
  MUX2_X1 U5270 ( .A(n10560), .B(n2560), .S(n1490), .Z(n8519) );
  MUX2_X1 U5271 ( .A(n10561), .B(n2549), .S(n1490), .Z(n8520) );
  MUX2_X1 U5272 ( .A(n10562), .B(n1834), .S(n1490), .Z(n8521) );
  MUX2_X1 U5273 ( .A(n10563), .B(n1823), .S(n1490), .Z(n8522) );
  MUX2_X1 U5274 ( .A(n10564), .B(n1812), .S(n1490), .Z(n8523) );
  MUX2_X1 U5275 ( .A(n10565), .B(n1801), .S(n1490), .Z(n8524) );
  MUX2_X1 U5276 ( .A(n10502), .B(n2948), .S(n1491), .Z(n8461) );
  MUX2_X1 U5277 ( .A(n10503), .B(n2937), .S(n1491), .Z(n8462) );
  MUX2_X1 U5278 ( .A(n10504), .B(n2926), .S(n1491), .Z(n8463) );
  MUX2_X1 U5279 ( .A(n10505), .B(n2910), .S(n1491), .Z(n8464) );
  MUX2_X1 U5280 ( .A(n10506), .B(n2899), .S(n1491), .Z(n8465) );
  MUX2_X1 U5281 ( .A(n10507), .B(n2887), .S(n1491), .Z(n8466) );
  MUX2_X1 U5282 ( .A(n10508), .B(n2876), .S(n1491), .Z(n8467) );
  MUX2_X1 U5283 ( .A(n10509), .B(n2865), .S(n1491), .Z(n8468) );
  MUX2_X1 U5284 ( .A(n10510), .B(n2854), .S(n1491), .Z(n8469) );
  MUX2_X1 U5285 ( .A(n10511), .B(n2843), .S(n1491), .Z(n8470) );
  MUX2_X1 U5286 ( .A(n10512), .B(n2832), .S(n1491), .Z(n8471) );
  MUX2_X1 U5287 ( .A(n10513), .B(n2821), .S(n1491), .Z(n8472) );
  MUX2_X1 U5288 ( .A(n10514), .B(n2810), .S(n1492), .Z(n8473) );
  MUX2_X1 U5289 ( .A(n10515), .B(n2799), .S(n1492), .Z(n8474) );
  MUX2_X1 U5290 ( .A(n10516), .B(n2788), .S(n1492), .Z(n8475) );
  MUX2_X1 U5291 ( .A(n10517), .B(n2777), .S(n1492), .Z(n8476) );
  MUX2_X1 U5292 ( .A(n10518), .B(n2766), .S(n1492), .Z(n8477) );
  MUX2_X1 U5293 ( .A(n10519), .B(n2755), .S(n1492), .Z(n8478) );
  MUX2_X1 U5294 ( .A(n10520), .B(n2744), .S(n1492), .Z(n8479) );
  MUX2_X1 U5295 ( .A(n10521), .B(n2733), .S(n1492), .Z(n8480) );
  MUX2_X1 U5296 ( .A(n10522), .B(n2722), .S(n1492), .Z(n8481) );
  MUX2_X1 U5297 ( .A(n10523), .B(n2711), .S(n1492), .Z(n8482) );
  MUX2_X1 U5298 ( .A(n10524), .B(n2604), .S(n1492), .Z(n8483) );
  MUX2_X1 U5299 ( .A(n10525), .B(n2593), .S(n1492), .Z(n8484) );
  MUX2_X1 U5300 ( .A(n10526), .B(n2582), .S(n1493), .Z(n8485) );
  MUX2_X1 U5301 ( .A(n10527), .B(n2571), .S(n1493), .Z(n8486) );
  MUX2_X1 U5302 ( .A(n10528), .B(n2560), .S(n1493), .Z(n8487) );
  MUX2_X1 U5303 ( .A(n10529), .B(n2549), .S(n1493), .Z(n8488) );
  MUX2_X1 U5304 ( .A(n10530), .B(n1834), .S(n1493), .Z(n8489) );
  MUX2_X1 U5305 ( .A(n10531), .B(n1823), .S(n1493), .Z(n8490) );
  MUX2_X1 U5306 ( .A(n10532), .B(n1812), .S(n1493), .Z(n8491) );
  MUX2_X1 U5307 ( .A(n10533), .B(n1801), .S(n1493), .Z(n8492) );
  MUX2_X1 U5308 ( .A(n10470), .B(n2948), .S(n1494), .Z(n8429) );
  MUX2_X1 U5309 ( .A(n10471), .B(n2937), .S(n1494), .Z(n8430) );
  MUX2_X1 U5310 ( .A(n10472), .B(n2926), .S(n1494), .Z(n8431) );
  MUX2_X1 U5311 ( .A(n10473), .B(n2910), .S(n1494), .Z(n8432) );
  MUX2_X1 U5312 ( .A(n10474), .B(n2899), .S(n1494), .Z(n8433) );
  MUX2_X1 U5313 ( .A(n10475), .B(n2887), .S(n1494), .Z(n8434) );
  MUX2_X1 U5314 ( .A(n10476), .B(n2876), .S(n1494), .Z(n8435) );
  MUX2_X1 U5315 ( .A(n10477), .B(n2865), .S(n1494), .Z(n8436) );
  MUX2_X1 U5316 ( .A(n10478), .B(n2854), .S(n1494), .Z(n8437) );
  MUX2_X1 U5317 ( .A(n10479), .B(n2843), .S(n1494), .Z(n8438) );
  MUX2_X1 U5318 ( .A(n10480), .B(n2832), .S(n1494), .Z(n8439) );
  MUX2_X1 U5319 ( .A(n10481), .B(n2821), .S(n1494), .Z(n8440) );
  MUX2_X1 U5320 ( .A(n10482), .B(n2810), .S(n1495), .Z(n8441) );
  MUX2_X1 U5321 ( .A(n10483), .B(n2799), .S(n1495), .Z(n8442) );
  MUX2_X1 U5322 ( .A(n10484), .B(n2788), .S(n1495), .Z(n8443) );
  MUX2_X1 U5323 ( .A(n10485), .B(n2777), .S(n1495), .Z(n8444) );
  MUX2_X1 U5324 ( .A(n10486), .B(n2766), .S(n1495), .Z(n8445) );
  MUX2_X1 U5325 ( .A(n10487), .B(n2755), .S(n1495), .Z(n8446) );
  MUX2_X1 U5326 ( .A(n10488), .B(n2744), .S(n1495), .Z(n8447) );
  MUX2_X1 U5327 ( .A(n10489), .B(n2733), .S(n1495), .Z(n8448) );
  MUX2_X1 U5328 ( .A(n10490), .B(n2722), .S(n1495), .Z(n8449) );
  MUX2_X1 U5329 ( .A(n10491), .B(n2711), .S(n1495), .Z(n8450) );
  MUX2_X1 U5330 ( .A(n10492), .B(n2604), .S(n1495), .Z(n8451) );
  MUX2_X1 U5331 ( .A(n10493), .B(n2593), .S(n1495), .Z(n8452) );
  MUX2_X1 U5332 ( .A(n10494), .B(n2582), .S(n1496), .Z(n8453) );
  MUX2_X1 U5333 ( .A(n10495), .B(n2571), .S(n1496), .Z(n8454) );
  MUX2_X1 U5334 ( .A(n10496), .B(n2560), .S(n1496), .Z(n8455) );
  MUX2_X1 U5335 ( .A(n10497), .B(n2549), .S(n1496), .Z(n8456) );
  MUX2_X1 U5336 ( .A(n10498), .B(n1834), .S(n1496), .Z(n8457) );
  MUX2_X1 U5337 ( .A(n10499), .B(n1823), .S(n1496), .Z(n8458) );
  MUX2_X1 U5338 ( .A(n10500), .B(n1812), .S(n1496), .Z(n8459) );
  MUX2_X1 U5339 ( .A(n10501), .B(n1801), .S(n1496), .Z(n8460) );
  MUX2_X1 U5340 ( .A(n10438), .B(n2949), .S(n1497), .Z(n8397) );
  MUX2_X1 U5341 ( .A(n10439), .B(n2938), .S(n1497), .Z(n8398) );
  MUX2_X1 U5342 ( .A(n10440), .B(n2927), .S(n1497), .Z(n8399) );
  MUX2_X1 U5343 ( .A(n10441), .B(n2911), .S(n1497), .Z(n8400) );
  MUX2_X1 U5344 ( .A(n10442), .B(n2900), .S(n1497), .Z(n8401) );
  MUX2_X1 U5345 ( .A(n10443), .B(n2888), .S(n1497), .Z(n8402) );
  MUX2_X1 U5346 ( .A(n10444), .B(n2877), .S(n1497), .Z(n8403) );
  MUX2_X1 U5347 ( .A(n10445), .B(n2866), .S(n1497), .Z(n8404) );
  MUX2_X1 U5348 ( .A(n10446), .B(n2855), .S(n1497), .Z(n8405) );
  MUX2_X1 U5349 ( .A(n10447), .B(n2844), .S(n1497), .Z(n8406) );
  MUX2_X1 U5350 ( .A(n10448), .B(n2833), .S(n1497), .Z(n8407) );
  MUX2_X1 U5351 ( .A(n10449), .B(n2822), .S(n1497), .Z(n8408) );
  MUX2_X1 U5352 ( .A(n10450), .B(n2811), .S(n1498), .Z(n8409) );
  MUX2_X1 U5353 ( .A(n10451), .B(n2800), .S(n1498), .Z(n8410) );
  MUX2_X1 U5354 ( .A(n10452), .B(n2789), .S(n1498), .Z(n8411) );
  MUX2_X1 U5355 ( .A(n10453), .B(n2778), .S(n1498), .Z(n8412) );
  MUX2_X1 U5356 ( .A(n10454), .B(n2767), .S(n1498), .Z(n8413) );
  MUX2_X1 U5357 ( .A(n10455), .B(n2756), .S(n1498), .Z(n8414) );
  MUX2_X1 U5358 ( .A(n10456), .B(n2745), .S(n1498), .Z(n8415) );
  MUX2_X1 U5359 ( .A(n10457), .B(n2734), .S(n1498), .Z(n8416) );
  MUX2_X1 U5360 ( .A(n10458), .B(n2723), .S(n1498), .Z(n8417) );
  MUX2_X1 U5361 ( .A(n10459), .B(n2712), .S(n1498), .Z(n8418) );
  MUX2_X1 U5362 ( .A(n10460), .B(n2605), .S(n1498), .Z(n8419) );
  MUX2_X1 U5363 ( .A(n10461), .B(n2594), .S(n1498), .Z(n8420) );
  MUX2_X1 U5364 ( .A(n10462), .B(n2583), .S(n1499), .Z(n8421) );
  MUX2_X1 U5365 ( .A(n10463), .B(n2572), .S(n1499), .Z(n8422) );
  MUX2_X1 U5366 ( .A(n10464), .B(n2561), .S(n1499), .Z(n8423) );
  MUX2_X1 U5367 ( .A(n10465), .B(n2550), .S(n1499), .Z(n8424) );
  MUX2_X1 U5368 ( .A(n10466), .B(n1835), .S(n1499), .Z(n8425) );
  MUX2_X1 U5369 ( .A(n10467), .B(n1824), .S(n1499), .Z(n8426) );
  MUX2_X1 U5370 ( .A(n10468), .B(n1813), .S(n1499), .Z(n8427) );
  MUX2_X1 U5371 ( .A(n10469), .B(n1802), .S(n1499), .Z(n8428) );
  MUX2_X1 U5372 ( .A(n10406), .B(n2949), .S(n1500), .Z(n8365) );
  MUX2_X1 U5373 ( .A(n10407), .B(n2938), .S(n1500), .Z(n8366) );
  MUX2_X1 U5374 ( .A(n10408), .B(n2927), .S(n1500), .Z(n8367) );
  MUX2_X1 U5375 ( .A(n10409), .B(n2911), .S(n1500), .Z(n8368) );
  MUX2_X1 U5376 ( .A(n10410), .B(n2900), .S(n1500), .Z(n8369) );
  MUX2_X1 U5377 ( .A(n10411), .B(n2888), .S(n1500), .Z(n8370) );
  MUX2_X1 U5378 ( .A(n10412), .B(n2877), .S(n1500), .Z(n8371) );
  MUX2_X1 U5379 ( .A(n10413), .B(n2866), .S(n1500), .Z(n8372) );
  MUX2_X1 U5380 ( .A(n10414), .B(n2855), .S(n1500), .Z(n8373) );
  MUX2_X1 U5381 ( .A(n10415), .B(n2844), .S(n1500), .Z(n8374) );
  MUX2_X1 U5382 ( .A(n10416), .B(n2833), .S(n1500), .Z(n8375) );
  MUX2_X1 U5383 ( .A(n10417), .B(n2822), .S(n1500), .Z(n8376) );
  MUX2_X1 U5384 ( .A(n10418), .B(n2811), .S(n1501), .Z(n8377) );
  MUX2_X1 U5385 ( .A(n10419), .B(n2800), .S(n1501), .Z(n8378) );
  MUX2_X1 U5386 ( .A(n10420), .B(n2789), .S(n1501), .Z(n8379) );
  MUX2_X1 U5387 ( .A(n10421), .B(n2778), .S(n1501), .Z(n8380) );
  MUX2_X1 U5388 ( .A(n10422), .B(n2767), .S(n1501), .Z(n8381) );
  MUX2_X1 U5389 ( .A(n10423), .B(n2756), .S(n1501), .Z(n8382) );
  MUX2_X1 U5390 ( .A(n10424), .B(n2745), .S(n1501), .Z(n8383) );
  MUX2_X1 U5391 ( .A(n10425), .B(n2734), .S(n1501), .Z(n8384) );
  MUX2_X1 U5392 ( .A(n10426), .B(n2723), .S(n1501), .Z(n8385) );
  MUX2_X1 U5393 ( .A(n10427), .B(n2712), .S(n1501), .Z(n8386) );
  MUX2_X1 U5394 ( .A(n10428), .B(n2605), .S(n1501), .Z(n8387) );
  MUX2_X1 U5395 ( .A(n10429), .B(n2594), .S(n1501), .Z(n8388) );
  MUX2_X1 U5396 ( .A(n10430), .B(n2583), .S(n1502), .Z(n8389) );
  MUX2_X1 U5397 ( .A(n10431), .B(n2572), .S(n1502), .Z(n8390) );
  MUX2_X1 U5398 ( .A(n10432), .B(n2561), .S(n1502), .Z(n8391) );
  MUX2_X1 U5399 ( .A(n10433), .B(n2550), .S(n1502), .Z(n8392) );
  MUX2_X1 U5400 ( .A(n10434), .B(n1835), .S(n1502), .Z(n8393) );
  MUX2_X1 U5401 ( .A(n10435), .B(n1824), .S(n1502), .Z(n8394) );
  MUX2_X1 U5402 ( .A(n10436), .B(n1813), .S(n1502), .Z(n8395) );
  MUX2_X1 U5403 ( .A(n10437), .B(n1802), .S(n1502), .Z(n8396) );
  MUX2_X1 U5404 ( .A(n10374), .B(n2949), .S(n1503), .Z(n8333) );
  MUX2_X1 U5405 ( .A(n10375), .B(n2938), .S(n1503), .Z(n8334) );
  MUX2_X1 U5406 ( .A(n10376), .B(n2927), .S(n1503), .Z(n8335) );
  MUX2_X1 U5407 ( .A(n10377), .B(n2911), .S(n1503), .Z(n8336) );
  MUX2_X1 U5408 ( .A(n10378), .B(n2900), .S(n1503), .Z(n8337) );
  MUX2_X1 U5409 ( .A(n10379), .B(n2888), .S(n1503), .Z(n8338) );
  MUX2_X1 U5410 ( .A(n10380), .B(n2877), .S(n1503), .Z(n8339) );
  MUX2_X1 U5411 ( .A(n10381), .B(n2866), .S(n1503), .Z(n8340) );
  MUX2_X1 U5412 ( .A(n10382), .B(n2855), .S(n1503), .Z(n8341) );
  MUX2_X1 U5413 ( .A(n10383), .B(n2844), .S(n1503), .Z(n8342) );
  MUX2_X1 U5414 ( .A(n10384), .B(n2833), .S(n1503), .Z(n8343) );
  MUX2_X1 U5415 ( .A(n10385), .B(n2822), .S(n1503), .Z(n8344) );
  MUX2_X1 U5416 ( .A(n10386), .B(n2811), .S(n1504), .Z(n8345) );
  MUX2_X1 U5417 ( .A(n10387), .B(n2800), .S(n1504), .Z(n8346) );
  MUX2_X1 U5418 ( .A(n10388), .B(n2789), .S(n1504), .Z(n8347) );
  MUX2_X1 U5419 ( .A(n10389), .B(n2778), .S(n1504), .Z(n8348) );
  MUX2_X1 U5420 ( .A(n10390), .B(n2767), .S(n1504), .Z(n8349) );
  MUX2_X1 U5421 ( .A(n10391), .B(n2756), .S(n1504), .Z(n8350) );
  MUX2_X1 U5422 ( .A(n10392), .B(n2745), .S(n1504), .Z(n8351) );
  MUX2_X1 U5423 ( .A(n10393), .B(n2734), .S(n1504), .Z(n8352) );
  MUX2_X1 U5424 ( .A(n10394), .B(n2723), .S(n1504), .Z(n8353) );
  MUX2_X1 U5425 ( .A(n10395), .B(n2712), .S(n1504), .Z(n8354) );
  MUX2_X1 U5426 ( .A(n10396), .B(n2605), .S(n1504), .Z(n8355) );
  MUX2_X1 U5427 ( .A(n10397), .B(n2594), .S(n1504), .Z(n8356) );
  MUX2_X1 U5428 ( .A(n10398), .B(n2583), .S(n1505), .Z(n8357) );
  MUX2_X1 U5429 ( .A(n10399), .B(n2572), .S(n1505), .Z(n8358) );
  MUX2_X1 U5430 ( .A(n10400), .B(n2561), .S(n1505), .Z(n8359) );
  MUX2_X1 U5431 ( .A(n10401), .B(n2550), .S(n1505), .Z(n8360) );
  MUX2_X1 U5432 ( .A(n10402), .B(n1835), .S(n1505), .Z(n8361) );
  MUX2_X1 U5433 ( .A(n10403), .B(n1824), .S(n1505), .Z(n8362) );
  MUX2_X1 U5434 ( .A(n10404), .B(n1813), .S(n1505), .Z(n8363) );
  MUX2_X1 U5435 ( .A(n10405), .B(n1802), .S(n1505), .Z(n8364) );
  MUX2_X1 U5436 ( .A(n10342), .B(n2949), .S(n1506), .Z(n8301) );
  MUX2_X1 U5437 ( .A(n10343), .B(n2938), .S(n1506), .Z(n8302) );
  MUX2_X1 U5438 ( .A(n10344), .B(n2927), .S(n1506), .Z(n8303) );
  MUX2_X1 U5439 ( .A(n10345), .B(n2911), .S(n1506), .Z(n8304) );
  MUX2_X1 U5440 ( .A(n10346), .B(n2900), .S(n1506), .Z(n8305) );
  MUX2_X1 U5441 ( .A(n10347), .B(n2888), .S(n1506), .Z(n8306) );
  MUX2_X1 U5442 ( .A(n10348), .B(n2877), .S(n1506), .Z(n8307) );
  MUX2_X1 U5443 ( .A(n10349), .B(n2866), .S(n1506), .Z(n8308) );
  MUX2_X1 U5444 ( .A(n10350), .B(n2855), .S(n1506), .Z(n8309) );
  MUX2_X1 U5445 ( .A(n10351), .B(n2844), .S(n1506), .Z(n8310) );
  MUX2_X1 U5446 ( .A(n10352), .B(n2833), .S(n1506), .Z(n8311) );
  MUX2_X1 U5447 ( .A(n10353), .B(n2822), .S(n1506), .Z(n8312) );
  MUX2_X1 U5448 ( .A(n10354), .B(n2811), .S(n1507), .Z(n8313) );
  MUX2_X1 U5449 ( .A(n10355), .B(n2800), .S(n1507), .Z(n8314) );
  MUX2_X1 U5450 ( .A(n10356), .B(n2789), .S(n1507), .Z(n8315) );
  MUX2_X1 U5451 ( .A(n10357), .B(n2778), .S(n1507), .Z(n8316) );
  MUX2_X1 U5452 ( .A(n10358), .B(n2767), .S(n1507), .Z(n8317) );
  MUX2_X1 U5453 ( .A(n10359), .B(n2756), .S(n1507), .Z(n8318) );
  MUX2_X1 U5454 ( .A(n10360), .B(n2745), .S(n1507), .Z(n8319) );
  MUX2_X1 U5455 ( .A(n10361), .B(n2734), .S(n1507), .Z(n8320) );
  MUX2_X1 U5456 ( .A(n10362), .B(n2723), .S(n1507), .Z(n8321) );
  MUX2_X1 U5457 ( .A(n10363), .B(n2712), .S(n1507), .Z(n8322) );
  MUX2_X1 U5458 ( .A(n10364), .B(n2605), .S(n1507), .Z(n8323) );
  MUX2_X1 U5459 ( .A(n10365), .B(n2594), .S(n1507), .Z(n8324) );
  MUX2_X1 U5460 ( .A(n10366), .B(n2583), .S(n1508), .Z(n8325) );
  MUX2_X1 U5461 ( .A(n10367), .B(n2572), .S(n1508), .Z(n8326) );
  MUX2_X1 U5462 ( .A(n10368), .B(n2561), .S(n1508), .Z(n8327) );
  MUX2_X1 U5463 ( .A(n10369), .B(n2550), .S(n1508), .Z(n8328) );
  MUX2_X1 U5464 ( .A(n10370), .B(n1835), .S(n1508), .Z(n8329) );
  MUX2_X1 U5465 ( .A(n10371), .B(n1824), .S(n1508), .Z(n8330) );
  MUX2_X1 U5466 ( .A(n10372), .B(n1813), .S(n1508), .Z(n8331) );
  MUX2_X1 U5467 ( .A(n10373), .B(n1802), .S(n1508), .Z(n8332) );
  MUX2_X1 U5468 ( .A(n10310), .B(n2949), .S(n1509), .Z(n8269) );
  MUX2_X1 U5469 ( .A(n10311), .B(n2938), .S(n1509), .Z(n8270) );
  MUX2_X1 U5470 ( .A(n10312), .B(n2927), .S(n1509), .Z(n8271) );
  MUX2_X1 U5471 ( .A(n10313), .B(n2911), .S(n1509), .Z(n8272) );
  MUX2_X1 U5472 ( .A(n10314), .B(n2900), .S(n1509), .Z(n8273) );
  MUX2_X1 U5473 ( .A(n10315), .B(n2888), .S(n1509), .Z(n8274) );
  MUX2_X1 U5474 ( .A(n10316), .B(n2877), .S(n1509), .Z(n8275) );
  MUX2_X1 U5475 ( .A(n10317), .B(n2866), .S(n1509), .Z(n8276) );
  MUX2_X1 U5476 ( .A(n10318), .B(n2855), .S(n1509), .Z(n8277) );
  MUX2_X1 U5477 ( .A(n10319), .B(n2844), .S(n1509), .Z(n8278) );
  MUX2_X1 U5478 ( .A(n10320), .B(n2833), .S(n1509), .Z(n8279) );
  MUX2_X1 U5479 ( .A(n10321), .B(n2822), .S(n1509), .Z(n8280) );
  MUX2_X1 U5480 ( .A(n10322), .B(n2811), .S(n1510), .Z(n8281) );
  MUX2_X1 U5481 ( .A(n10323), .B(n2800), .S(n1510), .Z(n8282) );
  MUX2_X1 U5482 ( .A(n10324), .B(n2789), .S(n1510), .Z(n8283) );
  MUX2_X1 U5483 ( .A(n10325), .B(n2778), .S(n1510), .Z(n8284) );
  MUX2_X1 U5484 ( .A(n10326), .B(n2767), .S(n1510), .Z(n8285) );
  MUX2_X1 U5485 ( .A(n10327), .B(n2756), .S(n1510), .Z(n8286) );
  MUX2_X1 U5486 ( .A(n10328), .B(n2745), .S(n1510), .Z(n8287) );
  MUX2_X1 U5487 ( .A(n10329), .B(n2734), .S(n1510), .Z(n8288) );
  MUX2_X1 U5488 ( .A(n10330), .B(n2723), .S(n1510), .Z(n8289) );
  MUX2_X1 U5489 ( .A(n10331), .B(n2712), .S(n1510), .Z(n8290) );
  MUX2_X1 U5490 ( .A(n10332), .B(n2605), .S(n1510), .Z(n8291) );
  MUX2_X1 U5491 ( .A(n10333), .B(n2594), .S(n1510), .Z(n8292) );
  MUX2_X1 U5492 ( .A(n10334), .B(n2583), .S(n1511), .Z(n8293) );
  MUX2_X1 U5493 ( .A(n10335), .B(n2572), .S(n1511), .Z(n8294) );
  MUX2_X1 U5494 ( .A(n10336), .B(n2561), .S(n1511), .Z(n8295) );
  MUX2_X1 U5495 ( .A(n10337), .B(n2550), .S(n1511), .Z(n8296) );
  MUX2_X1 U5496 ( .A(n10338), .B(n1835), .S(n1511), .Z(n8297) );
  MUX2_X1 U5497 ( .A(n10339), .B(n1824), .S(n1511), .Z(n8298) );
  MUX2_X1 U5498 ( .A(n10340), .B(n1813), .S(n1511), .Z(n8299) );
  MUX2_X1 U5499 ( .A(n10341), .B(n1802), .S(n1511), .Z(n8300) );
  MUX2_X1 U5500 ( .A(n10278), .B(n2949), .S(n1512), .Z(n8237) );
  MUX2_X1 U5501 ( .A(n10279), .B(n2938), .S(n1512), .Z(n8238) );
  MUX2_X1 U5502 ( .A(n10280), .B(n2927), .S(n1512), .Z(n8239) );
  MUX2_X1 U5503 ( .A(n10281), .B(n2911), .S(n1512), .Z(n8240) );
  MUX2_X1 U5504 ( .A(n10282), .B(n2900), .S(n1512), .Z(n8241) );
  MUX2_X1 U5505 ( .A(n10283), .B(n2888), .S(n1512), .Z(n8242) );
  MUX2_X1 U5506 ( .A(n10284), .B(n2877), .S(n1512), .Z(n8243) );
  MUX2_X1 U5507 ( .A(n10285), .B(n2866), .S(n1512), .Z(n8244) );
  MUX2_X1 U5508 ( .A(n10286), .B(n2855), .S(n1512), .Z(n8245) );
  MUX2_X1 U5509 ( .A(n10287), .B(n2844), .S(n1512), .Z(n8246) );
  MUX2_X1 U5510 ( .A(n10288), .B(n2833), .S(n1512), .Z(n8247) );
  MUX2_X1 U5511 ( .A(n10289), .B(n2822), .S(n1512), .Z(n8248) );
  MUX2_X1 U5512 ( .A(n10290), .B(n2811), .S(n1513), .Z(n8249) );
  MUX2_X1 U5513 ( .A(n10291), .B(n2800), .S(n1513), .Z(n8250) );
  MUX2_X1 U5514 ( .A(n10292), .B(n2789), .S(n1513), .Z(n8251) );
  MUX2_X1 U5515 ( .A(n10293), .B(n2778), .S(n1513), .Z(n8252) );
  MUX2_X1 U5516 ( .A(n10294), .B(n2767), .S(n1513), .Z(n8253) );
  MUX2_X1 U5517 ( .A(n10295), .B(n2756), .S(n1513), .Z(n8254) );
  MUX2_X1 U5518 ( .A(n10296), .B(n2745), .S(n1513), .Z(n8255) );
  MUX2_X1 U5519 ( .A(n10297), .B(n2734), .S(n1513), .Z(n8256) );
  MUX2_X1 U5520 ( .A(n10298), .B(n2723), .S(n1513), .Z(n8257) );
  MUX2_X1 U5521 ( .A(n10299), .B(n2712), .S(n1513), .Z(n8258) );
  MUX2_X1 U5522 ( .A(n10300), .B(n2605), .S(n1513), .Z(n8259) );
  MUX2_X1 U5523 ( .A(n10301), .B(n2594), .S(n1513), .Z(n8260) );
  MUX2_X1 U5524 ( .A(n10302), .B(n2583), .S(n1514), .Z(n8261) );
  MUX2_X1 U5525 ( .A(n10303), .B(n2572), .S(n1514), .Z(n8262) );
  MUX2_X1 U5526 ( .A(n10304), .B(n2561), .S(n1514), .Z(n8263) );
  MUX2_X1 U5527 ( .A(n10305), .B(n2550), .S(n1514), .Z(n8264) );
  MUX2_X1 U5528 ( .A(n10306), .B(n1835), .S(n1514), .Z(n8265) );
  MUX2_X1 U5529 ( .A(n10307), .B(n1824), .S(n1514), .Z(n8266) );
  MUX2_X1 U5530 ( .A(n10308), .B(n1813), .S(n1514), .Z(n8267) );
  MUX2_X1 U5531 ( .A(n10309), .B(n1802), .S(n1514), .Z(n8268) );
  MUX2_X1 U5532 ( .A(n10246), .B(n2949), .S(n1515), .Z(n8205) );
  MUX2_X1 U5533 ( .A(n10247), .B(n2938), .S(n1515), .Z(n8206) );
  MUX2_X1 U5534 ( .A(n10248), .B(n2927), .S(n1515), .Z(n8207) );
  MUX2_X1 U5535 ( .A(n10249), .B(n2911), .S(n1515), .Z(n8208) );
  MUX2_X1 U5536 ( .A(n10250), .B(n2900), .S(n1515), .Z(n8209) );
  MUX2_X1 U5537 ( .A(n10251), .B(n2888), .S(n1515), .Z(n8210) );
  MUX2_X1 U5538 ( .A(n10252), .B(n2877), .S(n1515), .Z(n8211) );
  MUX2_X1 U5539 ( .A(n10253), .B(n2866), .S(n1515), .Z(n8212) );
  MUX2_X1 U5540 ( .A(n10254), .B(n2855), .S(n1515), .Z(n8213) );
  MUX2_X1 U5541 ( .A(n10255), .B(n2844), .S(n1515), .Z(n8214) );
  MUX2_X1 U5542 ( .A(n10256), .B(n2833), .S(n1515), .Z(n8215) );
  MUX2_X1 U5543 ( .A(n10257), .B(n2822), .S(n1515), .Z(n8216) );
  MUX2_X1 U5544 ( .A(n10258), .B(n2811), .S(n1516), .Z(n8217) );
  MUX2_X1 U5545 ( .A(n10259), .B(n2800), .S(n1516), .Z(n8218) );
  MUX2_X1 U5546 ( .A(n10260), .B(n2789), .S(n1516), .Z(n8219) );
  MUX2_X1 U5547 ( .A(n10261), .B(n2778), .S(n1516), .Z(n8220) );
  MUX2_X1 U5548 ( .A(n10262), .B(n2767), .S(n1516), .Z(n8221) );
  MUX2_X1 U5549 ( .A(n10263), .B(n2756), .S(n1516), .Z(n8222) );
  MUX2_X1 U5550 ( .A(n10264), .B(n2745), .S(n1516), .Z(n8223) );
  MUX2_X1 U5551 ( .A(n10265), .B(n2734), .S(n1516), .Z(n8224) );
  MUX2_X1 U5552 ( .A(n10266), .B(n2723), .S(n1516), .Z(n8225) );
  MUX2_X1 U5553 ( .A(n10267), .B(n2712), .S(n1516), .Z(n8226) );
  MUX2_X1 U5554 ( .A(n10268), .B(n2605), .S(n1516), .Z(n8227) );
  MUX2_X1 U5555 ( .A(n10269), .B(n2594), .S(n1516), .Z(n8228) );
  MUX2_X1 U5556 ( .A(n10270), .B(n2583), .S(n1517), .Z(n8229) );
  MUX2_X1 U5557 ( .A(n10271), .B(n2572), .S(n1517), .Z(n8230) );
  MUX2_X1 U5558 ( .A(n10272), .B(n2561), .S(n1517), .Z(n8231) );
  MUX2_X1 U5559 ( .A(n10273), .B(n2550), .S(n1517), .Z(n8232) );
  MUX2_X1 U5560 ( .A(n10274), .B(n1835), .S(n1517), .Z(n8233) );
  MUX2_X1 U5561 ( .A(n10275), .B(n1824), .S(n1517), .Z(n8234) );
  MUX2_X1 U5562 ( .A(n10276), .B(n1813), .S(n1517), .Z(n8235) );
  MUX2_X1 U5563 ( .A(n10277), .B(n1802), .S(n1517), .Z(n8236) );
  MUX2_X1 U5564 ( .A(n10214), .B(n2949), .S(n1518), .Z(n8173) );
  MUX2_X1 U5565 ( .A(n10215), .B(n2938), .S(n1518), .Z(n8174) );
  MUX2_X1 U5566 ( .A(n10216), .B(n2927), .S(n1518), .Z(n8175) );
  MUX2_X1 U5567 ( .A(n10217), .B(n2911), .S(n1518), .Z(n8176) );
  MUX2_X1 U5568 ( .A(n10218), .B(n2900), .S(n1518), .Z(n8177) );
  MUX2_X1 U5569 ( .A(n10219), .B(n2888), .S(n1518), .Z(n8178) );
  MUX2_X1 U5570 ( .A(n10220), .B(n2877), .S(n1518), .Z(n8179) );
  MUX2_X1 U5571 ( .A(n10221), .B(n2866), .S(n1518), .Z(n8180) );
  MUX2_X1 U5572 ( .A(n10222), .B(n2855), .S(n1518), .Z(n8181) );
  MUX2_X1 U5573 ( .A(n10223), .B(n2844), .S(n1518), .Z(n8182) );
  MUX2_X1 U5574 ( .A(n10224), .B(n2833), .S(n1518), .Z(n8183) );
  MUX2_X1 U5575 ( .A(n10225), .B(n2822), .S(n1518), .Z(n8184) );
  MUX2_X1 U5576 ( .A(n10226), .B(n2811), .S(n1519), .Z(n8185) );
  MUX2_X1 U5577 ( .A(n10227), .B(n2800), .S(n1519), .Z(n8186) );
  MUX2_X1 U5578 ( .A(n10228), .B(n2789), .S(n1519), .Z(n8187) );
  MUX2_X1 U5579 ( .A(n10229), .B(n2778), .S(n1519), .Z(n8188) );
  MUX2_X1 U5580 ( .A(n10230), .B(n2767), .S(n1519), .Z(n8189) );
  MUX2_X1 U5581 ( .A(n10231), .B(n2756), .S(n1519), .Z(n8190) );
  MUX2_X1 U5582 ( .A(n10232), .B(n2745), .S(n1519), .Z(n8191) );
  MUX2_X1 U5583 ( .A(n10233), .B(n2734), .S(n1519), .Z(n8192) );
  MUX2_X1 U5584 ( .A(n10234), .B(n2723), .S(n1519), .Z(n8193) );
  MUX2_X1 U5585 ( .A(n10235), .B(n2712), .S(n1519), .Z(n8194) );
  MUX2_X1 U5586 ( .A(n10236), .B(n2605), .S(n1519), .Z(n8195) );
  MUX2_X1 U5587 ( .A(n10237), .B(n2594), .S(n1519), .Z(n8196) );
  MUX2_X1 U5588 ( .A(n10238), .B(n2583), .S(n1520), .Z(n8197) );
  MUX2_X1 U5589 ( .A(n10239), .B(n2572), .S(n1520), .Z(n8198) );
  MUX2_X1 U5590 ( .A(n10240), .B(n2561), .S(n1520), .Z(n8199) );
  MUX2_X1 U5591 ( .A(n10241), .B(n2550), .S(n1520), .Z(n8200) );
  MUX2_X1 U5592 ( .A(n10242), .B(n1835), .S(n1520), .Z(n8201) );
  MUX2_X1 U5593 ( .A(n10243), .B(n1824), .S(n1520), .Z(n8202) );
  MUX2_X1 U5594 ( .A(n10244), .B(n1813), .S(n1520), .Z(n8203) );
  MUX2_X1 U5595 ( .A(n10245), .B(n1802), .S(n1520), .Z(n8204) );
  MUX2_X1 U5596 ( .A(n10182), .B(n2949), .S(n1521), .Z(n8141) );
  MUX2_X1 U5597 ( .A(n10183), .B(n2938), .S(n1521), .Z(n8142) );
  MUX2_X1 U5598 ( .A(n10184), .B(n2927), .S(n1521), .Z(n8143) );
  MUX2_X1 U5599 ( .A(n10185), .B(n2911), .S(n1521), .Z(n8144) );
  MUX2_X1 U5600 ( .A(n10186), .B(n2900), .S(n1521), .Z(n8145) );
  MUX2_X1 U5601 ( .A(n10187), .B(n2888), .S(n1521), .Z(n8146) );
  MUX2_X1 U5602 ( .A(n10188), .B(n2877), .S(n1521), .Z(n8147) );
  MUX2_X1 U5603 ( .A(n10189), .B(n2866), .S(n1521), .Z(n8148) );
  MUX2_X1 U5604 ( .A(n10190), .B(n2855), .S(n1521), .Z(n8149) );
  MUX2_X1 U5605 ( .A(n10191), .B(n2844), .S(n1521), .Z(n8150) );
  MUX2_X1 U5606 ( .A(n10192), .B(n2833), .S(n1521), .Z(n8151) );
  MUX2_X1 U5607 ( .A(n10193), .B(n2822), .S(n1521), .Z(n8152) );
  MUX2_X1 U5608 ( .A(n10194), .B(n2811), .S(n1522), .Z(n8153) );
  MUX2_X1 U5609 ( .A(n10195), .B(n2800), .S(n1522), .Z(n8154) );
  MUX2_X1 U5610 ( .A(n10196), .B(n2789), .S(n1522), .Z(n8155) );
  MUX2_X1 U5611 ( .A(n10197), .B(n2778), .S(n1522), .Z(n8156) );
  MUX2_X1 U5612 ( .A(n10198), .B(n2767), .S(n1522), .Z(n8157) );
  MUX2_X1 U5613 ( .A(n10199), .B(n2756), .S(n1522), .Z(n8158) );
  MUX2_X1 U5614 ( .A(n10200), .B(n2745), .S(n1522), .Z(n8159) );
  MUX2_X1 U5615 ( .A(n10201), .B(n2734), .S(n1522), .Z(n8160) );
  MUX2_X1 U5616 ( .A(n10202), .B(n2723), .S(n1522), .Z(n8161) );
  MUX2_X1 U5617 ( .A(n10203), .B(n2712), .S(n1522), .Z(n8162) );
  MUX2_X1 U5618 ( .A(n10204), .B(n2605), .S(n1522), .Z(n8163) );
  MUX2_X1 U5619 ( .A(n10205), .B(n2594), .S(n1522), .Z(n8164) );
  MUX2_X1 U5620 ( .A(n10206), .B(n2583), .S(n1523), .Z(n8165) );
  MUX2_X1 U5621 ( .A(n10207), .B(n2572), .S(n1523), .Z(n8166) );
  MUX2_X1 U5622 ( .A(n10208), .B(n2561), .S(n1523), .Z(n8167) );
  MUX2_X1 U5623 ( .A(n10209), .B(n2550), .S(n1523), .Z(n8168) );
  MUX2_X1 U5624 ( .A(n10210), .B(n1835), .S(n1523), .Z(n8169) );
  MUX2_X1 U5625 ( .A(n10211), .B(n1824), .S(n1523), .Z(n8170) );
  MUX2_X1 U5626 ( .A(n10212), .B(n1813), .S(n1523), .Z(n8171) );
  MUX2_X1 U5627 ( .A(n10213), .B(n1802), .S(n1523), .Z(n8172) );
  MUX2_X1 U5628 ( .A(n10150), .B(n2949), .S(n1524), .Z(n8109) );
  MUX2_X1 U5629 ( .A(n10151), .B(n2938), .S(n1524), .Z(n8110) );
  MUX2_X1 U5630 ( .A(n10152), .B(n2927), .S(n1524), .Z(n8111) );
  MUX2_X1 U5631 ( .A(n10153), .B(n2911), .S(n1524), .Z(n8112) );
  MUX2_X1 U5632 ( .A(n10154), .B(n2900), .S(n1524), .Z(n8113) );
  MUX2_X1 U5633 ( .A(n10155), .B(n2888), .S(n1524), .Z(n8114) );
  MUX2_X1 U5634 ( .A(n10156), .B(n2877), .S(n1524), .Z(n8115) );
  MUX2_X1 U5635 ( .A(n10157), .B(n2866), .S(n1524), .Z(n8116) );
  MUX2_X1 U5636 ( .A(n10158), .B(n2855), .S(n1524), .Z(n8117) );
  MUX2_X1 U5637 ( .A(n10159), .B(n2844), .S(n1524), .Z(n8118) );
  MUX2_X1 U5638 ( .A(n10160), .B(n2833), .S(n1524), .Z(n8119) );
  MUX2_X1 U5639 ( .A(n10161), .B(n2822), .S(n1524), .Z(n8120) );
  MUX2_X1 U5640 ( .A(n10162), .B(n2811), .S(n1525), .Z(n8121) );
  MUX2_X1 U5641 ( .A(n10163), .B(n2800), .S(n1525), .Z(n8122) );
  MUX2_X1 U5642 ( .A(n10164), .B(n2789), .S(n1525), .Z(n8123) );
  MUX2_X1 U5643 ( .A(n10165), .B(n2778), .S(n1525), .Z(n8124) );
  MUX2_X1 U5644 ( .A(n10166), .B(n2767), .S(n1525), .Z(n8125) );
  MUX2_X1 U5645 ( .A(n10167), .B(n2756), .S(n1525), .Z(n8126) );
  MUX2_X1 U5646 ( .A(n10168), .B(n2745), .S(n1525), .Z(n8127) );
  MUX2_X1 U5647 ( .A(n10169), .B(n2734), .S(n1525), .Z(n8128) );
  MUX2_X1 U5648 ( .A(n10170), .B(n2723), .S(n1525), .Z(n8129) );
  MUX2_X1 U5649 ( .A(n10171), .B(n2712), .S(n1525), .Z(n8130) );
  MUX2_X1 U5650 ( .A(n10172), .B(n2605), .S(n1525), .Z(n8131) );
  MUX2_X1 U5651 ( .A(n10173), .B(n2594), .S(n1525), .Z(n8132) );
  MUX2_X1 U5652 ( .A(n10174), .B(n2583), .S(n1526), .Z(n8133) );
  MUX2_X1 U5653 ( .A(n10175), .B(n2572), .S(n1526), .Z(n8134) );
  MUX2_X1 U5654 ( .A(n10176), .B(n2561), .S(n1526), .Z(n8135) );
  MUX2_X1 U5655 ( .A(n10177), .B(n2550), .S(n1526), .Z(n8136) );
  MUX2_X1 U5656 ( .A(n10178), .B(n1835), .S(n1526), .Z(n8137) );
  MUX2_X1 U5657 ( .A(n10179), .B(n1824), .S(n1526), .Z(n8138) );
  MUX2_X1 U5658 ( .A(n10180), .B(n1813), .S(n1526), .Z(n8139) );
  MUX2_X1 U5659 ( .A(n10181), .B(n1802), .S(n1526), .Z(n8140) );
  MUX2_X1 U5660 ( .A(n10118), .B(n2949), .S(n1527), .Z(n8077) );
  MUX2_X1 U5661 ( .A(n10119), .B(n2938), .S(n1527), .Z(n8078) );
  MUX2_X1 U5662 ( .A(n10120), .B(n2927), .S(n1527), .Z(n8079) );
  MUX2_X1 U5663 ( .A(n10121), .B(n2911), .S(n1527), .Z(n8080) );
  MUX2_X1 U5664 ( .A(n10122), .B(n2900), .S(n1527), .Z(n8081) );
  MUX2_X1 U5665 ( .A(n10123), .B(n2888), .S(n1527), .Z(n8082) );
  MUX2_X1 U5666 ( .A(n10124), .B(n2877), .S(n1527), .Z(n8083) );
  MUX2_X1 U5667 ( .A(n10125), .B(n2866), .S(n1527), .Z(n8084) );
  MUX2_X1 U5668 ( .A(n10126), .B(n2855), .S(n1527), .Z(n8085) );
  MUX2_X1 U5669 ( .A(n10127), .B(n2844), .S(n1527), .Z(n8086) );
  MUX2_X1 U5670 ( .A(n10128), .B(n2833), .S(n1527), .Z(n8087) );
  MUX2_X1 U5671 ( .A(n10129), .B(n2822), .S(n1527), .Z(n8088) );
  MUX2_X1 U5672 ( .A(n10130), .B(n2811), .S(n1528), .Z(n8089) );
  MUX2_X1 U5673 ( .A(n10131), .B(n2800), .S(n1528), .Z(n8090) );
  MUX2_X1 U5674 ( .A(n10132), .B(n2789), .S(n1528), .Z(n8091) );
  MUX2_X1 U5675 ( .A(n10133), .B(n2778), .S(n1528), .Z(n8092) );
  MUX2_X1 U5676 ( .A(n10134), .B(n2767), .S(n1528), .Z(n8093) );
  MUX2_X1 U5677 ( .A(n10135), .B(n2756), .S(n1528), .Z(n8094) );
  MUX2_X1 U5678 ( .A(n10136), .B(n2745), .S(n1528), .Z(n8095) );
  MUX2_X1 U5679 ( .A(n10137), .B(n2734), .S(n1528), .Z(n8096) );
  MUX2_X1 U5680 ( .A(n10138), .B(n2723), .S(n1528), .Z(n8097) );
  MUX2_X1 U5681 ( .A(n10139), .B(n2712), .S(n1528), .Z(n8098) );
  MUX2_X1 U5682 ( .A(n10140), .B(n2605), .S(n1528), .Z(n8099) );
  MUX2_X1 U5683 ( .A(n10141), .B(n2594), .S(n1528), .Z(n8100) );
  MUX2_X1 U5684 ( .A(n10142), .B(n2583), .S(n1529), .Z(n8101) );
  MUX2_X1 U5685 ( .A(n10143), .B(n2572), .S(n1529), .Z(n8102) );
  MUX2_X1 U5686 ( .A(n10144), .B(n2561), .S(n1529), .Z(n8103) );
  MUX2_X1 U5687 ( .A(n10145), .B(n2550), .S(n1529), .Z(n8104) );
  MUX2_X1 U5688 ( .A(n10146), .B(n1835), .S(n1529), .Z(n8105) );
  MUX2_X1 U5689 ( .A(n10147), .B(n1824), .S(n1529), .Z(n8106) );
  MUX2_X1 U5690 ( .A(n10148), .B(n1813), .S(n1529), .Z(n8107) );
  MUX2_X1 U5691 ( .A(n10149), .B(n1802), .S(n1529), .Z(n8108) );
  MUX2_X1 U5692 ( .A(\REGISTERS[54][31] ), .B(n2950), .S(n1530), .Z(n8045) );
  MUX2_X1 U5693 ( .A(\REGISTERS[54][30] ), .B(n2939), .S(n1530), .Z(n8046) );
  MUX2_X1 U5694 ( .A(\REGISTERS[54][29] ), .B(n2928), .S(n1530), .Z(n8047) );
  MUX2_X1 U5695 ( .A(\REGISTERS[54][28] ), .B(n2912), .S(n1530), .Z(n8048) );
  MUX2_X1 U5696 ( .A(\REGISTERS[54][27] ), .B(n2901), .S(n1530), .Z(n8049) );
  MUX2_X1 U5697 ( .A(\REGISTERS[54][26] ), .B(n2889), .S(n1530), .Z(n8050) );
  MUX2_X1 U5698 ( .A(\REGISTERS[54][25] ), .B(n2878), .S(n1530), .Z(n8051) );
  MUX2_X1 U5699 ( .A(\REGISTERS[54][24] ), .B(n2867), .S(n1530), .Z(n8052) );
  MUX2_X1 U5700 ( .A(\REGISTERS[54][23] ), .B(n2856), .S(n1530), .Z(n8053) );
  MUX2_X1 U5701 ( .A(\REGISTERS[54][22] ), .B(n2845), .S(n1530), .Z(n8054) );
  MUX2_X1 U5702 ( .A(\REGISTERS[54][21] ), .B(n2834), .S(n1530), .Z(n8055) );
  MUX2_X1 U5703 ( .A(\REGISTERS[54][20] ), .B(n2823), .S(n1530), .Z(n8056) );
  MUX2_X1 U5704 ( .A(\REGISTERS[54][19] ), .B(n2812), .S(n1531), .Z(n8057) );
  MUX2_X1 U5705 ( .A(\REGISTERS[54][18] ), .B(n2801), .S(n1531), .Z(n8058) );
  MUX2_X1 U5706 ( .A(\REGISTERS[54][17] ), .B(n2790), .S(n1531), .Z(n8059) );
  MUX2_X1 U5707 ( .A(\REGISTERS[54][16] ), .B(n2779), .S(n1531), .Z(n8060) );
  MUX2_X1 U5708 ( .A(\REGISTERS[54][15] ), .B(n2768), .S(n1531), .Z(n8061) );
  MUX2_X1 U5709 ( .A(\REGISTERS[54][14] ), .B(n2757), .S(n1531), .Z(n8062) );
  MUX2_X1 U5710 ( .A(\REGISTERS[54][13] ), .B(n2746), .S(n1531), .Z(n8063) );
  MUX2_X1 U5711 ( .A(\REGISTERS[54][12] ), .B(n2735), .S(n1531), .Z(n8064) );
  MUX2_X1 U5712 ( .A(\REGISTERS[54][11] ), .B(n2724), .S(n1531), .Z(n8065) );
  MUX2_X1 U5713 ( .A(\REGISTERS[54][10] ), .B(n2713), .S(n1531), .Z(n8066) );
  MUX2_X1 U5714 ( .A(\REGISTERS[54][9] ), .B(n2606), .S(n1531), .Z(n8067) );
  MUX2_X1 U5715 ( .A(\REGISTERS[54][8] ), .B(n2595), .S(n1531), .Z(n8068) );
  MUX2_X1 U5716 ( .A(\REGISTERS[54][7] ), .B(n2584), .S(n1532), .Z(n8069) );
  MUX2_X1 U5717 ( .A(\REGISTERS[54][6] ), .B(n2573), .S(n1532), .Z(n8070) );
  MUX2_X1 U5718 ( .A(\REGISTERS[54][5] ), .B(n2562), .S(n1532), .Z(n8071) );
  MUX2_X1 U5719 ( .A(\REGISTERS[54][4] ), .B(n2551), .S(n1532), .Z(n8072) );
  MUX2_X1 U5720 ( .A(\REGISTERS[54][3] ), .B(n1836), .S(n1532), .Z(n8073) );
  MUX2_X1 U5721 ( .A(\REGISTERS[54][2] ), .B(n1825), .S(n1532), .Z(n8074) );
  MUX2_X1 U5722 ( .A(\REGISTERS[54][1] ), .B(n1814), .S(n1532), .Z(n8075) );
  MUX2_X1 U5723 ( .A(\REGISTERS[54][0] ), .B(n1803), .S(n1532), .Z(n8076) );
  MUX2_X1 U5724 ( .A(\REGISTERS[53][31] ), .B(n2950), .S(n1533), .Z(n8013) );
  MUX2_X1 U5725 ( .A(\REGISTERS[53][30] ), .B(n2939), .S(n1533), .Z(n8014) );
  MUX2_X1 U5726 ( .A(\REGISTERS[53][29] ), .B(n2928), .S(n1533), .Z(n8015) );
  MUX2_X1 U5727 ( .A(\REGISTERS[53][28] ), .B(n2912), .S(n1533), .Z(n8016) );
  MUX2_X1 U5728 ( .A(\REGISTERS[53][27] ), .B(n2901), .S(n1533), .Z(n8017) );
  MUX2_X1 U5729 ( .A(\REGISTERS[53][26] ), .B(n2889), .S(n1533), .Z(n8018) );
  MUX2_X1 U5730 ( .A(\REGISTERS[53][25] ), .B(n2878), .S(n1533), .Z(n8019) );
  MUX2_X1 U5731 ( .A(\REGISTERS[53][24] ), .B(n2867), .S(n1533), .Z(n8020) );
  MUX2_X1 U5732 ( .A(\REGISTERS[53][23] ), .B(n2856), .S(n1533), .Z(n8021) );
  MUX2_X1 U5733 ( .A(\REGISTERS[53][22] ), .B(n2845), .S(n1533), .Z(n8022) );
  MUX2_X1 U5734 ( .A(\REGISTERS[53][21] ), .B(n2834), .S(n1533), .Z(n8023) );
  MUX2_X1 U5735 ( .A(\REGISTERS[53][20] ), .B(n2823), .S(n1533), .Z(n8024) );
  MUX2_X1 U5736 ( .A(\REGISTERS[53][19] ), .B(n2812), .S(n1534), .Z(n8025) );
  MUX2_X1 U5737 ( .A(\REGISTERS[53][18] ), .B(n2801), .S(n1534), .Z(n8026) );
  MUX2_X1 U5738 ( .A(\REGISTERS[53][17] ), .B(n2790), .S(n1534), .Z(n8027) );
  MUX2_X1 U5739 ( .A(\REGISTERS[53][16] ), .B(n2779), .S(n1534), .Z(n8028) );
  MUX2_X1 U5740 ( .A(\REGISTERS[53][15] ), .B(n2768), .S(n1534), .Z(n8029) );
  MUX2_X1 U5741 ( .A(\REGISTERS[53][14] ), .B(n2757), .S(n1534), .Z(n8030) );
  MUX2_X1 U5742 ( .A(\REGISTERS[53][13] ), .B(n2746), .S(n1534), .Z(n8031) );
  MUX2_X1 U5743 ( .A(\REGISTERS[53][12] ), .B(n2735), .S(n1534), .Z(n8032) );
  MUX2_X1 U5744 ( .A(\REGISTERS[53][11] ), .B(n2724), .S(n1534), .Z(n8033) );
  MUX2_X1 U5745 ( .A(\REGISTERS[53][10] ), .B(n2713), .S(n1534), .Z(n8034) );
  MUX2_X1 U5746 ( .A(\REGISTERS[53][9] ), .B(n2606), .S(n1534), .Z(n8035) );
  MUX2_X1 U5747 ( .A(\REGISTERS[53][8] ), .B(n2595), .S(n1534), .Z(n8036) );
  MUX2_X1 U5748 ( .A(\REGISTERS[53][7] ), .B(n2584), .S(n1535), .Z(n8037) );
  MUX2_X1 U5749 ( .A(\REGISTERS[53][6] ), .B(n2573), .S(n1535), .Z(n8038) );
  MUX2_X1 U5750 ( .A(\REGISTERS[53][5] ), .B(n2562), .S(n1535), .Z(n8039) );
  MUX2_X1 U5751 ( .A(\REGISTERS[53][4] ), .B(n2551), .S(n1535), .Z(n8040) );
  MUX2_X1 U5752 ( .A(\REGISTERS[53][3] ), .B(n1836), .S(n1535), .Z(n8041) );
  MUX2_X1 U5753 ( .A(\REGISTERS[53][2] ), .B(n1825), .S(n1535), .Z(n8042) );
  MUX2_X1 U5754 ( .A(\REGISTERS[53][1] ), .B(n1814), .S(n1535), .Z(n8043) );
  MUX2_X1 U5755 ( .A(\REGISTERS[53][0] ), .B(n1803), .S(n1535), .Z(n8044) );
  MUX2_X1 U5756 ( .A(\REGISTERS[52][31] ), .B(n2950), .S(n1536), .Z(n7981) );
  MUX2_X1 U5757 ( .A(\REGISTERS[52][30] ), .B(n2939), .S(n1536), .Z(n7982) );
  MUX2_X1 U5758 ( .A(\REGISTERS[52][29] ), .B(n2928), .S(n1536), .Z(n7983) );
  MUX2_X1 U5759 ( .A(\REGISTERS[52][28] ), .B(n2912), .S(n1536), .Z(n7984) );
  MUX2_X1 U5760 ( .A(\REGISTERS[52][27] ), .B(n2901), .S(n1536), .Z(n7985) );
  MUX2_X1 U5761 ( .A(\REGISTERS[52][26] ), .B(n2889), .S(n1536), .Z(n7986) );
  MUX2_X1 U5762 ( .A(\REGISTERS[52][25] ), .B(n2878), .S(n1536), .Z(n7987) );
  MUX2_X1 U5763 ( .A(\REGISTERS[52][24] ), .B(n2867), .S(n1536), .Z(n7988) );
  MUX2_X1 U5764 ( .A(\REGISTERS[52][23] ), .B(n2856), .S(n1536), .Z(n7989) );
  MUX2_X1 U5765 ( .A(\REGISTERS[52][22] ), .B(n2845), .S(n1536), .Z(n7990) );
  MUX2_X1 U5766 ( .A(\REGISTERS[52][21] ), .B(n2834), .S(n1536), .Z(n7991) );
  MUX2_X1 U5767 ( .A(\REGISTERS[52][20] ), .B(n2823), .S(n1536), .Z(n7992) );
  MUX2_X1 U5768 ( .A(\REGISTERS[52][19] ), .B(n2812), .S(n1537), .Z(n7993) );
  MUX2_X1 U5769 ( .A(\REGISTERS[52][18] ), .B(n2801), .S(n1537), .Z(n7994) );
  MUX2_X1 U5770 ( .A(\REGISTERS[52][17] ), .B(n2790), .S(n1537), .Z(n7995) );
  MUX2_X1 U5771 ( .A(\REGISTERS[52][16] ), .B(n2779), .S(n1537), .Z(n7996) );
  MUX2_X1 U5772 ( .A(\REGISTERS[52][15] ), .B(n2768), .S(n1537), .Z(n7997) );
  MUX2_X1 U5773 ( .A(\REGISTERS[52][14] ), .B(n2757), .S(n1537), .Z(n7998) );
  MUX2_X1 U5774 ( .A(\REGISTERS[52][13] ), .B(n2746), .S(n1537), .Z(n7999) );
  MUX2_X1 U5775 ( .A(\REGISTERS[52][12] ), .B(n2735), .S(n1537), .Z(n8000) );
  MUX2_X1 U5776 ( .A(\REGISTERS[52][11] ), .B(n2724), .S(n1537), .Z(n8001) );
  MUX2_X1 U5777 ( .A(\REGISTERS[52][10] ), .B(n2713), .S(n1537), .Z(n8002) );
  MUX2_X1 U5778 ( .A(\REGISTERS[52][9] ), .B(n2606), .S(n1537), .Z(n8003) );
  MUX2_X1 U5779 ( .A(\REGISTERS[52][8] ), .B(n2595), .S(n1537), .Z(n8004) );
  MUX2_X1 U5780 ( .A(\REGISTERS[52][7] ), .B(n2584), .S(n1538), .Z(n8005) );
  MUX2_X1 U5781 ( .A(\REGISTERS[52][6] ), .B(n2573), .S(n1538), .Z(n8006) );
  MUX2_X1 U5782 ( .A(\REGISTERS[52][5] ), .B(n2562), .S(n1538), .Z(n8007) );
  MUX2_X1 U5783 ( .A(\REGISTERS[52][4] ), .B(n2551), .S(n1538), .Z(n8008) );
  MUX2_X1 U5784 ( .A(\REGISTERS[52][3] ), .B(n1836), .S(n1538), .Z(n8009) );
  MUX2_X1 U5785 ( .A(\REGISTERS[52][2] ), .B(n1825), .S(n1538), .Z(n8010) );
  MUX2_X1 U5786 ( .A(\REGISTERS[52][1] ), .B(n1814), .S(n1538), .Z(n8011) );
  MUX2_X1 U5787 ( .A(\REGISTERS[52][0] ), .B(n1803), .S(n1538), .Z(n8012) );
  MUX2_X1 U5788 ( .A(\REGISTERS[51][31] ), .B(n2950), .S(n1539), .Z(n7949) );
  MUX2_X1 U5789 ( .A(\REGISTERS[51][30] ), .B(n2939), .S(n1539), .Z(n7950) );
  MUX2_X1 U5790 ( .A(\REGISTERS[51][29] ), .B(n2928), .S(n1539), .Z(n7951) );
  MUX2_X1 U5791 ( .A(\REGISTERS[51][28] ), .B(n2912), .S(n1539), .Z(n7952) );
  MUX2_X1 U5792 ( .A(\REGISTERS[51][27] ), .B(n2901), .S(n1539), .Z(n7953) );
  MUX2_X1 U5793 ( .A(\REGISTERS[51][26] ), .B(n2889), .S(n1539), .Z(n7954) );
  MUX2_X1 U5794 ( .A(\REGISTERS[51][25] ), .B(n2878), .S(n1539), .Z(n7955) );
  MUX2_X1 U5795 ( .A(\REGISTERS[51][24] ), .B(n2867), .S(n1539), .Z(n7956) );
  MUX2_X1 U5796 ( .A(\REGISTERS[51][23] ), .B(n2856), .S(n1539), .Z(n7957) );
  MUX2_X1 U5797 ( .A(\REGISTERS[51][22] ), .B(n2845), .S(n1539), .Z(n7958) );
  MUX2_X1 U5798 ( .A(\REGISTERS[51][21] ), .B(n2834), .S(n1539), .Z(n7959) );
  MUX2_X1 U5799 ( .A(\REGISTERS[51][20] ), .B(n2823), .S(n1539), .Z(n7960) );
  MUX2_X1 U5800 ( .A(\REGISTERS[51][19] ), .B(n2812), .S(n1540), .Z(n7961) );
  MUX2_X1 U5801 ( .A(\REGISTERS[51][18] ), .B(n2801), .S(n1540), .Z(n7962) );
  MUX2_X1 U5802 ( .A(\REGISTERS[51][17] ), .B(n2790), .S(n1540), .Z(n7963) );
  MUX2_X1 U5803 ( .A(\REGISTERS[51][16] ), .B(n2779), .S(n1540), .Z(n7964) );
  MUX2_X1 U5804 ( .A(\REGISTERS[51][15] ), .B(n2768), .S(n1540), .Z(n7965) );
  MUX2_X1 U5805 ( .A(\REGISTERS[51][14] ), .B(n2757), .S(n1540), .Z(n7966) );
  MUX2_X1 U5806 ( .A(\REGISTERS[51][13] ), .B(n2746), .S(n1540), .Z(n7967) );
  MUX2_X1 U5807 ( .A(\REGISTERS[51][12] ), .B(n2735), .S(n1540), .Z(n7968) );
  MUX2_X1 U5808 ( .A(\REGISTERS[51][11] ), .B(n2724), .S(n1540), .Z(n7969) );
  MUX2_X1 U5809 ( .A(\REGISTERS[51][10] ), .B(n2713), .S(n1540), .Z(n7970) );
  MUX2_X1 U5810 ( .A(\REGISTERS[51][9] ), .B(n2606), .S(n1540), .Z(n7971) );
  MUX2_X1 U5811 ( .A(\REGISTERS[51][8] ), .B(n2595), .S(n1540), .Z(n7972) );
  MUX2_X1 U5812 ( .A(\REGISTERS[51][7] ), .B(n2584), .S(n1541), .Z(n7973) );
  MUX2_X1 U5813 ( .A(\REGISTERS[51][6] ), .B(n2573), .S(n1541), .Z(n7974) );
  MUX2_X1 U5814 ( .A(\REGISTERS[51][5] ), .B(n2562), .S(n1541), .Z(n7975) );
  MUX2_X1 U5815 ( .A(\REGISTERS[51][4] ), .B(n2551), .S(n1541), .Z(n7976) );
  MUX2_X1 U5816 ( .A(\REGISTERS[51][3] ), .B(n1836), .S(n1541), .Z(n7977) );
  MUX2_X1 U5817 ( .A(\REGISTERS[51][2] ), .B(n1825), .S(n1541), .Z(n7978) );
  MUX2_X1 U5818 ( .A(\REGISTERS[51][1] ), .B(n1814), .S(n1541), .Z(n7979) );
  MUX2_X1 U5819 ( .A(\REGISTERS[51][0] ), .B(n1803), .S(n1541), .Z(n7980) );
  MUX2_X1 U5820 ( .A(\REGISTERS[50][31] ), .B(n2950), .S(n1542), .Z(n7917) );
  MUX2_X1 U5821 ( .A(\REGISTERS[50][30] ), .B(n2939), .S(n1542), .Z(n7918) );
  MUX2_X1 U5822 ( .A(\REGISTERS[50][29] ), .B(n2928), .S(n1542), .Z(n7919) );
  MUX2_X1 U5823 ( .A(\REGISTERS[50][28] ), .B(n2912), .S(n1542), .Z(n7920) );
  MUX2_X1 U5824 ( .A(\REGISTERS[50][27] ), .B(n2901), .S(n1542), .Z(n7921) );
  MUX2_X1 U5825 ( .A(\REGISTERS[50][26] ), .B(n2889), .S(n1542), .Z(n7922) );
  MUX2_X1 U5826 ( .A(\REGISTERS[50][25] ), .B(n2878), .S(n1542), .Z(n7923) );
  MUX2_X1 U5827 ( .A(\REGISTERS[50][24] ), .B(n2867), .S(n1542), .Z(n7924) );
  MUX2_X1 U5828 ( .A(\REGISTERS[50][23] ), .B(n2856), .S(n1542), .Z(n7925) );
  MUX2_X1 U5829 ( .A(\REGISTERS[50][22] ), .B(n2845), .S(n1542), .Z(n7926) );
  MUX2_X1 U5830 ( .A(\REGISTERS[50][21] ), .B(n2834), .S(n1542), .Z(n7927) );
  MUX2_X1 U5831 ( .A(\REGISTERS[50][20] ), .B(n2823), .S(n1542), .Z(n7928) );
  MUX2_X1 U5832 ( .A(\REGISTERS[50][19] ), .B(n2812), .S(n1543), .Z(n7929) );
  MUX2_X1 U5833 ( .A(\REGISTERS[50][18] ), .B(n2801), .S(n1543), .Z(n7930) );
  MUX2_X1 U5834 ( .A(\REGISTERS[50][17] ), .B(n2790), .S(n1543), .Z(n7931) );
  MUX2_X1 U5835 ( .A(\REGISTERS[50][16] ), .B(n2779), .S(n1543), .Z(n7932) );
  MUX2_X1 U5836 ( .A(\REGISTERS[50][15] ), .B(n2768), .S(n1543), .Z(n7933) );
  MUX2_X1 U5837 ( .A(\REGISTERS[50][14] ), .B(n2757), .S(n1543), .Z(n7934) );
  MUX2_X1 U5838 ( .A(\REGISTERS[50][13] ), .B(n2746), .S(n1543), .Z(n7935) );
  MUX2_X1 U5839 ( .A(\REGISTERS[50][12] ), .B(n2735), .S(n1543), .Z(n7936) );
  MUX2_X1 U5840 ( .A(\REGISTERS[50][11] ), .B(n2724), .S(n1543), .Z(n7937) );
  MUX2_X1 U5841 ( .A(\REGISTERS[50][10] ), .B(n2713), .S(n1543), .Z(n7938) );
  MUX2_X1 U5842 ( .A(\REGISTERS[50][9] ), .B(n2606), .S(n1543), .Z(n7939) );
  MUX2_X1 U5843 ( .A(\REGISTERS[50][8] ), .B(n2595), .S(n1543), .Z(n7940) );
  MUX2_X1 U5844 ( .A(\REGISTERS[50][7] ), .B(n2584), .S(n1544), .Z(n7941) );
  MUX2_X1 U5845 ( .A(\REGISTERS[50][6] ), .B(n2573), .S(n1544), .Z(n7942) );
  MUX2_X1 U5846 ( .A(\REGISTERS[50][5] ), .B(n2562), .S(n1544), .Z(n7943) );
  MUX2_X1 U5847 ( .A(\REGISTERS[50][4] ), .B(n2551), .S(n1544), .Z(n7944) );
  MUX2_X1 U5848 ( .A(\REGISTERS[50][3] ), .B(n1836), .S(n1544), .Z(n7945) );
  MUX2_X1 U5849 ( .A(\REGISTERS[50][2] ), .B(n1825), .S(n1544), .Z(n7946) );
  MUX2_X1 U5850 ( .A(\REGISTERS[50][1] ), .B(n1814), .S(n1544), .Z(n7947) );
  MUX2_X1 U5851 ( .A(\REGISTERS[50][0] ), .B(n1803), .S(n1544), .Z(n7948) );
  MUX2_X1 U5852 ( .A(\REGISTERS[49][31] ), .B(n2950), .S(n1545), .Z(n7885) );
  MUX2_X1 U5853 ( .A(\REGISTERS[49][30] ), .B(n2939), .S(n1545), .Z(n7886) );
  MUX2_X1 U5854 ( .A(\REGISTERS[49][29] ), .B(n2928), .S(n1545), .Z(n7887) );
  MUX2_X1 U5855 ( .A(\REGISTERS[49][28] ), .B(n2912), .S(n1545), .Z(n7888) );
  MUX2_X1 U5856 ( .A(\REGISTERS[49][27] ), .B(n2901), .S(n1545), .Z(n7889) );
  MUX2_X1 U5857 ( .A(\REGISTERS[49][26] ), .B(n2889), .S(n1545), .Z(n7890) );
  MUX2_X1 U5858 ( .A(\REGISTERS[49][25] ), .B(n2878), .S(n1545), .Z(n7891) );
  MUX2_X1 U5859 ( .A(\REGISTERS[49][24] ), .B(n2867), .S(n1545), .Z(n7892) );
  MUX2_X1 U5860 ( .A(\REGISTERS[49][23] ), .B(n2856), .S(n1545), .Z(n7893) );
  MUX2_X1 U5861 ( .A(\REGISTERS[49][22] ), .B(n2845), .S(n1545), .Z(n7894) );
  MUX2_X1 U5862 ( .A(\REGISTERS[49][21] ), .B(n2834), .S(n1545), .Z(n7895) );
  MUX2_X1 U5863 ( .A(\REGISTERS[49][20] ), .B(n2823), .S(n1545), .Z(n7896) );
  MUX2_X1 U5864 ( .A(\REGISTERS[49][19] ), .B(n2812), .S(n1546), .Z(n7897) );
  MUX2_X1 U5865 ( .A(\REGISTERS[49][18] ), .B(n2801), .S(n1546), .Z(n7898) );
  MUX2_X1 U5866 ( .A(\REGISTERS[49][17] ), .B(n2790), .S(n1546), .Z(n7899) );
  MUX2_X1 U5867 ( .A(\REGISTERS[49][16] ), .B(n2779), .S(n1546), .Z(n7900) );
  MUX2_X1 U5868 ( .A(\REGISTERS[49][15] ), .B(n2768), .S(n1546), .Z(n7901) );
  MUX2_X1 U5869 ( .A(\REGISTERS[49][14] ), .B(n2757), .S(n1546), .Z(n7902) );
  MUX2_X1 U5870 ( .A(\REGISTERS[49][13] ), .B(n2746), .S(n1546), .Z(n7903) );
  MUX2_X1 U5871 ( .A(\REGISTERS[49][12] ), .B(n2735), .S(n1546), .Z(n7904) );
  MUX2_X1 U5872 ( .A(\REGISTERS[49][11] ), .B(n2724), .S(n1546), .Z(n7905) );
  MUX2_X1 U5873 ( .A(\REGISTERS[49][10] ), .B(n2713), .S(n1546), .Z(n7906) );
  MUX2_X1 U5874 ( .A(\REGISTERS[49][9] ), .B(n2606), .S(n1546), .Z(n7907) );
  MUX2_X1 U5875 ( .A(\REGISTERS[49][8] ), .B(n2595), .S(n1546), .Z(n7908) );
  MUX2_X1 U5876 ( .A(\REGISTERS[49][7] ), .B(n2584), .S(n1547), .Z(n7909) );
  MUX2_X1 U5877 ( .A(\REGISTERS[49][6] ), .B(n2573), .S(n1547), .Z(n7910) );
  MUX2_X1 U5878 ( .A(\REGISTERS[49][5] ), .B(n2562), .S(n1547), .Z(n7911) );
  MUX2_X1 U5879 ( .A(\REGISTERS[49][4] ), .B(n2551), .S(n1547), .Z(n7912) );
  MUX2_X1 U5880 ( .A(\REGISTERS[49][3] ), .B(n1836), .S(n1547), .Z(n7913) );
  MUX2_X1 U5881 ( .A(\REGISTERS[49][2] ), .B(n1825), .S(n1547), .Z(n7914) );
  MUX2_X1 U5882 ( .A(\REGISTERS[49][1] ), .B(n1814), .S(n1547), .Z(n7915) );
  MUX2_X1 U5883 ( .A(\REGISTERS[49][0] ), .B(n1803), .S(n1547), .Z(n7916) );
  MUX2_X1 U5884 ( .A(n10086), .B(n2950), .S(n1548), .Z(n7853) );
  MUX2_X1 U5885 ( .A(n10087), .B(n2939), .S(n1548), .Z(n7854) );
  MUX2_X1 U5886 ( .A(n10088), .B(n2928), .S(n1548), .Z(n7855) );
  MUX2_X1 U5887 ( .A(n10089), .B(n2912), .S(n1548), .Z(n7856) );
  MUX2_X1 U5888 ( .A(n10090), .B(n2901), .S(n1548), .Z(n7857) );
  MUX2_X1 U5889 ( .A(n10091), .B(n2889), .S(n1548), .Z(n7858) );
  MUX2_X1 U5890 ( .A(n10092), .B(n2878), .S(n1548), .Z(n7859) );
  MUX2_X1 U5891 ( .A(n10093), .B(n2867), .S(n1548), .Z(n7860) );
  MUX2_X1 U5892 ( .A(n10094), .B(n2856), .S(n1548), .Z(n7861) );
  MUX2_X1 U5893 ( .A(n10095), .B(n2845), .S(n1548), .Z(n7862) );
  MUX2_X1 U5894 ( .A(n10096), .B(n2834), .S(n1548), .Z(n7863) );
  MUX2_X1 U5895 ( .A(n10097), .B(n2823), .S(n1548), .Z(n7864) );
  MUX2_X1 U5896 ( .A(n10098), .B(n2812), .S(n1549), .Z(n7865) );
  MUX2_X1 U5897 ( .A(n10099), .B(n2801), .S(n1549), .Z(n7866) );
  MUX2_X1 U5898 ( .A(n10100), .B(n2790), .S(n1549), .Z(n7867) );
  MUX2_X1 U5899 ( .A(n10101), .B(n2779), .S(n1549), .Z(n7868) );
  MUX2_X1 U5900 ( .A(n10102), .B(n2768), .S(n1549), .Z(n7869) );
  MUX2_X1 U5901 ( .A(n10103), .B(n2757), .S(n1549), .Z(n7870) );
  MUX2_X1 U5902 ( .A(n10104), .B(n2746), .S(n1549), .Z(n7871) );
  MUX2_X1 U5903 ( .A(n10105), .B(n2735), .S(n1549), .Z(n7872) );
  MUX2_X1 U5904 ( .A(n10106), .B(n2724), .S(n1549), .Z(n7873) );
  MUX2_X1 U5905 ( .A(n10107), .B(n2713), .S(n1549), .Z(n7874) );
  MUX2_X1 U5906 ( .A(n10108), .B(n2606), .S(n1549), .Z(n7875) );
  MUX2_X1 U5907 ( .A(n10109), .B(n2595), .S(n1549), .Z(n7876) );
  MUX2_X1 U5908 ( .A(n10110), .B(n2584), .S(n1550), .Z(n7877) );
  MUX2_X1 U5909 ( .A(n10111), .B(n2573), .S(n1550), .Z(n7878) );
  MUX2_X1 U5910 ( .A(n10112), .B(n2562), .S(n1550), .Z(n7879) );
  MUX2_X1 U5911 ( .A(n10113), .B(n2551), .S(n1550), .Z(n7880) );
  MUX2_X1 U5912 ( .A(n10114), .B(n1836), .S(n1550), .Z(n7881) );
  MUX2_X1 U5913 ( .A(n10115), .B(n1825), .S(n1550), .Z(n7882) );
  MUX2_X1 U5914 ( .A(n10116), .B(n1814), .S(n1550), .Z(n7883) );
  MUX2_X1 U5915 ( .A(n10117), .B(n1803), .S(n1550), .Z(n7884) );
  MUX2_X1 U5916 ( .A(n10054), .B(n2950), .S(n1551), .Z(n7821) );
  MUX2_X1 U5917 ( .A(n10055), .B(n2939), .S(n1551), .Z(n7822) );
  MUX2_X1 U5918 ( .A(n10056), .B(n2928), .S(n1551), .Z(n7823) );
  MUX2_X1 U5919 ( .A(n10057), .B(n2912), .S(n1551), .Z(n7824) );
  MUX2_X1 U5920 ( .A(n10058), .B(n2901), .S(n1551), .Z(n7825) );
  MUX2_X1 U5921 ( .A(n10059), .B(n2889), .S(n1551), .Z(n7826) );
  MUX2_X1 U5922 ( .A(n10060), .B(n2878), .S(n1551), .Z(n7827) );
  MUX2_X1 U5923 ( .A(n10061), .B(n2867), .S(n1551), .Z(n7828) );
  MUX2_X1 U5924 ( .A(n10062), .B(n2856), .S(n1551), .Z(n7829) );
  MUX2_X1 U5925 ( .A(n10063), .B(n2845), .S(n1551), .Z(n7830) );
  MUX2_X1 U5926 ( .A(n10064), .B(n2834), .S(n1551), .Z(n7831) );
  MUX2_X1 U5927 ( .A(n10065), .B(n2823), .S(n1551), .Z(n7832) );
  MUX2_X1 U5928 ( .A(n10066), .B(n2812), .S(n1648), .Z(n7833) );
  MUX2_X1 U5929 ( .A(n10067), .B(n2801), .S(n1648), .Z(n7834) );
  MUX2_X1 U5930 ( .A(n10068), .B(n2790), .S(n1648), .Z(n7835) );
  MUX2_X1 U5931 ( .A(n10069), .B(n2779), .S(n1648), .Z(n7836) );
  MUX2_X1 U5932 ( .A(n10070), .B(n2768), .S(n1648), .Z(n7837) );
  MUX2_X1 U5933 ( .A(n10071), .B(n2757), .S(n1648), .Z(n7838) );
  MUX2_X1 U5934 ( .A(n10072), .B(n2746), .S(n1648), .Z(n7839) );
  MUX2_X1 U5935 ( .A(n10073), .B(n2735), .S(n1648), .Z(n7840) );
  MUX2_X1 U5936 ( .A(n10074), .B(n2724), .S(n1648), .Z(n7841) );
  MUX2_X1 U5937 ( .A(n10075), .B(n2713), .S(n1648), .Z(n7842) );
  MUX2_X1 U5938 ( .A(n10076), .B(n2606), .S(n1648), .Z(n7843) );
  MUX2_X1 U5939 ( .A(n10077), .B(n2595), .S(n1648), .Z(n7844) );
  MUX2_X1 U5940 ( .A(n10078), .B(n2584), .S(n1649), .Z(n7845) );
  MUX2_X1 U5941 ( .A(n10079), .B(n2573), .S(n1649), .Z(n7846) );
  MUX2_X1 U5942 ( .A(n10080), .B(n2562), .S(n1649), .Z(n7847) );
  MUX2_X1 U5943 ( .A(n10081), .B(n2551), .S(n1649), .Z(n7848) );
  MUX2_X1 U5944 ( .A(n10082), .B(n1836), .S(n1649), .Z(n7849) );
  MUX2_X1 U5945 ( .A(n10083), .B(n1825), .S(n1649), .Z(n7850) );
  MUX2_X1 U5946 ( .A(n10084), .B(n1814), .S(n1649), .Z(n7851) );
  MUX2_X1 U5947 ( .A(n10085), .B(n1803), .S(n1649), .Z(n7852) );
  MUX2_X1 U5948 ( .A(n10022), .B(n2950), .S(n1650), .Z(n7789) );
  MUX2_X1 U5949 ( .A(n10023), .B(n2939), .S(n1650), .Z(n7790) );
  MUX2_X1 U5950 ( .A(n10024), .B(n2928), .S(n1650), .Z(n7791) );
  MUX2_X1 U5951 ( .A(n10025), .B(n2912), .S(n1650), .Z(n7792) );
  MUX2_X1 U5952 ( .A(n10026), .B(n2901), .S(n1650), .Z(n7793) );
  MUX2_X1 U5953 ( .A(n10027), .B(n2889), .S(n1650), .Z(n7794) );
  MUX2_X1 U5954 ( .A(n10028), .B(n2878), .S(n1650), .Z(n7795) );
  MUX2_X1 U5955 ( .A(n10029), .B(n2867), .S(n1650), .Z(n7796) );
  MUX2_X1 U5956 ( .A(n10030), .B(n2856), .S(n1650), .Z(n7797) );
  MUX2_X1 U5957 ( .A(n10031), .B(n2845), .S(n1650), .Z(n7798) );
  MUX2_X1 U5958 ( .A(n10032), .B(n2834), .S(n1650), .Z(n7799) );
  MUX2_X1 U5959 ( .A(n10033), .B(n2823), .S(n1650), .Z(n7800) );
  MUX2_X1 U5960 ( .A(n10034), .B(n2812), .S(n1651), .Z(n7801) );
  MUX2_X1 U5961 ( .A(n10035), .B(n2801), .S(n1651), .Z(n7802) );
  MUX2_X1 U5962 ( .A(n10036), .B(n2790), .S(n1651), .Z(n7803) );
  MUX2_X1 U5963 ( .A(n10037), .B(n2779), .S(n1651), .Z(n7804) );
  MUX2_X1 U5964 ( .A(n10038), .B(n2768), .S(n1651), .Z(n7805) );
  MUX2_X1 U5965 ( .A(n10039), .B(n2757), .S(n1651), .Z(n7806) );
  MUX2_X1 U5966 ( .A(n10040), .B(n2746), .S(n1651), .Z(n7807) );
  MUX2_X1 U5967 ( .A(n10041), .B(n2735), .S(n1651), .Z(n7808) );
  MUX2_X1 U5968 ( .A(n10042), .B(n2724), .S(n1651), .Z(n7809) );
  MUX2_X1 U5969 ( .A(n10043), .B(n2713), .S(n1651), .Z(n7810) );
  MUX2_X1 U5970 ( .A(n10044), .B(n2606), .S(n1651), .Z(n7811) );
  MUX2_X1 U5971 ( .A(n10045), .B(n2595), .S(n1651), .Z(n7812) );
  MUX2_X1 U5972 ( .A(n10046), .B(n2584), .S(n1652), .Z(n7813) );
  MUX2_X1 U5973 ( .A(n10047), .B(n2573), .S(n1652), .Z(n7814) );
  MUX2_X1 U5974 ( .A(n10048), .B(n2562), .S(n1652), .Z(n7815) );
  MUX2_X1 U5975 ( .A(n10049), .B(n2551), .S(n1652), .Z(n7816) );
  MUX2_X1 U5976 ( .A(n10050), .B(n1836), .S(n1652), .Z(n7817) );
  MUX2_X1 U5977 ( .A(n10051), .B(n1825), .S(n1652), .Z(n7818) );
  MUX2_X1 U5978 ( .A(n10052), .B(n1814), .S(n1652), .Z(n7819) );
  MUX2_X1 U5979 ( .A(n10053), .B(n1803), .S(n1652), .Z(n7820) );
  MUX2_X1 U5980 ( .A(\REGISTERS[45][31] ), .B(n2950), .S(n1653), .Z(n7757) );
  MUX2_X1 U5981 ( .A(\REGISTERS[45][30] ), .B(n2939), .S(n1653), .Z(n7758) );
  MUX2_X1 U5982 ( .A(\REGISTERS[45][29] ), .B(n2928), .S(n1653), .Z(n7759) );
  MUX2_X1 U5983 ( .A(\REGISTERS[45][28] ), .B(n2912), .S(n1653), .Z(n7760) );
  MUX2_X1 U5984 ( .A(\REGISTERS[45][27] ), .B(n2901), .S(n1653), .Z(n7761) );
  MUX2_X1 U5985 ( .A(\REGISTERS[45][26] ), .B(n2889), .S(n1653), .Z(n7762) );
  MUX2_X1 U5986 ( .A(\REGISTERS[45][25] ), .B(n2878), .S(n1653), .Z(n7763) );
  MUX2_X1 U5987 ( .A(\REGISTERS[45][24] ), .B(n2867), .S(n1653), .Z(n7764) );
  MUX2_X1 U5988 ( .A(\REGISTERS[45][23] ), .B(n2856), .S(n1653), .Z(n7765) );
  MUX2_X1 U5989 ( .A(\REGISTERS[45][22] ), .B(n2845), .S(n1653), .Z(n7766) );
  MUX2_X1 U5990 ( .A(\REGISTERS[45][21] ), .B(n2834), .S(n1653), .Z(n7767) );
  MUX2_X1 U5991 ( .A(\REGISTERS[45][20] ), .B(n2823), .S(n1653), .Z(n7768) );
  MUX2_X1 U5992 ( .A(\REGISTERS[45][19] ), .B(n2812), .S(n1654), .Z(n7769) );
  MUX2_X1 U5993 ( .A(\REGISTERS[45][18] ), .B(n2801), .S(n1654), .Z(n7770) );
  MUX2_X1 U5994 ( .A(\REGISTERS[45][17] ), .B(n2790), .S(n1654), .Z(n7771) );
  MUX2_X1 U5995 ( .A(\REGISTERS[45][16] ), .B(n2779), .S(n1654), .Z(n7772) );
  MUX2_X1 U5996 ( .A(\REGISTERS[45][15] ), .B(n2768), .S(n1654), .Z(n7773) );
  MUX2_X1 U5997 ( .A(\REGISTERS[45][14] ), .B(n2757), .S(n1654), .Z(n7774) );
  MUX2_X1 U5998 ( .A(\REGISTERS[45][13] ), .B(n2746), .S(n1654), .Z(n7775) );
  MUX2_X1 U5999 ( .A(\REGISTERS[45][12] ), .B(n2735), .S(n1654), .Z(n7776) );
  MUX2_X1 U6000 ( .A(\REGISTERS[45][11] ), .B(n2724), .S(n1654), .Z(n7777) );
  MUX2_X1 U6001 ( .A(\REGISTERS[45][10] ), .B(n2713), .S(n1654), .Z(n7778) );
  MUX2_X1 U6002 ( .A(\REGISTERS[45][9] ), .B(n2606), .S(n1654), .Z(n7779) );
  MUX2_X1 U6003 ( .A(\REGISTERS[45][8] ), .B(n2595), .S(n1654), .Z(n7780) );
  MUX2_X1 U6004 ( .A(\REGISTERS[45][7] ), .B(n2584), .S(n1655), .Z(n7781) );
  MUX2_X1 U6005 ( .A(\REGISTERS[45][6] ), .B(n2573), .S(n1655), .Z(n7782) );
  MUX2_X1 U6006 ( .A(\REGISTERS[45][5] ), .B(n2562), .S(n1655), .Z(n7783) );
  MUX2_X1 U6007 ( .A(\REGISTERS[45][4] ), .B(n2551), .S(n1655), .Z(n7784) );
  MUX2_X1 U6008 ( .A(\REGISTERS[45][3] ), .B(n1836), .S(n1655), .Z(n7785) );
  MUX2_X1 U6009 ( .A(\REGISTERS[45][2] ), .B(n1825), .S(n1655), .Z(n7786) );
  MUX2_X1 U6010 ( .A(\REGISTERS[45][1] ), .B(n1814), .S(n1655), .Z(n7787) );
  MUX2_X1 U6011 ( .A(\REGISTERS[45][0] ), .B(n1803), .S(n1655), .Z(n7788) );
  MUX2_X1 U6012 ( .A(\REGISTERS[44][31] ), .B(n2950), .S(n1656), .Z(n7725) );
  MUX2_X1 U6013 ( .A(\REGISTERS[44][30] ), .B(n2939), .S(n1656), .Z(n7726) );
  MUX2_X1 U6014 ( .A(\REGISTERS[44][29] ), .B(n2928), .S(n1656), .Z(n7727) );
  MUX2_X1 U6015 ( .A(\REGISTERS[44][28] ), .B(n2912), .S(n1656), .Z(n7728) );
  MUX2_X1 U6016 ( .A(\REGISTERS[44][27] ), .B(n2901), .S(n1656), .Z(n7729) );
  MUX2_X1 U6017 ( .A(\REGISTERS[44][26] ), .B(n2889), .S(n1656), .Z(n7730) );
  MUX2_X1 U6018 ( .A(\REGISTERS[44][25] ), .B(n2878), .S(n1656), .Z(n7731) );
  MUX2_X1 U6019 ( .A(\REGISTERS[44][24] ), .B(n2867), .S(n1656), .Z(n7732) );
  MUX2_X1 U6020 ( .A(\REGISTERS[44][23] ), .B(n2856), .S(n1656), .Z(n7733) );
  MUX2_X1 U6021 ( .A(\REGISTERS[44][22] ), .B(n2845), .S(n1656), .Z(n7734) );
  MUX2_X1 U6022 ( .A(\REGISTERS[44][21] ), .B(n2834), .S(n1656), .Z(n7735) );
  MUX2_X1 U6023 ( .A(\REGISTERS[44][20] ), .B(n2823), .S(n1656), .Z(n7736) );
  MUX2_X1 U6024 ( .A(\REGISTERS[44][19] ), .B(n2812), .S(n1657), .Z(n7737) );
  MUX2_X1 U6025 ( .A(\REGISTERS[44][18] ), .B(n2801), .S(n1657), .Z(n7738) );
  MUX2_X1 U6026 ( .A(\REGISTERS[44][17] ), .B(n2790), .S(n1657), .Z(n7739) );
  MUX2_X1 U6027 ( .A(\REGISTERS[44][16] ), .B(n2779), .S(n1657), .Z(n7740) );
  MUX2_X1 U6028 ( .A(\REGISTERS[44][15] ), .B(n2768), .S(n1657), .Z(n7741) );
  MUX2_X1 U6029 ( .A(\REGISTERS[44][14] ), .B(n2757), .S(n1657), .Z(n7742) );
  MUX2_X1 U6030 ( .A(\REGISTERS[44][13] ), .B(n2746), .S(n1657), .Z(n7743) );
  MUX2_X1 U6031 ( .A(\REGISTERS[44][12] ), .B(n2735), .S(n1657), .Z(n7744) );
  MUX2_X1 U6032 ( .A(\REGISTERS[44][11] ), .B(n2724), .S(n1657), .Z(n7745) );
  MUX2_X1 U6033 ( .A(\REGISTERS[44][10] ), .B(n2713), .S(n1657), .Z(n7746) );
  MUX2_X1 U6034 ( .A(\REGISTERS[44][9] ), .B(n2606), .S(n1657), .Z(n7747) );
  MUX2_X1 U6035 ( .A(\REGISTERS[44][8] ), .B(n2595), .S(n1657), .Z(n7748) );
  MUX2_X1 U6036 ( .A(\REGISTERS[44][7] ), .B(n2584), .S(n1658), .Z(n7749) );
  MUX2_X1 U6037 ( .A(\REGISTERS[44][6] ), .B(n2573), .S(n1658), .Z(n7750) );
  MUX2_X1 U6038 ( .A(\REGISTERS[44][5] ), .B(n2562), .S(n1658), .Z(n7751) );
  MUX2_X1 U6039 ( .A(\REGISTERS[44][4] ), .B(n2551), .S(n1658), .Z(n7752) );
  MUX2_X1 U6040 ( .A(\REGISTERS[44][3] ), .B(n1836), .S(n1658), .Z(n7753) );
  MUX2_X1 U6041 ( .A(\REGISTERS[44][2] ), .B(n1825), .S(n1658), .Z(n7754) );
  MUX2_X1 U6042 ( .A(\REGISTERS[44][1] ), .B(n1814), .S(n1658), .Z(n7755) );
  MUX2_X1 U6043 ( .A(\REGISTERS[44][0] ), .B(n1803), .S(n1658), .Z(n7756) );
  MUX2_X1 U6044 ( .A(\REGISTERS[43][31] ), .B(n2951), .S(n1659), .Z(n7693) );
  MUX2_X1 U6045 ( .A(\REGISTERS[43][30] ), .B(n2940), .S(n1659), .Z(n7694) );
  MUX2_X1 U6046 ( .A(\REGISTERS[43][29] ), .B(n2929), .S(n1659), .Z(n7695) );
  MUX2_X1 U6047 ( .A(\REGISTERS[43][28] ), .B(n2913), .S(n1659), .Z(n7696) );
  MUX2_X1 U6048 ( .A(\REGISTERS[43][27] ), .B(n2902), .S(n1659), .Z(n7697) );
  MUX2_X1 U6049 ( .A(\REGISTERS[43][26] ), .B(n2890), .S(n1659), .Z(n7698) );
  MUX2_X1 U6050 ( .A(\REGISTERS[43][25] ), .B(n2879), .S(n1659), .Z(n7699) );
  MUX2_X1 U6051 ( .A(\REGISTERS[43][24] ), .B(n2868), .S(n1659), .Z(n7700) );
  MUX2_X1 U6052 ( .A(\REGISTERS[43][23] ), .B(n2857), .S(n1659), .Z(n7701) );
  MUX2_X1 U6053 ( .A(\REGISTERS[43][22] ), .B(n2846), .S(n1659), .Z(n7702) );
  MUX2_X1 U6054 ( .A(\REGISTERS[43][21] ), .B(n2835), .S(n1659), .Z(n7703) );
  MUX2_X1 U6055 ( .A(\REGISTERS[43][20] ), .B(n2824), .S(n1659), .Z(n7704) );
  MUX2_X1 U6056 ( .A(\REGISTERS[43][19] ), .B(n2813), .S(n1660), .Z(n7705) );
  MUX2_X1 U6057 ( .A(\REGISTERS[43][18] ), .B(n2802), .S(n1660), .Z(n7706) );
  MUX2_X1 U6058 ( .A(\REGISTERS[43][17] ), .B(n2791), .S(n1660), .Z(n7707) );
  MUX2_X1 U6059 ( .A(\REGISTERS[43][16] ), .B(n2780), .S(n1660), .Z(n7708) );
  MUX2_X1 U6060 ( .A(\REGISTERS[43][15] ), .B(n2769), .S(n1660), .Z(n7709) );
  MUX2_X1 U6061 ( .A(\REGISTERS[43][14] ), .B(n2758), .S(n1660), .Z(n7710) );
  MUX2_X1 U6062 ( .A(\REGISTERS[43][13] ), .B(n2747), .S(n1660), .Z(n7711) );
  MUX2_X1 U6063 ( .A(\REGISTERS[43][12] ), .B(n2736), .S(n1660), .Z(n7712) );
  MUX2_X1 U6064 ( .A(\REGISTERS[43][11] ), .B(n2725), .S(n1660), .Z(n7713) );
  MUX2_X1 U6065 ( .A(\REGISTERS[43][10] ), .B(n2714), .S(n1660), .Z(n7714) );
  MUX2_X1 U6066 ( .A(\REGISTERS[43][9] ), .B(n2607), .S(n1660), .Z(n7715) );
  MUX2_X1 U6067 ( .A(\REGISTERS[43][8] ), .B(n2596), .S(n1660), .Z(n7716) );
  MUX2_X1 U6068 ( .A(\REGISTERS[43][7] ), .B(n2585), .S(n1661), .Z(n7717) );
  MUX2_X1 U6069 ( .A(\REGISTERS[43][6] ), .B(n2574), .S(n1661), .Z(n7718) );
  MUX2_X1 U6070 ( .A(\REGISTERS[43][5] ), .B(n2563), .S(n1661), .Z(n7719) );
  MUX2_X1 U6071 ( .A(\REGISTERS[43][4] ), .B(n2552), .S(n1661), .Z(n7720) );
  MUX2_X1 U6072 ( .A(\REGISTERS[43][3] ), .B(n1837), .S(n1661), .Z(n7721) );
  MUX2_X1 U6073 ( .A(\REGISTERS[43][2] ), .B(n1826), .S(n1661), .Z(n7722) );
  MUX2_X1 U6074 ( .A(\REGISTERS[43][1] ), .B(n1815), .S(n1661), .Z(n7723) );
  MUX2_X1 U6075 ( .A(\REGISTERS[43][0] ), .B(n1804), .S(n1661), .Z(n7724) );
  MUX2_X1 U6076 ( .A(\REGISTERS[42][31] ), .B(n2951), .S(n1662), .Z(n7661) );
  MUX2_X1 U6077 ( .A(\REGISTERS[42][30] ), .B(n2940), .S(n1662), .Z(n7662) );
  MUX2_X1 U6078 ( .A(\REGISTERS[42][29] ), .B(n2929), .S(n1662), .Z(n7663) );
  MUX2_X1 U6079 ( .A(\REGISTERS[42][28] ), .B(n2913), .S(n1662), .Z(n7664) );
  MUX2_X1 U6080 ( .A(\REGISTERS[42][27] ), .B(n2902), .S(n1662), .Z(n7665) );
  MUX2_X1 U6081 ( .A(\REGISTERS[42][26] ), .B(n2890), .S(n1662), .Z(n7666) );
  MUX2_X1 U6082 ( .A(\REGISTERS[42][25] ), .B(n2879), .S(n1662), .Z(n7667) );
  MUX2_X1 U6083 ( .A(\REGISTERS[42][24] ), .B(n2868), .S(n1662), .Z(n7668) );
  MUX2_X1 U6084 ( .A(\REGISTERS[42][23] ), .B(n2857), .S(n1662), .Z(n7669) );
  MUX2_X1 U6085 ( .A(\REGISTERS[42][22] ), .B(n2846), .S(n1662), .Z(n7670) );
  MUX2_X1 U6086 ( .A(\REGISTERS[42][21] ), .B(n2835), .S(n1662), .Z(n7671) );
  MUX2_X1 U6087 ( .A(\REGISTERS[42][20] ), .B(n2824), .S(n1662), .Z(n7672) );
  MUX2_X1 U6088 ( .A(\REGISTERS[42][19] ), .B(n2813), .S(n1663), .Z(n7673) );
  MUX2_X1 U6089 ( .A(\REGISTERS[42][18] ), .B(n2802), .S(n1663), .Z(n7674) );
  MUX2_X1 U6090 ( .A(\REGISTERS[42][17] ), .B(n2791), .S(n1663), .Z(n7675) );
  MUX2_X1 U6091 ( .A(\REGISTERS[42][16] ), .B(n2780), .S(n1663), .Z(n7676) );
  MUX2_X1 U6092 ( .A(\REGISTERS[42][15] ), .B(n2769), .S(n1663), .Z(n7677) );
  MUX2_X1 U6093 ( .A(\REGISTERS[42][14] ), .B(n2758), .S(n1663), .Z(n7678) );
  MUX2_X1 U6094 ( .A(\REGISTERS[42][13] ), .B(n2747), .S(n1663), .Z(n7679) );
  MUX2_X1 U6095 ( .A(\REGISTERS[42][12] ), .B(n2736), .S(n1663), .Z(n7680) );
  MUX2_X1 U6096 ( .A(\REGISTERS[42][11] ), .B(n2725), .S(n1663), .Z(n7681) );
  MUX2_X1 U6097 ( .A(\REGISTERS[42][10] ), .B(n2714), .S(n1663), .Z(n7682) );
  MUX2_X1 U6098 ( .A(\REGISTERS[42][9] ), .B(n2607), .S(n1663), .Z(n7683) );
  MUX2_X1 U6099 ( .A(\REGISTERS[42][8] ), .B(n2596), .S(n1663), .Z(n7684) );
  MUX2_X1 U6100 ( .A(\REGISTERS[42][7] ), .B(n2585), .S(n1664), .Z(n7685) );
  MUX2_X1 U6101 ( .A(\REGISTERS[42][6] ), .B(n2574), .S(n1664), .Z(n7686) );
  MUX2_X1 U6102 ( .A(\REGISTERS[42][5] ), .B(n2563), .S(n1664), .Z(n7687) );
  MUX2_X1 U6103 ( .A(\REGISTERS[42][4] ), .B(n2552), .S(n1664), .Z(n7688) );
  MUX2_X1 U6104 ( .A(\REGISTERS[42][3] ), .B(n1837), .S(n1664), .Z(n7689) );
  MUX2_X1 U6105 ( .A(\REGISTERS[42][2] ), .B(n1826), .S(n1664), .Z(n7690) );
  MUX2_X1 U6106 ( .A(\REGISTERS[42][1] ), .B(n1815), .S(n1664), .Z(n7691) );
  MUX2_X1 U6107 ( .A(\REGISTERS[42][0] ), .B(n1804), .S(n1664), .Z(n7692) );
  MUX2_X1 U6108 ( .A(\REGISTERS[41][31] ), .B(n2951), .S(n1665), .Z(n7629) );
  MUX2_X1 U6109 ( .A(\REGISTERS[41][30] ), .B(n2940), .S(n1665), .Z(n7630) );
  MUX2_X1 U6110 ( .A(\REGISTERS[41][29] ), .B(n2929), .S(n1665), .Z(n7631) );
  MUX2_X1 U6111 ( .A(\REGISTERS[41][28] ), .B(n2913), .S(n1665), .Z(n7632) );
  MUX2_X1 U6112 ( .A(\REGISTERS[41][27] ), .B(n2902), .S(n1665), .Z(n7633) );
  MUX2_X1 U6113 ( .A(\REGISTERS[41][26] ), .B(n2890), .S(n1665), .Z(n7634) );
  MUX2_X1 U6114 ( .A(\REGISTERS[41][25] ), .B(n2879), .S(n1665), .Z(n7635) );
  MUX2_X1 U6115 ( .A(\REGISTERS[41][24] ), .B(n2868), .S(n1665), .Z(n7636) );
  MUX2_X1 U6116 ( .A(\REGISTERS[41][23] ), .B(n2857), .S(n1665), .Z(n7637) );
  MUX2_X1 U6117 ( .A(\REGISTERS[41][22] ), .B(n2846), .S(n1665), .Z(n7638) );
  MUX2_X1 U6118 ( .A(\REGISTERS[41][21] ), .B(n2835), .S(n1665), .Z(n7639) );
  MUX2_X1 U6119 ( .A(\REGISTERS[41][20] ), .B(n2824), .S(n1665), .Z(n7640) );
  MUX2_X1 U6120 ( .A(\REGISTERS[41][19] ), .B(n2813), .S(n1666), .Z(n7641) );
  MUX2_X1 U6121 ( .A(\REGISTERS[41][18] ), .B(n2802), .S(n1666), .Z(n7642) );
  MUX2_X1 U6122 ( .A(\REGISTERS[41][17] ), .B(n2791), .S(n1666), .Z(n7643) );
  MUX2_X1 U6123 ( .A(\REGISTERS[41][16] ), .B(n2780), .S(n1666), .Z(n7644) );
  MUX2_X1 U6124 ( .A(\REGISTERS[41][15] ), .B(n2769), .S(n1666), .Z(n7645) );
  MUX2_X1 U6125 ( .A(\REGISTERS[41][14] ), .B(n2758), .S(n1666), .Z(n7646) );
  MUX2_X1 U6126 ( .A(\REGISTERS[41][13] ), .B(n2747), .S(n1666), .Z(n7647) );
  MUX2_X1 U6127 ( .A(\REGISTERS[41][12] ), .B(n2736), .S(n1666), .Z(n7648) );
  MUX2_X1 U6128 ( .A(\REGISTERS[41][11] ), .B(n2725), .S(n1666), .Z(n7649) );
  MUX2_X1 U6129 ( .A(\REGISTERS[41][10] ), .B(n2714), .S(n1666), .Z(n7650) );
  MUX2_X1 U6130 ( .A(\REGISTERS[41][9] ), .B(n2607), .S(n1666), .Z(n7651) );
  MUX2_X1 U6131 ( .A(\REGISTERS[41][8] ), .B(n2596), .S(n1666), .Z(n7652) );
  MUX2_X1 U6132 ( .A(\REGISTERS[41][7] ), .B(n2585), .S(n1667), .Z(n7653) );
  MUX2_X1 U6133 ( .A(\REGISTERS[41][6] ), .B(n2574), .S(n1667), .Z(n7654) );
  MUX2_X1 U6134 ( .A(\REGISTERS[41][5] ), .B(n2563), .S(n1667), .Z(n7655) );
  MUX2_X1 U6135 ( .A(\REGISTERS[41][4] ), .B(n2552), .S(n1667), .Z(n7656) );
  MUX2_X1 U6136 ( .A(\REGISTERS[41][3] ), .B(n1837), .S(n1667), .Z(n7657) );
  MUX2_X1 U6137 ( .A(\REGISTERS[41][2] ), .B(n1826), .S(n1667), .Z(n7658) );
  MUX2_X1 U6138 ( .A(\REGISTERS[41][1] ), .B(n1815), .S(n1667), .Z(n7659) );
  MUX2_X1 U6139 ( .A(\REGISTERS[41][0] ), .B(n1804), .S(n1667), .Z(n7660) );
  MUX2_X1 U6140 ( .A(\REGISTERS[40][31] ), .B(n2951), .S(n1668), .Z(n7597) );
  MUX2_X1 U6141 ( .A(\REGISTERS[40][30] ), .B(n2940), .S(n1668), .Z(n7598) );
  MUX2_X1 U6142 ( .A(\REGISTERS[40][29] ), .B(n2929), .S(n1668), .Z(n7599) );
  MUX2_X1 U6143 ( .A(\REGISTERS[40][28] ), .B(n2913), .S(n1668), .Z(n7600) );
  MUX2_X1 U6144 ( .A(\REGISTERS[40][27] ), .B(n2902), .S(n1668), .Z(n7601) );
  MUX2_X1 U6145 ( .A(\REGISTERS[40][26] ), .B(n2890), .S(n1668), .Z(n7602) );
  MUX2_X1 U6146 ( .A(\REGISTERS[40][25] ), .B(n2879), .S(n1668), .Z(n7603) );
  MUX2_X1 U6147 ( .A(\REGISTERS[40][24] ), .B(n2868), .S(n1668), .Z(n7604) );
  MUX2_X1 U6148 ( .A(\REGISTERS[40][23] ), .B(n2857), .S(n1668), .Z(n7605) );
  MUX2_X1 U6149 ( .A(\REGISTERS[40][22] ), .B(n2846), .S(n1668), .Z(n7606) );
  MUX2_X1 U6150 ( .A(\REGISTERS[40][21] ), .B(n2835), .S(n1668), .Z(n7607) );
  MUX2_X1 U6151 ( .A(\REGISTERS[40][20] ), .B(n2824), .S(n1668), .Z(n7608) );
  MUX2_X1 U6152 ( .A(\REGISTERS[40][19] ), .B(n2813), .S(n1669), .Z(n7609) );
  MUX2_X1 U6153 ( .A(\REGISTERS[40][18] ), .B(n2802), .S(n1669), .Z(n7610) );
  MUX2_X1 U6154 ( .A(\REGISTERS[40][17] ), .B(n2791), .S(n1669), .Z(n7611) );
  MUX2_X1 U6155 ( .A(\REGISTERS[40][16] ), .B(n2780), .S(n1669), .Z(n7612) );
  MUX2_X1 U6156 ( .A(\REGISTERS[40][15] ), .B(n2769), .S(n1669), .Z(n7613) );
  MUX2_X1 U6157 ( .A(\REGISTERS[40][14] ), .B(n2758), .S(n1669), .Z(n7614) );
  MUX2_X1 U6158 ( .A(\REGISTERS[40][13] ), .B(n2747), .S(n1669), .Z(n7615) );
  MUX2_X1 U6159 ( .A(\REGISTERS[40][12] ), .B(n2736), .S(n1669), .Z(n7616) );
  MUX2_X1 U6160 ( .A(\REGISTERS[40][11] ), .B(n2725), .S(n1669), .Z(n7617) );
  MUX2_X1 U6161 ( .A(\REGISTERS[40][10] ), .B(n2714), .S(n1669), .Z(n7618) );
  MUX2_X1 U6162 ( .A(\REGISTERS[40][9] ), .B(n2607), .S(n1669), .Z(n7619) );
  MUX2_X1 U6163 ( .A(\REGISTERS[40][8] ), .B(n2596), .S(n1669), .Z(n7620) );
  MUX2_X1 U6164 ( .A(\REGISTERS[40][7] ), .B(n2585), .S(n1670), .Z(n7621) );
  MUX2_X1 U6165 ( .A(\REGISTERS[40][6] ), .B(n2574), .S(n1670), .Z(n7622) );
  MUX2_X1 U6166 ( .A(\REGISTERS[40][5] ), .B(n2563), .S(n1670), .Z(n7623) );
  MUX2_X1 U6167 ( .A(\REGISTERS[40][4] ), .B(n2552), .S(n1670), .Z(n7624) );
  MUX2_X1 U6168 ( .A(\REGISTERS[40][3] ), .B(n1837), .S(n1670), .Z(n7625) );
  MUX2_X1 U6169 ( .A(\REGISTERS[40][2] ), .B(n1826), .S(n1670), .Z(n7626) );
  MUX2_X1 U6170 ( .A(\REGISTERS[40][1] ), .B(n1815), .S(n1670), .Z(n7627) );
  MUX2_X1 U6171 ( .A(\REGISTERS[40][0] ), .B(n1804), .S(n1670), .Z(n7628) );
  MUX2_X1 U6172 ( .A(\REGISTERS[39][31] ), .B(n2951), .S(n1671), .Z(n7565) );
  MUX2_X1 U6173 ( .A(\REGISTERS[39][30] ), .B(n2940), .S(n1671), .Z(n7566) );
  MUX2_X1 U6174 ( .A(\REGISTERS[39][29] ), .B(n2929), .S(n1671), .Z(n7567) );
  MUX2_X1 U6175 ( .A(\REGISTERS[39][28] ), .B(n2913), .S(n1671), .Z(n7568) );
  MUX2_X1 U6176 ( .A(\REGISTERS[39][27] ), .B(n2902), .S(n1671), .Z(n7569) );
  MUX2_X1 U6177 ( .A(\REGISTERS[39][26] ), .B(n2890), .S(n1671), .Z(n7570) );
  MUX2_X1 U6178 ( .A(\REGISTERS[39][25] ), .B(n2879), .S(n1671), .Z(n7571) );
  MUX2_X1 U6179 ( .A(\REGISTERS[39][24] ), .B(n2868), .S(n1671), .Z(n7572) );
  MUX2_X1 U6180 ( .A(\REGISTERS[39][23] ), .B(n2857), .S(n1671), .Z(n7573) );
  MUX2_X1 U6181 ( .A(\REGISTERS[39][22] ), .B(n2846), .S(n1671), .Z(n7574) );
  MUX2_X1 U6182 ( .A(\REGISTERS[39][21] ), .B(n2835), .S(n1671), .Z(n7575) );
  MUX2_X1 U6183 ( .A(\REGISTERS[39][20] ), .B(n2824), .S(n1671), .Z(n7576) );
  MUX2_X1 U6184 ( .A(\REGISTERS[39][19] ), .B(n2813), .S(n1672), .Z(n7577) );
  MUX2_X1 U6185 ( .A(\REGISTERS[39][18] ), .B(n2802), .S(n1672), .Z(n7578) );
  MUX2_X1 U6186 ( .A(\REGISTERS[39][17] ), .B(n2791), .S(n1672), .Z(n7579) );
  MUX2_X1 U6187 ( .A(\REGISTERS[39][16] ), .B(n2780), .S(n1672), .Z(n7580) );
  MUX2_X1 U6188 ( .A(\REGISTERS[39][15] ), .B(n2769), .S(n1672), .Z(n7581) );
  MUX2_X1 U6189 ( .A(\REGISTERS[39][14] ), .B(n2758), .S(n1672), .Z(n7582) );
  MUX2_X1 U6190 ( .A(\REGISTERS[39][13] ), .B(n2747), .S(n1672), .Z(n7583) );
  MUX2_X1 U6191 ( .A(\REGISTERS[39][12] ), .B(n2736), .S(n1672), .Z(n7584) );
  MUX2_X1 U6192 ( .A(\REGISTERS[39][11] ), .B(n2725), .S(n1672), .Z(n7585) );
  MUX2_X1 U6193 ( .A(\REGISTERS[39][10] ), .B(n2714), .S(n1672), .Z(n7586) );
  MUX2_X1 U6194 ( .A(\REGISTERS[39][9] ), .B(n2607), .S(n1672), .Z(n7587) );
  MUX2_X1 U6195 ( .A(\REGISTERS[39][8] ), .B(n2596), .S(n1672), .Z(n7588) );
  MUX2_X1 U6196 ( .A(\REGISTERS[39][7] ), .B(n2585), .S(n1673), .Z(n7589) );
  MUX2_X1 U6197 ( .A(\REGISTERS[39][6] ), .B(n2574), .S(n1673), .Z(n7590) );
  MUX2_X1 U6198 ( .A(\REGISTERS[39][5] ), .B(n2563), .S(n1673), .Z(n7591) );
  MUX2_X1 U6199 ( .A(\REGISTERS[39][4] ), .B(n2552), .S(n1673), .Z(n7592) );
  MUX2_X1 U6200 ( .A(\REGISTERS[39][3] ), .B(n1837), .S(n1673), .Z(n7593) );
  MUX2_X1 U6201 ( .A(\REGISTERS[39][2] ), .B(n1826), .S(n1673), .Z(n7594) );
  MUX2_X1 U6202 ( .A(\REGISTERS[39][1] ), .B(n1815), .S(n1673), .Z(n7595) );
  MUX2_X1 U6203 ( .A(\REGISTERS[39][0] ), .B(n1804), .S(n1673), .Z(n7596) );
  MUX2_X1 U6204 ( .A(\REGISTERS[38][31] ), .B(n2951), .S(n1674), .Z(n7533) );
  MUX2_X1 U6205 ( .A(\REGISTERS[38][30] ), .B(n2940), .S(n1674), .Z(n7534) );
  MUX2_X1 U6206 ( .A(\REGISTERS[38][29] ), .B(n2929), .S(n1674), .Z(n7535) );
  MUX2_X1 U6207 ( .A(\REGISTERS[38][28] ), .B(n2913), .S(n1674), .Z(n7536) );
  MUX2_X1 U6208 ( .A(\REGISTERS[38][27] ), .B(n2902), .S(n1674), .Z(n7537) );
  MUX2_X1 U6209 ( .A(\REGISTERS[38][26] ), .B(n2890), .S(n1674), .Z(n7538) );
  MUX2_X1 U6210 ( .A(\REGISTERS[38][25] ), .B(n2879), .S(n1674), .Z(n7539) );
  MUX2_X1 U6211 ( .A(\REGISTERS[38][24] ), .B(n2868), .S(n1674), .Z(n7540) );
  MUX2_X1 U6212 ( .A(\REGISTERS[38][23] ), .B(n2857), .S(n1674), .Z(n7541) );
  MUX2_X1 U6213 ( .A(\REGISTERS[38][22] ), .B(n2846), .S(n1674), .Z(n7542) );
  MUX2_X1 U6214 ( .A(\REGISTERS[38][21] ), .B(n2835), .S(n1674), .Z(n7543) );
  MUX2_X1 U6215 ( .A(\REGISTERS[38][20] ), .B(n2824), .S(n1674), .Z(n7544) );
  MUX2_X1 U6216 ( .A(\REGISTERS[38][19] ), .B(n2813), .S(n1675), .Z(n7545) );
  MUX2_X1 U6217 ( .A(\REGISTERS[38][18] ), .B(n2802), .S(n1675), .Z(n7546) );
  MUX2_X1 U6218 ( .A(\REGISTERS[38][17] ), .B(n2791), .S(n1675), .Z(n7547) );
  MUX2_X1 U6219 ( .A(\REGISTERS[38][16] ), .B(n2780), .S(n1675), .Z(n7548) );
  MUX2_X1 U6220 ( .A(\REGISTERS[38][15] ), .B(n2769), .S(n1675), .Z(n7549) );
  MUX2_X1 U6221 ( .A(\REGISTERS[38][14] ), .B(n2758), .S(n1675), .Z(n7550) );
  MUX2_X1 U6222 ( .A(\REGISTERS[38][13] ), .B(n2747), .S(n1675), .Z(n7551) );
  MUX2_X1 U6223 ( .A(\REGISTERS[38][12] ), .B(n2736), .S(n1675), .Z(n7552) );
  MUX2_X1 U6224 ( .A(\REGISTERS[38][11] ), .B(n2725), .S(n1675), .Z(n7553) );
  MUX2_X1 U6225 ( .A(\REGISTERS[38][10] ), .B(n2714), .S(n1675), .Z(n7554) );
  MUX2_X1 U6226 ( .A(\REGISTERS[38][9] ), .B(n2607), .S(n1675), .Z(n7555) );
  MUX2_X1 U6227 ( .A(\REGISTERS[38][8] ), .B(n2596), .S(n1675), .Z(n7556) );
  MUX2_X1 U6228 ( .A(\REGISTERS[38][7] ), .B(n2585), .S(n1676), .Z(n7557) );
  MUX2_X1 U6229 ( .A(\REGISTERS[38][6] ), .B(n2574), .S(n1676), .Z(n7558) );
  MUX2_X1 U6230 ( .A(\REGISTERS[38][5] ), .B(n2563), .S(n1676), .Z(n7559) );
  MUX2_X1 U6231 ( .A(\REGISTERS[38][4] ), .B(n2552), .S(n1676), .Z(n7560) );
  MUX2_X1 U6232 ( .A(\REGISTERS[38][3] ), .B(n1837), .S(n1676), .Z(n7561) );
  MUX2_X1 U6233 ( .A(\REGISTERS[38][2] ), .B(n1826), .S(n1676), .Z(n7562) );
  MUX2_X1 U6234 ( .A(\REGISTERS[38][1] ), .B(n1815), .S(n1676), .Z(n7563) );
  MUX2_X1 U6235 ( .A(\REGISTERS[38][0] ), .B(n1804), .S(n1676), .Z(n7564) );
  MUX2_X1 U6236 ( .A(n9990), .B(n2951), .S(n1677), .Z(n7501) );
  MUX2_X1 U6237 ( .A(n9991), .B(n2940), .S(n1677), .Z(n7502) );
  MUX2_X1 U6238 ( .A(n9992), .B(n2929), .S(n1677), .Z(n7503) );
  MUX2_X1 U6239 ( .A(n9993), .B(n2913), .S(n1677), .Z(n7504) );
  MUX2_X1 U6240 ( .A(n9994), .B(n2902), .S(n1677), .Z(n7505) );
  MUX2_X1 U6241 ( .A(n9995), .B(n2890), .S(n1677), .Z(n7506) );
  MUX2_X1 U6242 ( .A(n9996), .B(n2879), .S(n1677), .Z(n7507) );
  MUX2_X1 U6243 ( .A(n9997), .B(n2868), .S(n1677), .Z(n7508) );
  MUX2_X1 U6244 ( .A(n9998), .B(n2857), .S(n1677), .Z(n7509) );
  MUX2_X1 U6245 ( .A(n9999), .B(n2846), .S(n1677), .Z(n7510) );
  MUX2_X1 U6246 ( .A(n10000), .B(n2835), .S(n1677), .Z(n7511) );
  MUX2_X1 U6247 ( .A(n10001), .B(n2824), .S(n1677), .Z(n7512) );
  MUX2_X1 U6248 ( .A(n10002), .B(n2813), .S(n1678), .Z(n7513) );
  MUX2_X1 U6249 ( .A(n10003), .B(n2802), .S(n1678), .Z(n7514) );
  MUX2_X1 U6250 ( .A(n10004), .B(n2791), .S(n1678), .Z(n7515) );
  MUX2_X1 U6251 ( .A(n10005), .B(n2780), .S(n1678), .Z(n7516) );
  MUX2_X1 U6252 ( .A(n10006), .B(n2769), .S(n1678), .Z(n7517) );
  MUX2_X1 U6253 ( .A(n10007), .B(n2758), .S(n1678), .Z(n7518) );
  MUX2_X1 U6254 ( .A(n10008), .B(n2747), .S(n1678), .Z(n7519) );
  MUX2_X1 U6255 ( .A(n10009), .B(n2736), .S(n1678), .Z(n7520) );
  MUX2_X1 U6256 ( .A(n10010), .B(n2725), .S(n1678), .Z(n7521) );
  MUX2_X1 U6257 ( .A(n10011), .B(n2714), .S(n1678), .Z(n7522) );
  MUX2_X1 U6258 ( .A(n10012), .B(n2607), .S(n1678), .Z(n7523) );
  MUX2_X1 U6259 ( .A(n10013), .B(n2596), .S(n1678), .Z(n7524) );
  MUX2_X1 U6260 ( .A(n10014), .B(n2585), .S(n1679), .Z(n7525) );
  MUX2_X1 U6261 ( .A(n10015), .B(n2574), .S(n1679), .Z(n7526) );
  MUX2_X1 U6262 ( .A(n10016), .B(n2563), .S(n1679), .Z(n7527) );
  MUX2_X1 U6263 ( .A(n10017), .B(n2552), .S(n1679), .Z(n7528) );
  MUX2_X1 U6264 ( .A(n10018), .B(n1837), .S(n1679), .Z(n7529) );
  MUX2_X1 U6265 ( .A(n10019), .B(n1826), .S(n1679), .Z(n7530) );
  MUX2_X1 U6266 ( .A(n10020), .B(n1815), .S(n1679), .Z(n7531) );
  MUX2_X1 U6267 ( .A(n10021), .B(n1804), .S(n1679), .Z(n7532) );
  MUX2_X1 U6268 ( .A(n9958), .B(n2951), .S(n1680), .Z(n7469) );
  MUX2_X1 U6269 ( .A(n9959), .B(n2940), .S(n1680), .Z(n7470) );
  MUX2_X1 U6270 ( .A(n9960), .B(n2929), .S(n1680), .Z(n7471) );
  MUX2_X1 U6271 ( .A(n9961), .B(n2913), .S(n1680), .Z(n7472) );
  MUX2_X1 U6272 ( .A(n9962), .B(n2902), .S(n1680), .Z(n7473) );
  MUX2_X1 U6273 ( .A(n9963), .B(n2890), .S(n1680), .Z(n7474) );
  MUX2_X1 U6274 ( .A(n9964), .B(n2879), .S(n1680), .Z(n7475) );
  MUX2_X1 U6275 ( .A(n9965), .B(n2868), .S(n1680), .Z(n7476) );
  MUX2_X1 U6276 ( .A(n9966), .B(n2857), .S(n1680), .Z(n7477) );
  MUX2_X1 U6277 ( .A(n9967), .B(n2846), .S(n1680), .Z(n7478) );
  MUX2_X1 U6278 ( .A(n9968), .B(n2835), .S(n1680), .Z(n7479) );
  MUX2_X1 U6279 ( .A(n9969), .B(n2824), .S(n1680), .Z(n7480) );
  MUX2_X1 U6280 ( .A(n9970), .B(n2813), .S(n1681), .Z(n7481) );
  MUX2_X1 U6281 ( .A(n9971), .B(n2802), .S(n1681), .Z(n7482) );
  MUX2_X1 U6282 ( .A(n9972), .B(n2791), .S(n1681), .Z(n7483) );
  MUX2_X1 U6283 ( .A(n9973), .B(n2780), .S(n1681), .Z(n7484) );
  MUX2_X1 U6284 ( .A(n9974), .B(n2769), .S(n1681), .Z(n7485) );
  MUX2_X1 U6285 ( .A(n9975), .B(n2758), .S(n1681), .Z(n7486) );
  MUX2_X1 U6286 ( .A(n9976), .B(n2747), .S(n1681), .Z(n7487) );
  MUX2_X1 U6287 ( .A(n9977), .B(n2736), .S(n1681), .Z(n7488) );
  MUX2_X1 U6288 ( .A(n9978), .B(n2725), .S(n1681), .Z(n7489) );
  MUX2_X1 U6289 ( .A(n9979), .B(n2714), .S(n1681), .Z(n7490) );
  MUX2_X1 U6290 ( .A(n9980), .B(n2607), .S(n1681), .Z(n7491) );
  MUX2_X1 U6291 ( .A(n9981), .B(n2596), .S(n1681), .Z(n7492) );
  MUX2_X1 U6292 ( .A(n9982), .B(n2585), .S(n1682), .Z(n7493) );
  MUX2_X1 U6293 ( .A(n9983), .B(n2574), .S(n1682), .Z(n7494) );
  MUX2_X1 U6294 ( .A(n9984), .B(n2563), .S(n1682), .Z(n7495) );
  MUX2_X1 U6295 ( .A(n9985), .B(n2552), .S(n1682), .Z(n7496) );
  MUX2_X1 U6296 ( .A(n9986), .B(n1837), .S(n1682), .Z(n7497) );
  MUX2_X1 U6297 ( .A(n9987), .B(n1826), .S(n1682), .Z(n7498) );
  MUX2_X1 U6298 ( .A(n9988), .B(n1815), .S(n1682), .Z(n7499) );
  MUX2_X1 U6299 ( .A(n9989), .B(n1804), .S(n1682), .Z(n7500) );
  MUX2_X1 U6300 ( .A(n9926), .B(n2951), .S(n1683), .Z(n7437) );
  MUX2_X1 U6301 ( .A(n9927), .B(n2940), .S(n1683), .Z(n7438) );
  MUX2_X1 U6302 ( .A(n9928), .B(n2929), .S(n1683), .Z(n7439) );
  MUX2_X1 U6303 ( .A(n9929), .B(n2913), .S(n1683), .Z(n7440) );
  MUX2_X1 U6304 ( .A(n9930), .B(n2902), .S(n1683), .Z(n7441) );
  MUX2_X1 U6305 ( .A(n9931), .B(n2890), .S(n1683), .Z(n7442) );
  MUX2_X1 U6306 ( .A(n9932), .B(n2879), .S(n1683), .Z(n7443) );
  MUX2_X1 U6307 ( .A(n9933), .B(n2868), .S(n1683), .Z(n7444) );
  MUX2_X1 U6308 ( .A(n9934), .B(n2857), .S(n1683), .Z(n7445) );
  MUX2_X1 U6309 ( .A(n9935), .B(n2846), .S(n1683), .Z(n7446) );
  MUX2_X1 U6310 ( .A(n9936), .B(n2835), .S(n1683), .Z(n7447) );
  MUX2_X1 U6311 ( .A(n9937), .B(n2824), .S(n1683), .Z(n7448) );
  MUX2_X1 U6312 ( .A(n9938), .B(n2813), .S(n1684), .Z(n7449) );
  MUX2_X1 U6313 ( .A(n9939), .B(n2802), .S(n1684), .Z(n7450) );
  MUX2_X1 U6314 ( .A(n9940), .B(n2791), .S(n1684), .Z(n7451) );
  MUX2_X1 U6315 ( .A(n9941), .B(n2780), .S(n1684), .Z(n7452) );
  MUX2_X1 U6316 ( .A(n9942), .B(n2769), .S(n1684), .Z(n7453) );
  MUX2_X1 U6317 ( .A(n9943), .B(n2758), .S(n1684), .Z(n7454) );
  MUX2_X1 U6318 ( .A(n9944), .B(n2747), .S(n1684), .Z(n7455) );
  MUX2_X1 U6319 ( .A(n9945), .B(n2736), .S(n1684), .Z(n7456) );
  MUX2_X1 U6320 ( .A(n9946), .B(n2725), .S(n1684), .Z(n7457) );
  MUX2_X1 U6321 ( .A(n9947), .B(n2714), .S(n1684), .Z(n7458) );
  MUX2_X1 U6322 ( .A(n9948), .B(n2607), .S(n1684), .Z(n7459) );
  MUX2_X1 U6323 ( .A(n9949), .B(n2596), .S(n1684), .Z(n7460) );
  MUX2_X1 U6324 ( .A(n9950), .B(n2585), .S(n1685), .Z(n7461) );
  MUX2_X1 U6325 ( .A(n9951), .B(n2574), .S(n1685), .Z(n7462) );
  MUX2_X1 U6326 ( .A(n9952), .B(n2563), .S(n1685), .Z(n7463) );
  MUX2_X1 U6327 ( .A(n9953), .B(n2552), .S(n1685), .Z(n7464) );
  MUX2_X1 U6328 ( .A(n9954), .B(n1837), .S(n1685), .Z(n7465) );
  MUX2_X1 U6329 ( .A(n9955), .B(n1826), .S(n1685), .Z(n7466) );
  MUX2_X1 U6330 ( .A(n9956), .B(n1815), .S(n1685), .Z(n7467) );
  MUX2_X1 U6331 ( .A(n9957), .B(n1804), .S(n1685), .Z(n7468) );
  MUX2_X1 U6332 ( .A(\REGISTERS[34][31] ), .B(n2951), .S(n1686), .Z(n7405) );
  MUX2_X1 U6333 ( .A(\REGISTERS[34][30] ), .B(n2940), .S(n1686), .Z(n7406) );
  MUX2_X1 U6334 ( .A(\REGISTERS[34][29] ), .B(n2929), .S(n1686), .Z(n7407) );
  MUX2_X1 U6335 ( .A(\REGISTERS[34][28] ), .B(n2913), .S(n1686), .Z(n7408) );
  MUX2_X1 U6336 ( .A(\REGISTERS[34][27] ), .B(n2902), .S(n1686), .Z(n7409) );
  MUX2_X1 U6337 ( .A(\REGISTERS[34][26] ), .B(n2890), .S(n1686), .Z(n7410) );
  MUX2_X1 U6338 ( .A(\REGISTERS[34][25] ), .B(n2879), .S(n1686), .Z(n7411) );
  MUX2_X1 U6339 ( .A(\REGISTERS[34][24] ), .B(n2868), .S(n1686), .Z(n7412) );
  MUX2_X1 U6340 ( .A(\REGISTERS[34][23] ), .B(n2857), .S(n1686), .Z(n7413) );
  MUX2_X1 U6341 ( .A(\REGISTERS[34][22] ), .B(n2846), .S(n1686), .Z(n7414) );
  MUX2_X1 U6342 ( .A(\REGISTERS[34][21] ), .B(n2835), .S(n1686), .Z(n7415) );
  MUX2_X1 U6343 ( .A(\REGISTERS[34][20] ), .B(n2824), .S(n1686), .Z(n7416) );
  MUX2_X1 U6344 ( .A(\REGISTERS[34][19] ), .B(n2813), .S(n1687), .Z(n7417) );
  MUX2_X1 U6345 ( .A(\REGISTERS[34][18] ), .B(n2802), .S(n1687), .Z(n7418) );
  MUX2_X1 U6346 ( .A(\REGISTERS[34][17] ), .B(n2791), .S(n1687), .Z(n7419) );
  MUX2_X1 U6347 ( .A(\REGISTERS[34][16] ), .B(n2780), .S(n1687), .Z(n7420) );
  MUX2_X1 U6348 ( .A(\REGISTERS[34][15] ), .B(n2769), .S(n1687), .Z(n7421) );
  MUX2_X1 U6349 ( .A(\REGISTERS[34][14] ), .B(n2758), .S(n1687), .Z(n7422) );
  MUX2_X1 U6350 ( .A(\REGISTERS[34][13] ), .B(n2747), .S(n1687), .Z(n7423) );
  MUX2_X1 U6351 ( .A(\REGISTERS[34][12] ), .B(n2736), .S(n1687), .Z(n7424) );
  MUX2_X1 U6352 ( .A(\REGISTERS[34][11] ), .B(n2725), .S(n1687), .Z(n7425) );
  MUX2_X1 U6353 ( .A(\REGISTERS[34][10] ), .B(n2714), .S(n1687), .Z(n7426) );
  MUX2_X1 U6354 ( .A(\REGISTERS[34][9] ), .B(n2607), .S(n1687), .Z(n7427) );
  MUX2_X1 U6355 ( .A(\REGISTERS[34][8] ), .B(n2596), .S(n1687), .Z(n7428) );
  MUX2_X1 U6356 ( .A(\REGISTERS[34][7] ), .B(n2585), .S(n1688), .Z(n7429) );
  MUX2_X1 U6357 ( .A(\REGISTERS[34][6] ), .B(n2574), .S(n1688), .Z(n7430) );
  MUX2_X1 U6358 ( .A(\REGISTERS[34][5] ), .B(n2563), .S(n1688), .Z(n7431) );
  MUX2_X1 U6359 ( .A(\REGISTERS[34][4] ), .B(n2552), .S(n1688), .Z(n7432) );
  MUX2_X1 U6360 ( .A(\REGISTERS[34][3] ), .B(n1837), .S(n1688), .Z(n7433) );
  MUX2_X1 U6361 ( .A(\REGISTERS[34][2] ), .B(n1826), .S(n1688), .Z(n7434) );
  MUX2_X1 U6362 ( .A(\REGISTERS[34][1] ), .B(n1815), .S(n1688), .Z(n7435) );
  MUX2_X1 U6363 ( .A(\REGISTERS[34][0] ), .B(n1804), .S(n1688), .Z(n7436) );
  MUX2_X1 U6364 ( .A(\REGISTERS[33][31] ), .B(n2951), .S(n1689), .Z(n7373) );
  MUX2_X1 U6365 ( .A(\REGISTERS[33][30] ), .B(n2940), .S(n1689), .Z(n7374) );
  MUX2_X1 U6366 ( .A(\REGISTERS[33][29] ), .B(n2929), .S(n1689), .Z(n7375) );
  MUX2_X1 U6367 ( .A(\REGISTERS[33][28] ), .B(n2913), .S(n1689), .Z(n7376) );
  MUX2_X1 U6368 ( .A(\REGISTERS[33][27] ), .B(n2902), .S(n1689), .Z(n7377) );
  MUX2_X1 U6369 ( .A(\REGISTERS[33][26] ), .B(n2890), .S(n1689), .Z(n7378) );
  MUX2_X1 U6370 ( .A(\REGISTERS[33][25] ), .B(n2879), .S(n1689), .Z(n7379) );
  MUX2_X1 U6371 ( .A(\REGISTERS[33][24] ), .B(n2868), .S(n1689), .Z(n7380) );
  MUX2_X1 U6372 ( .A(\REGISTERS[33][23] ), .B(n2857), .S(n1689), .Z(n7381) );
  MUX2_X1 U6373 ( .A(\REGISTERS[33][22] ), .B(n2846), .S(n1689), .Z(n7382) );
  MUX2_X1 U6374 ( .A(\REGISTERS[33][21] ), .B(n2835), .S(n1689), .Z(n7383) );
  MUX2_X1 U6375 ( .A(\REGISTERS[33][20] ), .B(n2824), .S(n1689), .Z(n7384) );
  MUX2_X1 U6376 ( .A(\REGISTERS[33][19] ), .B(n2813), .S(n1690), .Z(n7385) );
  MUX2_X1 U6377 ( .A(\REGISTERS[33][18] ), .B(n2802), .S(n1690), .Z(n7386) );
  MUX2_X1 U6378 ( .A(\REGISTERS[33][17] ), .B(n2791), .S(n1690), .Z(n7387) );
  MUX2_X1 U6379 ( .A(\REGISTERS[33][16] ), .B(n2780), .S(n1690), .Z(n7388) );
  MUX2_X1 U6380 ( .A(\REGISTERS[33][15] ), .B(n2769), .S(n1690), .Z(n7389) );
  MUX2_X1 U6381 ( .A(\REGISTERS[33][14] ), .B(n2758), .S(n1690), .Z(n7390) );
  MUX2_X1 U6382 ( .A(\REGISTERS[33][13] ), .B(n2747), .S(n1690), .Z(n7391) );
  MUX2_X1 U6383 ( .A(\REGISTERS[33][12] ), .B(n2736), .S(n1690), .Z(n7392) );
  MUX2_X1 U6384 ( .A(\REGISTERS[33][11] ), .B(n2725), .S(n1690), .Z(n7393) );
  MUX2_X1 U6385 ( .A(\REGISTERS[33][10] ), .B(n2714), .S(n1690), .Z(n7394) );
  MUX2_X1 U6386 ( .A(\REGISTERS[33][9] ), .B(n2607), .S(n1690), .Z(n7395) );
  MUX2_X1 U6387 ( .A(\REGISTERS[33][8] ), .B(n2596), .S(n1690), .Z(n7396) );
  MUX2_X1 U6388 ( .A(\REGISTERS[33][7] ), .B(n2585), .S(n1691), .Z(n7397) );
  MUX2_X1 U6389 ( .A(\REGISTERS[33][6] ), .B(n2574), .S(n1691), .Z(n7398) );
  MUX2_X1 U6390 ( .A(\REGISTERS[33][5] ), .B(n2563), .S(n1691), .Z(n7399) );
  MUX2_X1 U6391 ( .A(\REGISTERS[33][4] ), .B(n2552), .S(n1691), .Z(n7400) );
  MUX2_X1 U6392 ( .A(\REGISTERS[33][3] ), .B(n1837), .S(n1691), .Z(n7401) );
  MUX2_X1 U6393 ( .A(\REGISTERS[33][2] ), .B(n1826), .S(n1691), .Z(n7402) );
  MUX2_X1 U6394 ( .A(\REGISTERS[33][1] ), .B(n1815), .S(n1691), .Z(n7403) );
  MUX2_X1 U6395 ( .A(\REGISTERS[33][0] ), .B(n1804), .S(n1691), .Z(n7404) );
  MUX2_X1 U6396 ( .A(n9894), .B(n2952), .S(n1692), .Z(n7341) );
  MUX2_X1 U6397 ( .A(n9895), .B(n2941), .S(n1692), .Z(n7342) );
  MUX2_X1 U6398 ( .A(n9896), .B(n2930), .S(n1692), .Z(n7343) );
  MUX2_X1 U6399 ( .A(n9897), .B(n2914), .S(n1692), .Z(n7344) );
  MUX2_X1 U6400 ( .A(n9898), .B(n2903), .S(n1692), .Z(n7345) );
  MUX2_X1 U6401 ( .A(n9899), .B(n2891), .S(n1692), .Z(n7346) );
  MUX2_X1 U6402 ( .A(n9900), .B(n2880), .S(n1692), .Z(n7347) );
  MUX2_X1 U6403 ( .A(n9901), .B(n2869), .S(n1692), .Z(n7348) );
  MUX2_X1 U6404 ( .A(n9902), .B(n2858), .S(n1692), .Z(n7349) );
  MUX2_X1 U6405 ( .A(n9903), .B(n2847), .S(n1692), .Z(n7350) );
  MUX2_X1 U6406 ( .A(n9904), .B(n2836), .S(n1692), .Z(n7351) );
  MUX2_X1 U6407 ( .A(n9905), .B(n2825), .S(n1692), .Z(n7352) );
  MUX2_X1 U6408 ( .A(n9906), .B(n2814), .S(n1693), .Z(n7353) );
  MUX2_X1 U6409 ( .A(n9907), .B(n2803), .S(n1693), .Z(n7354) );
  MUX2_X1 U6410 ( .A(n9908), .B(n2792), .S(n1693), .Z(n7355) );
  MUX2_X1 U6411 ( .A(n9909), .B(n2781), .S(n1693), .Z(n7356) );
  MUX2_X1 U6412 ( .A(n9910), .B(n2770), .S(n1693), .Z(n7357) );
  MUX2_X1 U6413 ( .A(n9911), .B(n2759), .S(n1693), .Z(n7358) );
  MUX2_X1 U6414 ( .A(n9912), .B(n2748), .S(n1693), .Z(n7359) );
  MUX2_X1 U6415 ( .A(n9913), .B(n2737), .S(n1693), .Z(n7360) );
  MUX2_X1 U6416 ( .A(n9914), .B(n2726), .S(n1693), .Z(n7361) );
  MUX2_X1 U6417 ( .A(n9915), .B(n2715), .S(n1693), .Z(n7362) );
  MUX2_X1 U6418 ( .A(n9916), .B(n2704), .S(n1693), .Z(n7363) );
  MUX2_X1 U6419 ( .A(n9917), .B(n2597), .S(n1693), .Z(n7364) );
  MUX2_X1 U6420 ( .A(n9918), .B(n2586), .S(n1694), .Z(n7365) );
  MUX2_X1 U6421 ( .A(n9919), .B(n2575), .S(n1694), .Z(n7366) );
  MUX2_X1 U6422 ( .A(n9920), .B(n2564), .S(n1694), .Z(n7367) );
  MUX2_X1 U6423 ( .A(n9921), .B(n2553), .S(n1694), .Z(n7368) );
  MUX2_X1 U6424 ( .A(n9922), .B(n1838), .S(n1694), .Z(n7369) );
  MUX2_X1 U6425 ( .A(n9923), .B(n1827), .S(n1694), .Z(n7370) );
  MUX2_X1 U6426 ( .A(n9924), .B(n1816), .S(n1694), .Z(n7371) );
  MUX2_X1 U6427 ( .A(n9925), .B(n1805), .S(n1694), .Z(n7372) );
  MUX2_X1 U6428 ( .A(n9862), .B(n2952), .S(n1695), .Z(n7309) );
  MUX2_X1 U6429 ( .A(n9863), .B(n2941), .S(n1695), .Z(n7310) );
  MUX2_X1 U6430 ( .A(n9864), .B(n2930), .S(n1695), .Z(n7311) );
  MUX2_X1 U6431 ( .A(n9865), .B(n2914), .S(n1695), .Z(n7312) );
  MUX2_X1 U6432 ( .A(n9866), .B(n2903), .S(n1695), .Z(n7313) );
  MUX2_X1 U6433 ( .A(n9867), .B(n2891), .S(n1695), .Z(n7314) );
  MUX2_X1 U6434 ( .A(n9868), .B(n2880), .S(n1695), .Z(n7315) );
  MUX2_X1 U6435 ( .A(n9869), .B(n2869), .S(n1695), .Z(n7316) );
  MUX2_X1 U6436 ( .A(n9870), .B(n2858), .S(n1695), .Z(n7317) );
  MUX2_X1 U6437 ( .A(n9871), .B(n2847), .S(n1695), .Z(n7318) );
  MUX2_X1 U6438 ( .A(n9872), .B(n2836), .S(n1695), .Z(n7319) );
  MUX2_X1 U6439 ( .A(n9873), .B(n2825), .S(n1695), .Z(n7320) );
  MUX2_X1 U6440 ( .A(n9874), .B(n2814), .S(n1696), .Z(n7321) );
  MUX2_X1 U6441 ( .A(n9875), .B(n2803), .S(n1696), .Z(n7322) );
  MUX2_X1 U6442 ( .A(n9876), .B(n2792), .S(n1696), .Z(n7323) );
  MUX2_X1 U6443 ( .A(n9877), .B(n2781), .S(n1696), .Z(n7324) );
  MUX2_X1 U6444 ( .A(n9878), .B(n2770), .S(n1696), .Z(n7325) );
  MUX2_X1 U6445 ( .A(n9879), .B(n2759), .S(n1696), .Z(n7326) );
  MUX2_X1 U6446 ( .A(n9880), .B(n2748), .S(n1696), .Z(n7327) );
  MUX2_X1 U6447 ( .A(n9881), .B(n2737), .S(n1696), .Z(n7328) );
  MUX2_X1 U6448 ( .A(n9882), .B(n2726), .S(n1696), .Z(n7329) );
  MUX2_X1 U6449 ( .A(n9883), .B(n2715), .S(n1696), .Z(n7330) );
  MUX2_X1 U6450 ( .A(n9884), .B(n2704), .S(n1696), .Z(n7331) );
  MUX2_X1 U6451 ( .A(n9885), .B(n2597), .S(n1696), .Z(n7332) );
  MUX2_X1 U6452 ( .A(n9886), .B(n2586), .S(n1697), .Z(n7333) );
  MUX2_X1 U6453 ( .A(n9887), .B(n2575), .S(n1697), .Z(n7334) );
  MUX2_X1 U6454 ( .A(n9888), .B(n2564), .S(n1697), .Z(n7335) );
  MUX2_X1 U6455 ( .A(n9889), .B(n2553), .S(n1697), .Z(n7336) );
  MUX2_X1 U6456 ( .A(n9890), .B(n1838), .S(n1697), .Z(n7337) );
  MUX2_X1 U6457 ( .A(n9891), .B(n1827), .S(n1697), .Z(n7338) );
  MUX2_X1 U6458 ( .A(n9892), .B(n1816), .S(n1697), .Z(n7339) );
  MUX2_X1 U6459 ( .A(n9893), .B(n1805), .S(n1697), .Z(n7340) );
  MUX2_X1 U6460 ( .A(n9830), .B(n2952), .S(n1698), .Z(n7277) );
  MUX2_X1 U6461 ( .A(n9831), .B(n2941), .S(n1698), .Z(n7278) );
  MUX2_X1 U6462 ( .A(n9832), .B(n2930), .S(n1698), .Z(n7279) );
  MUX2_X1 U6463 ( .A(n9833), .B(n2914), .S(n1698), .Z(n7280) );
  MUX2_X1 U6464 ( .A(n9834), .B(n2903), .S(n1698), .Z(n7281) );
  MUX2_X1 U6465 ( .A(n9835), .B(n2891), .S(n1698), .Z(n7282) );
  MUX2_X1 U6466 ( .A(n9836), .B(n2880), .S(n1698), .Z(n7283) );
  MUX2_X1 U6467 ( .A(n9837), .B(n2869), .S(n1698), .Z(n7284) );
  MUX2_X1 U6468 ( .A(n9838), .B(n2858), .S(n1698), .Z(n7285) );
  MUX2_X1 U6469 ( .A(n9839), .B(n2847), .S(n1698), .Z(n7286) );
  MUX2_X1 U6470 ( .A(n9840), .B(n2836), .S(n1698), .Z(n7287) );
  MUX2_X1 U6471 ( .A(n9841), .B(n2825), .S(n1698), .Z(n7288) );
  MUX2_X1 U6472 ( .A(n9842), .B(n2814), .S(n1699), .Z(n7289) );
  MUX2_X1 U6473 ( .A(n9843), .B(n2803), .S(n1699), .Z(n7290) );
  MUX2_X1 U6474 ( .A(n9844), .B(n2792), .S(n1699), .Z(n7291) );
  MUX2_X1 U6475 ( .A(n9845), .B(n2781), .S(n1699), .Z(n7292) );
  MUX2_X1 U6476 ( .A(n9846), .B(n2770), .S(n1699), .Z(n7293) );
  MUX2_X1 U6477 ( .A(n9847), .B(n2759), .S(n1699), .Z(n7294) );
  MUX2_X1 U6478 ( .A(n9848), .B(n2748), .S(n1699), .Z(n7295) );
  MUX2_X1 U6479 ( .A(n9849), .B(n2737), .S(n1699), .Z(n7296) );
  MUX2_X1 U6480 ( .A(n9850), .B(n2726), .S(n1699), .Z(n7297) );
  MUX2_X1 U6481 ( .A(n9851), .B(n2715), .S(n1699), .Z(n7298) );
  MUX2_X1 U6482 ( .A(n9852), .B(n2704), .S(n1699), .Z(n7299) );
  MUX2_X1 U6483 ( .A(n9853), .B(n2597), .S(n1699), .Z(n7300) );
  MUX2_X1 U6484 ( .A(n9854), .B(n2586), .S(n1700), .Z(n7301) );
  MUX2_X1 U6485 ( .A(n9855), .B(n2575), .S(n1700), .Z(n7302) );
  MUX2_X1 U6486 ( .A(n9856), .B(n2564), .S(n1700), .Z(n7303) );
  MUX2_X1 U6487 ( .A(n9857), .B(n2553), .S(n1700), .Z(n7304) );
  MUX2_X1 U6488 ( .A(n9858), .B(n1838), .S(n1700), .Z(n7305) );
  MUX2_X1 U6489 ( .A(n9859), .B(n1827), .S(n1700), .Z(n7306) );
  MUX2_X1 U6490 ( .A(n9860), .B(n1816), .S(n1700), .Z(n7307) );
  MUX2_X1 U6491 ( .A(n9861), .B(n1805), .S(n1700), .Z(n7308) );
  MUX2_X1 U6492 ( .A(n9798), .B(n2952), .S(n1701), .Z(n7245) );
  MUX2_X1 U6493 ( .A(n9799), .B(n2941), .S(n1701), .Z(n7246) );
  MUX2_X1 U6494 ( .A(n9800), .B(n2930), .S(n1701), .Z(n7247) );
  MUX2_X1 U6495 ( .A(n9801), .B(n2914), .S(n1701), .Z(n7248) );
  MUX2_X1 U6496 ( .A(n9802), .B(n2903), .S(n1701), .Z(n7249) );
  MUX2_X1 U6497 ( .A(n9803), .B(n2891), .S(n1701), .Z(n7250) );
  MUX2_X1 U6498 ( .A(n9804), .B(n2880), .S(n1701), .Z(n7251) );
  MUX2_X1 U6499 ( .A(n9805), .B(n2869), .S(n1701), .Z(n7252) );
  MUX2_X1 U6500 ( .A(n9806), .B(n2858), .S(n1701), .Z(n7253) );
  MUX2_X1 U6501 ( .A(n9807), .B(n2847), .S(n1701), .Z(n7254) );
  MUX2_X1 U6502 ( .A(n9808), .B(n2836), .S(n1701), .Z(n7255) );
  MUX2_X1 U6503 ( .A(n9809), .B(n2825), .S(n1701), .Z(n7256) );
  MUX2_X1 U6504 ( .A(n9810), .B(n2814), .S(n1702), .Z(n7257) );
  MUX2_X1 U6505 ( .A(n9811), .B(n2803), .S(n1702), .Z(n7258) );
  MUX2_X1 U6506 ( .A(n9812), .B(n2792), .S(n1702), .Z(n7259) );
  MUX2_X1 U6507 ( .A(n9813), .B(n2781), .S(n1702), .Z(n7260) );
  MUX2_X1 U6508 ( .A(n9814), .B(n2770), .S(n1702), .Z(n7261) );
  MUX2_X1 U6509 ( .A(n9815), .B(n2759), .S(n1702), .Z(n7262) );
  MUX2_X1 U6510 ( .A(n9816), .B(n2748), .S(n1702), .Z(n7263) );
  MUX2_X1 U6511 ( .A(n9817), .B(n2737), .S(n1702), .Z(n7264) );
  MUX2_X1 U6512 ( .A(n9818), .B(n2726), .S(n1702), .Z(n7265) );
  MUX2_X1 U6513 ( .A(n9819), .B(n2715), .S(n1702), .Z(n7266) );
  MUX2_X1 U6514 ( .A(n9820), .B(n2704), .S(n1702), .Z(n7267) );
  MUX2_X1 U6515 ( .A(n9821), .B(n2597), .S(n1702), .Z(n7268) );
  MUX2_X1 U6516 ( .A(n9822), .B(n2586), .S(n1703), .Z(n7269) );
  MUX2_X1 U6517 ( .A(n9823), .B(n2575), .S(n1703), .Z(n7270) );
  MUX2_X1 U6518 ( .A(n9824), .B(n2564), .S(n1703), .Z(n7271) );
  MUX2_X1 U6519 ( .A(n9825), .B(n2553), .S(n1703), .Z(n7272) );
  MUX2_X1 U6520 ( .A(n9826), .B(n1838), .S(n1703), .Z(n7273) );
  MUX2_X1 U6521 ( .A(n9827), .B(n1827), .S(n1703), .Z(n7274) );
  MUX2_X1 U6522 ( .A(n9828), .B(n1816), .S(n1703), .Z(n7275) );
  MUX2_X1 U6523 ( .A(n9829), .B(n1805), .S(n1703), .Z(n7276) );
  MUX2_X1 U6524 ( .A(n9766), .B(n2952), .S(n1704), .Z(n7213) );
  MUX2_X1 U6525 ( .A(n9767), .B(n2941), .S(n1704), .Z(n7214) );
  MUX2_X1 U6526 ( .A(n9768), .B(n2930), .S(n1704), .Z(n7215) );
  MUX2_X1 U6527 ( .A(n9769), .B(n2914), .S(n1704), .Z(n7216) );
  MUX2_X1 U6528 ( .A(n9770), .B(n2903), .S(n1704), .Z(n7217) );
  MUX2_X1 U6529 ( .A(n9771), .B(n2891), .S(n1704), .Z(n7218) );
  MUX2_X1 U6530 ( .A(n9772), .B(n2880), .S(n1704), .Z(n7219) );
  MUX2_X1 U6531 ( .A(n9773), .B(n2869), .S(n1704), .Z(n7220) );
  MUX2_X1 U6532 ( .A(n9774), .B(n2858), .S(n1704), .Z(n7221) );
  MUX2_X1 U6533 ( .A(n9775), .B(n2847), .S(n1704), .Z(n7222) );
  MUX2_X1 U6534 ( .A(n9776), .B(n2836), .S(n1704), .Z(n7223) );
  MUX2_X1 U6535 ( .A(n9777), .B(n2825), .S(n1704), .Z(n7224) );
  MUX2_X1 U6536 ( .A(n9778), .B(n2814), .S(n1705), .Z(n7225) );
  MUX2_X1 U6537 ( .A(n9779), .B(n2803), .S(n1705), .Z(n7226) );
  MUX2_X1 U6538 ( .A(n9780), .B(n2792), .S(n1705), .Z(n7227) );
  MUX2_X1 U6539 ( .A(n9781), .B(n2781), .S(n1705), .Z(n7228) );
  MUX2_X1 U6540 ( .A(n9782), .B(n2770), .S(n1705), .Z(n7229) );
  MUX2_X1 U6541 ( .A(n9783), .B(n2759), .S(n1705), .Z(n7230) );
  MUX2_X1 U6542 ( .A(n9784), .B(n2748), .S(n1705), .Z(n7231) );
  MUX2_X1 U6543 ( .A(n9785), .B(n2737), .S(n1705), .Z(n7232) );
  MUX2_X1 U6544 ( .A(n9786), .B(n2726), .S(n1705), .Z(n7233) );
  MUX2_X1 U6545 ( .A(n9787), .B(n2715), .S(n1705), .Z(n7234) );
  MUX2_X1 U6546 ( .A(n9788), .B(n2704), .S(n1705), .Z(n7235) );
  MUX2_X1 U6547 ( .A(n9789), .B(n2597), .S(n1705), .Z(n7236) );
  MUX2_X1 U6548 ( .A(n9790), .B(n2586), .S(n1706), .Z(n7237) );
  MUX2_X1 U6549 ( .A(n9791), .B(n2575), .S(n1706), .Z(n7238) );
  MUX2_X1 U6550 ( .A(n9792), .B(n2564), .S(n1706), .Z(n7239) );
  MUX2_X1 U6551 ( .A(n9793), .B(n2553), .S(n1706), .Z(n7240) );
  MUX2_X1 U6552 ( .A(n9794), .B(n1838), .S(n1706), .Z(n7241) );
  MUX2_X1 U6553 ( .A(n9795), .B(n1827), .S(n1706), .Z(n7242) );
  MUX2_X1 U6554 ( .A(n9796), .B(n1816), .S(n1706), .Z(n7243) );
  MUX2_X1 U6555 ( .A(n9797), .B(n1805), .S(n1706), .Z(n7244) );
  MUX2_X1 U6556 ( .A(n9734), .B(n2952), .S(n1707), .Z(n7181) );
  MUX2_X1 U6557 ( .A(n9735), .B(n2941), .S(n1707), .Z(n7182) );
  MUX2_X1 U6558 ( .A(n9736), .B(n2930), .S(n1707), .Z(n7183) );
  MUX2_X1 U6559 ( .A(n9737), .B(n2914), .S(n1707), .Z(n7184) );
  MUX2_X1 U6560 ( .A(n9738), .B(n2903), .S(n1707), .Z(n7185) );
  MUX2_X1 U6561 ( .A(n9739), .B(n2891), .S(n1707), .Z(n7186) );
  MUX2_X1 U6562 ( .A(n9740), .B(n2880), .S(n1707), .Z(n7187) );
  MUX2_X1 U6563 ( .A(n9741), .B(n2869), .S(n1707), .Z(n7188) );
  MUX2_X1 U6564 ( .A(n9742), .B(n2858), .S(n1707), .Z(n7189) );
  MUX2_X1 U6565 ( .A(n9743), .B(n2847), .S(n1707), .Z(n7190) );
  MUX2_X1 U6566 ( .A(n9744), .B(n2836), .S(n1707), .Z(n7191) );
  MUX2_X1 U6567 ( .A(n9745), .B(n2825), .S(n1707), .Z(n7192) );
  MUX2_X1 U6568 ( .A(n9746), .B(n2814), .S(n1708), .Z(n7193) );
  MUX2_X1 U6569 ( .A(n9747), .B(n2803), .S(n1708), .Z(n7194) );
  MUX2_X1 U6570 ( .A(n9748), .B(n2792), .S(n1708), .Z(n7195) );
  MUX2_X1 U6571 ( .A(n9749), .B(n2781), .S(n1708), .Z(n7196) );
  MUX2_X1 U6572 ( .A(n9750), .B(n2770), .S(n1708), .Z(n7197) );
  MUX2_X1 U6573 ( .A(n9751), .B(n2759), .S(n1708), .Z(n7198) );
  MUX2_X1 U6574 ( .A(n9752), .B(n2748), .S(n1708), .Z(n7199) );
  MUX2_X1 U6575 ( .A(n9753), .B(n2737), .S(n1708), .Z(n7200) );
  MUX2_X1 U6576 ( .A(n9754), .B(n2726), .S(n1708), .Z(n7201) );
  MUX2_X1 U6577 ( .A(n9755), .B(n2715), .S(n1708), .Z(n7202) );
  MUX2_X1 U6578 ( .A(n9756), .B(n2704), .S(n1708), .Z(n7203) );
  MUX2_X1 U6579 ( .A(n9757), .B(n2597), .S(n1708), .Z(n7204) );
  MUX2_X1 U6580 ( .A(n9758), .B(n2586), .S(n1709), .Z(n7205) );
  MUX2_X1 U6581 ( .A(n9759), .B(n2575), .S(n1709), .Z(n7206) );
  MUX2_X1 U6582 ( .A(n9760), .B(n2564), .S(n1709), .Z(n7207) );
  MUX2_X1 U6583 ( .A(n9761), .B(n2553), .S(n1709), .Z(n7208) );
  MUX2_X1 U6584 ( .A(n9762), .B(n1838), .S(n1709), .Z(n7209) );
  MUX2_X1 U6585 ( .A(n9763), .B(n1827), .S(n1709), .Z(n7210) );
  MUX2_X1 U6586 ( .A(n9764), .B(n1816), .S(n1709), .Z(n7211) );
  MUX2_X1 U6587 ( .A(n9765), .B(n1805), .S(n1709), .Z(n7212) );
  MUX2_X1 U6588 ( .A(n9702), .B(n2952), .S(n1710), .Z(n7149) );
  MUX2_X1 U6589 ( .A(n9703), .B(n2941), .S(n1710), .Z(n7150) );
  MUX2_X1 U6590 ( .A(n9704), .B(n2930), .S(n1710), .Z(n7151) );
  MUX2_X1 U6591 ( .A(n9705), .B(n2914), .S(n1710), .Z(n7152) );
  MUX2_X1 U6592 ( .A(n9706), .B(n2903), .S(n1710), .Z(n7153) );
  MUX2_X1 U6593 ( .A(n9707), .B(n2891), .S(n1710), .Z(n7154) );
  MUX2_X1 U6594 ( .A(n9708), .B(n2880), .S(n1710), .Z(n7155) );
  MUX2_X1 U6595 ( .A(n9709), .B(n2869), .S(n1710), .Z(n7156) );
  MUX2_X1 U6596 ( .A(n9710), .B(n2858), .S(n1710), .Z(n7157) );
  MUX2_X1 U6597 ( .A(n9711), .B(n2847), .S(n1710), .Z(n7158) );
  MUX2_X1 U6598 ( .A(n9712), .B(n2836), .S(n1710), .Z(n7159) );
  MUX2_X1 U6599 ( .A(n9713), .B(n2825), .S(n1710), .Z(n7160) );
  MUX2_X1 U6600 ( .A(n9714), .B(n2814), .S(n1711), .Z(n7161) );
  MUX2_X1 U6601 ( .A(n9715), .B(n2803), .S(n1711), .Z(n7162) );
  MUX2_X1 U6602 ( .A(n9716), .B(n2792), .S(n1711), .Z(n7163) );
  MUX2_X1 U6603 ( .A(n9717), .B(n2781), .S(n1711), .Z(n7164) );
  MUX2_X1 U6604 ( .A(n9718), .B(n2770), .S(n1711), .Z(n7165) );
  MUX2_X1 U6605 ( .A(n9719), .B(n2759), .S(n1711), .Z(n7166) );
  MUX2_X1 U6606 ( .A(n9720), .B(n2748), .S(n1711), .Z(n7167) );
  MUX2_X1 U6607 ( .A(n9721), .B(n2737), .S(n1711), .Z(n7168) );
  MUX2_X1 U6608 ( .A(n9722), .B(n2726), .S(n1711), .Z(n7169) );
  MUX2_X1 U6609 ( .A(n9723), .B(n2715), .S(n1711), .Z(n7170) );
  MUX2_X1 U6610 ( .A(n9724), .B(n2704), .S(n1711), .Z(n7171) );
  MUX2_X1 U6611 ( .A(n9725), .B(n2597), .S(n1711), .Z(n7172) );
  MUX2_X1 U6612 ( .A(n9726), .B(n2586), .S(n1712), .Z(n7173) );
  MUX2_X1 U6613 ( .A(n9727), .B(n2575), .S(n1712), .Z(n7174) );
  MUX2_X1 U6614 ( .A(n9728), .B(n2564), .S(n1712), .Z(n7175) );
  MUX2_X1 U6615 ( .A(n9729), .B(n2553), .S(n1712), .Z(n7176) );
  MUX2_X1 U6616 ( .A(n9730), .B(n1838), .S(n1712), .Z(n7177) );
  MUX2_X1 U6617 ( .A(n9731), .B(n1827), .S(n1712), .Z(n7178) );
  MUX2_X1 U6618 ( .A(n9732), .B(n1816), .S(n1712), .Z(n7179) );
  MUX2_X1 U6619 ( .A(n9733), .B(n1805), .S(n1712), .Z(n7180) );
  MUX2_X1 U6620 ( .A(n9670), .B(n2952), .S(n1713), .Z(n7117) );
  MUX2_X1 U6621 ( .A(n9671), .B(n2941), .S(n1713), .Z(n7118) );
  MUX2_X1 U6622 ( .A(n9672), .B(n2930), .S(n1713), .Z(n7119) );
  MUX2_X1 U6623 ( .A(n9673), .B(n2914), .S(n1713), .Z(n7120) );
  MUX2_X1 U6624 ( .A(n9674), .B(n2903), .S(n1713), .Z(n7121) );
  MUX2_X1 U6625 ( .A(n9675), .B(n2891), .S(n1713), .Z(n7122) );
  MUX2_X1 U6626 ( .A(n9676), .B(n2880), .S(n1713), .Z(n7123) );
  MUX2_X1 U6627 ( .A(n9677), .B(n2869), .S(n1713), .Z(n7124) );
  MUX2_X1 U6628 ( .A(n9678), .B(n2858), .S(n1713), .Z(n7125) );
  MUX2_X1 U6629 ( .A(n9679), .B(n2847), .S(n1713), .Z(n7126) );
  MUX2_X1 U6630 ( .A(n9680), .B(n2836), .S(n1713), .Z(n7127) );
  MUX2_X1 U6631 ( .A(n9681), .B(n2825), .S(n1713), .Z(n7128) );
  MUX2_X1 U6632 ( .A(n9682), .B(n2814), .S(n1714), .Z(n7129) );
  MUX2_X1 U6633 ( .A(n9683), .B(n2803), .S(n1714), .Z(n7130) );
  MUX2_X1 U6634 ( .A(n9684), .B(n2792), .S(n1714), .Z(n7131) );
  MUX2_X1 U6635 ( .A(n9685), .B(n2781), .S(n1714), .Z(n7132) );
  MUX2_X1 U6636 ( .A(n9686), .B(n2770), .S(n1714), .Z(n7133) );
  MUX2_X1 U6637 ( .A(n9687), .B(n2759), .S(n1714), .Z(n7134) );
  MUX2_X1 U6638 ( .A(n9688), .B(n2748), .S(n1714), .Z(n7135) );
  MUX2_X1 U6639 ( .A(n9689), .B(n2737), .S(n1714), .Z(n7136) );
  MUX2_X1 U6640 ( .A(n9690), .B(n2726), .S(n1714), .Z(n7137) );
  MUX2_X1 U6641 ( .A(n9691), .B(n2715), .S(n1714), .Z(n7138) );
  MUX2_X1 U6642 ( .A(n9692), .B(n2704), .S(n1714), .Z(n7139) );
  MUX2_X1 U6643 ( .A(n9693), .B(n2597), .S(n1714), .Z(n7140) );
  MUX2_X1 U6644 ( .A(n9694), .B(n2586), .S(n1715), .Z(n7141) );
  MUX2_X1 U6645 ( .A(n9695), .B(n2575), .S(n1715), .Z(n7142) );
  MUX2_X1 U6646 ( .A(n9696), .B(n2564), .S(n1715), .Z(n7143) );
  MUX2_X1 U6647 ( .A(n9697), .B(n2553), .S(n1715), .Z(n7144) );
  MUX2_X1 U6648 ( .A(n9698), .B(n1838), .S(n1715), .Z(n7145) );
  MUX2_X1 U6649 ( .A(n9699), .B(n1827), .S(n1715), .Z(n7146) );
  MUX2_X1 U6650 ( .A(n9700), .B(n1816), .S(n1715), .Z(n7147) );
  MUX2_X1 U6651 ( .A(n9701), .B(n1805), .S(n1715), .Z(n7148) );
  MUX2_X1 U6652 ( .A(n9638), .B(n2952), .S(n1716), .Z(n7085) );
  MUX2_X1 U6653 ( .A(n9639), .B(n2941), .S(n1716), .Z(n7086) );
  MUX2_X1 U6654 ( .A(n9640), .B(n2930), .S(n1716), .Z(n7087) );
  MUX2_X1 U6655 ( .A(n9641), .B(n2914), .S(n1716), .Z(n7088) );
  MUX2_X1 U6656 ( .A(n9642), .B(n2903), .S(n1716), .Z(n7089) );
  MUX2_X1 U6657 ( .A(n9643), .B(n2891), .S(n1716), .Z(n7090) );
  MUX2_X1 U6658 ( .A(n9644), .B(n2880), .S(n1716), .Z(n7091) );
  MUX2_X1 U6659 ( .A(n9645), .B(n2869), .S(n1716), .Z(n7092) );
  MUX2_X1 U6660 ( .A(n9646), .B(n2858), .S(n1716), .Z(n7093) );
  MUX2_X1 U6661 ( .A(n9647), .B(n2847), .S(n1716), .Z(n7094) );
  MUX2_X1 U6662 ( .A(n9648), .B(n2836), .S(n1716), .Z(n7095) );
  MUX2_X1 U6663 ( .A(n9649), .B(n2825), .S(n1716), .Z(n7096) );
  MUX2_X1 U6664 ( .A(n9650), .B(n2814), .S(n1717), .Z(n7097) );
  MUX2_X1 U6665 ( .A(n9651), .B(n2803), .S(n1717), .Z(n7098) );
  MUX2_X1 U6666 ( .A(n9652), .B(n2792), .S(n1717), .Z(n7099) );
  MUX2_X1 U6667 ( .A(n9653), .B(n2781), .S(n1717), .Z(n7100) );
  MUX2_X1 U6668 ( .A(n9654), .B(n2770), .S(n1717), .Z(n7101) );
  MUX2_X1 U6669 ( .A(n9655), .B(n2759), .S(n1717), .Z(n7102) );
  MUX2_X1 U6670 ( .A(n9656), .B(n2748), .S(n1717), .Z(n7103) );
  MUX2_X1 U6671 ( .A(n9657), .B(n2737), .S(n1717), .Z(n7104) );
  MUX2_X1 U6672 ( .A(n9658), .B(n2726), .S(n1717), .Z(n7105) );
  MUX2_X1 U6673 ( .A(n9659), .B(n2715), .S(n1717), .Z(n7106) );
  MUX2_X1 U6674 ( .A(n9660), .B(n2704), .S(n1717), .Z(n7107) );
  MUX2_X1 U6675 ( .A(n9661), .B(n2597), .S(n1717), .Z(n7108) );
  MUX2_X1 U6676 ( .A(n9662), .B(n2586), .S(n1718), .Z(n7109) );
  MUX2_X1 U6677 ( .A(n9663), .B(n2575), .S(n1718), .Z(n7110) );
  MUX2_X1 U6678 ( .A(n9664), .B(n2564), .S(n1718), .Z(n7111) );
  MUX2_X1 U6679 ( .A(n9665), .B(n2553), .S(n1718), .Z(n7112) );
  MUX2_X1 U6680 ( .A(n9666), .B(n1838), .S(n1718), .Z(n7113) );
  MUX2_X1 U6681 ( .A(n9667), .B(n1827), .S(n1718), .Z(n7114) );
  MUX2_X1 U6682 ( .A(n9668), .B(n1816), .S(n1718), .Z(n7115) );
  MUX2_X1 U6683 ( .A(n9669), .B(n1805), .S(n1718), .Z(n7116) );
  MUX2_X1 U6684 ( .A(n9606), .B(n2952), .S(n1719), .Z(n7053) );
  MUX2_X1 U6685 ( .A(n9607), .B(n2941), .S(n1719), .Z(n7054) );
  MUX2_X1 U6686 ( .A(n9608), .B(n2930), .S(n1719), .Z(n7055) );
  MUX2_X1 U6687 ( .A(n9609), .B(n2914), .S(n1719), .Z(n7056) );
  MUX2_X1 U6688 ( .A(n9610), .B(n2903), .S(n1719), .Z(n7057) );
  MUX2_X1 U6689 ( .A(n9611), .B(n2891), .S(n1719), .Z(n7058) );
  MUX2_X1 U6690 ( .A(n9612), .B(n2880), .S(n1719), .Z(n7059) );
  MUX2_X1 U6691 ( .A(n9613), .B(n2869), .S(n1719), .Z(n7060) );
  MUX2_X1 U6692 ( .A(n9614), .B(n2858), .S(n1719), .Z(n7061) );
  MUX2_X1 U6693 ( .A(n9615), .B(n2847), .S(n1719), .Z(n7062) );
  MUX2_X1 U6694 ( .A(n9616), .B(n2836), .S(n1719), .Z(n7063) );
  MUX2_X1 U6695 ( .A(n9617), .B(n2825), .S(n1719), .Z(n7064) );
  MUX2_X1 U6696 ( .A(n9618), .B(n2814), .S(n1720), .Z(n7065) );
  MUX2_X1 U6697 ( .A(n9619), .B(n2803), .S(n1720), .Z(n7066) );
  MUX2_X1 U6698 ( .A(n9620), .B(n2792), .S(n1720), .Z(n7067) );
  MUX2_X1 U6699 ( .A(n9621), .B(n2781), .S(n1720), .Z(n7068) );
  MUX2_X1 U6700 ( .A(n9622), .B(n2770), .S(n1720), .Z(n7069) );
  MUX2_X1 U6701 ( .A(n9623), .B(n2759), .S(n1720), .Z(n7070) );
  MUX2_X1 U6702 ( .A(n9624), .B(n2748), .S(n1720), .Z(n7071) );
  MUX2_X1 U6703 ( .A(n9625), .B(n2737), .S(n1720), .Z(n7072) );
  MUX2_X1 U6704 ( .A(n9626), .B(n2726), .S(n1720), .Z(n7073) );
  MUX2_X1 U6705 ( .A(n9627), .B(n2715), .S(n1720), .Z(n7074) );
  MUX2_X1 U6706 ( .A(n9628), .B(n2704), .S(n1720), .Z(n7075) );
  MUX2_X1 U6707 ( .A(n9629), .B(n2597), .S(n1720), .Z(n7076) );
  MUX2_X1 U6708 ( .A(n9630), .B(n2586), .S(n1721), .Z(n7077) );
  MUX2_X1 U6709 ( .A(n9631), .B(n2575), .S(n1721), .Z(n7078) );
  MUX2_X1 U6710 ( .A(n9632), .B(n2564), .S(n1721), .Z(n7079) );
  MUX2_X1 U6711 ( .A(n9633), .B(n2553), .S(n1721), .Z(n7080) );
  MUX2_X1 U6712 ( .A(n9634), .B(n1838), .S(n1721), .Z(n7081) );
  MUX2_X1 U6713 ( .A(n9635), .B(n1827), .S(n1721), .Z(n7082) );
  MUX2_X1 U6714 ( .A(n9636), .B(n1816), .S(n1721), .Z(n7083) );
  MUX2_X1 U6715 ( .A(n9637), .B(n1805), .S(n1721), .Z(n7084) );
  MUX2_X1 U6716 ( .A(n9574), .B(n2952), .S(n1722), .Z(n7021) );
  MUX2_X1 U6717 ( .A(n9575), .B(n2941), .S(n1722), .Z(n7022) );
  MUX2_X1 U6718 ( .A(n9576), .B(n2930), .S(n1722), .Z(n7023) );
  MUX2_X1 U6719 ( .A(n9577), .B(n2914), .S(n1722), .Z(n7024) );
  MUX2_X1 U6720 ( .A(n9578), .B(n2903), .S(n1722), .Z(n7025) );
  MUX2_X1 U6721 ( .A(n9579), .B(n2891), .S(n1722), .Z(n7026) );
  MUX2_X1 U6722 ( .A(n9580), .B(n2880), .S(n1722), .Z(n7027) );
  MUX2_X1 U6723 ( .A(n9581), .B(n2869), .S(n1722), .Z(n7028) );
  MUX2_X1 U6724 ( .A(n9582), .B(n2858), .S(n1722), .Z(n7029) );
  MUX2_X1 U6725 ( .A(n9583), .B(n2847), .S(n1722), .Z(n7030) );
  MUX2_X1 U6726 ( .A(n9584), .B(n2836), .S(n1722), .Z(n7031) );
  MUX2_X1 U6727 ( .A(n9585), .B(n2825), .S(n1722), .Z(n7032) );
  MUX2_X1 U6728 ( .A(n9586), .B(n2814), .S(n1723), .Z(n7033) );
  MUX2_X1 U6729 ( .A(n9587), .B(n2803), .S(n1723), .Z(n7034) );
  MUX2_X1 U6730 ( .A(n9588), .B(n2792), .S(n1723), .Z(n7035) );
  MUX2_X1 U6731 ( .A(n9589), .B(n2781), .S(n1723), .Z(n7036) );
  MUX2_X1 U6732 ( .A(n9590), .B(n2770), .S(n1723), .Z(n7037) );
  MUX2_X1 U6733 ( .A(n9591), .B(n2759), .S(n1723), .Z(n7038) );
  MUX2_X1 U6734 ( .A(n9592), .B(n2748), .S(n1723), .Z(n7039) );
  MUX2_X1 U6735 ( .A(n9593), .B(n2737), .S(n1723), .Z(n7040) );
  MUX2_X1 U6736 ( .A(n9594), .B(n2726), .S(n1723), .Z(n7041) );
  MUX2_X1 U6737 ( .A(n9595), .B(n2715), .S(n1723), .Z(n7042) );
  MUX2_X1 U6738 ( .A(n9596), .B(n2704), .S(n1723), .Z(n7043) );
  MUX2_X1 U6739 ( .A(n9597), .B(n2597), .S(n1723), .Z(n7044) );
  MUX2_X1 U6740 ( .A(n9598), .B(n2586), .S(n1724), .Z(n7045) );
  MUX2_X1 U6741 ( .A(n9599), .B(n2575), .S(n1724), .Z(n7046) );
  MUX2_X1 U6742 ( .A(n9600), .B(n2564), .S(n1724), .Z(n7047) );
  MUX2_X1 U6743 ( .A(n9601), .B(n2553), .S(n1724), .Z(n7048) );
  MUX2_X1 U6744 ( .A(n9602), .B(n1838), .S(n1724), .Z(n7049) );
  MUX2_X1 U6745 ( .A(n9603), .B(n1827), .S(n1724), .Z(n7050) );
  MUX2_X1 U6746 ( .A(n9604), .B(n1816), .S(n1724), .Z(n7051) );
  MUX2_X1 U6747 ( .A(n9605), .B(n1805), .S(n1724), .Z(n7052) );
  MUX2_X1 U6748 ( .A(\REGISTERS[21][31] ), .B(n2953), .S(n1725), .Z(n6989) );
  MUX2_X1 U6749 ( .A(\REGISTERS[21][30] ), .B(n2942), .S(n1725), .Z(n6990) );
  MUX2_X1 U6750 ( .A(\REGISTERS[21][29] ), .B(n2931), .S(n1725), .Z(n6991) );
  MUX2_X1 U6751 ( .A(\REGISTERS[21][28] ), .B(n2915), .S(n1725), .Z(n6992) );
  MUX2_X1 U6752 ( .A(\REGISTERS[21][27] ), .B(n2904), .S(n1725), .Z(n6993) );
  MUX2_X1 U6753 ( .A(\REGISTERS[21][26] ), .B(n2892), .S(n1725), .Z(n6994) );
  MUX2_X1 U6754 ( .A(\REGISTERS[21][25] ), .B(n2881), .S(n1725), .Z(n6995) );
  MUX2_X1 U6755 ( .A(\REGISTERS[21][24] ), .B(n2870), .S(n1725), .Z(n6996) );
  MUX2_X1 U6756 ( .A(\REGISTERS[21][23] ), .B(n2859), .S(n1725), .Z(n6997) );
  MUX2_X1 U6757 ( .A(\REGISTERS[21][22] ), .B(n2848), .S(n1725), .Z(n6998) );
  MUX2_X1 U6758 ( .A(\REGISTERS[21][21] ), .B(n2837), .S(n1725), .Z(n6999) );
  MUX2_X1 U6759 ( .A(\REGISTERS[21][20] ), .B(n2826), .S(n1725), .Z(n7000) );
  MUX2_X1 U6760 ( .A(\REGISTERS[21][19] ), .B(n2815), .S(n1726), .Z(n7001) );
  MUX2_X1 U6761 ( .A(\REGISTERS[21][18] ), .B(n2804), .S(n1726), .Z(n7002) );
  MUX2_X1 U6762 ( .A(\REGISTERS[21][17] ), .B(n2793), .S(n1726), .Z(n7003) );
  MUX2_X1 U6763 ( .A(\REGISTERS[21][16] ), .B(n2782), .S(n1726), .Z(n7004) );
  MUX2_X1 U6764 ( .A(\REGISTERS[21][15] ), .B(n2771), .S(n1726), .Z(n7005) );
  MUX2_X1 U6765 ( .A(\REGISTERS[21][14] ), .B(n2760), .S(n1726), .Z(n7006) );
  MUX2_X1 U6766 ( .A(\REGISTERS[21][13] ), .B(n2749), .S(n1726), .Z(n7007) );
  MUX2_X1 U6767 ( .A(\REGISTERS[21][12] ), .B(n2738), .S(n1726), .Z(n7008) );
  MUX2_X1 U6768 ( .A(\REGISTERS[21][11] ), .B(n2727), .S(n1726), .Z(n7009) );
  MUX2_X1 U6769 ( .A(\REGISTERS[21][10] ), .B(n2716), .S(n1726), .Z(n7010) );
  MUX2_X1 U6770 ( .A(\REGISTERS[21][9] ), .B(n2705), .S(n1726), .Z(n7011) );
  MUX2_X1 U6771 ( .A(\REGISTERS[21][8] ), .B(n2598), .S(n1726), .Z(n7012) );
  MUX2_X1 U6772 ( .A(\REGISTERS[21][7] ), .B(n2587), .S(n1727), .Z(n7013) );
  MUX2_X1 U6773 ( .A(\REGISTERS[21][6] ), .B(n2576), .S(n1727), .Z(n7014) );
  MUX2_X1 U6774 ( .A(\REGISTERS[21][5] ), .B(n2565), .S(n1727), .Z(n7015) );
  MUX2_X1 U6775 ( .A(\REGISTERS[21][4] ), .B(n2554), .S(n1727), .Z(n7016) );
  MUX2_X1 U6776 ( .A(\REGISTERS[21][3] ), .B(n1839), .S(n1727), .Z(n7017) );
  MUX2_X1 U6777 ( .A(\REGISTERS[21][2] ), .B(n1828), .S(n1727), .Z(n7018) );
  MUX2_X1 U6778 ( .A(\REGISTERS[21][1] ), .B(n1817), .S(n1727), .Z(n7019) );
  MUX2_X1 U6779 ( .A(\REGISTERS[21][0] ), .B(n1806), .S(n1727), .Z(n7020) );
  MUX2_X1 U6780 ( .A(\REGISTERS[20][31] ), .B(n2953), .S(n1728), .Z(n6957) );
  MUX2_X1 U6781 ( .A(\REGISTERS[20][30] ), .B(n2942), .S(n1728), .Z(n6958) );
  MUX2_X1 U6782 ( .A(\REGISTERS[20][29] ), .B(n2931), .S(n1728), .Z(n6959) );
  MUX2_X1 U6783 ( .A(\REGISTERS[20][28] ), .B(n2915), .S(n1728), .Z(n6960) );
  MUX2_X1 U6784 ( .A(\REGISTERS[20][27] ), .B(n2904), .S(n1728), .Z(n6961) );
  MUX2_X1 U6785 ( .A(\REGISTERS[20][26] ), .B(n2892), .S(n1728), .Z(n6962) );
  MUX2_X1 U6786 ( .A(\REGISTERS[20][25] ), .B(n2881), .S(n1728), .Z(n6963) );
  MUX2_X1 U6787 ( .A(\REGISTERS[20][24] ), .B(n2870), .S(n1728), .Z(n6964) );
  MUX2_X1 U6788 ( .A(\REGISTERS[20][23] ), .B(n2859), .S(n1728), .Z(n6965) );
  MUX2_X1 U6789 ( .A(\REGISTERS[20][22] ), .B(n2848), .S(n1728), .Z(n6966) );
  MUX2_X1 U6790 ( .A(\REGISTERS[20][21] ), .B(n2837), .S(n1728), .Z(n6967) );
  MUX2_X1 U6791 ( .A(\REGISTERS[20][20] ), .B(n2826), .S(n1728), .Z(n6968) );
  MUX2_X1 U6792 ( .A(\REGISTERS[20][19] ), .B(n2815), .S(n1729), .Z(n6969) );
  MUX2_X1 U6793 ( .A(\REGISTERS[20][18] ), .B(n2804), .S(n1729), .Z(n6970) );
  MUX2_X1 U6794 ( .A(\REGISTERS[20][17] ), .B(n2793), .S(n1729), .Z(n6971) );
  MUX2_X1 U6795 ( .A(\REGISTERS[20][16] ), .B(n2782), .S(n1729), .Z(n6972) );
  MUX2_X1 U6796 ( .A(\REGISTERS[20][15] ), .B(n2771), .S(n1729), .Z(n6973) );
  MUX2_X1 U6797 ( .A(\REGISTERS[20][14] ), .B(n2760), .S(n1729), .Z(n6974) );
  MUX2_X1 U6798 ( .A(\REGISTERS[20][13] ), .B(n2749), .S(n1729), .Z(n6975) );
  MUX2_X1 U6799 ( .A(\REGISTERS[20][12] ), .B(n2738), .S(n1729), .Z(n6976) );
  MUX2_X1 U6800 ( .A(\REGISTERS[20][11] ), .B(n2727), .S(n1729), .Z(n6977) );
  MUX2_X1 U6801 ( .A(\REGISTERS[20][10] ), .B(n2716), .S(n1729), .Z(n6978) );
  MUX2_X1 U6802 ( .A(\REGISTERS[20][9] ), .B(n2705), .S(n1729), .Z(n6979) );
  MUX2_X1 U6803 ( .A(\REGISTERS[20][8] ), .B(n2598), .S(n1729), .Z(n6980) );
  MUX2_X1 U6804 ( .A(\REGISTERS[20][7] ), .B(n2587), .S(n1730), .Z(n6981) );
  MUX2_X1 U6805 ( .A(\REGISTERS[20][6] ), .B(n2576), .S(n1730), .Z(n6982) );
  MUX2_X1 U6806 ( .A(\REGISTERS[20][5] ), .B(n2565), .S(n1730), .Z(n6983) );
  MUX2_X1 U6807 ( .A(\REGISTERS[20][4] ), .B(n2554), .S(n1730), .Z(n6984) );
  MUX2_X1 U6808 ( .A(\REGISTERS[20][3] ), .B(n1839), .S(n1730), .Z(n6985) );
  MUX2_X1 U6809 ( .A(\REGISTERS[20][2] ), .B(n1828), .S(n1730), .Z(n6986) );
  MUX2_X1 U6810 ( .A(\REGISTERS[20][1] ), .B(n1817), .S(n1730), .Z(n6987) );
  MUX2_X1 U6811 ( .A(\REGISTERS[20][0] ), .B(n1806), .S(n1730), .Z(n6988) );
  MUX2_X1 U6812 ( .A(\REGISTERS[19][31] ), .B(n2953), .S(n1731), .Z(n6925) );
  MUX2_X1 U6813 ( .A(\REGISTERS[19][30] ), .B(n2942), .S(n1731), .Z(n6926) );
  MUX2_X1 U6814 ( .A(\REGISTERS[19][29] ), .B(n2931), .S(n1731), .Z(n6927) );
  MUX2_X1 U6815 ( .A(\REGISTERS[19][28] ), .B(n2915), .S(n1731), .Z(n6928) );
  MUX2_X1 U6816 ( .A(\REGISTERS[19][27] ), .B(n2904), .S(n1731), .Z(n6929) );
  MUX2_X1 U6817 ( .A(\REGISTERS[19][26] ), .B(n2892), .S(n1731), .Z(n6930) );
  MUX2_X1 U6818 ( .A(\REGISTERS[19][25] ), .B(n2881), .S(n1731), .Z(n6931) );
  MUX2_X1 U6819 ( .A(\REGISTERS[19][24] ), .B(n2870), .S(n1731), .Z(n6932) );
  MUX2_X1 U6820 ( .A(\REGISTERS[19][23] ), .B(n2859), .S(n1731), .Z(n6933) );
  MUX2_X1 U6821 ( .A(\REGISTERS[19][22] ), .B(n2848), .S(n1731), .Z(n6934) );
  MUX2_X1 U6822 ( .A(\REGISTERS[19][21] ), .B(n2837), .S(n1731), .Z(n6935) );
  MUX2_X1 U6823 ( .A(\REGISTERS[19][20] ), .B(n2826), .S(n1731), .Z(n6936) );
  MUX2_X1 U6824 ( .A(\REGISTERS[19][19] ), .B(n2815), .S(n1732), .Z(n6937) );
  MUX2_X1 U6825 ( .A(\REGISTERS[19][18] ), .B(n2804), .S(n1732), .Z(n6938) );
  MUX2_X1 U6826 ( .A(\REGISTERS[19][17] ), .B(n2793), .S(n1732), .Z(n6939) );
  MUX2_X1 U6827 ( .A(\REGISTERS[19][16] ), .B(n2782), .S(n1732), .Z(n6940) );
  MUX2_X1 U6828 ( .A(\REGISTERS[19][15] ), .B(n2771), .S(n1732), .Z(n6941) );
  MUX2_X1 U6829 ( .A(\REGISTERS[19][14] ), .B(n2760), .S(n1732), .Z(n6942) );
  MUX2_X1 U6830 ( .A(\REGISTERS[19][13] ), .B(n2749), .S(n1732), .Z(n6943) );
  MUX2_X1 U6831 ( .A(\REGISTERS[19][12] ), .B(n2738), .S(n1732), .Z(n6944) );
  MUX2_X1 U6832 ( .A(\REGISTERS[19][11] ), .B(n2727), .S(n1732), .Z(n6945) );
  MUX2_X1 U6833 ( .A(\REGISTERS[19][10] ), .B(n2716), .S(n1732), .Z(n6946) );
  MUX2_X1 U6834 ( .A(\REGISTERS[19][9] ), .B(n2705), .S(n1732), .Z(n6947) );
  MUX2_X1 U6835 ( .A(\REGISTERS[19][8] ), .B(n2598), .S(n1732), .Z(n6948) );
  MUX2_X1 U6836 ( .A(\REGISTERS[19][7] ), .B(n2587), .S(n1733), .Z(n6949) );
  MUX2_X1 U6837 ( .A(\REGISTERS[19][6] ), .B(n2576), .S(n1733), .Z(n6950) );
  MUX2_X1 U6838 ( .A(\REGISTERS[19][5] ), .B(n2565), .S(n1733), .Z(n6951) );
  MUX2_X1 U6839 ( .A(\REGISTERS[19][4] ), .B(n2554), .S(n1733), .Z(n6952) );
  MUX2_X1 U6840 ( .A(\REGISTERS[19][3] ), .B(n1839), .S(n1733), .Z(n6953) );
  MUX2_X1 U6841 ( .A(\REGISTERS[19][2] ), .B(n1828), .S(n1733), .Z(n6954) );
  MUX2_X1 U6842 ( .A(\REGISTERS[19][1] ), .B(n1817), .S(n1733), .Z(n6955) );
  MUX2_X1 U6843 ( .A(\REGISTERS[19][0] ), .B(n1806), .S(n1733), .Z(n6956) );
  MUX2_X1 U6844 ( .A(\REGISTERS[18][31] ), .B(n2953), .S(n1734), .Z(n6893) );
  MUX2_X1 U6845 ( .A(\REGISTERS[18][30] ), .B(n2942), .S(n1734), .Z(n6894) );
  MUX2_X1 U6846 ( .A(\REGISTERS[18][29] ), .B(n2931), .S(n1734), .Z(n6895) );
  MUX2_X1 U6847 ( .A(\REGISTERS[18][28] ), .B(n2915), .S(n1734), .Z(n6896) );
  MUX2_X1 U6848 ( .A(\REGISTERS[18][27] ), .B(n2904), .S(n1734), .Z(n6897) );
  MUX2_X1 U6849 ( .A(\REGISTERS[18][26] ), .B(n2892), .S(n1734), .Z(n6898) );
  MUX2_X1 U6850 ( .A(\REGISTERS[18][25] ), .B(n2881), .S(n1734), .Z(n6899) );
  MUX2_X1 U6851 ( .A(\REGISTERS[18][24] ), .B(n2870), .S(n1734), .Z(n6900) );
  MUX2_X1 U6852 ( .A(\REGISTERS[18][23] ), .B(n2859), .S(n1734), .Z(n6901) );
  MUX2_X1 U6853 ( .A(\REGISTERS[18][22] ), .B(n2848), .S(n1734), .Z(n6902) );
  MUX2_X1 U6854 ( .A(\REGISTERS[18][21] ), .B(n2837), .S(n1734), .Z(n6903) );
  MUX2_X1 U6855 ( .A(\REGISTERS[18][20] ), .B(n2826), .S(n1734), .Z(n6904) );
  MUX2_X1 U6856 ( .A(\REGISTERS[18][19] ), .B(n2815), .S(n1735), .Z(n6905) );
  MUX2_X1 U6857 ( .A(\REGISTERS[18][18] ), .B(n2804), .S(n1735), .Z(n6906) );
  MUX2_X1 U6858 ( .A(\REGISTERS[18][17] ), .B(n2793), .S(n1735), .Z(n6907) );
  MUX2_X1 U6859 ( .A(\REGISTERS[18][16] ), .B(n2782), .S(n1735), .Z(n6908) );
  MUX2_X1 U6860 ( .A(\REGISTERS[18][15] ), .B(n2771), .S(n1735), .Z(n6909) );
  MUX2_X1 U6861 ( .A(\REGISTERS[18][14] ), .B(n2760), .S(n1735), .Z(n6910) );
  MUX2_X1 U6862 ( .A(\REGISTERS[18][13] ), .B(n2749), .S(n1735), .Z(n6911) );
  MUX2_X1 U6863 ( .A(\REGISTERS[18][12] ), .B(n2738), .S(n1735), .Z(n6912) );
  MUX2_X1 U6864 ( .A(\REGISTERS[18][11] ), .B(n2727), .S(n1735), .Z(n6913) );
  MUX2_X1 U6865 ( .A(\REGISTERS[18][10] ), .B(n2716), .S(n1735), .Z(n6914) );
  MUX2_X1 U6866 ( .A(\REGISTERS[18][9] ), .B(n2705), .S(n1735), .Z(n6915) );
  MUX2_X1 U6867 ( .A(\REGISTERS[18][8] ), .B(n2598), .S(n1735), .Z(n6916) );
  MUX2_X1 U6868 ( .A(\REGISTERS[18][7] ), .B(n2587), .S(n1736), .Z(n6917) );
  MUX2_X1 U6869 ( .A(\REGISTERS[18][6] ), .B(n2576), .S(n1736), .Z(n6918) );
  MUX2_X1 U6870 ( .A(\REGISTERS[18][5] ), .B(n2565), .S(n1736), .Z(n6919) );
  MUX2_X1 U6871 ( .A(\REGISTERS[18][4] ), .B(n2554), .S(n1736), .Z(n6920) );
  MUX2_X1 U6872 ( .A(\REGISTERS[18][3] ), .B(n1839), .S(n1736), .Z(n6921) );
  MUX2_X1 U6873 ( .A(\REGISTERS[18][2] ), .B(n1828), .S(n1736), .Z(n6922) );
  MUX2_X1 U6874 ( .A(\REGISTERS[18][1] ), .B(n1817), .S(n1736), .Z(n6923) );
  MUX2_X1 U6875 ( .A(\REGISTERS[18][0] ), .B(n1806), .S(n1736), .Z(n6924) );
  MUX2_X1 U6876 ( .A(\REGISTERS[17][31] ), .B(n2953), .S(n1737), .Z(n6861) );
  MUX2_X1 U6877 ( .A(\REGISTERS[17][30] ), .B(n2942), .S(n1737), .Z(n6862) );
  MUX2_X1 U6878 ( .A(\REGISTERS[17][29] ), .B(n2931), .S(n1737), .Z(n6863) );
  MUX2_X1 U6879 ( .A(\REGISTERS[17][28] ), .B(n2915), .S(n1737), .Z(n6864) );
  MUX2_X1 U6880 ( .A(\REGISTERS[17][27] ), .B(n2904), .S(n1737), .Z(n6865) );
  MUX2_X1 U6881 ( .A(\REGISTERS[17][26] ), .B(n2892), .S(n1737), .Z(n6866) );
  MUX2_X1 U6882 ( .A(\REGISTERS[17][25] ), .B(n2881), .S(n1737), .Z(n6867) );
  MUX2_X1 U6883 ( .A(\REGISTERS[17][24] ), .B(n2870), .S(n1737), .Z(n6868) );
  MUX2_X1 U6884 ( .A(\REGISTERS[17][23] ), .B(n2859), .S(n1737), .Z(n6869) );
  MUX2_X1 U6885 ( .A(\REGISTERS[17][22] ), .B(n2848), .S(n1737), .Z(n6870) );
  MUX2_X1 U6886 ( .A(\REGISTERS[17][21] ), .B(n2837), .S(n1737), .Z(n6871) );
  MUX2_X1 U6887 ( .A(\REGISTERS[17][20] ), .B(n2826), .S(n1737), .Z(n6872) );
  MUX2_X1 U6888 ( .A(\REGISTERS[17][19] ), .B(n2815), .S(n1738), .Z(n6873) );
  MUX2_X1 U6889 ( .A(\REGISTERS[17][18] ), .B(n2804), .S(n1738), .Z(n6874) );
  MUX2_X1 U6890 ( .A(\REGISTERS[17][17] ), .B(n2793), .S(n1738), .Z(n6875) );
  MUX2_X1 U6891 ( .A(\REGISTERS[17][16] ), .B(n2782), .S(n1738), .Z(n6876) );
  MUX2_X1 U6892 ( .A(\REGISTERS[17][15] ), .B(n2771), .S(n1738), .Z(n6877) );
  MUX2_X1 U6893 ( .A(\REGISTERS[17][14] ), .B(n2760), .S(n1738), .Z(n6878) );
  MUX2_X1 U6894 ( .A(\REGISTERS[17][13] ), .B(n2749), .S(n1738), .Z(n6879) );
  MUX2_X1 U6895 ( .A(\REGISTERS[17][12] ), .B(n2738), .S(n1738), .Z(n6880) );
  MUX2_X1 U6896 ( .A(\REGISTERS[17][11] ), .B(n2727), .S(n1738), .Z(n6881) );
  MUX2_X1 U6897 ( .A(\REGISTERS[17][10] ), .B(n2716), .S(n1738), .Z(n6882) );
  MUX2_X1 U6898 ( .A(\REGISTERS[17][9] ), .B(n2705), .S(n1738), .Z(n6883) );
  MUX2_X1 U6899 ( .A(\REGISTERS[17][8] ), .B(n2598), .S(n1738), .Z(n6884) );
  MUX2_X1 U6900 ( .A(\REGISTERS[17][7] ), .B(n2587), .S(n1739), .Z(n6885) );
  MUX2_X1 U6901 ( .A(\REGISTERS[17][6] ), .B(n2576), .S(n1739), .Z(n6886) );
  MUX2_X1 U6902 ( .A(\REGISTERS[17][5] ), .B(n2565), .S(n1739), .Z(n6887) );
  MUX2_X1 U6903 ( .A(\REGISTERS[17][4] ), .B(n2554), .S(n1739), .Z(n6888) );
  MUX2_X1 U6904 ( .A(\REGISTERS[17][3] ), .B(n1839), .S(n1739), .Z(n6889) );
  MUX2_X1 U6905 ( .A(\REGISTERS[17][2] ), .B(n1828), .S(n1739), .Z(n6890) );
  MUX2_X1 U6906 ( .A(\REGISTERS[17][1] ), .B(n1817), .S(n1739), .Z(n6891) );
  MUX2_X1 U6907 ( .A(\REGISTERS[17][0] ), .B(n1806), .S(n1739), .Z(n6892) );
  MUX2_X1 U6908 ( .A(\REGISTERS[16][31] ), .B(n2953), .S(n1740), .Z(n6829) );
  MUX2_X1 U6909 ( .A(\REGISTERS[16][30] ), .B(n2942), .S(n1740), .Z(n6830) );
  MUX2_X1 U6910 ( .A(\REGISTERS[16][29] ), .B(n2931), .S(n1740), .Z(n6831) );
  MUX2_X1 U6911 ( .A(\REGISTERS[16][28] ), .B(n2915), .S(n1740), .Z(n6832) );
  MUX2_X1 U6912 ( .A(\REGISTERS[16][27] ), .B(n2904), .S(n1740), .Z(n6833) );
  MUX2_X1 U6913 ( .A(\REGISTERS[16][26] ), .B(n2892), .S(n1740), .Z(n6834) );
  MUX2_X1 U6914 ( .A(\REGISTERS[16][25] ), .B(n2881), .S(n1740), .Z(n6835) );
  MUX2_X1 U6915 ( .A(\REGISTERS[16][24] ), .B(n2870), .S(n1740), .Z(n6836) );
  MUX2_X1 U6916 ( .A(\REGISTERS[16][23] ), .B(n2859), .S(n1740), .Z(n6837) );
  MUX2_X1 U6917 ( .A(\REGISTERS[16][22] ), .B(n2848), .S(n1740), .Z(n6838) );
  MUX2_X1 U6918 ( .A(\REGISTERS[16][21] ), .B(n2837), .S(n1740), .Z(n6839) );
  MUX2_X1 U6919 ( .A(\REGISTERS[16][20] ), .B(n2826), .S(n1740), .Z(n6840) );
  MUX2_X1 U6920 ( .A(\REGISTERS[16][19] ), .B(n2815), .S(n1741), .Z(n6841) );
  MUX2_X1 U6921 ( .A(\REGISTERS[16][18] ), .B(n2804), .S(n1741), .Z(n6842) );
  MUX2_X1 U6922 ( .A(\REGISTERS[16][17] ), .B(n2793), .S(n1741), .Z(n6843) );
  MUX2_X1 U6923 ( .A(\REGISTERS[16][16] ), .B(n2782), .S(n1741), .Z(n6844) );
  MUX2_X1 U6924 ( .A(\REGISTERS[16][15] ), .B(n2771), .S(n1741), .Z(n6845) );
  MUX2_X1 U6925 ( .A(\REGISTERS[16][14] ), .B(n2760), .S(n1741), .Z(n6846) );
  MUX2_X1 U6926 ( .A(\REGISTERS[16][13] ), .B(n2749), .S(n1741), .Z(n6847) );
  MUX2_X1 U6927 ( .A(\REGISTERS[16][12] ), .B(n2738), .S(n1741), .Z(n6848) );
  MUX2_X1 U6928 ( .A(\REGISTERS[16][11] ), .B(n2727), .S(n1741), .Z(n6849) );
  MUX2_X1 U6929 ( .A(\REGISTERS[16][10] ), .B(n2716), .S(n1741), .Z(n6850) );
  MUX2_X1 U6930 ( .A(\REGISTERS[16][9] ), .B(n2705), .S(n1741), .Z(n6851) );
  MUX2_X1 U6931 ( .A(\REGISTERS[16][8] ), .B(n2598), .S(n1741), .Z(n6852) );
  MUX2_X1 U6932 ( .A(\REGISTERS[16][7] ), .B(n2587), .S(n1742), .Z(n6853) );
  MUX2_X1 U6933 ( .A(\REGISTERS[16][6] ), .B(n2576), .S(n1742), .Z(n6854) );
  MUX2_X1 U6934 ( .A(\REGISTERS[16][5] ), .B(n2565), .S(n1742), .Z(n6855) );
  MUX2_X1 U6935 ( .A(\REGISTERS[16][4] ), .B(n2554), .S(n1742), .Z(n6856) );
  MUX2_X1 U6936 ( .A(\REGISTERS[16][3] ), .B(n1839), .S(n1742), .Z(n6857) );
  MUX2_X1 U6937 ( .A(\REGISTERS[16][2] ), .B(n1828), .S(n1742), .Z(n6858) );
  MUX2_X1 U6938 ( .A(\REGISTERS[16][1] ), .B(n1817), .S(n1742), .Z(n6859) );
  MUX2_X1 U6939 ( .A(\REGISTERS[16][0] ), .B(n1806), .S(n1742), .Z(n6860) );
  MUX2_X1 U6940 ( .A(n9542), .B(n2953), .S(n1743), .Z(n6797) );
  MUX2_X1 U6941 ( .A(n9543), .B(n2942), .S(n1743), .Z(n6798) );
  MUX2_X1 U6942 ( .A(n9544), .B(n2931), .S(n1743), .Z(n6799) );
  MUX2_X1 U6943 ( .A(n9545), .B(n2915), .S(n1743), .Z(n6800) );
  MUX2_X1 U6944 ( .A(n9546), .B(n2904), .S(n1743), .Z(n6801) );
  MUX2_X1 U6945 ( .A(n9547), .B(n2892), .S(n1743), .Z(n6802) );
  MUX2_X1 U6946 ( .A(n9548), .B(n2881), .S(n1743), .Z(n6803) );
  MUX2_X1 U6947 ( .A(n9549), .B(n2870), .S(n1743), .Z(n6804) );
  MUX2_X1 U6948 ( .A(n9550), .B(n2859), .S(n1743), .Z(n6805) );
  MUX2_X1 U6949 ( .A(n9551), .B(n2848), .S(n1743), .Z(n6806) );
  MUX2_X1 U6950 ( .A(n9552), .B(n2837), .S(n1743), .Z(n6807) );
  MUX2_X1 U6951 ( .A(n9553), .B(n2826), .S(n1743), .Z(n6808) );
  MUX2_X1 U6952 ( .A(n9554), .B(n2815), .S(n1744), .Z(n6809) );
  MUX2_X1 U6953 ( .A(n9555), .B(n2804), .S(n1744), .Z(n6810) );
  MUX2_X1 U6954 ( .A(n9556), .B(n2793), .S(n1744), .Z(n6811) );
  MUX2_X1 U6955 ( .A(n9557), .B(n2782), .S(n1744), .Z(n6812) );
  MUX2_X1 U6956 ( .A(n9558), .B(n2771), .S(n1744), .Z(n6813) );
  MUX2_X1 U6957 ( .A(n9559), .B(n2760), .S(n1744), .Z(n6814) );
  MUX2_X1 U6958 ( .A(n9560), .B(n2749), .S(n1744), .Z(n6815) );
  MUX2_X1 U6959 ( .A(n9561), .B(n2738), .S(n1744), .Z(n6816) );
  MUX2_X1 U6960 ( .A(n9562), .B(n2727), .S(n1744), .Z(n6817) );
  MUX2_X1 U6961 ( .A(n9563), .B(n2716), .S(n1744), .Z(n6818) );
  MUX2_X1 U6962 ( .A(n9564), .B(n2705), .S(n1744), .Z(n6819) );
  MUX2_X1 U6963 ( .A(n9565), .B(n2598), .S(n1744), .Z(n6820) );
  MUX2_X1 U6964 ( .A(n9566), .B(n2587), .S(n1745), .Z(n6821) );
  MUX2_X1 U6965 ( .A(n9567), .B(n2576), .S(n1745), .Z(n6822) );
  MUX2_X1 U6966 ( .A(n9568), .B(n2565), .S(n1745), .Z(n6823) );
  MUX2_X1 U6967 ( .A(n9569), .B(n2554), .S(n1745), .Z(n6824) );
  MUX2_X1 U6968 ( .A(n9570), .B(n1839), .S(n1745), .Z(n6825) );
  MUX2_X1 U6969 ( .A(n9571), .B(n1828), .S(n1745), .Z(n6826) );
  MUX2_X1 U6970 ( .A(n9572), .B(n1817), .S(n1745), .Z(n6827) );
  MUX2_X1 U6971 ( .A(n9573), .B(n1806), .S(n1745), .Z(n6828) );
  MUX2_X1 U6972 ( .A(n9510), .B(n2953), .S(n1746), .Z(n6765) );
  MUX2_X1 U6973 ( .A(n9511), .B(n2942), .S(n1746), .Z(n6766) );
  MUX2_X1 U6974 ( .A(n9512), .B(n2931), .S(n1746), .Z(n6767) );
  MUX2_X1 U6975 ( .A(n9513), .B(n2915), .S(n1746), .Z(n6768) );
  MUX2_X1 U6976 ( .A(n9514), .B(n2904), .S(n1746), .Z(n6769) );
  MUX2_X1 U6977 ( .A(n9515), .B(n2892), .S(n1746), .Z(n6770) );
  MUX2_X1 U6978 ( .A(n9516), .B(n2881), .S(n1746), .Z(n6771) );
  MUX2_X1 U6979 ( .A(n9517), .B(n2870), .S(n1746), .Z(n6772) );
  MUX2_X1 U6980 ( .A(n9518), .B(n2859), .S(n1746), .Z(n6773) );
  MUX2_X1 U6981 ( .A(n9519), .B(n2848), .S(n1746), .Z(n6774) );
  MUX2_X1 U6982 ( .A(n9520), .B(n2837), .S(n1746), .Z(n6775) );
  MUX2_X1 U6983 ( .A(n9521), .B(n2826), .S(n1746), .Z(n6776) );
  MUX2_X1 U6984 ( .A(n9522), .B(n2815), .S(n1747), .Z(n6777) );
  MUX2_X1 U6985 ( .A(n9523), .B(n2804), .S(n1747), .Z(n6778) );
  MUX2_X1 U6986 ( .A(n9524), .B(n2793), .S(n1747), .Z(n6779) );
  MUX2_X1 U6987 ( .A(n9525), .B(n2782), .S(n1747), .Z(n6780) );
  MUX2_X1 U6988 ( .A(n9526), .B(n2771), .S(n1747), .Z(n6781) );
  MUX2_X1 U6989 ( .A(n9527), .B(n2760), .S(n1747), .Z(n6782) );
  MUX2_X1 U6990 ( .A(n9528), .B(n2749), .S(n1747), .Z(n6783) );
  MUX2_X1 U6991 ( .A(n9529), .B(n2738), .S(n1747), .Z(n6784) );
  MUX2_X1 U6992 ( .A(n9530), .B(n2727), .S(n1747), .Z(n6785) );
  MUX2_X1 U6993 ( .A(n9531), .B(n2716), .S(n1747), .Z(n6786) );
  MUX2_X1 U6994 ( .A(n9532), .B(n2705), .S(n1747), .Z(n6787) );
  MUX2_X1 U6995 ( .A(n9533), .B(n2598), .S(n1747), .Z(n6788) );
  MUX2_X1 U6996 ( .A(n9534), .B(n2587), .S(n1748), .Z(n6789) );
  MUX2_X1 U6997 ( .A(n9535), .B(n2576), .S(n1748), .Z(n6790) );
  MUX2_X1 U6998 ( .A(n9536), .B(n2565), .S(n1748), .Z(n6791) );
  MUX2_X1 U6999 ( .A(n9537), .B(n2554), .S(n1748), .Z(n6792) );
  MUX2_X1 U7000 ( .A(n9538), .B(n1839), .S(n1748), .Z(n6793) );
  MUX2_X1 U7001 ( .A(n9539), .B(n1828), .S(n1748), .Z(n6794) );
  MUX2_X1 U7002 ( .A(n9540), .B(n1817), .S(n1748), .Z(n6795) );
  MUX2_X1 U7003 ( .A(n9541), .B(n1806), .S(n1748), .Z(n6796) );
  MUX2_X1 U7004 ( .A(n9478), .B(n2953), .S(n1749), .Z(n6733) );
  MUX2_X1 U7005 ( .A(n9479), .B(n2942), .S(n1749), .Z(n6734) );
  MUX2_X1 U7006 ( .A(n9480), .B(n2931), .S(n1749), .Z(n6735) );
  MUX2_X1 U7007 ( .A(n9481), .B(n2915), .S(n1749), .Z(n6736) );
  MUX2_X1 U7008 ( .A(n9482), .B(n2904), .S(n1749), .Z(n6737) );
  MUX2_X1 U7009 ( .A(n9483), .B(n2892), .S(n1749), .Z(n6738) );
  MUX2_X1 U7010 ( .A(n9484), .B(n2881), .S(n1749), .Z(n6739) );
  MUX2_X1 U7011 ( .A(n9485), .B(n2870), .S(n1749), .Z(n6740) );
  MUX2_X1 U7012 ( .A(n9486), .B(n2859), .S(n1749), .Z(n6741) );
  MUX2_X1 U7013 ( .A(n9487), .B(n2848), .S(n1749), .Z(n6742) );
  MUX2_X1 U7014 ( .A(n9488), .B(n2837), .S(n1749), .Z(n6743) );
  MUX2_X1 U7015 ( .A(n9489), .B(n2826), .S(n1749), .Z(n6744) );
  MUX2_X1 U7016 ( .A(n9490), .B(n2815), .S(n1750), .Z(n6745) );
  MUX2_X1 U7017 ( .A(n9491), .B(n2804), .S(n1750), .Z(n6746) );
  MUX2_X1 U7018 ( .A(n9492), .B(n2793), .S(n1750), .Z(n6747) );
  MUX2_X1 U7019 ( .A(n9493), .B(n2782), .S(n1750), .Z(n6748) );
  MUX2_X1 U7020 ( .A(n9494), .B(n2771), .S(n1750), .Z(n6749) );
  MUX2_X1 U7021 ( .A(n9495), .B(n2760), .S(n1750), .Z(n6750) );
  MUX2_X1 U7022 ( .A(n9496), .B(n2749), .S(n1750), .Z(n6751) );
  MUX2_X1 U7023 ( .A(n9497), .B(n2738), .S(n1750), .Z(n6752) );
  MUX2_X1 U7024 ( .A(n9498), .B(n2727), .S(n1750), .Z(n6753) );
  MUX2_X1 U7025 ( .A(n9499), .B(n2716), .S(n1750), .Z(n6754) );
  MUX2_X1 U7026 ( .A(n9500), .B(n2705), .S(n1750), .Z(n6755) );
  MUX2_X1 U7027 ( .A(n9501), .B(n2598), .S(n1750), .Z(n6756) );
  MUX2_X1 U7028 ( .A(n9502), .B(n2587), .S(n1751), .Z(n6757) );
  MUX2_X1 U7029 ( .A(n9503), .B(n2576), .S(n1751), .Z(n6758) );
  MUX2_X1 U7030 ( .A(n9504), .B(n2565), .S(n1751), .Z(n6759) );
  MUX2_X1 U7031 ( .A(n9505), .B(n2554), .S(n1751), .Z(n6760) );
  MUX2_X1 U7032 ( .A(n9506), .B(n1839), .S(n1751), .Z(n6761) );
  MUX2_X1 U7033 ( .A(n9507), .B(n1828), .S(n1751), .Z(n6762) );
  MUX2_X1 U7034 ( .A(n9508), .B(n1817), .S(n1751), .Z(n6763) );
  MUX2_X1 U7035 ( .A(n9509), .B(n1806), .S(n1751), .Z(n6764) );
  MUX2_X1 U7036 ( .A(\REGISTERS[12][31] ), .B(n2953), .S(n1752), .Z(n6701) );
  MUX2_X1 U7037 ( .A(\REGISTERS[12][30] ), .B(n2942), .S(n1752), .Z(n6702) );
  MUX2_X1 U7038 ( .A(\REGISTERS[12][29] ), .B(n2931), .S(n1752), .Z(n6703) );
  MUX2_X1 U7039 ( .A(\REGISTERS[12][28] ), .B(n2915), .S(n1752), .Z(n6704) );
  MUX2_X1 U7040 ( .A(\REGISTERS[12][27] ), .B(n2904), .S(n1752), .Z(n6705) );
  MUX2_X1 U7041 ( .A(\REGISTERS[12][26] ), .B(n2892), .S(n1752), .Z(n6706) );
  MUX2_X1 U7042 ( .A(\REGISTERS[12][25] ), .B(n2881), .S(n1752), .Z(n6707) );
  MUX2_X1 U7043 ( .A(\REGISTERS[12][24] ), .B(n2870), .S(n1752), .Z(n6708) );
  MUX2_X1 U7044 ( .A(\REGISTERS[12][23] ), .B(n2859), .S(n1752), .Z(n6709) );
  MUX2_X1 U7045 ( .A(\REGISTERS[12][22] ), .B(n2848), .S(n1752), .Z(n6710) );
  MUX2_X1 U7046 ( .A(\REGISTERS[12][21] ), .B(n2837), .S(n1752), .Z(n6711) );
  MUX2_X1 U7047 ( .A(\REGISTERS[12][20] ), .B(n2826), .S(n1752), .Z(n6712) );
  MUX2_X1 U7048 ( .A(\REGISTERS[12][19] ), .B(n2815), .S(n1753), .Z(n6713) );
  MUX2_X1 U7049 ( .A(\REGISTERS[12][18] ), .B(n2804), .S(n1753), .Z(n6714) );
  MUX2_X1 U7050 ( .A(\REGISTERS[12][17] ), .B(n2793), .S(n1753), .Z(n6715) );
  MUX2_X1 U7051 ( .A(\REGISTERS[12][16] ), .B(n2782), .S(n1753), .Z(n6716) );
  MUX2_X1 U7052 ( .A(\REGISTERS[12][15] ), .B(n2771), .S(n1753), .Z(n6717) );
  MUX2_X1 U7053 ( .A(\REGISTERS[12][14] ), .B(n2760), .S(n1753), .Z(n6718) );
  MUX2_X1 U7054 ( .A(\REGISTERS[12][13] ), .B(n2749), .S(n1753), .Z(n6719) );
  MUX2_X1 U7055 ( .A(\REGISTERS[12][12] ), .B(n2738), .S(n1753), .Z(n6720) );
  MUX2_X1 U7056 ( .A(\REGISTERS[12][11] ), .B(n2727), .S(n1753), .Z(n6721) );
  MUX2_X1 U7057 ( .A(\REGISTERS[12][10] ), .B(n2716), .S(n1753), .Z(n6722) );
  MUX2_X1 U7058 ( .A(\REGISTERS[12][9] ), .B(n2705), .S(n1753), .Z(n6723) );
  MUX2_X1 U7059 ( .A(\REGISTERS[12][8] ), .B(n2598), .S(n1753), .Z(n6724) );
  MUX2_X1 U7060 ( .A(\REGISTERS[12][7] ), .B(n2587), .S(n1754), .Z(n6725) );
  MUX2_X1 U7061 ( .A(\REGISTERS[12][6] ), .B(n2576), .S(n1754), .Z(n6726) );
  MUX2_X1 U7062 ( .A(\REGISTERS[12][5] ), .B(n2565), .S(n1754), .Z(n6727) );
  MUX2_X1 U7063 ( .A(\REGISTERS[12][4] ), .B(n2554), .S(n1754), .Z(n6728) );
  MUX2_X1 U7064 ( .A(\REGISTERS[12][3] ), .B(n1839), .S(n1754), .Z(n6729) );
  MUX2_X1 U7065 ( .A(\REGISTERS[12][2] ), .B(n1828), .S(n1754), .Z(n6730) );
  MUX2_X1 U7066 ( .A(\REGISTERS[12][1] ), .B(n1817), .S(n1754), .Z(n6731) );
  MUX2_X1 U7067 ( .A(\REGISTERS[12][0] ), .B(n1806), .S(n1754), .Z(n6732) );
  MUX2_X1 U7068 ( .A(\REGISTERS[11][31] ), .B(n2953), .S(n1755), .Z(n6669) );
  MUX2_X1 U7069 ( .A(\REGISTERS[11][30] ), .B(n2942), .S(n1755), .Z(n6670) );
  MUX2_X1 U7070 ( .A(\REGISTERS[11][29] ), .B(n2931), .S(n1755), .Z(n6671) );
  MUX2_X1 U7071 ( .A(\REGISTERS[11][28] ), .B(n2915), .S(n1755), .Z(n6672) );
  MUX2_X1 U7072 ( .A(\REGISTERS[11][27] ), .B(n2904), .S(n1755), .Z(n6673) );
  MUX2_X1 U7073 ( .A(\REGISTERS[11][26] ), .B(n2892), .S(n1755), .Z(n6674) );
  MUX2_X1 U7074 ( .A(\REGISTERS[11][25] ), .B(n2881), .S(n1755), .Z(n6675) );
  MUX2_X1 U7075 ( .A(\REGISTERS[11][24] ), .B(n2870), .S(n1755), .Z(n6676) );
  MUX2_X1 U7076 ( .A(\REGISTERS[11][23] ), .B(n2859), .S(n1755), .Z(n6677) );
  MUX2_X1 U7077 ( .A(\REGISTERS[11][22] ), .B(n2848), .S(n1755), .Z(n6678) );
  MUX2_X1 U7078 ( .A(\REGISTERS[11][21] ), .B(n2837), .S(n1755), .Z(n6679) );
  MUX2_X1 U7079 ( .A(\REGISTERS[11][20] ), .B(n2826), .S(n1755), .Z(n6680) );
  MUX2_X1 U7080 ( .A(\REGISTERS[11][19] ), .B(n2815), .S(n1756), .Z(n6681) );
  MUX2_X1 U7081 ( .A(\REGISTERS[11][18] ), .B(n2804), .S(n1756), .Z(n6682) );
  MUX2_X1 U7082 ( .A(\REGISTERS[11][17] ), .B(n2793), .S(n1756), .Z(n6683) );
  MUX2_X1 U7083 ( .A(\REGISTERS[11][16] ), .B(n2782), .S(n1756), .Z(n6684) );
  MUX2_X1 U7084 ( .A(\REGISTERS[11][15] ), .B(n2771), .S(n1756), .Z(n6685) );
  MUX2_X1 U7085 ( .A(\REGISTERS[11][14] ), .B(n2760), .S(n1756), .Z(n6686) );
  MUX2_X1 U7086 ( .A(\REGISTERS[11][13] ), .B(n2749), .S(n1756), .Z(n6687) );
  MUX2_X1 U7087 ( .A(\REGISTERS[11][12] ), .B(n2738), .S(n1756), .Z(n6688) );
  MUX2_X1 U7088 ( .A(\REGISTERS[11][11] ), .B(n2727), .S(n1756), .Z(n6689) );
  MUX2_X1 U7089 ( .A(\REGISTERS[11][10] ), .B(n2716), .S(n1756), .Z(n6690) );
  MUX2_X1 U7090 ( .A(\REGISTERS[11][9] ), .B(n2705), .S(n1756), .Z(n6691) );
  MUX2_X1 U7091 ( .A(\REGISTERS[11][8] ), .B(n2598), .S(n1756), .Z(n6692) );
  MUX2_X1 U7092 ( .A(\REGISTERS[11][7] ), .B(n2587), .S(n1757), .Z(n6693) );
  MUX2_X1 U7093 ( .A(\REGISTERS[11][6] ), .B(n2576), .S(n1757), .Z(n6694) );
  MUX2_X1 U7094 ( .A(\REGISTERS[11][5] ), .B(n2565), .S(n1757), .Z(n6695) );
  MUX2_X1 U7095 ( .A(\REGISTERS[11][4] ), .B(n2554), .S(n1757), .Z(n6696) );
  MUX2_X1 U7096 ( .A(\REGISTERS[11][3] ), .B(n1839), .S(n1757), .Z(n6697) );
  MUX2_X1 U7097 ( .A(\REGISTERS[11][2] ), .B(n1828), .S(n1757), .Z(n6698) );
  MUX2_X1 U7098 ( .A(\REGISTERS[11][1] ), .B(n1817), .S(n1757), .Z(n6699) );
  MUX2_X1 U7099 ( .A(\REGISTERS[11][0] ), .B(n1806), .S(n1757), .Z(n6700) );
  MUX2_X1 U7100 ( .A(n9446), .B(n2954), .S(n1758), .Z(n6637) );
  MUX2_X1 U7101 ( .A(n9447), .B(n2943), .S(n1758), .Z(n6638) );
  MUX2_X1 U7102 ( .A(n9448), .B(n2932), .S(n1758), .Z(n6639) );
  MUX2_X1 U7103 ( .A(n9449), .B(n2917), .S(n1758), .Z(n6640) );
  MUX2_X1 U7104 ( .A(n9450), .B(n2905), .S(n1758), .Z(n6641) );
  MUX2_X1 U7105 ( .A(n9451), .B(n2893), .S(n1758), .Z(n6642) );
  MUX2_X1 U7106 ( .A(n9452), .B(n2882), .S(n1758), .Z(n6643) );
  MUX2_X1 U7107 ( .A(n9453), .B(n2871), .S(n1758), .Z(n6644) );
  MUX2_X1 U7108 ( .A(n9454), .B(n2860), .S(n1758), .Z(n6645) );
  MUX2_X1 U7109 ( .A(n9455), .B(n2849), .S(n1758), .Z(n6646) );
  MUX2_X1 U7110 ( .A(n9456), .B(n2838), .S(n1758), .Z(n6647) );
  MUX2_X1 U7111 ( .A(n9457), .B(n2827), .S(n1758), .Z(n6648) );
  MUX2_X1 U7112 ( .A(n9458), .B(n2816), .S(n1759), .Z(n6649) );
  MUX2_X1 U7113 ( .A(n9459), .B(n2805), .S(n1759), .Z(n6650) );
  MUX2_X1 U7114 ( .A(n9460), .B(n2794), .S(n1759), .Z(n6651) );
  MUX2_X1 U7115 ( .A(n9461), .B(n2783), .S(n1759), .Z(n6652) );
  MUX2_X1 U7116 ( .A(n9462), .B(n2772), .S(n1759), .Z(n6653) );
  MUX2_X1 U7117 ( .A(n9463), .B(n2761), .S(n1759), .Z(n6654) );
  MUX2_X1 U7118 ( .A(n9464), .B(n2750), .S(n1759), .Z(n6655) );
  MUX2_X1 U7119 ( .A(n9465), .B(n2739), .S(n1759), .Z(n6656) );
  MUX2_X1 U7120 ( .A(n9466), .B(n2728), .S(n1759), .Z(n6657) );
  MUX2_X1 U7121 ( .A(n9467), .B(n2717), .S(n1759), .Z(n6658) );
  MUX2_X1 U7122 ( .A(n9468), .B(n2706), .S(n1759), .Z(n6659) );
  MUX2_X1 U7123 ( .A(n9469), .B(n2599), .S(n1759), .Z(n6660) );
  MUX2_X1 U7124 ( .A(n9470), .B(n2588), .S(n1760), .Z(n6661) );
  MUX2_X1 U7125 ( .A(n9471), .B(n2577), .S(n1760), .Z(n6662) );
  MUX2_X1 U7126 ( .A(n9472), .B(n2566), .S(n1760), .Z(n6663) );
  MUX2_X1 U7127 ( .A(n9473), .B(n2555), .S(n1760), .Z(n6664) );
  MUX2_X1 U7128 ( .A(n9474), .B(n2544), .S(n1760), .Z(n6665) );
  MUX2_X1 U7129 ( .A(n9475), .B(n1829), .S(n1760), .Z(n6666) );
  MUX2_X1 U7130 ( .A(n9476), .B(n1818), .S(n1760), .Z(n6667) );
  MUX2_X1 U7131 ( .A(n9477), .B(n1807), .S(n1760), .Z(n6668) );
  MUX2_X1 U7132 ( .A(n9414), .B(n2954), .S(n1761), .Z(n6605) );
  MUX2_X1 U7133 ( .A(n9415), .B(n2943), .S(n1761), .Z(n6606) );
  MUX2_X1 U7134 ( .A(n9416), .B(n2932), .S(n1761), .Z(n6607) );
  MUX2_X1 U7135 ( .A(n9417), .B(n2917), .S(n1761), .Z(n6608) );
  MUX2_X1 U7136 ( .A(n9418), .B(n2905), .S(n1761), .Z(n6609) );
  MUX2_X1 U7137 ( .A(n9419), .B(n2893), .S(n1761), .Z(n6610) );
  MUX2_X1 U7138 ( .A(n9420), .B(n2882), .S(n1761), .Z(n6611) );
  MUX2_X1 U7139 ( .A(n9421), .B(n2871), .S(n1761), .Z(n6612) );
  MUX2_X1 U7140 ( .A(n9422), .B(n2860), .S(n1761), .Z(n6613) );
  MUX2_X1 U7141 ( .A(n9423), .B(n2849), .S(n1761), .Z(n6614) );
  MUX2_X1 U7142 ( .A(n9424), .B(n2838), .S(n1761), .Z(n6615) );
  MUX2_X1 U7143 ( .A(n9425), .B(n2827), .S(n1761), .Z(n6616) );
  MUX2_X1 U7144 ( .A(n9426), .B(n2816), .S(n1762), .Z(n6617) );
  MUX2_X1 U7145 ( .A(n9427), .B(n2805), .S(n1762), .Z(n6618) );
  MUX2_X1 U7146 ( .A(n9428), .B(n2794), .S(n1762), .Z(n6619) );
  MUX2_X1 U7147 ( .A(n9429), .B(n2783), .S(n1762), .Z(n6620) );
  MUX2_X1 U7148 ( .A(n9430), .B(n2772), .S(n1762), .Z(n6621) );
  MUX2_X1 U7149 ( .A(n9431), .B(n2761), .S(n1762), .Z(n6622) );
  MUX2_X1 U7150 ( .A(n9432), .B(n2750), .S(n1762), .Z(n6623) );
  MUX2_X1 U7151 ( .A(n9433), .B(n2739), .S(n1762), .Z(n6624) );
  MUX2_X1 U7152 ( .A(n9434), .B(n2728), .S(n1762), .Z(n6625) );
  MUX2_X1 U7153 ( .A(n9435), .B(n2717), .S(n1762), .Z(n6626) );
  MUX2_X1 U7154 ( .A(n9436), .B(n2706), .S(n1762), .Z(n6627) );
  MUX2_X1 U7155 ( .A(n9437), .B(n2599), .S(n1762), .Z(n6628) );
  MUX2_X1 U7156 ( .A(n9438), .B(n2588), .S(n1763), .Z(n6629) );
  MUX2_X1 U7157 ( .A(n9439), .B(n2577), .S(n1763), .Z(n6630) );
  MUX2_X1 U7158 ( .A(n9440), .B(n2566), .S(n1763), .Z(n6631) );
  MUX2_X1 U7159 ( .A(n9441), .B(n2555), .S(n1763), .Z(n6632) );
  MUX2_X1 U7160 ( .A(n9442), .B(n2544), .S(n1763), .Z(n6633) );
  MUX2_X1 U7161 ( .A(n9443), .B(n1829), .S(n1763), .Z(n6634) );
  MUX2_X1 U7162 ( .A(n9444), .B(n1818), .S(n1763), .Z(n6635) );
  MUX2_X1 U7163 ( .A(n9445), .B(n1807), .S(n1763), .Z(n6636) );
  MUX2_X1 U7164 ( .A(n9382), .B(n2954), .S(n1764), .Z(n6573) );
  MUX2_X1 U7165 ( .A(n9383), .B(n2943), .S(n1764), .Z(n6574) );
  MUX2_X1 U7166 ( .A(n9384), .B(n2932), .S(n1764), .Z(n6575) );
  MUX2_X1 U7167 ( .A(n9385), .B(n2917), .S(n1764), .Z(n6576) );
  MUX2_X1 U7168 ( .A(n9386), .B(n2905), .S(n1764), .Z(n6577) );
  MUX2_X1 U7169 ( .A(n9387), .B(n2893), .S(n1764), .Z(n6578) );
  MUX2_X1 U7170 ( .A(n9388), .B(n2882), .S(n1764), .Z(n6579) );
  MUX2_X1 U7171 ( .A(n9389), .B(n2871), .S(n1764), .Z(n6580) );
  MUX2_X1 U7172 ( .A(n9390), .B(n2860), .S(n1764), .Z(n6581) );
  MUX2_X1 U7173 ( .A(n9391), .B(n2849), .S(n1764), .Z(n6582) );
  MUX2_X1 U7174 ( .A(n9392), .B(n2838), .S(n1764), .Z(n6583) );
  MUX2_X1 U7175 ( .A(n9393), .B(n2827), .S(n1764), .Z(n6584) );
  MUX2_X1 U7176 ( .A(n9394), .B(n2816), .S(n1765), .Z(n6585) );
  MUX2_X1 U7177 ( .A(n9395), .B(n2805), .S(n1765), .Z(n6586) );
  MUX2_X1 U7178 ( .A(n9396), .B(n2794), .S(n1765), .Z(n6587) );
  MUX2_X1 U7179 ( .A(n9397), .B(n2783), .S(n1765), .Z(n6588) );
  MUX2_X1 U7180 ( .A(n9398), .B(n2772), .S(n1765), .Z(n6589) );
  MUX2_X1 U7181 ( .A(n9399), .B(n2761), .S(n1765), .Z(n6590) );
  MUX2_X1 U7182 ( .A(n9400), .B(n2750), .S(n1765), .Z(n6591) );
  MUX2_X1 U7183 ( .A(n9401), .B(n2739), .S(n1765), .Z(n6592) );
  MUX2_X1 U7184 ( .A(n9402), .B(n2728), .S(n1765), .Z(n6593) );
  MUX2_X1 U7185 ( .A(n9403), .B(n2717), .S(n1765), .Z(n6594) );
  MUX2_X1 U7186 ( .A(n9404), .B(n2706), .S(n1765), .Z(n6595) );
  MUX2_X1 U7187 ( .A(n9405), .B(n2599), .S(n1765), .Z(n6596) );
  MUX2_X1 U7188 ( .A(n9406), .B(n2588), .S(n1766), .Z(n6597) );
  MUX2_X1 U7189 ( .A(n9407), .B(n2577), .S(n1766), .Z(n6598) );
  MUX2_X1 U7190 ( .A(n9408), .B(n2566), .S(n1766), .Z(n6599) );
  MUX2_X1 U7191 ( .A(n9409), .B(n2555), .S(n1766), .Z(n6600) );
  MUX2_X1 U7192 ( .A(n9410), .B(n2544), .S(n1766), .Z(n6601) );
  MUX2_X1 U7193 ( .A(n9411), .B(n1829), .S(n1766), .Z(n6602) );
  MUX2_X1 U7194 ( .A(n9412), .B(n1818), .S(n1766), .Z(n6603) );
  MUX2_X1 U7195 ( .A(n9413), .B(n1807), .S(n1766), .Z(n6604) );
  MUX2_X1 U7196 ( .A(n9350), .B(n2954), .S(n1767), .Z(n6541) );
  MUX2_X1 U7197 ( .A(n9351), .B(n2943), .S(n1767), .Z(n6542) );
  MUX2_X1 U7198 ( .A(n9352), .B(n2932), .S(n1767), .Z(n6543) );
  MUX2_X1 U7199 ( .A(n9353), .B(n2917), .S(n1767), .Z(n6544) );
  MUX2_X1 U7200 ( .A(n9354), .B(n2905), .S(n1767), .Z(n6545) );
  MUX2_X1 U7201 ( .A(n9355), .B(n2893), .S(n1767), .Z(n6546) );
  MUX2_X1 U7202 ( .A(n9356), .B(n2882), .S(n1767), .Z(n6547) );
  MUX2_X1 U7203 ( .A(n9357), .B(n2871), .S(n1767), .Z(n6548) );
  MUX2_X1 U7204 ( .A(n9358), .B(n2860), .S(n1767), .Z(n6549) );
  MUX2_X1 U7205 ( .A(n9359), .B(n2849), .S(n1767), .Z(n6550) );
  MUX2_X1 U7206 ( .A(n9360), .B(n2838), .S(n1767), .Z(n6551) );
  MUX2_X1 U7207 ( .A(n9361), .B(n2827), .S(n1767), .Z(n6552) );
  MUX2_X1 U7208 ( .A(n9362), .B(n2816), .S(n1768), .Z(n6553) );
  MUX2_X1 U7209 ( .A(n9363), .B(n2805), .S(n1768), .Z(n6554) );
  MUX2_X1 U7210 ( .A(n9364), .B(n2794), .S(n1768), .Z(n6555) );
  MUX2_X1 U7211 ( .A(n9365), .B(n2783), .S(n1768), .Z(n6556) );
  MUX2_X1 U7212 ( .A(n9366), .B(n2772), .S(n1768), .Z(n6557) );
  MUX2_X1 U7213 ( .A(n9367), .B(n2761), .S(n1768), .Z(n6558) );
  MUX2_X1 U7214 ( .A(n9368), .B(n2750), .S(n1768), .Z(n6559) );
  MUX2_X1 U7215 ( .A(n9369), .B(n2739), .S(n1768), .Z(n6560) );
  MUX2_X1 U7216 ( .A(n9370), .B(n2728), .S(n1768), .Z(n6561) );
  MUX2_X1 U7217 ( .A(n9371), .B(n2717), .S(n1768), .Z(n6562) );
  MUX2_X1 U7218 ( .A(n9372), .B(n2706), .S(n1768), .Z(n6563) );
  MUX2_X1 U7219 ( .A(n9373), .B(n2599), .S(n1768), .Z(n6564) );
  MUX2_X1 U7220 ( .A(n9374), .B(n2588), .S(n1769), .Z(n6565) );
  MUX2_X1 U7221 ( .A(n9375), .B(n2577), .S(n1769), .Z(n6566) );
  MUX2_X1 U7222 ( .A(n9376), .B(n2566), .S(n1769), .Z(n6567) );
  MUX2_X1 U7223 ( .A(n9377), .B(n2555), .S(n1769), .Z(n6568) );
  MUX2_X1 U7224 ( .A(n9378), .B(n2544), .S(n1769), .Z(n6569) );
  MUX2_X1 U7225 ( .A(n9379), .B(n1829), .S(n1769), .Z(n6570) );
  MUX2_X1 U7226 ( .A(n9380), .B(n1818), .S(n1769), .Z(n6571) );
  MUX2_X1 U7227 ( .A(n9381), .B(n1807), .S(n1769), .Z(n6572) );
  MUX2_X1 U7228 ( .A(n9318), .B(n2954), .S(n1770), .Z(n6509) );
  MUX2_X1 U7229 ( .A(n9319), .B(n2943), .S(n1770), .Z(n6510) );
  MUX2_X1 U7230 ( .A(n9320), .B(n2932), .S(n1770), .Z(n6511) );
  MUX2_X1 U7231 ( .A(n9321), .B(n2917), .S(n1770), .Z(n6512) );
  MUX2_X1 U7232 ( .A(n9322), .B(n2905), .S(n1770), .Z(n6513) );
  MUX2_X1 U7233 ( .A(n9323), .B(n2893), .S(n1770), .Z(n6514) );
  MUX2_X1 U7234 ( .A(n9324), .B(n2882), .S(n1770), .Z(n6515) );
  MUX2_X1 U7235 ( .A(n9325), .B(n2871), .S(n1770), .Z(n6516) );
  MUX2_X1 U7236 ( .A(n9326), .B(n2860), .S(n1770), .Z(n6517) );
  MUX2_X1 U7237 ( .A(n9327), .B(n2849), .S(n1770), .Z(n6518) );
  MUX2_X1 U7238 ( .A(n9328), .B(n2838), .S(n1770), .Z(n6519) );
  MUX2_X1 U7239 ( .A(n9329), .B(n2827), .S(n1770), .Z(n6520) );
  MUX2_X1 U7240 ( .A(n9330), .B(n2816), .S(n1771), .Z(n6521) );
  MUX2_X1 U7241 ( .A(n9331), .B(n2805), .S(n1771), .Z(n6522) );
  MUX2_X1 U7242 ( .A(n9332), .B(n2794), .S(n1771), .Z(n6523) );
  MUX2_X1 U7243 ( .A(n9333), .B(n2783), .S(n1771), .Z(n6524) );
  MUX2_X1 U7244 ( .A(n9334), .B(n2772), .S(n1771), .Z(n6525) );
  MUX2_X1 U7245 ( .A(n9335), .B(n2761), .S(n1771), .Z(n6526) );
  MUX2_X1 U7246 ( .A(n9336), .B(n2750), .S(n1771), .Z(n6527) );
  MUX2_X1 U7247 ( .A(n9337), .B(n2739), .S(n1771), .Z(n6528) );
  MUX2_X1 U7248 ( .A(n9338), .B(n2728), .S(n1771), .Z(n6529) );
  MUX2_X1 U7249 ( .A(n9339), .B(n2717), .S(n1771), .Z(n6530) );
  MUX2_X1 U7250 ( .A(n9340), .B(n2706), .S(n1771), .Z(n6531) );
  MUX2_X1 U7251 ( .A(n9341), .B(n2599), .S(n1771), .Z(n6532) );
  MUX2_X1 U7252 ( .A(n9342), .B(n2588), .S(n1772), .Z(n6533) );
  MUX2_X1 U7253 ( .A(n9343), .B(n2577), .S(n1772), .Z(n6534) );
  MUX2_X1 U7254 ( .A(n9344), .B(n2566), .S(n1772), .Z(n6535) );
  MUX2_X1 U7255 ( .A(n9345), .B(n2555), .S(n1772), .Z(n6536) );
  MUX2_X1 U7256 ( .A(n9346), .B(n2544), .S(n1772), .Z(n6537) );
  MUX2_X1 U7257 ( .A(n9347), .B(n1829), .S(n1772), .Z(n6538) );
  MUX2_X1 U7258 ( .A(n9348), .B(n1818), .S(n1772), .Z(n6539) );
  MUX2_X1 U7259 ( .A(n9349), .B(n1807), .S(n1772), .Z(n6540) );
  MUX2_X1 U7260 ( .A(n9286), .B(n2954), .S(n1773), .Z(n6477) );
  MUX2_X1 U7261 ( .A(n9287), .B(n2943), .S(n1773), .Z(n6478) );
  MUX2_X1 U7262 ( .A(n9288), .B(n2932), .S(n1773), .Z(n6479) );
  MUX2_X1 U7263 ( .A(n9289), .B(n2917), .S(n1773), .Z(n6480) );
  MUX2_X1 U7264 ( .A(n9290), .B(n2905), .S(n1773), .Z(n6481) );
  MUX2_X1 U7265 ( .A(n9291), .B(n2893), .S(n1773), .Z(n6482) );
  MUX2_X1 U7266 ( .A(n9292), .B(n2882), .S(n1773), .Z(n6483) );
  MUX2_X1 U7267 ( .A(n9293), .B(n2871), .S(n1773), .Z(n6484) );
  MUX2_X1 U7268 ( .A(n9294), .B(n2860), .S(n1773), .Z(n6485) );
  MUX2_X1 U7269 ( .A(n9295), .B(n2849), .S(n1773), .Z(n6486) );
  MUX2_X1 U7270 ( .A(n9296), .B(n2838), .S(n1773), .Z(n6487) );
  MUX2_X1 U7271 ( .A(n9297), .B(n2827), .S(n1773), .Z(n6488) );
  MUX2_X1 U7272 ( .A(n9298), .B(n2816), .S(n1774), .Z(n6489) );
  MUX2_X1 U7273 ( .A(n9299), .B(n2805), .S(n1774), .Z(n6490) );
  MUX2_X1 U7274 ( .A(n9300), .B(n2794), .S(n1774), .Z(n6491) );
  MUX2_X1 U7275 ( .A(n9301), .B(n2783), .S(n1774), .Z(n6492) );
  MUX2_X1 U7276 ( .A(n9302), .B(n2772), .S(n1774), .Z(n6493) );
  MUX2_X1 U7277 ( .A(n9303), .B(n2761), .S(n1774), .Z(n6494) );
  MUX2_X1 U7278 ( .A(n9304), .B(n2750), .S(n1774), .Z(n6495) );
  MUX2_X1 U7279 ( .A(n9305), .B(n2739), .S(n1774), .Z(n6496) );
  MUX2_X1 U7280 ( .A(n9306), .B(n2728), .S(n1774), .Z(n6497) );
  MUX2_X1 U7281 ( .A(n9307), .B(n2717), .S(n1774), .Z(n6498) );
  MUX2_X1 U7282 ( .A(n9308), .B(n2706), .S(n1774), .Z(n6499) );
  MUX2_X1 U7283 ( .A(n9309), .B(n2599), .S(n1774), .Z(n6500) );
  MUX2_X1 U7284 ( .A(n9310), .B(n2588), .S(n1775), .Z(n6501) );
  MUX2_X1 U7285 ( .A(n9311), .B(n2577), .S(n1775), .Z(n6502) );
  MUX2_X1 U7286 ( .A(n9312), .B(n2566), .S(n1775), .Z(n6503) );
  MUX2_X1 U7287 ( .A(n9313), .B(n2555), .S(n1775), .Z(n6504) );
  MUX2_X1 U7288 ( .A(n9314), .B(n2544), .S(n1775), .Z(n6505) );
  MUX2_X1 U7289 ( .A(n9315), .B(n1829), .S(n1775), .Z(n6506) );
  MUX2_X1 U7290 ( .A(n9316), .B(n1818), .S(n1775), .Z(n6507) );
  MUX2_X1 U7291 ( .A(n9317), .B(n1807), .S(n1775), .Z(n6508) );
  MUX2_X1 U7292 ( .A(n9254), .B(n2954), .S(n1776), .Z(n6445) );
  MUX2_X1 U7293 ( .A(n9255), .B(n2943), .S(n1776), .Z(n6446) );
  MUX2_X1 U7294 ( .A(n9256), .B(n2932), .S(n1776), .Z(n6447) );
  MUX2_X1 U7295 ( .A(n9257), .B(n2917), .S(n1776), .Z(n6448) );
  MUX2_X1 U7296 ( .A(n9258), .B(n2905), .S(n1776), .Z(n6449) );
  MUX2_X1 U7297 ( .A(n9259), .B(n2893), .S(n1776), .Z(n6450) );
  MUX2_X1 U7298 ( .A(n9260), .B(n2882), .S(n1776), .Z(n6451) );
  MUX2_X1 U7299 ( .A(n9261), .B(n2871), .S(n1776), .Z(n6452) );
  MUX2_X1 U7300 ( .A(n9262), .B(n2860), .S(n1776), .Z(n6453) );
  MUX2_X1 U7301 ( .A(n9263), .B(n2849), .S(n1776), .Z(n6454) );
  MUX2_X1 U7302 ( .A(n9264), .B(n2838), .S(n1776), .Z(n6455) );
  MUX2_X1 U7303 ( .A(n9265), .B(n2827), .S(n1776), .Z(n6456) );
  MUX2_X1 U7304 ( .A(n9266), .B(n2816), .S(n1777), .Z(n6457) );
  MUX2_X1 U7305 ( .A(n9267), .B(n2805), .S(n1777), .Z(n6458) );
  MUX2_X1 U7306 ( .A(n9268), .B(n2794), .S(n1777), .Z(n6459) );
  MUX2_X1 U7307 ( .A(n9269), .B(n2783), .S(n1777), .Z(n6460) );
  MUX2_X1 U7308 ( .A(n9270), .B(n2772), .S(n1777), .Z(n6461) );
  MUX2_X1 U7309 ( .A(n9271), .B(n2761), .S(n1777), .Z(n6462) );
  MUX2_X1 U7310 ( .A(n9272), .B(n2750), .S(n1777), .Z(n6463) );
  MUX2_X1 U7311 ( .A(n9273), .B(n2739), .S(n1777), .Z(n6464) );
  MUX2_X1 U7312 ( .A(n9274), .B(n2728), .S(n1777), .Z(n6465) );
  MUX2_X1 U7313 ( .A(n9275), .B(n2717), .S(n1777), .Z(n6466) );
  MUX2_X1 U7314 ( .A(n9276), .B(n2706), .S(n1777), .Z(n6467) );
  MUX2_X1 U7315 ( .A(n9277), .B(n2599), .S(n1777), .Z(n6468) );
  MUX2_X1 U7316 ( .A(n9278), .B(n2588), .S(n1778), .Z(n6469) );
  MUX2_X1 U7317 ( .A(n9279), .B(n2577), .S(n1778), .Z(n6470) );
  MUX2_X1 U7318 ( .A(n9280), .B(n2566), .S(n1778), .Z(n6471) );
  MUX2_X1 U7319 ( .A(n9281), .B(n2555), .S(n1778), .Z(n6472) );
  MUX2_X1 U7320 ( .A(n9282), .B(n2544), .S(n1778), .Z(n6473) );
  MUX2_X1 U7321 ( .A(n9283), .B(n1829), .S(n1778), .Z(n6474) );
  MUX2_X1 U7322 ( .A(n9284), .B(n1818), .S(n1778), .Z(n6475) );
  MUX2_X1 U7323 ( .A(n9285), .B(n1807), .S(n1778), .Z(n6476) );
  MUX2_X1 U7324 ( .A(n9222), .B(n2954), .S(n1779), .Z(n6413) );
  MUX2_X1 U7325 ( .A(n9223), .B(n2943), .S(n1779), .Z(n6414) );
  MUX2_X1 U7326 ( .A(n9224), .B(n2932), .S(n1779), .Z(n6415) );
  MUX2_X1 U7327 ( .A(n9225), .B(n2917), .S(n1779), .Z(n6416) );
  MUX2_X1 U7328 ( .A(n9226), .B(n2905), .S(n1779), .Z(n6417) );
  MUX2_X1 U7329 ( .A(n9227), .B(n2893), .S(n1779), .Z(n6418) );
  MUX2_X1 U7330 ( .A(n9228), .B(n2882), .S(n1779), .Z(n6419) );
  MUX2_X1 U7331 ( .A(n9229), .B(n2871), .S(n1779), .Z(n6420) );
  MUX2_X1 U7332 ( .A(n9230), .B(n2860), .S(n1779), .Z(n6421) );
  MUX2_X1 U7333 ( .A(n9231), .B(n2849), .S(n1779), .Z(n6422) );
  MUX2_X1 U7334 ( .A(n9232), .B(n2838), .S(n1779), .Z(n6423) );
  MUX2_X1 U7335 ( .A(n9233), .B(n2827), .S(n1779), .Z(n6424) );
  MUX2_X1 U7336 ( .A(n9234), .B(n2816), .S(n1780), .Z(n6425) );
  MUX2_X1 U7337 ( .A(n9235), .B(n2805), .S(n1780), .Z(n6426) );
  MUX2_X1 U7338 ( .A(n9236), .B(n2794), .S(n1780), .Z(n6427) );
  MUX2_X1 U7339 ( .A(n9237), .B(n2783), .S(n1780), .Z(n6428) );
  MUX2_X1 U7340 ( .A(n9238), .B(n2772), .S(n1780), .Z(n6429) );
  MUX2_X1 U7341 ( .A(n9239), .B(n2761), .S(n1780), .Z(n6430) );
  MUX2_X1 U7342 ( .A(n9240), .B(n2750), .S(n1780), .Z(n6431) );
  MUX2_X1 U7343 ( .A(n9241), .B(n2739), .S(n1780), .Z(n6432) );
  MUX2_X1 U7344 ( .A(n9242), .B(n2728), .S(n1780), .Z(n6433) );
  MUX2_X1 U7345 ( .A(n9243), .B(n2717), .S(n1780), .Z(n6434) );
  MUX2_X1 U7346 ( .A(n9244), .B(n2706), .S(n1780), .Z(n6435) );
  MUX2_X1 U7347 ( .A(n9245), .B(n2599), .S(n1780), .Z(n6436) );
  MUX2_X1 U7348 ( .A(n9246), .B(n2588), .S(n1781), .Z(n6437) );
  MUX2_X1 U7349 ( .A(n9247), .B(n2577), .S(n1781), .Z(n6438) );
  MUX2_X1 U7350 ( .A(n9248), .B(n2566), .S(n1781), .Z(n6439) );
  MUX2_X1 U7351 ( .A(n9249), .B(n2555), .S(n1781), .Z(n6440) );
  MUX2_X1 U7352 ( .A(n9250), .B(n2544), .S(n1781), .Z(n6441) );
  MUX2_X1 U7353 ( .A(n9251), .B(n1829), .S(n1781), .Z(n6442) );
  MUX2_X1 U7354 ( .A(n9252), .B(n1818), .S(n1781), .Z(n6443) );
  MUX2_X1 U7355 ( .A(n9253), .B(n1807), .S(n1781), .Z(n6444) );
  MUX2_X1 U7356 ( .A(n9190), .B(n2954), .S(n1782), .Z(n6381) );
  MUX2_X1 U7357 ( .A(n9191), .B(n2943), .S(n1782), .Z(n6382) );
  MUX2_X1 U7358 ( .A(n9192), .B(n2932), .S(n1782), .Z(n6383) );
  MUX2_X1 U7359 ( .A(n9193), .B(n2917), .S(n1782), .Z(n6384) );
  MUX2_X1 U7360 ( .A(n9194), .B(n2905), .S(n1782), .Z(n6385) );
  MUX2_X1 U7361 ( .A(n9195), .B(n2893), .S(n1782), .Z(n6386) );
  MUX2_X1 U7362 ( .A(n9196), .B(n2882), .S(n1782), .Z(n6387) );
  MUX2_X1 U7363 ( .A(n9197), .B(n2871), .S(n1782), .Z(n6388) );
  MUX2_X1 U7364 ( .A(n9198), .B(n2860), .S(n1782), .Z(n6389) );
  MUX2_X1 U7365 ( .A(n9199), .B(n2849), .S(n1782), .Z(n6390) );
  MUX2_X1 U7366 ( .A(n9200), .B(n2838), .S(n1782), .Z(n6391) );
  MUX2_X1 U7367 ( .A(n9201), .B(n2827), .S(n1782), .Z(n6392) );
  MUX2_X1 U7368 ( .A(n9202), .B(n2816), .S(n1783), .Z(n6393) );
  MUX2_X1 U7369 ( .A(n9203), .B(n2805), .S(n1783), .Z(n6394) );
  MUX2_X1 U7370 ( .A(n9204), .B(n2794), .S(n1783), .Z(n6395) );
  MUX2_X1 U7371 ( .A(n9205), .B(n2783), .S(n1783), .Z(n6396) );
  MUX2_X1 U7372 ( .A(n9206), .B(n2772), .S(n1783), .Z(n6397) );
  MUX2_X1 U7373 ( .A(n9207), .B(n2761), .S(n1783), .Z(n6398) );
  MUX2_X1 U7374 ( .A(n9208), .B(n2750), .S(n1783), .Z(n6399) );
  MUX2_X1 U7375 ( .A(n9209), .B(n2739), .S(n1783), .Z(n6400) );
  MUX2_X1 U7376 ( .A(n9210), .B(n2728), .S(n1783), .Z(n6401) );
  MUX2_X1 U7377 ( .A(n9211), .B(n2717), .S(n1783), .Z(n6402) );
  MUX2_X1 U7378 ( .A(n9212), .B(n2706), .S(n1783), .Z(n6403) );
  MUX2_X1 U7379 ( .A(n9213), .B(n2599), .S(n1783), .Z(n6404) );
  MUX2_X1 U7380 ( .A(n9214), .B(n2588), .S(n1784), .Z(n6405) );
  MUX2_X1 U7381 ( .A(n9215), .B(n2577), .S(n1784), .Z(n6406) );
  MUX2_X1 U7382 ( .A(n9216), .B(n2566), .S(n1784), .Z(n6407) );
  MUX2_X1 U7383 ( .A(n9217), .B(n2555), .S(n1784), .Z(n6408) );
  MUX2_X1 U7384 ( .A(n9218), .B(n2544), .S(n1784), .Z(n6409) );
  MUX2_X1 U7385 ( .A(n9219), .B(n1829), .S(n1784), .Z(n6410) );
  MUX2_X1 U7386 ( .A(n9220), .B(n1818), .S(n1784), .Z(n6411) );
  MUX2_X1 U7387 ( .A(n9221), .B(n1807), .S(n1784), .Z(n6412) );
  MUX2_X1 U7388 ( .A(n9158), .B(n2954), .S(n1785), .Z(n6349) );
  MUX2_X1 U7389 ( .A(n9159), .B(n2943), .S(n1785), .Z(n6350) );
  MUX2_X1 U7390 ( .A(n9160), .B(n2932), .S(n1785), .Z(n6351) );
  MUX2_X1 U7391 ( .A(n9161), .B(n2917), .S(n1785), .Z(n6352) );
  MUX2_X1 U7392 ( .A(n9162), .B(n2905), .S(n1785), .Z(n6353) );
  MUX2_X1 U7393 ( .A(n9163), .B(n2893), .S(n1785), .Z(n6354) );
  MUX2_X1 U7394 ( .A(n9164), .B(n2882), .S(n1785), .Z(n6355) );
  MUX2_X1 U7395 ( .A(n9165), .B(n2871), .S(n1785), .Z(n6356) );
  MUX2_X1 U7396 ( .A(n9166), .B(n2860), .S(n1785), .Z(n6357) );
  MUX2_X1 U7397 ( .A(n9167), .B(n2849), .S(n1785), .Z(n6358) );
  MUX2_X1 U7398 ( .A(n9168), .B(n2838), .S(n1785), .Z(n6359) );
  MUX2_X1 U7399 ( .A(n9169), .B(n2827), .S(n1785), .Z(n6360) );
  MUX2_X1 U7400 ( .A(n9170), .B(n2816), .S(n1786), .Z(n6361) );
  MUX2_X1 U7401 ( .A(n9171), .B(n2805), .S(n1786), .Z(n6362) );
  MUX2_X1 U7402 ( .A(n9172), .B(n2794), .S(n1786), .Z(n6363) );
  MUX2_X1 U7403 ( .A(n9173), .B(n2783), .S(n1786), .Z(n6364) );
  MUX2_X1 U7404 ( .A(n9174), .B(n2772), .S(n1786), .Z(n6365) );
  MUX2_X1 U7405 ( .A(n9175), .B(n2761), .S(n1786), .Z(n6366) );
  MUX2_X1 U7406 ( .A(n9176), .B(n2750), .S(n1786), .Z(n6367) );
  MUX2_X1 U7407 ( .A(n9177), .B(n2739), .S(n1786), .Z(n6368) );
  MUX2_X1 U7408 ( .A(n9178), .B(n2728), .S(n1786), .Z(n6369) );
  MUX2_X1 U7409 ( .A(n9179), .B(n2717), .S(n1786), .Z(n6370) );
  MUX2_X1 U7410 ( .A(n9180), .B(n2706), .S(n1786), .Z(n6371) );
  MUX2_X1 U7411 ( .A(n9181), .B(n2599), .S(n1786), .Z(n6372) );
  MUX2_X1 U7412 ( .A(n9182), .B(n2588), .S(n1787), .Z(n6373) );
  MUX2_X1 U7413 ( .A(n9183), .B(n2577), .S(n1787), .Z(n6374) );
  MUX2_X1 U7414 ( .A(n9184), .B(n2566), .S(n1787), .Z(n6375) );
  MUX2_X1 U7415 ( .A(n9185), .B(n2555), .S(n1787), .Z(n6376) );
  MUX2_X1 U7416 ( .A(n9186), .B(n2544), .S(n1787), .Z(n6377) );
  MUX2_X1 U7417 ( .A(n9187), .B(n1829), .S(n1787), .Z(n6378) );
  MUX2_X1 U7418 ( .A(n9188), .B(n1818), .S(n1787), .Z(n6379) );
  MUX2_X1 U7419 ( .A(n9189), .B(n1807), .S(n1787), .Z(n6380) );
  MUX2_X1 U7420 ( .A(n3393), .B(n2954), .S(n1788), .Z(n6317) );
  MUX2_X1 U7421 ( .A(n3395), .B(n2943), .S(n1788), .Z(n6318) );
  MUX2_X1 U7422 ( .A(n3396), .B(n2932), .S(n1788), .Z(n6319) );
  MUX2_X1 U7423 ( .A(n3397), .B(n2917), .S(n1788), .Z(n6320) );
  MUX2_X1 U7424 ( .A(n3399), .B(n2905), .S(n1788), .Z(n6321) );
  MUX2_X1 U7425 ( .A(n3401), .B(n2893), .S(n1788), .Z(n6322) );
  MUX2_X1 U7426 ( .A(n3402), .B(n2882), .S(n1788), .Z(n6323) );
  MUX2_X1 U7427 ( .A(n3404), .B(n2871), .S(n1788), .Z(n6324) );
  MUX2_X1 U7428 ( .A(n3407), .B(n2860), .S(n1788), .Z(n6325) );
  MUX2_X1 U7429 ( .A(n3408), .B(n2849), .S(n1788), .Z(n6326) );
  MUX2_X1 U7430 ( .A(n3410), .B(n2838), .S(n1788), .Z(n6327) );
  MUX2_X1 U7431 ( .A(n3411), .B(n2827), .S(n1788), .Z(n6328) );
  MUX2_X1 U7432 ( .A(n3412), .B(n2816), .S(n1789), .Z(n6329) );
  MUX2_X1 U7433 ( .A(n3414), .B(n2805), .S(n1789), .Z(n6330) );
  MUX2_X1 U7434 ( .A(n9140), .B(n2794), .S(n1789), .Z(n6331) );
  MUX2_X1 U7435 ( .A(n9141), .B(n2783), .S(n1789), .Z(n6332) );
  MUX2_X1 U7436 ( .A(n9142), .B(n2772), .S(n1789), .Z(n6333) );
  MUX2_X1 U7437 ( .A(n9143), .B(n2761), .S(n1789), .Z(n6334) );
  MUX2_X1 U7438 ( .A(n9144), .B(n2750), .S(n1789), .Z(n6335) );
  MUX2_X1 U7439 ( .A(n9145), .B(n2739), .S(n1789), .Z(n6336) );
  MUX2_X1 U7440 ( .A(n9146), .B(n2728), .S(n1789), .Z(n6337) );
  MUX2_X1 U7441 ( .A(n9147), .B(n2717), .S(n1789), .Z(n6338) );
  MUX2_X1 U7442 ( .A(n9148), .B(n2706), .S(n1789), .Z(n6339) );
  MUX2_X1 U7443 ( .A(n9149), .B(n2599), .S(n1789), .Z(n6340) );
  MUX2_X1 U7444 ( .A(n9150), .B(n2588), .S(n1790), .Z(n6341) );
  MUX2_X1 U7445 ( .A(n9151), .B(n2577), .S(n1790), .Z(n6342) );
  MUX2_X1 U7446 ( .A(n9152), .B(n2566), .S(n1790), .Z(n6343) );
  MUX2_X1 U7447 ( .A(n9153), .B(n2555), .S(n1790), .Z(n6344) );
  MUX2_X1 U7448 ( .A(n9154), .B(n2544), .S(n1790), .Z(n6345) );
  MUX2_X1 U7449 ( .A(n9155), .B(n1829), .S(n1790), .Z(n6346) );
  MUX2_X1 U7450 ( .A(n9156), .B(n1818), .S(n1790), .Z(n6347) );
  MUX2_X1 U7451 ( .A(n9157), .B(n1807), .S(n1790), .Z(n6348) );
endmodule


module FF_0 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n3, n4, n1, n2;

  DFF_X1 Q_reg ( .D(n4), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n3), .A2(n1), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n2), .ZN(n3) );
  INV_X1 U5 ( .A(EN), .ZN(n2) );
  INV_X1 U6 ( .A(RESET), .ZN(n1) );
endmodule


module regFFD_NBIT32_10 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_9 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_8 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_7 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT5_0 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  DFFR_X1 \Q_reg[2]  ( .D(n13), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n8) );
  DFFR_X1 \Q_reg[3]  ( .D(n14), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n9) );
  DFFR_X1 \Q_reg[0]  ( .D(n11), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n6) );
  DFFR_X1 \Q_reg[4]  ( .D(n15), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n10) );
  DFFR_X1 \Q_reg[1]  ( .D(n12), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n7) );
  OAI21_X1 U2 ( .B1(n7), .B2(ENABLE), .A(n2), .ZN(n12) );
  NAND2_X1 U3 ( .A1(D[1]), .A2(ENABLE), .ZN(n2) );
  OAI21_X1 U4 ( .B1(n8), .B2(ENABLE), .A(n3), .ZN(n13) );
  NAND2_X1 U5 ( .A1(D[2]), .A2(ENABLE), .ZN(n3) );
  OAI21_X1 U6 ( .B1(n9), .B2(ENABLE), .A(n4), .ZN(n14) );
  NAND2_X1 U7 ( .A1(D[3]), .A2(ENABLE), .ZN(n4) );
  OAI21_X1 U8 ( .B1(n10), .B2(ENABLE), .A(n5), .ZN(n15) );
  NAND2_X1 U9 ( .A1(D[4]), .A2(ENABLE), .ZN(n5) );
  OAI21_X1 U10 ( .B1(n6), .B2(ENABLE), .A(n1), .ZN(n11) );
  NAND2_X1 U11 ( .A1(ENABLE), .A2(D[0]), .ZN(n1) );
endmodule


module FF_7 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n1, n2, n5, n6;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n1), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n2), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n2) );
  INV_X1 U6 ( .A(RESET), .ZN(n1) );
endmodule


module regFFD_NBIT6_0 ( CK, RESET, ENABLE, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  DFFR_X1 \Q_reg[5]  ( .D(n18), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n12) );
  DFFR_X1 \Q_reg[2]  ( .D(n15), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n9) );
  DFFR_X1 \Q_reg[1]  ( .D(n14), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n8) );
  DFFR_X1 \Q_reg[0]  ( .D(n13), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n7) );
  DFFR_X1 \Q_reg[3]  ( .D(n16), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n10) );
  DFFR_X1 \Q_reg[4]  ( .D(n17), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n11) );
  OAI21_X1 U2 ( .B1(n9), .B2(ENABLE), .A(n3), .ZN(n15) );
  NAND2_X1 U3 ( .A1(D[2]), .A2(ENABLE), .ZN(n3) );
  OAI21_X1 U4 ( .B1(n8), .B2(ENABLE), .A(n2), .ZN(n14) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n2) );
  OAI21_X1 U6 ( .B1(n7), .B2(ENABLE), .A(n1), .ZN(n13) );
  NAND2_X1 U7 ( .A1(ENABLE), .A2(D[0]), .ZN(n1) );
  OAI21_X1 U8 ( .B1(n12), .B2(ENABLE), .A(n6), .ZN(n18) );
  NAND2_X1 U9 ( .A1(D[5]), .A2(ENABLE), .ZN(n6) );
  OAI21_X1 U10 ( .B1(n11), .B2(ENABLE), .A(n5), .ZN(n17) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n5) );
  OAI21_X1 U12 ( .B1(n10), .B2(ENABLE), .A(n4), .ZN(n16) );
  NAND2_X1 U13 ( .A1(D[3]), .A2(ENABLE), .ZN(n4) );
endmodule


module regFFD_NBIT32_6 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U6 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U7 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U8 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U9 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U10 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U11 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U12 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U13 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U14 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U15 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U16 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U17 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U18 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U19 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U20 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U21 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U22 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U23 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U24 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U25 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U26 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U27 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U28 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U29 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U30 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U31 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U32 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U33 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U34 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U35 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U36 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
  OAI21_X1 U37 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U38 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U39 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U40 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U41 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U42 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U43 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U44 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U45 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U46 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U47 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U48 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U49 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U50 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U51 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U52 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U53 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U54 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U55 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U56 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U57 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U58 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U59 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U60 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U61 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U62 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U63 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U64 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U65 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U66 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U67 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U68 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
endmodule


module IV_224 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_672 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_671 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_670 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_224 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_224 UIV ( .A(S), .Y(SB) );
  ND2_672 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_671 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_670 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_223 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_669 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_668 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_667 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_223 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_223 UIV ( .A(S), .Y(SB) );
  ND2_669 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_668 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_667 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_222 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_666 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_665 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_664 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_222 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_222 UIV ( .A(S), .Y(SB) );
  ND2_666 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_665 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_664 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_221 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_663 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_662 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_661 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_221 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_221 UIV ( .A(S), .Y(SB) );
  ND2_663 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_662 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_661 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_220 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_660 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_659 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_658 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_220 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_220 UIV ( .A(S), .Y(SB) );
  ND2_660 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_659 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_658 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_219 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_657 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_656 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_655 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_219 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_219 UIV ( .A(S), .Y(SB) );
  ND2_657 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_656 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_655 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_218 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_654 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_653 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_652 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_218 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_218 UIV ( .A(S), .Y(SB) );
  ND2_654 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_653 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_652 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_217 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_651 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_650 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_649 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_217 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_217 UIV ( .A(S), .Y(SB) );
  ND2_651 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_650 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_649 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_216 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_648 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_647 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_646 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_216 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_216 UIV ( .A(S), .Y(SB) );
  ND2_648 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_647 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_646 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_215 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_645 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_644 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_643 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_215 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_215 UIV ( .A(S), .Y(SB) );
  ND2_645 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_644 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_643 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_214 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_642 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_641 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_640 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_214 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_214 UIV ( .A(S), .Y(SB) );
  ND2_642 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_641 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_640 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_213 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_639 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_638 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_637 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_213 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_213 UIV ( .A(S), .Y(SB) );
  ND2_639 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_638 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_637 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_212 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_636 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_635 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_634 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_212 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_212 UIV ( .A(S), .Y(SB) );
  ND2_636 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_635 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_634 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_211 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_633 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_632 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_631 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_211 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_211 UIV ( .A(S), .Y(SB) );
  ND2_633 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_632 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_631 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_210 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_630 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_629 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_628 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_210 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_210 UIV ( .A(S), .Y(SB) );
  ND2_630 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_629 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_628 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_209 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_627 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_626 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_625 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_209 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_209 UIV ( .A(S), .Y(SB) );
  ND2_627 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_626 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_625 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_208 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_624 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_623 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_622 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_208 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_208 UIV ( .A(S), .Y(SB) );
  ND2_624 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_623 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_622 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_207 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_621 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_620 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_619 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_207 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_207 UIV ( .A(S), .Y(SB) );
  ND2_621 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_620 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_619 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_206 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_618 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_617 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_616 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_206 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_206 UIV ( .A(S), .Y(SB) );
  ND2_618 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_617 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_616 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_205 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_615 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_614 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_205 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_205 UIV ( .A(S), .Y(SB) );
  ND2_615 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_614 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_613 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_204 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_204 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_204 UIV ( .A(S), .Y(SB) );
  ND2_612 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_611 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_610 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_203 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_203 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_203 UIV ( .A(S), .Y(SB) );
  ND2_609 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_608 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_607 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_202 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_202 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_202 UIV ( .A(S), .Y(SB) );
  ND2_606 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_605 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_604 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_201 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_201 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_201 UIV ( .A(S), .Y(SB) );
  ND2_603 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_602 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_601 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_200 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_200 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_200 UIV ( .A(S), .Y(SB) );
  ND2_600 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_599 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_598 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_199 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_199 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_199 UIV ( .A(S), .Y(SB) );
  ND2_597 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_596 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_595 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_198 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_198 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_198 UIV ( .A(S), .Y(SB) );
  ND2_594 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_593 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_592 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_197 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_197 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_197 UIV ( .A(S), .Y(SB) );
  ND2_591 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_590 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_589 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_196 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_196 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_196 UIV ( .A(S), .Y(SB) );
  ND2_588 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_587 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_586 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_195 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_195 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_195 UIV ( .A(S), .Y(SB) );
  ND2_585 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_584 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_583 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_194 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_194 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_194 UIV ( .A(S), .Y(SB) );
  ND2_582 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_581 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_580 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_193 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_193 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_193 UIV ( .A(S), .Y(SB) );
  ND2_579 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_578 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_577 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_6 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_224 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_223 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_222 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_221 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_220 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_219 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_218 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_217 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_216 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_215 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_214 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_213 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_212 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_211 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_210 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_209 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_208 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_207 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_206 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_205 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_204 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_203 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_202 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_201 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_200 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_199 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_198 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_197 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_196 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_195 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_194 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_193 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_192 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_192 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_192 UIV ( .A(S), .Y(SB) );
  ND2_576 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_575 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_574 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_191 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_191 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_191 UIV ( .A(S), .Y(SB) );
  ND2_573 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_572 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_571 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_190 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_190 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_190 UIV ( .A(S), .Y(SB) );
  ND2_570 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_569 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_568 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_189 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_189 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_189 UIV ( .A(S), .Y(SB) );
  ND2_567 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_566 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_565 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_188 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_188 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_188 UIV ( .A(S), .Y(SB) );
  ND2_564 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_563 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_562 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_187 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_187 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_187 UIV ( .A(S), .Y(SB) );
  ND2_561 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_560 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_559 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_186 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_186 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_186 UIV ( .A(S), .Y(SB) );
  ND2_558 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_557 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_556 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_185 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_185 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_185 UIV ( .A(S), .Y(SB) );
  ND2_555 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_554 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_553 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_184 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_184 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_184 UIV ( .A(S), .Y(SB) );
  ND2_552 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_551 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_550 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_183 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_183 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_183 UIV ( .A(S), .Y(SB) );
  ND2_549 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_548 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_547 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_182 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_182 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_182 UIV ( .A(S), .Y(SB) );
  ND2_546 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_545 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_544 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_181 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_181 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_181 UIV ( .A(S), .Y(SB) );
  ND2_543 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_542 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_541 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_180 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_180 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_180 UIV ( .A(S), .Y(SB) );
  ND2_540 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_539 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_538 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_179 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_179 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_179 UIV ( .A(S), .Y(SB) );
  ND2_537 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_536 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_535 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_178 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_178 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_178 UIV ( .A(S), .Y(SB) );
  ND2_534 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_533 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_532 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_177 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_177 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_177 UIV ( .A(S), .Y(SB) );
  ND2_531 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_530 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_529 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_176 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_176 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_176 UIV ( .A(S), .Y(SB) );
  ND2_528 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_527 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_526 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_175 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_175 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_175 UIV ( .A(S), .Y(SB) );
  ND2_525 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_524 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_523 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_174 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_174 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_174 UIV ( .A(S), .Y(SB) );
  ND2_522 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_521 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_520 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_173 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_173 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_173 UIV ( .A(S), .Y(SB) );
  ND2_519 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_518 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_517 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_172 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_172 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_172 UIV ( .A(S), .Y(SB) );
  ND2_516 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_515 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_514 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_171 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_171 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_171 UIV ( .A(S), .Y(SB) );
  ND2_513 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_512 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_511 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_170 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_170 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_170 UIV ( .A(S), .Y(SB) );
  ND2_510 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_509 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_508 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_169 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_169 UIV ( .A(S), .Y(SB) );
  ND2_507 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_506 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_505 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_168 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_168 UIV ( .A(S), .Y(SB) );
  ND2_504 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_503 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_502 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_167 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_167 UIV ( .A(S), .Y(SB) );
  ND2_501 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_500 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_499 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_166 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_166 UIV ( .A(S), .Y(SB) );
  ND2_498 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_497 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_496 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_165 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_165 UIV ( .A(S), .Y(SB) );
  ND2_495 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_494 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_493 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_164 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_164 UIV ( .A(S), .Y(SB) );
  ND2_492 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_491 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_490 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_163 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_163 UIV ( .A(S), .Y(SB) );
  ND2_489 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_488 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_487 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_162 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_162 UIV ( .A(S), .Y(SB) );
  ND2_486 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_485 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_484 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_161 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_161 UIV ( .A(S), .Y(SB) );
  ND2_483 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_482 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_481 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_5 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_192 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_191 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_190 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_189 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_188 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_187 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_186 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_185 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_184 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_183 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_182 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_181 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_180 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_179 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_178 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_177 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_176 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_175 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_174 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_173 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_172 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_171 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_170 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_169 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_168 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_167 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_166 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_165 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_164 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_163 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_162 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_161 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module logic_N32 ( .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , 
        \FUNC[1] , \FUNC[0] }), DATA1, DATA2, OUT_ALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUT_ALU;
  input \FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155;
  wire   [5:0] FUNC;

  NAND3_X1 U173 ( .A1(n140), .A2(n154), .A3(FUNC[4]), .ZN(n136) );
  BUF_X1 U2 ( .A(n71), .Z(n12) );
  BUF_X1 U3 ( .A(n71), .Z(n13) );
  BUF_X1 U4 ( .A(n71), .Z(n14) );
  BUF_X1 U5 ( .A(n72), .Z(n5) );
  BUF_X1 U6 ( .A(n72), .Z(n4) );
  BUF_X1 U7 ( .A(n73), .Z(n2) );
  BUF_X1 U8 ( .A(n73), .Z(n1) );
  BUF_X1 U9 ( .A(n72), .Z(n7) );
  BUF_X1 U10 ( .A(n72), .Z(n8) );
  OAI22_X1 U11 ( .A1(n86), .A2(n53), .B1(n87), .B2(n21), .ZN(OUT_ALU[31]) );
  AOI21_X1 U12 ( .B1(n13), .B2(n53), .A(n7), .ZN(n87) );
  AOI221_X1 U13 ( .B1(n12), .B2(n21), .C1(DATA1[31]), .C2(n3), .A(n6), .ZN(n86) );
  INV_X1 U14 ( .A(DATA2[31]), .ZN(n53) );
  OAI22_X1 U15 ( .A1(n88), .A2(n54), .B1(n89), .B2(n22), .ZN(OUT_ALU[30]) );
  AOI21_X1 U16 ( .B1(n13), .B2(n54), .A(n7), .ZN(n89) );
  AOI221_X1 U17 ( .B1(n12), .B2(n22), .C1(DATA1[30]), .C2(n2), .A(n6), .ZN(n88) );
  INV_X1 U18 ( .A(DATA2[30]), .ZN(n54) );
  OAI22_X1 U19 ( .A1(n92), .A2(n55), .B1(n93), .B2(n23), .ZN(OUT_ALU[29]) );
  AOI21_X1 U20 ( .B1(n13), .B2(n55), .A(n7), .ZN(n93) );
  AOI221_X1 U21 ( .B1(n12), .B2(n23), .C1(DATA1[29]), .C2(n2), .A(n6), .ZN(n92) );
  INV_X1 U22 ( .A(DATA2[29]), .ZN(n55) );
  OAI22_X1 U23 ( .A1(n94), .A2(n56), .B1(n95), .B2(n24), .ZN(OUT_ALU[28]) );
  AOI21_X1 U24 ( .B1(n13), .B2(n56), .A(n7), .ZN(n95) );
  AOI221_X1 U25 ( .B1(n12), .B2(n24), .C1(DATA1[28]), .C2(n2), .A(n6), .ZN(n94) );
  INV_X1 U26 ( .A(DATA2[28]), .ZN(n56) );
  OAI22_X1 U27 ( .A1(n96), .A2(n57), .B1(n97), .B2(n25), .ZN(OUT_ALU[27]) );
  AOI21_X1 U28 ( .B1(n13), .B2(n57), .A(n7), .ZN(n97) );
  AOI221_X1 U29 ( .B1(n12), .B2(n25), .C1(DATA1[27]), .C2(n2), .A(n6), .ZN(n96) );
  INV_X1 U30 ( .A(DATA2[27]), .ZN(n57) );
  OAI22_X1 U31 ( .A1(n98), .A2(n58), .B1(n99), .B2(n26), .ZN(OUT_ALU[26]) );
  AOI21_X1 U32 ( .B1(n13), .B2(n58), .A(n7), .ZN(n99) );
  AOI221_X1 U33 ( .B1(n11), .B2(n26), .C1(DATA1[26]), .C2(n2), .A(n5), .ZN(n98) );
  INV_X1 U34 ( .A(DATA2[26]), .ZN(n58) );
  OAI22_X1 U35 ( .A1(n100), .A2(n59), .B1(n101), .B2(n27), .ZN(OUT_ALU[25]) );
  AOI21_X1 U36 ( .B1(n13), .B2(n59), .A(n7), .ZN(n101) );
  AOI221_X1 U37 ( .B1(n12), .B2(n27), .C1(DATA1[25]), .C2(n2), .A(n6), .ZN(
        n100) );
  INV_X1 U38 ( .A(DATA2[25]), .ZN(n59) );
  OAI22_X1 U39 ( .A1(n102), .A2(n60), .B1(n103), .B2(n28), .ZN(OUT_ALU[24]) );
  AOI21_X1 U40 ( .B1(n14), .B2(n60), .A(n7), .ZN(n103) );
  AOI221_X1 U41 ( .B1(n12), .B2(n28), .C1(DATA1[24]), .C2(n2), .A(n6), .ZN(
        n102) );
  INV_X1 U42 ( .A(DATA2[24]), .ZN(n60) );
  OAI22_X1 U43 ( .A1(n104), .A2(n61), .B1(n105), .B2(n29), .ZN(OUT_ALU[23]) );
  AOI21_X1 U44 ( .B1(n14), .B2(n61), .A(n8), .ZN(n105) );
  AOI221_X1 U45 ( .B1(n11), .B2(n29), .C1(DATA1[23]), .C2(n2), .A(n5), .ZN(
        n104) );
  INV_X1 U46 ( .A(DATA2[23]), .ZN(n61) );
  OAI22_X1 U47 ( .A1(n106), .A2(n62), .B1(n107), .B2(n30), .ZN(OUT_ALU[22]) );
  AOI21_X1 U48 ( .B1(n14), .B2(n62), .A(n8), .ZN(n107) );
  AOI221_X1 U49 ( .B1(n11), .B2(n30), .C1(DATA1[22]), .C2(n2), .A(n5), .ZN(
        n106) );
  INV_X1 U50 ( .A(DATA2[22]), .ZN(n62) );
  OAI22_X1 U51 ( .A1(n108), .A2(n63), .B1(n109), .B2(n31), .ZN(OUT_ALU[21]) );
  AOI21_X1 U52 ( .B1(n14), .B2(n63), .A(n8), .ZN(n109) );
  AOI221_X1 U53 ( .B1(n11), .B2(n31), .C1(DATA1[21]), .C2(n2), .A(n5), .ZN(
        n108) );
  INV_X1 U54 ( .A(DATA2[21]), .ZN(n63) );
  OAI22_X1 U55 ( .A1(n110), .A2(n64), .B1(n111), .B2(n32), .ZN(OUT_ALU[20]) );
  AOI21_X1 U56 ( .B1(n14), .B2(n64), .A(n8), .ZN(n111) );
  AOI221_X1 U57 ( .B1(n11), .B2(n32), .C1(DATA1[20]), .C2(n2), .A(n5), .ZN(
        n110) );
  INV_X1 U58 ( .A(DATA2[20]), .ZN(n64) );
  OAI22_X1 U59 ( .A1(n114), .A2(n65), .B1(n115), .B2(n33), .ZN(OUT_ALU[19]) );
  AOI21_X1 U60 ( .B1(n14), .B2(n65), .A(n8), .ZN(n115) );
  AOI221_X1 U61 ( .B1(n11), .B2(n33), .C1(DATA1[19]), .C2(n1), .A(n5), .ZN(
        n114) );
  INV_X1 U62 ( .A(DATA2[19]), .ZN(n65) );
  OAI22_X1 U63 ( .A1(n116), .A2(n66), .B1(n117), .B2(n34), .ZN(OUT_ALU[18]) );
  AOI21_X1 U64 ( .B1(n14), .B2(n66), .A(n8), .ZN(n117) );
  AOI221_X1 U65 ( .B1(n11), .B2(n34), .C1(DATA1[18]), .C2(n1), .A(n5), .ZN(
        n116) );
  INV_X1 U66 ( .A(DATA2[18]), .ZN(n66) );
  OAI22_X1 U67 ( .A1(n118), .A2(n67), .B1(n119), .B2(n35), .ZN(OUT_ALU[17]) );
  AOI21_X1 U68 ( .B1(n14), .B2(n67), .A(n8), .ZN(n119) );
  AOI221_X1 U69 ( .B1(n11), .B2(n35), .C1(DATA1[17]), .C2(n1), .A(n5), .ZN(
        n118) );
  INV_X1 U70 ( .A(DATA2[17]), .ZN(n67) );
  OAI22_X1 U71 ( .A1(n120), .A2(n68), .B1(n121), .B2(n36), .ZN(OUT_ALU[16]) );
  AOI21_X1 U72 ( .B1(n14), .B2(n68), .A(n8), .ZN(n121) );
  AOI221_X1 U73 ( .B1(n10), .B2(n36), .C1(DATA1[16]), .C2(n1), .A(n4), .ZN(
        n120) );
  INV_X1 U74 ( .A(DATA2[16]), .ZN(n68) );
  OAI22_X1 U75 ( .A1(n122), .A2(n141), .B1(n123), .B2(n37), .ZN(OUT_ALU[15])
         );
  AOI21_X1 U76 ( .B1(n14), .B2(n141), .A(n8), .ZN(n123) );
  AOI221_X1 U77 ( .B1(n10), .B2(n37), .C1(DATA1[15]), .C2(n1), .A(n4), .ZN(
        n122) );
  INV_X1 U78 ( .A(DATA2[15]), .ZN(n141) );
  OAI22_X1 U79 ( .A1(n124), .A2(n142), .B1(n125), .B2(n38), .ZN(OUT_ALU[14])
         );
  AOI21_X1 U80 ( .B1(n14), .B2(n142), .A(n8), .ZN(n125) );
  AOI221_X1 U81 ( .B1(n10), .B2(n38), .C1(DATA1[14]), .C2(n1), .A(n4), .ZN(
        n124) );
  INV_X1 U82 ( .A(DATA2[14]), .ZN(n142) );
  OAI22_X1 U83 ( .A1(n126), .A2(n143), .B1(n127), .B2(n39), .ZN(OUT_ALU[13])
         );
  AOI21_X1 U84 ( .B1(n15), .B2(n143), .A(n8), .ZN(n127) );
  AOI221_X1 U85 ( .B1(n10), .B2(n39), .C1(DATA1[13]), .C2(n1), .A(n4), .ZN(
        n126) );
  INV_X1 U86 ( .A(DATA2[13]), .ZN(n143) );
  OAI22_X1 U87 ( .A1(n128), .A2(n144), .B1(n129), .B2(n40), .ZN(OUT_ALU[12])
         );
  AOI21_X1 U88 ( .B1(n15), .B2(n144), .A(n8), .ZN(n129) );
  AOI221_X1 U89 ( .B1(n10), .B2(n40), .C1(DATA1[12]), .C2(n1), .A(n4), .ZN(
        n128) );
  INV_X1 U90 ( .A(DATA2[12]), .ZN(n144) );
  OAI22_X1 U91 ( .A1(n130), .A2(n145), .B1(n131), .B2(n41), .ZN(OUT_ALU[11])
         );
  AOI21_X1 U92 ( .B1(n15), .B2(n145), .A(n9), .ZN(n131) );
  AOI221_X1 U93 ( .B1(n10), .B2(n41), .C1(DATA1[11]), .C2(n1), .A(n4), .ZN(
        n130) );
  INV_X1 U94 ( .A(DATA2[11]), .ZN(n145) );
  OAI22_X1 U95 ( .A1(n132), .A2(n146), .B1(n133), .B2(n42), .ZN(OUT_ALU[10])
         );
  AOI21_X1 U96 ( .B1(n15), .B2(n146), .A(n9), .ZN(n133) );
  AOI221_X1 U97 ( .B1(n10), .B2(n42), .C1(DATA1[10]), .C2(n1), .A(n4), .ZN(
        n132) );
  INV_X1 U98 ( .A(DATA2[10]), .ZN(n146) );
  OAI22_X1 U99 ( .A1(n69), .A2(n147), .B1(n70), .B2(n43), .ZN(OUT_ALU[9]) );
  AOI21_X1 U100 ( .B1(n13), .B2(n147), .A(n7), .ZN(n70) );
  AOI221_X1 U101 ( .B1(n10), .B2(n43), .C1(n3), .C2(DATA1[9]), .A(n4), .ZN(n69) );
  INV_X1 U102 ( .A(DATA2[9]), .ZN(n147) );
  OAI22_X1 U103 ( .A1(n74), .A2(n148), .B1(n75), .B2(n44), .ZN(OUT_ALU[8]) );
  AOI21_X1 U104 ( .B1(n12), .B2(n148), .A(n6), .ZN(n75) );
  AOI221_X1 U105 ( .B1(n10), .B2(n44), .C1(DATA1[8]), .C2(n3), .A(n4), .ZN(n74) );
  INV_X1 U106 ( .A(DATA2[8]), .ZN(n148) );
  OAI22_X1 U107 ( .A1(n76), .A2(n149), .B1(n77), .B2(n45), .ZN(OUT_ALU[7]) );
  AOI21_X1 U108 ( .B1(n13), .B2(n149), .A(n7), .ZN(n77) );
  AOI221_X1 U109 ( .B1(n10), .B2(n45), .C1(DATA1[7]), .C2(n3), .A(n4), .ZN(n76) );
  INV_X1 U110 ( .A(DATA2[7]), .ZN(n149) );
  OAI22_X1 U111 ( .A1(n78), .A2(n150), .B1(n79), .B2(n46), .ZN(OUT_ALU[6]) );
  AOI21_X1 U112 ( .B1(n12), .B2(n150), .A(n6), .ZN(n79) );
  AOI221_X1 U113 ( .B1(n10), .B2(n46), .C1(DATA1[6]), .C2(n3), .A(n4), .ZN(n78) );
  INV_X1 U114 ( .A(DATA2[6]), .ZN(n150) );
  OAI22_X1 U115 ( .A1(n80), .A2(n151), .B1(n81), .B2(n47), .ZN(OUT_ALU[5]) );
  AOI21_X1 U116 ( .B1(n12), .B2(n151), .A(n6), .ZN(n81) );
  AOI221_X1 U117 ( .B1(n11), .B2(n47), .C1(DATA1[5]), .C2(n3), .A(n5), .ZN(n80) );
  INV_X1 U118 ( .A(DATA2[5]), .ZN(n151) );
  OAI22_X1 U119 ( .A1(n82), .A2(n20), .B1(n83), .B2(n48), .ZN(OUT_ALU[4]) );
  AOI21_X1 U120 ( .B1(n13), .B2(n20), .A(n7), .ZN(n83) );
  AOI221_X1 U121 ( .B1(n11), .B2(n48), .C1(DATA1[4]), .C2(n3), .A(n5), .ZN(n82) );
  OAI22_X1 U122 ( .A1(n84), .A2(n19), .B1(n85), .B2(n49), .ZN(OUT_ALU[3]) );
  AOI21_X1 U123 ( .B1(n13), .B2(n19), .A(n7), .ZN(n85) );
  AOI221_X1 U124 ( .B1(n11), .B2(n49), .C1(DATA1[3]), .C2(n3), .A(n5), .ZN(n84) );
  OAI22_X1 U125 ( .A1(n90), .A2(n18), .B1(n91), .B2(n50), .ZN(OUT_ALU[2]) );
  AOI21_X1 U126 ( .B1(n13), .B2(n18), .A(n7), .ZN(n91) );
  AOI221_X1 U127 ( .B1(n12), .B2(n50), .C1(DATA1[2]), .C2(n2), .A(n6), .ZN(n90) );
  OAI22_X1 U128 ( .A1(n112), .A2(n17), .B1(n113), .B2(n51), .ZN(OUT_ALU[1]) );
  AOI21_X1 U129 ( .B1(n14), .B2(n17), .A(n8), .ZN(n113) );
  AOI221_X1 U130 ( .B1(n11), .B2(n51), .C1(DATA1[1]), .C2(n1), .A(n5), .ZN(
        n112) );
  OAI22_X1 U131 ( .A1(n134), .A2(n16), .B1(n135), .B2(n52), .ZN(OUT_ALU[0]) );
  AOI21_X1 U132 ( .B1(n12), .B2(n16), .A(n6), .ZN(n135) );
  AOI221_X1 U133 ( .B1(n10), .B2(n52), .C1(DATA1[0]), .C2(n1), .A(n4), .ZN(
        n134) );
  BUF_X1 U134 ( .A(n72), .Z(n6) );
  BUF_X1 U135 ( .A(n71), .Z(n11) );
  BUF_X1 U136 ( .A(n71), .Z(n10) );
  BUF_X1 U137 ( .A(n73), .Z(n3) );
  INV_X1 U138 ( .A(DATA1[12]), .ZN(n40) );
  INV_X1 U139 ( .A(DATA1[23]), .ZN(n29) );
  INV_X1 U140 ( .A(DATA1[14]), .ZN(n38) );
  INV_X1 U141 ( .A(DATA1[17]), .ZN(n35) );
  INV_X1 U142 ( .A(DATA1[21]), .ZN(n31) );
  INV_X1 U143 ( .A(DATA1[13]), .ZN(n39) );
  INV_X1 U144 ( .A(DATA1[22]), .ZN(n30) );
  INV_X1 U145 ( .A(DATA1[16]), .ZN(n36) );
  INV_X1 U146 ( .A(DATA1[15]), .ZN(n37) );
  INV_X1 U147 ( .A(DATA1[9]), .ZN(n43) );
  INV_X1 U148 ( .A(DATA1[11]), .ZN(n41) );
  INV_X1 U149 ( .A(DATA1[10]), .ZN(n42) );
  INV_X1 U150 ( .A(DATA1[8]), .ZN(n44) );
  INV_X1 U151 ( .A(DATA1[7]), .ZN(n45) );
  INV_X1 U152 ( .A(DATA1[2]), .ZN(n50) );
  INV_X1 U153 ( .A(DATA1[3]), .ZN(n49) );
  INV_X1 U154 ( .A(DATA1[28]), .ZN(n24) );
  INV_X1 U155 ( .A(DATA1[27]), .ZN(n25) );
  INV_X1 U156 ( .A(DATA1[26]), .ZN(n26) );
  INV_X1 U157 ( .A(DATA1[25]), .ZN(n27) );
  INV_X1 U158 ( .A(DATA1[24]), .ZN(n28) );
  INV_X1 U159 ( .A(DATA1[18]), .ZN(n34) );
  INV_X1 U160 ( .A(DATA1[0]), .ZN(n52) );
  INV_X1 U161 ( .A(DATA1[29]), .ZN(n23) );
  INV_X1 U162 ( .A(DATA1[4]), .ZN(n48) );
  INV_X1 U163 ( .A(DATA1[6]), .ZN(n46) );
  INV_X1 U164 ( .A(DATA1[31]), .ZN(n21) );
  INV_X1 U165 ( .A(DATA1[19]), .ZN(n33) );
  INV_X1 U166 ( .A(DATA1[20]), .ZN(n32) );
  INV_X1 U167 ( .A(DATA1[1]), .ZN(n51) );
  INV_X1 U168 ( .A(DATA1[5]), .ZN(n47) );
  INV_X1 U169 ( .A(DATA1[30]), .ZN(n22) );
  OAI21_X1 U170 ( .B1(FUNC[0]), .B2(n136), .A(n137), .ZN(n72) );
  OR3_X1 U171 ( .A1(n138), .A2(FUNC[3]), .A3(n155), .ZN(n137) );
  NAND4_X1 U172 ( .A1(FUNC[2]), .A2(FUNC[1]), .A3(n153), .A4(n152), .ZN(n138)
         );
  INV_X1 U174 ( .A(FUNC[5]), .ZN(n152) );
  NOR3_X1 U175 ( .A1(FUNC[2]), .A2(FUNC[5]), .A3(FUNC[1]), .ZN(n140) );
  AOI21_X1 U176 ( .B1(n155), .B2(FUNC[3]), .A(n138), .ZN(n73) );
  INV_X1 U177 ( .A(FUNC[3]), .ZN(n154) );
  NAND2_X1 U178 ( .A1(n136), .A2(n139), .ZN(n71) );
  NAND4_X1 U179 ( .A1(FUNC[3]), .A2(n140), .A3(n155), .A4(n153), .ZN(n139) );
  INV_X1 U180 ( .A(FUNC[0]), .ZN(n155) );
  INV_X1 U181 ( .A(FUNC[4]), .ZN(n153) );
  CLKBUF_X1 U182 ( .A(n72), .Z(n9) );
  CLKBUF_X1 U183 ( .A(n71), .Z(n15) );
  INV_X1 U184 ( .A(DATA2[0]), .ZN(n16) );
  INV_X1 U185 ( .A(DATA2[1]), .ZN(n17) );
  INV_X1 U186 ( .A(DATA2[2]), .ZN(n18) );
  INV_X1 U187 ( .A(DATA2[3]), .ZN(n19) );
  INV_X1 U188 ( .A(DATA2[4]), .ZN(n20) );
endmodule


module comparator ( DATA1, DATA2i, .tipo({\tipo[5] , \tipo[4] , \tipo[3] , 
        \tipo[2] , \tipo[1] , \tipo[0] }), OUTALU );
  input [31:0] DATA1;
  output [31:0] OUTALU;
  input DATA2i, \tipo[5] , \tipo[4] , \tipo[3] , \tipo[2] , \tipo[1] ,
         \tipo[0] ;
  wire   N57, N58, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [5:0] tipo;
  assign OUTALU[31] = 1'b0;
  assign OUTALU[30] = 1'b0;
  assign OUTALU[29] = 1'b0;
  assign OUTALU[28] = 1'b0;
  assign OUTALU[27] = 1'b0;
  assign OUTALU[26] = 1'b0;
  assign OUTALU[25] = 1'b0;
  assign OUTALU[24] = 1'b0;
  assign OUTALU[23] = 1'b0;
  assign OUTALU[22] = 1'b0;
  assign OUTALU[21] = 1'b0;
  assign OUTALU[20] = 1'b0;
  assign OUTALU[19] = 1'b0;
  assign OUTALU[18] = 1'b0;
  assign OUTALU[17] = 1'b0;
  assign OUTALU[16] = 1'b0;
  assign OUTALU[15] = 1'b0;
  assign OUTALU[14] = 1'b0;
  assign OUTALU[13] = 1'b0;
  assign OUTALU[12] = 1'b0;
  assign OUTALU[11] = 1'b0;
  assign OUTALU[10] = 1'b0;
  assign OUTALU[9] = 1'b0;
  assign OUTALU[8] = 1'b0;
  assign OUTALU[7] = 1'b0;
  assign OUTALU[6] = 1'b0;
  assign OUTALU[5] = 1'b0;
  assign OUTALU[4] = 1'b0;
  assign OUTALU[3] = 1'b0;
  assign OUTALU[2] = 1'b0;
  assign OUTALU[1] = 1'b0;

  DLH_X1 \OUTALU_reg[0]  ( .G(N57), .D(N58), .Q(OUTALU[0]) );
  NAND3_X1 U80 ( .A1(n48), .A2(n7), .A3(tipo[5]), .ZN(n37) );
  NAND3_X1 U81 ( .A1(tipo[3]), .A2(n48), .A3(tipo[5]), .ZN(n43) );
  NAND3_X1 U82 ( .A1(tipo[3]), .A2(n49), .A3(tipo[1]), .ZN(n46) );
  NAND3_X1 U83 ( .A1(n48), .A2(n5), .A3(tipo[3]), .ZN(n42) );
  INV_X1 U33 ( .A(n19), .ZN(n1) );
  NOR4_X1 U34 ( .A1(DATA1[23]), .A2(DATA1[22]), .A3(DATA1[21]), .A4(DATA1[20]), 
        .ZN(n27) );
  NOR4_X1 U35 ( .A1(DATA1[9]), .A2(DATA1[8]), .A3(DATA1[7]), .A4(DATA1[6]), 
        .ZN(n31) );
  NOR4_X1 U36 ( .A1(DATA1[16]), .A2(DATA1[15]), .A3(DATA1[14]), .A4(DATA1[13]), 
        .ZN(n25) );
  NOR2_X1 U37 ( .A1(n22), .A2(n23), .ZN(n19) );
  NAND4_X1 U38 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n22) );
  NAND4_X1 U39 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n23) );
  NOR4_X1 U40 ( .A1(DATA1[27]), .A2(DATA1[26]), .A3(DATA1[25]), .A4(DATA1[24]), 
        .ZN(n28) );
  INV_X1 U41 ( .A(DATA2i), .ZN(n2) );
  NOR4_X1 U42 ( .A1(DATA1[1]), .A2(DATA1[19]), .A3(DATA1[18]), .A4(DATA1[17]), 
        .ZN(n26) );
  NOR4_X1 U43 ( .A1(DATA1[5]), .A2(DATA1[4]), .A3(DATA1[3]), .A4(DATA1[31]), 
        .ZN(n30) );
  NOR4_X1 U44 ( .A1(DATA1[30]), .A2(DATA1[2]), .A3(DATA1[29]), .A4(DATA1[28]), 
        .ZN(n29) );
  OAI221_X1 U45 ( .B1(n39), .B2(n36), .C1(n34), .C2(n40), .A(n4), .ZN(n21) );
  INV_X1 U46 ( .A(n41), .ZN(n4) );
  AOI211_X1 U47 ( .C1(n37), .C2(n42), .A(n9), .B(n11), .ZN(n41) );
  NOR4_X1 U48 ( .A1(DATA1[12]), .A2(DATA1[11]), .A3(DATA1[10]), .A4(DATA1[0]), 
        .ZN(n24) );
  OAI22_X1 U49 ( .A1(n39), .A2(n40), .B1(n34), .B2(n42), .ZN(n18) );
  OAI22_X1 U50 ( .A1(n42), .A2(n39), .B1(n40), .B2(n38), .ZN(n16) );
  OAI21_X1 U51 ( .B1(n33), .B2(n34), .A(n6), .ZN(n20) );
  INV_X1 U52 ( .A(n35), .ZN(n6) );
  AOI21_X1 U53 ( .B1(n36), .B2(n37), .A(n38), .ZN(n35) );
  NAND2_X1 U54 ( .A1(n11), .A2(n9), .ZN(n38) );
  OAI211_X1 U55 ( .C1(n12), .C2(n2), .A(n13), .B(n14), .ZN(N58) );
  OAI21_X1 U56 ( .B1(n17), .B2(n18), .A(n19), .ZN(n13) );
  AOI21_X1 U57 ( .B1(n20), .B2(n1), .A(n21), .ZN(n12) );
  AOI22_X1 U58 ( .A1(n15), .A2(n2), .B1(n16), .B2(n1), .ZN(n14) );
  OR4_X1 U59 ( .A1(n16), .A2(n15), .A3(n32), .A4(n20), .ZN(N57) );
  OR2_X1 U60 ( .A1(n17), .A2(n21), .ZN(n32) );
  AND2_X1 U61 ( .A1(n43), .A2(n37), .ZN(n33) );
  NAND4_X1 U62 ( .A1(tipo[4]), .A2(tipo[2]), .A3(n7), .A4(n5), .ZN(n40) );
  OAI221_X1 U63 ( .B1(n46), .B2(n47), .C1(n33), .C2(n39), .A(n3), .ZN(n15) );
  INV_X1 U64 ( .A(n18), .ZN(n3) );
  NAND2_X1 U65 ( .A1(tipo[0]), .A2(tipo[2]), .ZN(n47) );
  NAND4_X1 U66 ( .A1(tipo[5]), .A2(tipo[4]), .A3(n8), .A4(n7), .ZN(n36) );
  INV_X1 U67 ( .A(tipo[2]), .ZN(n8) );
  NAND2_X1 U68 ( .A1(tipo[1]), .A2(n11), .ZN(n34) );
  NAND2_X1 U69 ( .A1(tipo[0]), .A2(n9), .ZN(n39) );
  INV_X1 U70 ( .A(tipo[3]), .ZN(n7) );
  NOR2_X1 U71 ( .A1(tipo[4]), .A2(tipo[2]), .ZN(n48) );
  OAI21_X1 U72 ( .B1(n43), .B2(n38), .A(n44), .ZN(n17) );
  NAND4_X1 U73 ( .A1(tipo[4]), .A2(tipo[2]), .A3(n45), .A4(n10), .ZN(n44) );
  INV_X1 U74 ( .A(n34), .ZN(n10) );
  NOR2_X1 U75 ( .A1(tipo[5]), .A2(n7), .ZN(n45) );
  XNOR2_X1 U76 ( .A(n5), .B(tipo[4]), .ZN(n49) );
  INV_X1 U77 ( .A(tipo[1]), .ZN(n9) );
  INV_X1 U78 ( .A(tipo[5]), .ZN(n5) );
  INV_X1 U79 ( .A(tipo[0]), .ZN(n11) );
endmodule


module SHIFTER_GENERIC_N32_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[5][31] , \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] ,
         \ML_int[5][15] , \ML_int[5][14] , \ML_int[5][13] , \ML_int[5][12] ,
         \ML_int[5][11] , \ML_int[5][10] , \ML_int[5][9] , \ML_int[5][8] ,
         \ML_int[5][7] , \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] ,
         \ML_int[5][3] , \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  assign B[31] = \ML_int[5][31] ;
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[8] = \ML_int[5][8] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n11), .Z(
        \ML_int[5][31] ) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n11), .Z(
        \ML_int[5][30] ) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n11), .Z(
        \ML_int[5][29] ) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n11), .Z(
        \ML_int[5][28] ) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n11), .Z(
        \ML_int[5][27] ) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n11), .Z(
        \ML_int[5][26] ) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n11), .Z(
        \ML_int[5][25] ) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n11), .Z(
        \ML_int[5][24] ) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(n13), .S(n11), .Z(\ML_int[5][23] )
         );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(n14), .S(n11), .Z(\ML_int[5][22] )
         );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(n15), .S(n11), .Z(\ML_int[5][21] )
         );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(n16), .S(n11), .Z(\ML_int[5][20] )
         );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(n17), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(n18), .S(n11), .Z(\ML_int[5][18] )
         );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(n19), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(n20), .S(SH[4]), .Z(
        \ML_int[5][16] ) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n9), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n9), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n9), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n9), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n9), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n9), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n9), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n9), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n9), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n9), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(SH[3]), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n9), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n9), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n9), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n9), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n9), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n9), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n9), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n9), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n9), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n9), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n9), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n9), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n9), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n7), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n7), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n7), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n7), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n7), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n7), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(SH[2]), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n7), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(SH[2]), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n7), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(SH[2]), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n7), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n7), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n7), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n7), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n7), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n7), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n7), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n7), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n7), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n7), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n7), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n7), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n7), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n7), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n7), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n5), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n4), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n5), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n4), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n5), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n4), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n5), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n5), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n5), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n5), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n5), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n5), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n5), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n5), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n5), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n5), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n5), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n5), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n4), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n4), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n4), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n4), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n4), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n4), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n4), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n4), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n4), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n4), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n4), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n4), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n2), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n1), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n2), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n1), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n2), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n1), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n2), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n2), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n2), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n2), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n2), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n2), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n2), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n2), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n2), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n2), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n2), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n2), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n2), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n1), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n1), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n1), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n1), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n1), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n1), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n1), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n1), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n1), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n1), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n1), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n1), .Z(\ML_int[1][1] ) );
  INV_X1 U3 ( .A(n12), .ZN(n11) );
  INV_X1 U4 ( .A(n21), .ZN(n13) );
  INV_X1 U5 ( .A(n22), .ZN(n14) );
  INV_X1 U6 ( .A(n23), .ZN(n15) );
  INV_X1 U7 ( .A(n24), .ZN(n16) );
  INV_X1 U8 ( .A(n25), .ZN(n17) );
  INV_X1 U9 ( .A(n26), .ZN(n18) );
  INV_X1 U10 ( .A(n27), .ZN(n19) );
  INV_X1 U11 ( .A(n28), .ZN(n20) );
  INV_X1 U12 ( .A(n8), .ZN(n7) );
  INV_X1 U13 ( .A(n6), .ZN(n5) );
  INV_X1 U14 ( .A(n6), .ZN(n4) );
  INV_X1 U15 ( .A(n3), .ZN(n2) );
  INV_X1 U16 ( .A(n3), .ZN(n1) );
  INV_X1 U17 ( .A(SH[1]), .ZN(n6) );
  INV_X1 U18 ( .A(SH[0]), .ZN(n3) );
  INV_X1 U19 ( .A(SH[3]), .ZN(n10) );
  INV_X1 U20 ( .A(SH[2]), .ZN(n8) );
  INV_X1 U21 ( .A(n10), .ZN(n9) );
  INV_X1 U22 ( .A(SH[4]), .ZN(n12) );
  AND2_X1 U23 ( .A1(\ML_int[4][9] ), .A2(n12), .ZN(\ML_int[5][9] ) );
  AND2_X1 U24 ( .A1(\ML_int[4][8] ), .A2(n12), .ZN(\ML_int[5][8] ) );
  NOR2_X1 U25 ( .A1(n11), .A2(n21), .ZN(\ML_int[5][7] ) );
  NOR2_X1 U26 ( .A1(SH[4]), .A2(n22), .ZN(\ML_int[5][6] ) );
  NOR2_X1 U27 ( .A1(n11), .A2(n23), .ZN(\ML_int[5][5] ) );
  NOR2_X1 U28 ( .A1(SH[4]), .A2(n24), .ZN(\ML_int[5][4] ) );
  NOR2_X1 U29 ( .A1(n11), .A2(n25), .ZN(\ML_int[5][3] ) );
  NOR2_X1 U30 ( .A1(SH[4]), .A2(n26), .ZN(\ML_int[5][2] ) );
  NOR2_X1 U31 ( .A1(n11), .A2(n27), .ZN(\ML_int[5][1] ) );
  AND2_X1 U32 ( .A1(\ML_int[4][15] ), .A2(n12), .ZN(\ML_int[5][15] ) );
  AND2_X1 U33 ( .A1(\ML_int[4][14] ), .A2(n12), .ZN(\ML_int[5][14] ) );
  AND2_X1 U34 ( .A1(\ML_int[4][13] ), .A2(n12), .ZN(\ML_int[5][13] ) );
  AND2_X1 U35 ( .A1(\ML_int[4][12] ), .A2(n12), .ZN(\ML_int[5][12] ) );
  AND2_X1 U36 ( .A1(\ML_int[4][11] ), .A2(n12), .ZN(\ML_int[5][11] ) );
  AND2_X1 U37 ( .A1(\ML_int[4][10] ), .A2(n12), .ZN(\ML_int[5][10] ) );
  NOR2_X1 U38 ( .A1(SH[4]), .A2(n28), .ZN(\ML_int[5][0] ) );
  NAND2_X1 U39 ( .A1(\ML_int[3][7] ), .A2(n10), .ZN(n21) );
  NAND2_X1 U40 ( .A1(\ML_int[3][6] ), .A2(n10), .ZN(n22) );
  NAND2_X1 U41 ( .A1(\ML_int[3][5] ), .A2(n10), .ZN(n23) );
  NAND2_X1 U42 ( .A1(\ML_int[3][4] ), .A2(n10), .ZN(n24) );
  NAND2_X1 U43 ( .A1(\ML_int[3][3] ), .A2(n10), .ZN(n25) );
  NAND2_X1 U44 ( .A1(\ML_int[3][2] ), .A2(n10), .ZN(n26) );
  NAND2_X1 U45 ( .A1(\ML_int[3][1] ), .A2(n10), .ZN(n27) );
  NAND2_X1 U46 ( .A1(\ML_int[3][0] ), .A2(n10), .ZN(n28) );
  AND2_X1 U47 ( .A1(\ML_int[2][3] ), .A2(n8), .ZN(\ML_int[3][3] ) );
  AND2_X1 U48 ( .A1(\ML_int[2][2] ), .A2(n8), .ZN(\ML_int[3][2] ) );
  AND2_X1 U49 ( .A1(\ML_int[2][1] ), .A2(n8), .ZN(\ML_int[3][1] ) );
  AND2_X1 U50 ( .A1(\ML_int[2][0] ), .A2(n8), .ZN(\ML_int[3][0] ) );
  AND2_X1 U51 ( .A1(\ML_int[1][1] ), .A2(n6), .ZN(\ML_int[2][1] ) );
  AND2_X1 U52 ( .A1(\ML_int[1][0] ), .A2(n6), .ZN(\ML_int[2][0] ) );
  AND2_X1 U53 ( .A1(A[0]), .A2(n3), .ZN(\ML_int[1][0] ) );
endmodule


module SHIFTER_GENERIC_N32_DW_sla_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188;
  assign B[0] = \A[0] ;
  assign \A[0]  = A[0];

  NOR2_X2 U2 ( .A1(SH[2]), .A2(SH[3]), .ZN(n130) );
  INV_X1 U3 ( .A(n82), .ZN(n72) );
  INV_X1 U4 ( .A(n15), .ZN(n18) );
  INV_X1 U5 ( .A(n114), .ZN(n73) );
  BUF_X1 U6 ( .A(n94), .Z(n10) );
  BUF_X1 U7 ( .A(n94), .Z(n11) );
  AND2_X1 U8 ( .A1(n166), .A2(n14), .ZN(n88) );
  BUF_X1 U9 ( .A(n93), .Z(n7) );
  BUF_X1 U10 ( .A(n93), .Z(n8) );
  BUF_X1 U11 ( .A(n90), .Z(n1) );
  BUF_X1 U12 ( .A(n90), .Z(n2) );
  BUF_X1 U13 ( .A(n91), .Z(n4) );
  BUF_X1 U14 ( .A(n91), .Z(n5) );
  BUF_X1 U15 ( .A(SH[4]), .Z(n15) );
  BUF_X1 U16 ( .A(SH[4]), .Z(n16) );
  BUF_X1 U17 ( .A(n93), .Z(n9) );
  BUF_X1 U18 ( .A(n94), .Z(n12) );
  BUF_X1 U19 ( .A(n90), .Z(n3) );
  BUF_X1 U20 ( .A(n91), .Z(n6) );
  BUF_X1 U21 ( .A(SH[4]), .Z(n17) );
  INV_X1 U22 ( .A(n168), .ZN(n55) );
  INV_X1 U23 ( .A(n171), .ZN(n58) );
  INV_X1 U24 ( .A(n177), .ZN(n60) );
  INV_X1 U25 ( .A(n181), .ZN(n62) );
  INV_X1 U26 ( .A(n185), .ZN(n65) );
  INV_X1 U27 ( .A(n131), .ZN(n67) );
  INV_X1 U28 ( .A(n173), .ZN(n48) );
  INV_X1 U29 ( .A(n75), .ZN(n70) );
  INV_X1 U30 ( .A(n153), .ZN(n69) );
  INV_X1 U31 ( .A(n86), .ZN(n38) );
  INV_X1 U32 ( .A(n97), .ZN(n40) );
  INV_X1 U33 ( .A(n104), .ZN(n42) );
  INV_X1 U34 ( .A(n110), .ZN(n44) );
  INV_X1 U35 ( .A(n138), .ZN(n50) );
  INV_X1 U36 ( .A(n89), .ZN(n30) );
  INV_X1 U37 ( .A(n99), .ZN(n32) );
  INV_X1 U38 ( .A(n106), .ZN(n34) );
  INV_X1 U39 ( .A(n112), .ZN(n36) );
  NAND2_X1 U40 ( .A1(n17), .A2(\A[0] ), .ZN(n75) );
  INV_X1 U41 ( .A(A[29]), .ZN(n19) );
  INV_X1 U42 ( .A(n186), .ZN(n66) );
  INV_X1 U43 ( .A(A[12]), .ZN(n49) );
  INV_X1 U44 ( .A(A[23]), .ZN(n29) );
  INV_X1 U45 ( .A(A[14]), .ZN(n46) );
  INV_X1 U46 ( .A(A[17]), .ZN(n41) );
  INV_X1 U47 ( .A(A[21]), .ZN(n33) );
  INV_X1 U48 ( .A(A[13]), .ZN(n47) );
  INV_X1 U49 ( .A(A[22]), .ZN(n31) );
  INV_X1 U50 ( .A(A[16]), .ZN(n43) );
  INV_X1 U51 ( .A(A[15]), .ZN(n45) );
  INV_X1 U52 ( .A(A[9]), .ZN(n53) );
  INV_X1 U53 ( .A(A[7]), .ZN(n56) );
  INV_X1 U54 ( .A(A[10]), .ZN(n52) );
  INV_X1 U55 ( .A(A[11]), .ZN(n51) );
  INV_X1 U56 ( .A(A[8]), .ZN(n54) );
  INV_X1 U57 ( .A(A[2]), .ZN(n64) );
  INV_X1 U58 ( .A(A[28]), .ZN(n20) );
  INV_X1 U59 ( .A(A[27]), .ZN(n21) );
  INV_X1 U60 ( .A(A[26]), .ZN(n23) );
  INV_X1 U61 ( .A(A[25]), .ZN(n25) );
  INV_X1 U62 ( .A(A[24]), .ZN(n27) );
  INV_X1 U63 ( .A(A[3]), .ZN(n63) );
  INV_X1 U64 ( .A(A[18]), .ZN(n39) );
  INV_X1 U65 ( .A(\A[0] ), .ZN(n71) );
  INV_X1 U66 ( .A(A[4]), .ZN(n61) );
  INV_X1 U67 ( .A(A[6]), .ZN(n57) );
  INV_X1 U68 ( .A(A[19]), .ZN(n37) );
  INV_X1 U69 ( .A(A[20]), .ZN(n35) );
  INV_X1 U70 ( .A(A[1]), .ZN(n68) );
  INV_X1 U71 ( .A(A[5]), .ZN(n59) );
  INV_X1 U72 ( .A(n118), .ZN(n22) );
  INV_X1 U73 ( .A(n123), .ZN(n24) );
  INV_X1 U74 ( .A(n135), .ZN(n26) );
  INV_X1 U75 ( .A(n141), .ZN(n28) );
  INV_X1 U76 ( .A(SH[0]), .ZN(n13) );
  INV_X1 U77 ( .A(SH[2]), .ZN(n14) );
  OAI21_X1 U78 ( .B1(n15), .B2(n74), .A(n75), .ZN(B[9]) );
  OAI21_X1 U79 ( .B1(n15), .B2(n76), .A(n75), .ZN(B[8]) );
  OAI21_X1 U80 ( .B1(n15), .B2(n77), .A(n75), .ZN(B[7]) );
  OAI21_X1 U81 ( .B1(n15), .B2(n78), .A(n75), .ZN(B[6]) );
  OAI21_X1 U82 ( .B1(n15), .B2(n79), .A(n75), .ZN(B[5]) );
  OAI21_X1 U83 ( .B1(n16), .B2(n80), .A(n75), .ZN(B[4]) );
  OAI21_X1 U84 ( .B1(n16), .B2(n81), .A(n75), .ZN(B[3]) );
  OAI221_X1 U85 ( .B1(n22), .B2(n82), .C1(n83), .C2(n18), .A(n84), .ZN(B[31])
         );
  AOI222_X1 U86 ( .A1(n85), .A2(n86), .B1(n73), .B2(n87), .C1(n88), .C2(n89), 
        .ZN(n84) );
  OAI221_X1 U87 ( .B1(n2), .B2(n19), .C1(n5), .C2(n20), .A(n92), .ZN(n87) );
  AOI22_X1 U88 ( .A1(A[30]), .A2(n8), .B1(A[31]), .B2(n11), .ZN(n92) );
  OAI221_X1 U89 ( .B1(n24), .B2(n82), .C1(n95), .C2(n18), .A(n96), .ZN(B[30])
         );
  AOI222_X1 U90 ( .A1(n85), .A2(n97), .B1(n73), .B2(n98), .C1(n88), .C2(n99), 
        .ZN(n96) );
  OAI221_X1 U91 ( .B1(n1), .B2(n20), .C1(n4), .C2(n21), .A(n100), .ZN(n98) );
  AOI22_X1 U92 ( .A1(A[29]), .A2(n7), .B1(A[30]), .B2(n10), .ZN(n100) );
  OAI21_X1 U93 ( .B1(n16), .B2(n101), .A(n75), .ZN(B[2]) );
  OAI221_X1 U94 ( .B1(n26), .B2(n82), .C1(n102), .C2(n18), .A(n103), .ZN(B[29]) );
  AOI222_X1 U95 ( .A1(n85), .A2(n104), .B1(n73), .B2(n105), .C1(n88), .C2(n106), .ZN(n103) );
  OAI221_X1 U96 ( .B1(n1), .B2(n21), .C1(n4), .C2(n23), .A(n107), .ZN(n105) );
  AOI22_X1 U97 ( .A1(A[28]), .A2(n7), .B1(A[29]), .B2(n10), .ZN(n107) );
  OAI221_X1 U98 ( .B1(n28), .B2(n82), .C1(n108), .C2(n18), .A(n109), .ZN(B[28]) );
  AOI222_X1 U99 ( .A1(n85), .A2(n110), .B1(n73), .B2(n111), .C1(n88), .C2(n112), .ZN(n109) );
  OAI221_X1 U100 ( .B1(n1), .B2(n23), .C1(n4), .C2(n25), .A(n113), .ZN(n111)
         );
  AOI22_X1 U101 ( .A1(A[27]), .A2(n7), .B1(A[28]), .B2(n10), .ZN(n113) );
  OAI221_X1 U102 ( .B1(n22), .B2(n114), .C1(n115), .C2(n18), .A(n116), .ZN(
        B[27]) );
  AOI222_X1 U103 ( .A1(n72), .A2(n89), .B1(n88), .B2(n86), .C1(n85), .C2(n117), 
        .ZN(n116) );
  OAI221_X1 U104 ( .B1(n1), .B2(n25), .C1(n4), .C2(n27), .A(n119), .ZN(n118)
         );
  AOI22_X1 U105 ( .A1(A[26]), .A2(n7), .B1(A[27]), .B2(n10), .ZN(n119) );
  OAI221_X1 U106 ( .B1(n24), .B2(n114), .C1(n120), .C2(n18), .A(n121), .ZN(
        B[26]) );
  AOI222_X1 U107 ( .A1(n72), .A2(n99), .B1(n88), .B2(n97), .C1(n85), .C2(n122), 
        .ZN(n121) );
  OAI221_X1 U108 ( .B1(n1), .B2(n27), .C1(n4), .C2(n29), .A(n124), .ZN(n123)
         );
  AOI22_X1 U109 ( .A1(A[25]), .A2(n7), .B1(A[26]), .B2(n10), .ZN(n124) );
  OAI221_X1 U110 ( .B1(n26), .B2(n114), .C1(n74), .C2(n18), .A(n125), .ZN(
        B[25]) );
  AOI222_X1 U111 ( .A1(n72), .A2(n106), .B1(n88), .B2(n104), .C1(n85), .C2(
        n126), .ZN(n125) );
  AOI221_X1 U112 ( .B1(n127), .B2(n128), .C1(n129), .C2(n130), .A(n67), .ZN(
        n74) );
  AOI21_X1 U113 ( .B1(n132), .B2(n133), .A(n134), .ZN(n131) );
  OAI221_X1 U114 ( .B1(n1), .B2(n29), .C1(n4), .C2(n31), .A(n136), .ZN(n135)
         );
  AOI22_X1 U115 ( .A1(A[24]), .A2(n7), .B1(A[25]), .B2(n10), .ZN(n136) );
  OAI221_X1 U116 ( .B1(n28), .B2(n114), .C1(n76), .C2(n18), .A(n137), .ZN(
        B[24]) );
  AOI222_X1 U117 ( .A1(n72), .A2(n112), .B1(n88), .B2(n110), .C1(n85), .C2(
        n138), .ZN(n137) );
  AOI221_X1 U118 ( .B1(n139), .B2(n128), .C1(n140), .C2(n130), .A(n69), .ZN(
        n76) );
  OAI221_X1 U119 ( .B1(n1), .B2(n31), .C1(n4), .C2(n33), .A(n142), .ZN(n141)
         );
  AOI22_X1 U120 ( .A1(A[23]), .A2(n7), .B1(A[24]), .B2(n10), .ZN(n142) );
  OAI221_X1 U121 ( .B1(n30), .B2(n114), .C1(n77), .C2(n18), .A(n143), .ZN(
        B[23]) );
  AOI222_X1 U122 ( .A1(n72), .A2(n86), .B1(n88), .B2(n117), .C1(n85), .C2(n144), .ZN(n143) );
  AOI221_X1 U123 ( .B1(n145), .B2(n128), .C1(n146), .C2(n130), .A(n69), .ZN(
        n77) );
  OAI221_X1 U124 ( .B1(n1), .B2(n33), .C1(n4), .C2(n35), .A(n147), .ZN(n89) );
  AOI22_X1 U125 ( .A1(A[22]), .A2(n7), .B1(A[23]), .B2(n10), .ZN(n147) );
  OAI221_X1 U126 ( .B1(n32), .B2(n114), .C1(n78), .C2(n18), .A(n148), .ZN(
        B[22]) );
  AOI222_X1 U127 ( .A1(n72), .A2(n97), .B1(n88), .B2(n122), .C1(n85), .C2(n149), .ZN(n148) );
  AOI221_X1 U128 ( .B1(n66), .B2(n128), .C1(n150), .C2(n130), .A(n69), .ZN(n78) );
  OAI221_X1 U129 ( .B1(n1), .B2(n35), .C1(n5), .C2(n37), .A(n151), .ZN(n99) );
  AOI22_X1 U130 ( .A1(A[21]), .A2(n7), .B1(A[22]), .B2(n10), .ZN(n151) );
  OAI221_X1 U131 ( .B1(n34), .B2(n114), .C1(n79), .C2(n18), .A(n152), .ZN(
        B[21]) );
  AOI222_X1 U132 ( .A1(n72), .A2(n104), .B1(n88), .B2(n126), .C1(n85), .C2(
        n129), .ZN(n152) );
  AOI221_X1 U133 ( .B1(n133), .B2(n128), .C1(n127), .C2(n130), .A(n69), .ZN(
        n79) );
  OAI221_X1 U134 ( .B1(n1), .B2(n37), .C1(n5), .C2(n39), .A(n154), .ZN(n106)
         );
  AOI22_X1 U135 ( .A1(A[20]), .A2(n7), .B1(A[21]), .B2(n10), .ZN(n154) );
  OAI221_X1 U136 ( .B1(n36), .B2(n114), .C1(n80), .C2(n18), .A(n155), .ZN(
        B[20]) );
  AOI222_X1 U137 ( .A1(n72), .A2(n110), .B1(n88), .B2(n138), .C1(n85), .C2(
        n140), .ZN(n155) );
  AOI21_X1 U138 ( .B1(n139), .B2(n130), .A(n156), .ZN(n80) );
  OAI221_X1 U139 ( .B1(n1), .B2(n39), .C1(n5), .C2(n41), .A(n157), .ZN(n112)
         );
  AOI22_X1 U140 ( .A1(A[19]), .A2(n7), .B1(A[20]), .B2(n11), .ZN(n157) );
  OAI21_X1 U141 ( .B1(n16), .B2(n158), .A(n75), .ZN(B[1]) );
  OAI221_X1 U142 ( .B1(n38), .B2(n114), .C1(n81), .C2(n18), .A(n159), .ZN(
        B[19]) );
  AOI222_X1 U143 ( .A1(n72), .A2(n117), .B1(n88), .B2(n144), .C1(n85), .C2(
        n146), .ZN(n159) );
  AOI21_X1 U144 ( .B1(n145), .B2(n130), .A(n156), .ZN(n81) );
  OAI221_X1 U145 ( .B1(n2), .B2(n41), .C1(n5), .C2(n43), .A(n160), .ZN(n86) );
  AOI22_X1 U146 ( .A1(A[18]), .A2(n8), .B1(A[19]), .B2(n11), .ZN(n160) );
  OAI221_X1 U147 ( .B1(n40), .B2(n114), .C1(n101), .C2(n18), .A(n161), .ZN(
        B[18]) );
  AOI222_X1 U148 ( .A1(n72), .A2(n122), .B1(n88), .B2(n149), .C1(n85), .C2(
        n150), .ZN(n161) );
  AOI21_X1 U149 ( .B1(n66), .B2(n130), .A(n156), .ZN(n101) );
  OAI221_X1 U150 ( .B1(n2), .B2(n43), .C1(n5), .C2(n45), .A(n162), .ZN(n97) );
  AOI22_X1 U151 ( .A1(A[17]), .A2(n8), .B1(A[18]), .B2(n11), .ZN(n162) );
  OAI221_X1 U152 ( .B1(n42), .B2(n114), .C1(n158), .C2(n18), .A(n163), .ZN(
        B[17]) );
  AOI222_X1 U153 ( .A1(n72), .A2(n126), .B1(n88), .B2(n129), .C1(n85), .C2(
        n127), .ZN(n163) );
  AOI21_X1 U154 ( .B1(n133), .B2(n130), .A(n156), .ZN(n158) );
  OAI21_X1 U155 ( .B1(n71), .B2(n14), .A(n153), .ZN(n156) );
  OAI221_X1 U156 ( .B1(n2), .B2(n45), .C1(n5), .C2(n46), .A(n164), .ZN(n104)
         );
  AOI22_X1 U157 ( .A1(A[16]), .A2(n8), .B1(A[17]), .B2(n11), .ZN(n164) );
  OAI221_X1 U158 ( .B1(n50), .B2(n82), .C1(n44), .C2(n114), .A(n165), .ZN(
        B[16]) );
  AOI221_X1 U159 ( .B1(n85), .B2(n139), .C1(n88), .C2(n140), .A(n70), .ZN(n165) );
  AND2_X1 U160 ( .A1(n166), .A2(SH[2]), .ZN(n85) );
  AND2_X1 U161 ( .A1(SH[3]), .A2(n18), .ZN(n166) );
  NAND2_X1 U162 ( .A1(n130), .A2(n18), .ZN(n114) );
  OAI221_X1 U163 ( .B1(n2), .B2(n46), .C1(n5), .C2(n47), .A(n167), .ZN(n110)
         );
  AOI22_X1 U164 ( .A1(A[15]), .A2(n8), .B1(A[16]), .B2(n11), .ZN(n167) );
  NAND2_X1 U165 ( .A1(n128), .A2(n18), .ZN(n82) );
  OAI21_X1 U166 ( .B1(n16), .B2(n83), .A(n75), .ZN(B[15]) );
  AOI221_X1 U167 ( .B1(n144), .B2(n128), .C1(n117), .C2(n130), .A(n55), .ZN(
        n83) );
  AOI22_X1 U168 ( .A1(n169), .A2(n145), .B1(n132), .B2(n146), .ZN(n168) );
  OAI221_X1 U169 ( .B1(n2), .B2(n47), .C1(n5), .C2(n49), .A(n170), .ZN(n117)
         );
  AOI22_X1 U170 ( .A1(A[14]), .A2(n8), .B1(A[15]), .B2(n11), .ZN(n170) );
  OAI21_X1 U171 ( .B1(n16), .B2(n95), .A(n75), .ZN(B[14]) );
  AOI221_X1 U172 ( .B1(n149), .B2(n128), .C1(n122), .C2(n130), .A(n58), .ZN(
        n95) );
  AOI22_X1 U173 ( .A1(n169), .A2(n66), .B1(n132), .B2(n150), .ZN(n171) );
  OAI221_X1 U174 ( .B1(n2), .B2(n49), .C1(n5), .C2(n51), .A(n172), .ZN(n122)
         );
  AOI22_X1 U175 ( .A1(A[13]), .A2(n8), .B1(A[14]), .B2(n11), .ZN(n172) );
  OAI21_X1 U176 ( .B1(n16), .B2(n102), .A(n75), .ZN(B[13]) );
  AOI221_X1 U177 ( .B1(n133), .B2(n169), .C1(n127), .C2(n132), .A(n48), .ZN(
        n102) );
  AOI22_X1 U178 ( .A1(n128), .A2(n129), .B1(n130), .B2(n126), .ZN(n173) );
  OAI221_X1 U179 ( .B1(n2), .B2(n51), .C1(n5), .C2(n52), .A(n174), .ZN(n126)
         );
  AOI22_X1 U180 ( .A1(A[12]), .A2(n8), .B1(A[13]), .B2(n11), .ZN(n174) );
  OAI221_X1 U181 ( .B1(n2), .B2(n56), .C1(n5), .C2(n57), .A(n175), .ZN(n129)
         );
  AOI22_X1 U182 ( .A1(A[8]), .A2(n8), .B1(A[9]), .B2(n11), .ZN(n175) );
  OAI221_X1 U183 ( .B1(n2), .B2(n63), .C1(n6), .C2(n64), .A(n176), .ZN(n127)
         );
  AOI22_X1 U184 ( .A1(A[4]), .A2(n8), .B1(A[5]), .B2(n11), .ZN(n176) );
  AND2_X1 U185 ( .A1(SH[2]), .A2(SH[3]), .ZN(n169) );
  MUX2_X1 U186 ( .A(\A[0] ), .B(A[1]), .S(n10), .Z(n133) );
  OAI21_X1 U187 ( .B1(n17), .B2(n108), .A(n75), .ZN(B[12]) );
  AOI221_X1 U188 ( .B1(n140), .B2(n128), .C1(n138), .C2(n130), .A(n60), .ZN(
        n108) );
  AOI21_X1 U189 ( .B1(n132), .B2(n139), .A(n134), .ZN(n177) );
  OAI221_X1 U190 ( .B1(n2), .B2(n64), .C1(n68), .C2(n4), .A(n178), .ZN(n139)
         );
  AOI22_X1 U191 ( .A1(n9), .A2(A[3]), .B1(A[4]), .B2(n11), .ZN(n178) );
  OAI221_X1 U192 ( .B1(n2), .B2(n52), .C1(n6), .C2(n53), .A(n179), .ZN(n138)
         );
  AOI22_X1 U193 ( .A1(A[11]), .A2(n8), .B1(A[12]), .B2(n11), .ZN(n179) );
  OAI221_X1 U194 ( .B1(n3), .B2(n57), .C1(n6), .C2(n59), .A(n180), .ZN(n140)
         );
  AOI22_X1 U195 ( .A1(A[7]), .A2(n8), .B1(A[8]), .B2(n12), .ZN(n180) );
  OAI21_X1 U196 ( .B1(n17), .B2(n115), .A(n75), .ZN(B[11]) );
  AOI221_X1 U197 ( .B1(n146), .B2(n128), .C1(n144), .C2(n130), .A(n62), .ZN(
        n115) );
  AOI21_X1 U198 ( .B1(n132), .B2(n145), .A(n134), .ZN(n181) );
  OAI221_X1 U199 ( .B1(n68), .B2(n3), .C1(n71), .C2(n4), .A(n182), .ZN(n145)
         );
  AOI22_X1 U200 ( .A1(n9), .A2(A[2]), .B1(A[3]), .B2(n12), .ZN(n182) );
  OAI221_X1 U201 ( .B1(n3), .B2(n53), .C1(n6), .C2(n54), .A(n183), .ZN(n144)
         );
  AOI22_X1 U202 ( .A1(A[10]), .A2(n9), .B1(A[11]), .B2(n12), .ZN(n183) );
  OAI221_X1 U203 ( .B1(n3), .B2(n59), .C1(n6), .C2(n61), .A(n184), .ZN(n146)
         );
  AOI22_X1 U204 ( .A1(A[6]), .A2(n9), .B1(A[7]), .B2(n12), .ZN(n184) );
  OAI21_X1 U205 ( .B1(n17), .B2(n120), .A(n75), .ZN(B[10]) );
  AOI221_X1 U206 ( .B1(n150), .B2(n128), .C1(n149), .C2(n130), .A(n65), .ZN(
        n120) );
  AOI21_X1 U207 ( .B1(n132), .B2(n66), .A(n134), .ZN(n185) );
  NOR2_X1 U208 ( .A1(n14), .A2(n153), .ZN(n134) );
  NAND2_X1 U209 ( .A1(SH[3]), .A2(\A[0] ), .ZN(n153) );
  AOI222_X1 U210 ( .A1(n10), .A2(A[2]), .B1(A[1]), .B2(n9), .C1(\A[0] ), .C2(
        SH[1]), .ZN(n186) );
  AND2_X1 U211 ( .A1(SH[3]), .A2(n14), .ZN(n132) );
  OAI221_X1 U212 ( .B1(n3), .B2(n54), .C1(n4), .C2(n56), .A(n187), .ZN(n149)
         );
  AOI22_X1 U213 ( .A1(A[9]), .A2(n9), .B1(A[10]), .B2(n12), .ZN(n187) );
  NOR2_X1 U214 ( .A1(n14), .A2(SH[3]), .ZN(n128) );
  OAI221_X1 U215 ( .B1(n1), .B2(n61), .C1(n63), .C2(n4), .A(n188), .ZN(n150)
         );
  AOI22_X1 U216 ( .A1(A[5]), .A2(n7), .B1(A[6]), .B2(n10), .ZN(n188) );
  NOR2_X1 U217 ( .A1(SH[0]), .A2(SH[1]), .ZN(n94) );
  NOR2_X1 U218 ( .A1(n13), .A2(SH[1]), .ZN(n93) );
  NAND2_X1 U219 ( .A1(SH[0]), .A2(SH[1]), .ZN(n91) );
  NAND2_X1 U220 ( .A1(SH[1]), .A2(n13), .ZN(n90) );
endmodule


module SHIFTER_GENERIC_N32_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168;

  INV_X1 U3 ( .A(n62), .ZN(n55) );
  INV_X1 U4 ( .A(n143), .ZN(n56) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  INV_X1 U6 ( .A(n92), .ZN(n54) );
  INV_X1 U7 ( .A(n97), .ZN(n60) );
  INV_X1 U8 ( .A(n101), .ZN(n57) );
  INV_X1 U9 ( .A(n100), .ZN(n58) );
  INV_X1 U10 ( .A(n98), .ZN(n59) );
  AND2_X1 U11 ( .A1(n160), .A2(n4), .ZN(n66) );
  BUF_X1 U12 ( .A(SH[4]), .Z(n8) );
  BUF_X1 U13 ( .A(SH[4]), .Z(n6) );
  BUF_X1 U14 ( .A(SH[4]), .Z(n7) );
  BUF_X1 U15 ( .A(n98), .Z(n1) );
  BUF_X1 U16 ( .A(n98), .Z(n2) );
  INV_X1 U17 ( .A(n128), .ZN(n14) );
  NOR2_X2 U18 ( .A1(n3), .A2(SH[1]), .ZN(n100) );
  INV_X1 U19 ( .A(n129), .ZN(n13) );
  INV_X1 U20 ( .A(n131), .ZN(n15) );
  INV_X1 U21 ( .A(n163), .ZN(n10) );
  INV_X1 U22 ( .A(n142), .ZN(n12) );
  INV_X1 U23 ( .A(n141), .ZN(B[12]) );
  INV_X1 U24 ( .A(n61), .ZN(n41) );
  INV_X1 U25 ( .A(n79), .ZN(n31) );
  INV_X1 U26 ( .A(n108), .ZN(n40) );
  INV_X1 U27 ( .A(n70), .ZN(n44) );
  INV_X1 U28 ( .A(n96), .ZN(n38) );
  INV_X1 U29 ( .A(n84), .ZN(n33) );
  INV_X1 U30 ( .A(n65), .ZN(n35) );
  INV_X1 U31 ( .A(n85), .ZN(n26) );
  INV_X1 U32 ( .A(n67), .ZN(n28) );
  INV_X1 U33 ( .A(n80), .ZN(n25) );
  INV_X1 U34 ( .A(A[14]), .ZN(n39) );
  INV_X1 U35 ( .A(A[23]), .ZN(n24) );
  INV_X1 U36 ( .A(A[12]), .ZN(n42) );
  INV_X1 U37 ( .A(A[2]), .ZN(n53) );
  INV_X1 U38 ( .A(A[31]), .ZN(n16) );
  INV_X1 U39 ( .A(A[20]), .ZN(n29) );
  INV_X1 U40 ( .A(A[5]), .ZN(n50) );
  INV_X1 U41 ( .A(A[30]), .ZN(n17) );
  INV_X1 U42 ( .A(A[6]), .ZN(n49) );
  INV_X1 U43 ( .A(A[4]), .ZN(n51) );
  INV_X1 U44 ( .A(A[29]), .ZN(n18) );
  INV_X1 U45 ( .A(A[19]), .ZN(n30) );
  INV_X1 U46 ( .A(A[17]), .ZN(n34) );
  INV_X1 U47 ( .A(A[21]), .ZN(n27) );
  INV_X1 U48 ( .A(A[9]), .ZN(n46) );
  INV_X1 U49 ( .A(A[11]), .ZN(n43) );
  INV_X1 U50 ( .A(A[10]), .ZN(n45) );
  INV_X1 U51 ( .A(A[8]), .ZN(n47) );
  INV_X1 U52 ( .A(A[7]), .ZN(n48) );
  INV_X1 U53 ( .A(A[16]), .ZN(n36) );
  INV_X1 U54 ( .A(A[15]), .ZN(n37) );
  INV_X1 U55 ( .A(A[3]), .ZN(n52) );
  INV_X1 U56 ( .A(A[26]), .ZN(n21) );
  INV_X1 U57 ( .A(A[27]), .ZN(n20) );
  INV_X1 U58 ( .A(A[28]), .ZN(n19) );
  INV_X1 U59 ( .A(A[25]), .ZN(n22) );
  INV_X1 U60 ( .A(A[24]), .ZN(n23) );
  INV_X1 U61 ( .A(A[18]), .ZN(n32) );
  NOR2_X2 U62 ( .A1(SH[0]), .A2(SH[1]), .ZN(n101) );
  INV_X1 U63 ( .A(SH[0]), .ZN(n3) );
  INV_X1 U64 ( .A(SH[2]), .ZN(n4) );
  INV_X1 U65 ( .A(SH[3]), .ZN(n5) );
  OAI221_X1 U66 ( .B1(n61), .B2(n62), .C1(n63), .C2(n9), .A(n64), .ZN(B[9]) );
  AOI222_X1 U67 ( .A1(n54), .A2(n65), .B1(n66), .B2(n67), .C1(n68), .C2(n69), 
        .ZN(n64) );
  OAI221_X1 U68 ( .B1(n70), .B2(n62), .C1(n71), .C2(n9), .A(n72), .ZN(B[8]) );
  AOI222_X1 U69 ( .A1(n54), .A2(n73), .B1(n66), .B2(n74), .C1(n68), .C2(n75), 
        .ZN(n72) );
  OAI221_X1 U70 ( .B1(n76), .B2(n62), .C1(n77), .C2(n9), .A(n78), .ZN(B[7]) );
  AOI222_X1 U71 ( .A1(n54), .A2(n38), .B1(n66), .B2(n79), .C1(n68), .C2(n80), 
        .ZN(n78) );
  OAI221_X1 U72 ( .B1(n81), .B2(n62), .C1(n82), .C2(n9), .A(n83), .ZN(B[6]) );
  AOI222_X1 U73 ( .A1(n54), .A2(n40), .B1(n66), .B2(n84), .C1(n68), .C2(n85), 
        .ZN(n83) );
  OAI221_X1 U74 ( .B1(n86), .B2(n62), .C1(n87), .C2(n9), .A(n88), .ZN(B[5]) );
  AOI222_X1 U75 ( .A1(n54), .A2(n41), .B1(n66), .B2(n65), .C1(n68), .C2(n67), 
        .ZN(n88) );
  OAI221_X1 U76 ( .B1(n89), .B2(n62), .C1(n90), .C2(n9), .A(n91), .ZN(B[4]) );
  AOI222_X1 U77 ( .A1(n54), .A2(n44), .B1(n66), .B2(n73), .C1(n68), .C2(n74), 
        .ZN(n91) );
  OAI221_X1 U78 ( .B1(n76), .B2(n92), .C1(n93), .C2(n9), .A(n94), .ZN(B[3]) );
  AOI222_X1 U79 ( .A1(n68), .A2(n79), .B1(n55), .B2(n95), .C1(n66), .C2(n38), 
        .ZN(n94) );
  OAI221_X1 U80 ( .B1(n97), .B2(n49), .C1(n1), .C2(n50), .A(n99), .ZN(n95) );
  AOI22_X1 U81 ( .A1(A[4]), .A2(n100), .B1(A[3]), .B2(n101), .ZN(n99) );
  AOI221_X1 U82 ( .B1(n60), .B2(A[10]), .C1(n59), .C2(A[9]), .A(n102), .ZN(n76) );
  OAI22_X1 U83 ( .A1(n47), .A2(n58), .B1(n48), .B2(n57), .ZN(n102) );
  AND2_X1 U84 ( .A1(n55), .A2(n103), .ZN(B[31]) );
  AND2_X1 U85 ( .A1(n104), .A2(n55), .ZN(B[30]) );
  OAI221_X1 U86 ( .B1(n81), .B2(n92), .C1(n105), .C2(n9), .A(n106), .ZN(B[2])
         );
  AOI222_X1 U87 ( .A1(n68), .A2(n84), .B1(n55), .B2(n107), .C1(n66), .C2(n40), 
        .ZN(n106) );
  OAI221_X1 U88 ( .B1(n97), .B2(n50), .C1(n2), .C2(n51), .A(n109), .ZN(n107)
         );
  AOI22_X1 U89 ( .A1(A[3]), .A2(n100), .B1(A[2]), .B2(n101), .ZN(n109) );
  AOI221_X1 U90 ( .B1(n60), .B2(A[9]), .C1(n59), .C2(A[8]), .A(n110), .ZN(n81)
         );
  OAI22_X1 U91 ( .A1(n48), .A2(n58), .B1(n49), .B2(n57), .ZN(n110) );
  AND2_X1 U92 ( .A1(n111), .A2(n55), .ZN(B[29]) );
  AND2_X1 U93 ( .A1(n112), .A2(n55), .ZN(B[28]) );
  NOR3_X1 U94 ( .A1(n14), .A2(n8), .A3(SH[3]), .ZN(B[27]) );
  NOR2_X1 U95 ( .A1(n6), .A2(n113), .ZN(B[26]) );
  NOR2_X1 U96 ( .A1(n6), .A2(n63), .ZN(B[25]) );
  AOI22_X1 U97 ( .A1(n114), .A2(n56), .B1(n111), .B2(n115), .ZN(n63) );
  NOR2_X1 U98 ( .A1(n6), .A2(n71), .ZN(B[24]) );
  AOI22_X1 U99 ( .A1(n116), .A2(n56), .B1(n112), .B2(n115), .ZN(n71) );
  NOR2_X1 U100 ( .A1(n6), .A2(n77), .ZN(B[23]) );
  AOI222_X1 U101 ( .A1(n117), .A2(n115), .B1(n103), .B2(n118), .C1(n119), .C2(
        n56), .ZN(n77) );
  NOR2_X1 U102 ( .A1(n6), .A2(n82), .ZN(B[22]) );
  AOI222_X1 U103 ( .A1(n120), .A2(n115), .B1(n104), .B2(n118), .C1(n121), .C2(
        n56), .ZN(n82) );
  NOR2_X1 U104 ( .A1(n7), .A2(n87), .ZN(B[21]) );
  AOI222_X1 U105 ( .A1(n114), .A2(n115), .B1(n111), .B2(n118), .C1(n69), .C2(
        n56), .ZN(n87) );
  NOR2_X1 U106 ( .A1(n7), .A2(n90), .ZN(B[20]) );
  AOI222_X1 U107 ( .A1(n116), .A2(n115), .B1(n112), .B2(n118), .C1(n75), .C2(
        n56), .ZN(n90) );
  OAI221_X1 U108 ( .B1(n86), .B2(n92), .C1(n122), .C2(n9), .A(n123), .ZN(B[1])
         );
  AOI222_X1 U109 ( .A1(n68), .A2(n65), .B1(n55), .B2(n124), .C1(n66), .C2(n41), 
        .ZN(n123) );
  AOI221_X1 U110 ( .B1(n60), .B2(A[12]), .C1(n59), .C2(A[11]), .A(n125), .ZN(
        n61) );
  OAI22_X1 U111 ( .A1(n45), .A2(n58), .B1(n46), .B2(n57), .ZN(n125) );
  OAI221_X1 U112 ( .B1(n97), .B2(n51), .C1(n2), .C2(n52), .A(n126), .ZN(n124)
         );
  AOI22_X1 U113 ( .A1(A[2]), .A2(n100), .B1(A[1]), .B2(n101), .ZN(n126) );
  AOI221_X1 U114 ( .B1(n60), .B2(A[8]), .C1(n59), .C2(A[7]), .A(n127), .ZN(n86) );
  OAI22_X1 U115 ( .A1(n49), .A2(n58), .B1(n50), .B2(n57), .ZN(n127) );
  NOR2_X1 U116 ( .A1(n7), .A2(n93), .ZN(B[19]) );
  AOI222_X1 U117 ( .A1(n80), .A2(n56), .B1(n119), .B2(n115), .C1(n128), .C2(
        SH[3]), .ZN(n93) );
  NOR2_X1 U118 ( .A1(n7), .A2(n105), .ZN(B[18]) );
  AOI221_X1 U119 ( .B1(n121), .B2(n115), .C1(n85), .C2(n56), .A(n13), .ZN(n105) );
  AOI22_X1 U120 ( .A1(n130), .A2(n104), .B1(n118), .B2(n120), .ZN(n129) );
  NOR2_X1 U121 ( .A1(n7), .A2(n122), .ZN(B[17]) );
  AOI221_X1 U122 ( .B1(n69), .B2(n115), .C1(n67), .C2(n56), .A(n15), .ZN(n122)
         );
  AOI22_X1 U123 ( .A1(n130), .A2(n111), .B1(n118), .B2(n114), .ZN(n131) );
  NOR2_X1 U124 ( .A1(n8), .A2(n132), .ZN(B[16]) );
  OAI221_X1 U125 ( .B1(n25), .B2(n92), .C1(n31), .C2(n62), .A(n133), .ZN(B[15]) );
  AOI222_X1 U126 ( .A1(n68), .A2(n117), .B1(n134), .B2(n103), .C1(n66), .C2(
        n119), .ZN(n133) );
  OAI221_X1 U127 ( .B1(n26), .B2(n92), .C1(n33), .C2(n62), .A(n135), .ZN(B[14]) );
  AOI222_X1 U128 ( .A1(n68), .A2(n120), .B1(n134), .B2(n104), .C1(n66), .C2(
        n121), .ZN(n135) );
  OAI221_X1 U129 ( .B1(n28), .B2(n92), .C1(n35), .C2(n62), .A(n136), .ZN(B[13]) );
  AOI222_X1 U130 ( .A1(n68), .A2(n114), .B1(n134), .B2(n111), .C1(n66), .C2(
        n69), .ZN(n136) );
  OAI221_X1 U131 ( .B1(n97), .B2(n23), .C1(n1), .C2(n24), .A(n137), .ZN(n69)
         );
  AOI22_X1 U132 ( .A1(A[22]), .A2(n100), .B1(A[21]), .B2(n101), .ZN(n137) );
  OAI222_X1 U133 ( .A1(n58), .A2(n17), .B1(n1), .B2(n16), .C1(n57), .C2(n18), 
        .ZN(n111) );
  OAI221_X1 U134 ( .B1(n97), .B2(n19), .C1(n1), .C2(n20), .A(n138), .ZN(n114)
         );
  AOI22_X1 U135 ( .A1(A[26]), .A2(n100), .B1(A[25]), .B2(n101), .ZN(n138) );
  OAI221_X1 U136 ( .B1(n97), .B2(n36), .C1(n2), .C2(n37), .A(n139), .ZN(n65)
         );
  AOI22_X1 U137 ( .A1(A[14]), .A2(n100), .B1(A[13]), .B2(n101), .ZN(n139) );
  OAI221_X1 U138 ( .B1(n97), .B2(n29), .C1(n2), .C2(n30), .A(n140), .ZN(n67)
         );
  AOI22_X1 U139 ( .A1(A[18]), .A2(n100), .B1(A[17]), .B2(n101), .ZN(n140) );
  AOI221_X1 U140 ( .B1(n74), .B2(n54), .C1(n73), .C2(n55), .A(n12), .ZN(n141)
         );
  AOI222_X1 U141 ( .A1(n68), .A2(n116), .B1(n134), .B2(n112), .C1(n66), .C2(
        n75), .ZN(n142) );
  NOR2_X1 U142 ( .A1(n9), .A2(n143), .ZN(n134) );
  OAI221_X1 U143 ( .B1(n31), .B2(n92), .C1(n96), .C2(n62), .A(n144), .ZN(B[11]) );
  AOI221_X1 U144 ( .B1(n68), .B2(n119), .C1(n66), .C2(n80), .A(n145), .ZN(n144) );
  NOR3_X1 U145 ( .A1(n9), .A2(SH[3]), .A3(n14), .ZN(n145) );
  MUX2_X1 U146 ( .A(n117), .B(n103), .S(SH[2]), .Z(n128) );
  NOR2_X1 U147 ( .A1(n16), .A2(n57), .ZN(n103) );
  OAI221_X1 U148 ( .B1(n97), .B2(n17), .C1(n1), .C2(n18), .A(n146), .ZN(n117)
         );
  AOI22_X1 U149 ( .A1(A[28]), .A2(n100), .B1(A[27]), .B2(n101), .ZN(n146) );
  OAI221_X1 U150 ( .B1(n29), .B2(n58), .C1(n30), .C2(n57), .A(n147), .ZN(n80)
         );
  AOI22_X1 U151 ( .A1(A[22]), .A2(n60), .B1(A[21]), .B2(n59), .ZN(n147) );
  OAI221_X1 U152 ( .B1(n97), .B2(n21), .C1(n1), .C2(n22), .A(n148), .ZN(n119)
         );
  AOI22_X1 U153 ( .A1(A[24]), .A2(n100), .B1(A[23]), .B2(n101), .ZN(n148) );
  AOI221_X1 U154 ( .B1(n60), .B2(A[14]), .C1(n59), .C2(A[13]), .A(n149), .ZN(
        n96) );
  OAI22_X1 U155 ( .A1(n42), .A2(n58), .B1(n43), .B2(n57), .ZN(n149) );
  OAI221_X1 U156 ( .B1(n97), .B2(n32), .C1(n2), .C2(n34), .A(n150), .ZN(n79)
         );
  AOI22_X1 U157 ( .A1(A[16]), .A2(n100), .B1(A[15]), .B2(n101), .ZN(n150) );
  OAI221_X1 U158 ( .B1(n108), .B2(n62), .C1(n113), .C2(n9), .A(n151), .ZN(
        B[10]) );
  AOI222_X1 U159 ( .A1(n54), .A2(n84), .B1(n66), .B2(n85), .C1(n68), .C2(n121), 
        .ZN(n151) );
  OAI221_X1 U160 ( .B1(n97), .B2(n22), .C1(n2), .C2(n23), .A(n152), .ZN(n121)
         );
  AOI22_X1 U161 ( .A1(A[23]), .A2(n100), .B1(A[22]), .B2(n101), .ZN(n152) );
  OAI221_X1 U162 ( .B1(n97), .B2(n27), .C1(n29), .C2(n2), .A(n153), .ZN(n85)
         );
  AOI22_X1 U163 ( .A1(n100), .A2(A[19]), .B1(n101), .B2(A[18]), .ZN(n153) );
  OAI221_X1 U164 ( .B1(n97), .B2(n34), .C1(n1), .C2(n36), .A(n154), .ZN(n84)
         );
  AOI22_X1 U165 ( .A1(A[15]), .A2(n100), .B1(A[14]), .B2(n101), .ZN(n154) );
  AOI22_X1 U166 ( .A1(n120), .A2(n56), .B1(n104), .B2(n115), .ZN(n113) );
  OAI22_X1 U167 ( .A1(n57), .A2(n17), .B1(n58), .B2(n16), .ZN(n104) );
  OAI221_X1 U168 ( .B1(n97), .B2(n18), .C1(n1), .C2(n19), .A(n155), .ZN(n120)
         );
  AOI22_X1 U169 ( .A1(A[27]), .A2(n100), .B1(A[26]), .B2(n101), .ZN(n155) );
  AOI221_X1 U170 ( .B1(n60), .B2(A[13]), .C1(n59), .C2(A[12]), .A(n156), .ZN(
        n108) );
  OAI22_X1 U171 ( .A1(n43), .A2(n58), .B1(n45), .B2(n57), .ZN(n156) );
  OAI221_X1 U172 ( .B1(n89), .B2(n92), .C1(n132), .C2(n9), .A(n157), .ZN(B[0])
         );
  AOI222_X1 U173 ( .A1(n68), .A2(n73), .B1(n55), .B2(n158), .C1(n66), .C2(n44), 
        .ZN(n157) );
  AOI221_X1 U174 ( .B1(n60), .B2(A[11]), .C1(n59), .C2(A[10]), .A(n159), .ZN(
        n70) );
  OAI22_X1 U175 ( .A1(n46), .A2(n58), .B1(n47), .B2(n57), .ZN(n159) );
  OAI221_X1 U176 ( .B1(n97), .B2(n52), .C1(n2), .C2(n53), .A(n161), .ZN(n158)
         );
  AOI22_X1 U177 ( .A1(A[1]), .A2(n100), .B1(A[0]), .B2(n101), .ZN(n161) );
  NAND2_X1 U178 ( .A1(n56), .A2(n9), .ZN(n62) );
  OAI221_X1 U179 ( .B1(n97), .B2(n37), .C1(n2), .C2(n39), .A(n162), .ZN(n73)
         );
  AOI22_X1 U180 ( .A1(A[13]), .A2(n100), .B1(A[12]), .B2(n101), .ZN(n162) );
  AND2_X1 U181 ( .A1(SH[2]), .A2(n160), .ZN(n68) );
  NOR2_X1 U182 ( .A1(n5), .A2(n8), .ZN(n160) );
  AOI221_X1 U183 ( .B1(n75), .B2(n115), .C1(n74), .C2(n56), .A(n10), .ZN(n132)
         );
  AOI22_X1 U184 ( .A1(n130), .A2(n112), .B1(n118), .B2(n116), .ZN(n163) );
  OAI221_X1 U185 ( .B1(n97), .B2(n20), .C1(n1), .C2(n21), .A(n164), .ZN(n116)
         );
  AOI22_X1 U186 ( .A1(A[25]), .A2(n100), .B1(A[24]), .B2(n101), .ZN(n164) );
  NOR2_X1 U187 ( .A1(n5), .A2(SH[2]), .ZN(n118) );
  OAI221_X1 U188 ( .B1(n97), .B2(n16), .C1(n1), .C2(n17), .A(n165), .ZN(n112)
         );
  AOI22_X1 U189 ( .A1(A[29]), .A2(n100), .B1(A[28]), .B2(n101), .ZN(n165) );
  NOR2_X1 U190 ( .A1(n4), .A2(n5), .ZN(n130) );
  NAND2_X1 U191 ( .A1(n4), .A2(n5), .ZN(n143) );
  OAI221_X1 U192 ( .B1(n97), .B2(n30), .C1(n2), .C2(n32), .A(n166), .ZN(n74)
         );
  AOI22_X1 U193 ( .A1(A[17]), .A2(n100), .B1(A[16]), .B2(n101), .ZN(n166) );
  OAI221_X1 U194 ( .B1(n58), .B2(n27), .C1(n29), .C2(n57), .A(n167), .ZN(n75)
         );
  AOI22_X1 U195 ( .A1(A[23]), .A2(n60), .B1(A[22]), .B2(n59), .ZN(n167) );
  NAND2_X1 U196 ( .A1(n115), .A2(n9), .ZN(n92) );
  NOR2_X1 U197 ( .A1(n4), .A2(SH[3]), .ZN(n115) );
  AOI221_X1 U198 ( .B1(n60), .B2(A[7]), .C1(n59), .C2(A[6]), .A(n168), .ZN(n89) );
  OAI22_X1 U199 ( .A1(n50), .A2(n58), .B1(n51), .B2(n57), .ZN(n168) );
  NAND2_X1 U200 ( .A1(SH[1]), .A2(n3), .ZN(n98) );
  NAND2_X1 U201 ( .A1(SH[1]), .A2(SH[0]), .ZN(n97) );
endmodule


module SHIFTER_GENERIC_N32_DW_sra_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  NOR2_X2 U2 ( .A1(n2), .A2(SH[0]), .ZN(n94) );
  NOR2_X2 U3 ( .A1(SH[2]), .A2(SH[3]), .ZN(n114) );
  INV_X1 U4 ( .A(n98), .ZN(n59) );
  INV_X1 U5 ( .A(n95), .ZN(n57) );
  INV_X1 U6 ( .A(n88), .ZN(n54) );
  INV_X1 U7 ( .A(n4), .ZN(n7) );
  INV_X1 U8 ( .A(n61), .ZN(n55) );
  INV_X1 U9 ( .A(n97), .ZN(n58) );
  INV_X1 U10 ( .A(n94), .ZN(n56) );
  NOR2_X2 U11 ( .A1(n1), .A2(n2), .ZN(n95) );
  NAND2_X1 U12 ( .A1(n1), .A2(n2), .ZN(n98) );
  AND2_X1 U13 ( .A1(n166), .A2(n3), .ZN(n64) );
  BUF_X1 U14 ( .A(SH[4]), .Z(n4) );
  BUF_X1 U15 ( .A(SH[4]), .Z(n5) );
  BUF_X1 U16 ( .A(SH[4]), .Z(n6) );
  INV_X1 U17 ( .A(n121), .ZN(n13) );
  INV_X1 U18 ( .A(n125), .ZN(n11) );
  INV_X1 U19 ( .A(n126), .ZN(n9) );
  INV_X1 U20 ( .A(n134), .ZN(n15) );
  INV_X1 U21 ( .A(n138), .ZN(n10) );
  INV_X1 U22 ( .A(n169), .ZN(n8) );
  INV_X1 U23 ( .A(n137), .ZN(n22) );
  INV_X1 U24 ( .A(n100), .ZN(n16) );
  INV_X1 U25 ( .A(n141), .ZN(n33) );
  INV_X1 U26 ( .A(n132), .ZN(n34) );
  INV_X1 U27 ( .A(n149), .ZN(n36) );
  INV_X1 U28 ( .A(n92), .ZN(n38) );
  INV_X1 U29 ( .A(n104), .ZN(n39) );
  INV_X1 U30 ( .A(n60), .ZN(n41) );
  INV_X1 U31 ( .A(n68), .ZN(n44) );
  INV_X1 U32 ( .A(n135), .ZN(n14) );
  INV_X1 U33 ( .A(n77), .ZN(n26) );
  INV_X1 U34 ( .A(n76), .ZN(n30) );
  INV_X1 U35 ( .A(A[17]), .ZN(n32) );
  INV_X1 U36 ( .A(n168), .ZN(n40) );
  INV_X1 U37 ( .A(A[12]), .ZN(n42) );
  INV_X1 U38 ( .A(n160), .ZN(n35) );
  INV_X1 U39 ( .A(n148), .ZN(n37) );
  INV_X1 U40 ( .A(A[21]), .ZN(n27) );
  INV_X1 U41 ( .A(A[23]), .ZN(n25) );
  NAND2_X1 U42 ( .A1(n6), .A2(\A[31] ), .ZN(n100) );
  INV_X1 U43 ( .A(A[2]), .ZN(n53) );
  INV_X1 U44 ( .A(A[19]), .ZN(n29) );
  INV_X1 U45 ( .A(A[5]), .ZN(n50) );
  INV_X1 U46 ( .A(A[18]), .ZN(n31) );
  INV_X1 U47 ( .A(A[6]), .ZN(n49) );
  INV_X1 U48 ( .A(A[4]), .ZN(n51) );
  INV_X1 U49 ( .A(A[29]), .ZN(n18) );
  INV_X1 U50 ( .A(\A[31] ), .ZN(n12) );
  INV_X1 U51 ( .A(A[20]), .ZN(n28) );
  INV_X1 U52 ( .A(A[9]), .ZN(n46) );
  INV_X1 U53 ( .A(A[11]), .ZN(n43) );
  INV_X1 U54 ( .A(A[10]), .ZN(n45) );
  INV_X1 U55 ( .A(A[8]), .ZN(n47) );
  INV_X1 U56 ( .A(A[7]), .ZN(n48) );
  INV_X1 U57 ( .A(A[3]), .ZN(n52) );
  INV_X1 U58 ( .A(A[27]), .ZN(n20) );
  INV_X1 U59 ( .A(A[26]), .ZN(n21) );
  INV_X1 U60 ( .A(A[25]), .ZN(n23) );
  INV_X1 U61 ( .A(A[28]), .ZN(n19) );
  INV_X1 U62 ( .A(A[24]), .ZN(n24) );
  INV_X1 U63 ( .A(A[30]), .ZN(n17) );
  INV_X1 U64 ( .A(SH[0]), .ZN(n1) );
  INV_X1 U65 ( .A(SH[1]), .ZN(n2) );
  INV_X1 U66 ( .A(SH[2]), .ZN(n3) );
  OAI221_X1 U67 ( .B1(n60), .B2(n61), .C1(n62), .C2(n7), .A(n63), .ZN(B[9]) );
  AOI222_X1 U68 ( .A1(n54), .A2(n34), .B1(n64), .B2(n65), .C1(n66), .C2(n67), 
        .ZN(n63) );
  OAI221_X1 U69 ( .B1(n68), .B2(n61), .C1(n69), .C2(n7), .A(n70), .ZN(B[8]) );
  AOI222_X1 U70 ( .A1(n54), .A2(n36), .B1(n64), .B2(n71), .C1(n66), .C2(n72), 
        .ZN(n70) );
  OAI221_X1 U71 ( .B1(n73), .B2(n61), .C1(n74), .C2(n7), .A(n75), .ZN(B[7]) );
  AOI222_X1 U72 ( .A1(n54), .A2(n38), .B1(n64), .B2(n76), .C1(n66), .C2(n77), 
        .ZN(n75) );
  OAI221_X1 U73 ( .B1(n78), .B2(n61), .C1(n79), .C2(n7), .A(n80), .ZN(B[6]) );
  AOI222_X1 U74 ( .A1(n54), .A2(n39), .B1(n64), .B2(n33), .C1(n66), .C2(n81), 
        .ZN(n80) );
  OAI221_X1 U75 ( .B1(n82), .B2(n61), .C1(n83), .C2(n7), .A(n84), .ZN(B[5]) );
  AOI222_X1 U76 ( .A1(n54), .A2(n41), .B1(n64), .B2(n34), .C1(n66), .C2(n65), 
        .ZN(n84) );
  OAI221_X1 U77 ( .B1(n85), .B2(n61), .C1(n86), .C2(n7), .A(n87), .ZN(B[4]) );
  AOI222_X1 U78 ( .A1(n54), .A2(n44), .B1(n64), .B2(n36), .C1(n66), .C2(n71), 
        .ZN(n87) );
  OAI221_X1 U79 ( .B1(n73), .B2(n88), .C1(n89), .C2(n7), .A(n90), .ZN(B[3]) );
  AOI222_X1 U80 ( .A1(n66), .A2(n76), .B1(n55), .B2(n91), .C1(n64), .C2(n38), 
        .ZN(n90) );
  OAI221_X1 U81 ( .B1(n56), .B2(n50), .C1(n57), .C2(n49), .A(n93), .ZN(n91) );
  AOI22_X1 U82 ( .A1(A[4]), .A2(n58), .B1(A[3]), .B2(n59), .ZN(n93) );
  AOI221_X1 U83 ( .B1(n94), .B2(A[9]), .C1(n95), .C2(A[10]), .A(n96), .ZN(n73)
         );
  OAI22_X1 U84 ( .A1(n47), .A2(n97), .B1(n48), .B2(n98), .ZN(n96) );
  OAI21_X1 U85 ( .B1(n4), .B2(n99), .A(n100), .ZN(B[30]) );
  OAI221_X1 U86 ( .B1(n78), .B2(n88), .C1(n101), .C2(n7), .A(n102), .ZN(B[2])
         );
  AOI222_X1 U87 ( .A1(n66), .A2(n33), .B1(n55), .B2(n103), .C1(n64), .C2(n39), 
        .ZN(n102) );
  OAI221_X1 U88 ( .B1(n56), .B2(n51), .C1(n57), .C2(n50), .A(n105), .ZN(n103)
         );
  AOI22_X1 U89 ( .A1(A[3]), .A2(n58), .B1(A[2]), .B2(n59), .ZN(n105) );
  AOI221_X1 U90 ( .B1(n94), .B2(A[8]), .C1(n95), .C2(A[9]), .A(n106), .ZN(n78)
         );
  OAI22_X1 U91 ( .A1(n48), .A2(n97), .B1(n49), .B2(n98), .ZN(n106) );
  OAI21_X1 U92 ( .B1(n4), .B2(n107), .A(n100), .ZN(B[29]) );
  OAI21_X1 U93 ( .B1(n4), .B2(n108), .A(n100), .ZN(B[28]) );
  OAI21_X1 U94 ( .B1(n4), .B2(n109), .A(n100), .ZN(B[27]) );
  OAI21_X1 U95 ( .B1(n4), .B2(n110), .A(n100), .ZN(B[26]) );
  OAI21_X1 U96 ( .B1(n5), .B2(n62), .A(n100), .ZN(B[25]) );
  AOI221_X1 U97 ( .B1(n111), .B2(n112), .C1(n113), .C2(n114), .A(n14), .ZN(n62) );
  OAI21_X1 U98 ( .B1(n5), .B2(n69), .A(n100), .ZN(B[24]) );
  AOI221_X1 U99 ( .B1(n115), .B2(n112), .C1(n116), .C2(n114), .A(n14), .ZN(n69) );
  OAI21_X1 U100 ( .B1(n5), .B2(n74), .A(n100), .ZN(B[23]) );
  AOI221_X1 U101 ( .B1(n117), .B2(n112), .C1(n118), .C2(n114), .A(n14), .ZN(
        n74) );
  OAI21_X1 U102 ( .B1(n5), .B2(n79), .A(n100), .ZN(B[22]) );
  AOI221_X1 U103 ( .B1(n119), .B2(n112), .C1(n120), .C2(n114), .A(n13), .ZN(
        n79) );
  AOI21_X1 U104 ( .B1(n122), .B2(n123), .A(n124), .ZN(n121) );
  OAI21_X1 U105 ( .B1(n5), .B2(n83), .A(n100), .ZN(B[21]) );
  AOI221_X1 U106 ( .B1(n113), .B2(n112), .C1(n67), .C2(n114), .A(n11), .ZN(n83) );
  AOI21_X1 U107 ( .B1(n122), .B2(n111), .A(n124), .ZN(n125) );
  OAI21_X1 U108 ( .B1(n5), .B2(n86), .A(n100), .ZN(B[20]) );
  AOI221_X1 U109 ( .B1(n116), .B2(n112), .C1(n72), .C2(n114), .A(n9), .ZN(n86)
         );
  AOI21_X1 U110 ( .B1(n122), .B2(n115), .A(n124), .ZN(n126) );
  OAI221_X1 U111 ( .B1(n82), .B2(n88), .C1(n127), .C2(n7), .A(n128), .ZN(B[1])
         );
  AOI222_X1 U112 ( .A1(n66), .A2(n34), .B1(n55), .B2(n129), .C1(n64), .C2(n41), 
        .ZN(n128) );
  AOI221_X1 U113 ( .B1(n94), .B2(A[11]), .C1(n95), .C2(A[12]), .A(n130), .ZN(
        n60) );
  OAI22_X1 U114 ( .A1(n45), .A2(n97), .B1(n46), .B2(n98), .ZN(n130) );
  OAI221_X1 U115 ( .B1(n56), .B2(n52), .C1(n57), .C2(n51), .A(n131), .ZN(n129)
         );
  AOI22_X1 U116 ( .A1(A[2]), .A2(n58), .B1(A[1]), .B2(n59), .ZN(n131) );
  AOI221_X1 U117 ( .B1(n94), .B2(A[7]), .C1(n95), .C2(A[8]), .A(n133), .ZN(n82) );
  OAI22_X1 U118 ( .A1(n49), .A2(n97), .B1(n50), .B2(n98), .ZN(n133) );
  OAI21_X1 U119 ( .B1(n5), .B2(n89), .A(n100), .ZN(B[19]) );
  AOI221_X1 U120 ( .B1(n118), .B2(n112), .C1(n77), .C2(n114), .A(n15), .ZN(n89) );
  AOI21_X1 U121 ( .B1(n122), .B2(n117), .A(n124), .ZN(n134) );
  NOR2_X1 U122 ( .A1(n135), .A2(n3), .ZN(n124) );
  OAI21_X1 U123 ( .B1(n6), .B2(n101), .A(n100), .ZN(B[18]) );
  AOI221_X1 U124 ( .B1(n123), .B2(n136), .C1(n119), .C2(n122), .A(n22), .ZN(
        n101) );
  AOI22_X1 U125 ( .A1(n112), .A2(n120), .B1(n114), .B2(n81), .ZN(n137) );
  OAI21_X1 U126 ( .B1(n6), .B2(n127), .A(n100), .ZN(B[17]) );
  AOI221_X1 U127 ( .B1(n67), .B2(n112), .C1(n65), .C2(n114), .A(n10), .ZN(n127) );
  AOI22_X1 U128 ( .A1(n136), .A2(n111), .B1(n122), .B2(n113), .ZN(n138) );
  OAI21_X1 U129 ( .B1(n6), .B2(n139), .A(n100), .ZN(B[16]) );
  OAI221_X1 U130 ( .B1(n26), .B2(n88), .C1(n30), .C2(n61), .A(n140), .ZN(B[15]) );
  AOI221_X1 U131 ( .B1(n66), .B2(n117), .C1(n64), .C2(n118), .A(n16), .ZN(n140) );
  OAI221_X1 U132 ( .B1(n141), .B2(n61), .C1(n99), .C2(n7), .A(n142), .ZN(B[14]) );
  AOI222_X1 U133 ( .A1(n54), .A2(n81), .B1(n64), .B2(n120), .C1(n66), .C2(n119), .ZN(n142) );
  AOI21_X1 U134 ( .B1(n123), .B2(n114), .A(n143), .ZN(n99) );
  OAI221_X1 U135 ( .B1(n132), .B2(n61), .C1(n107), .C2(n7), .A(n144), .ZN(
        B[13]) );
  AOI222_X1 U136 ( .A1(n54), .A2(n65), .B1(n64), .B2(n67), .C1(n66), .C2(n113), 
        .ZN(n144) );
  OAI221_X1 U137 ( .B1(n56), .B2(n20), .C1(n57), .C2(n19), .A(n145), .ZN(n113)
         );
  AOI22_X1 U138 ( .A1(A[26]), .A2(n58), .B1(A[25]), .B2(n59), .ZN(n145) );
  OAI221_X1 U139 ( .B1(n56), .B2(n25), .C1(n57), .C2(n24), .A(n146), .ZN(n67)
         );
  AOI22_X1 U140 ( .A1(A[22]), .A2(n58), .B1(A[21]), .B2(n59), .ZN(n146) );
  OAI221_X1 U141 ( .B1(n56), .B2(n29), .C1(n57), .C2(n28), .A(n147), .ZN(n65)
         );
  AOI22_X1 U142 ( .A1(A[18]), .A2(n58), .B1(A[17]), .B2(n59), .ZN(n147) );
  AOI21_X1 U143 ( .B1(n111), .B2(n114), .A(n143), .ZN(n107) );
  OAI222_X1 U144 ( .A1(n98), .A2(n18), .B1(n97), .B2(n17), .C1(n2), .C2(n12), 
        .ZN(n111) );
  AOI221_X1 U145 ( .B1(n94), .B2(A[15]), .C1(n95), .C2(A[16]), .A(n37), .ZN(
        n132) );
  AOI22_X1 U146 ( .A1(A[14]), .A2(n58), .B1(A[13]), .B2(n59), .ZN(n148) );
  OAI221_X1 U147 ( .B1(n149), .B2(n61), .C1(n108), .C2(n7), .A(n150), .ZN(
        B[12]) );
  AOI222_X1 U148 ( .A1(n54), .A2(n71), .B1(n64), .B2(n72), .C1(n66), .C2(n116), 
        .ZN(n150) );
  AOI21_X1 U149 ( .B1(n115), .B2(n114), .A(n143), .ZN(n108) );
  OAI221_X1 U150 ( .B1(n92), .B2(n61), .C1(n109), .C2(n7), .A(n151), .ZN(B[11]) );
  AOI222_X1 U151 ( .A1(n54), .A2(n76), .B1(n64), .B2(n77), .C1(n66), .C2(n118), 
        .ZN(n151) );
  OAI221_X1 U152 ( .B1(n56), .B2(n23), .C1(n57), .C2(n21), .A(n152), .ZN(n118)
         );
  AOI22_X1 U153 ( .A1(A[24]), .A2(n58), .B1(A[23]), .B2(n59), .ZN(n152) );
  OAI221_X1 U154 ( .B1(n28), .B2(n97), .C1(n29), .C2(n98), .A(n153), .ZN(n77)
         );
  AOI22_X1 U155 ( .A1(A[21]), .A2(n94), .B1(A[22]), .B2(n95), .ZN(n153) );
  OAI221_X1 U156 ( .B1(n56), .B2(n32), .C1(n57), .C2(n31), .A(n154), .ZN(n76)
         );
  AOI22_X1 U157 ( .A1(A[16]), .A2(n58), .B1(A[15]), .B2(n59), .ZN(n154) );
  AOI21_X1 U158 ( .B1(n117), .B2(n114), .A(n143), .ZN(n109) );
  OAI21_X1 U159 ( .B1(n3), .B2(n12), .A(n135), .ZN(n143) );
  OAI221_X1 U160 ( .B1(n56), .B2(n18), .C1(n57), .C2(n17), .A(n155), .ZN(n117)
         );
  AOI22_X1 U161 ( .A1(A[28]), .A2(n58), .B1(A[27]), .B2(n59), .ZN(n155) );
  AOI221_X1 U162 ( .B1(n94), .B2(A[13]), .C1(n95), .C2(A[14]), .A(n156), .ZN(
        n92) );
  OAI22_X1 U163 ( .A1(n42), .A2(n97), .B1(n43), .B2(n98), .ZN(n156) );
  OAI221_X1 U164 ( .B1(n104), .B2(n61), .C1(n110), .C2(n7), .A(n157), .ZN(
        B[10]) );
  AOI222_X1 U165 ( .A1(n54), .A2(n33), .B1(n64), .B2(n81), .C1(n66), .C2(n120), 
        .ZN(n157) );
  OAI221_X1 U166 ( .B1(n56), .B2(n24), .C1(n57), .C2(n23), .A(n158), .ZN(n120)
         );
  AOI22_X1 U167 ( .A1(A[23]), .A2(n58), .B1(A[22]), .B2(n59), .ZN(n158) );
  OAI221_X1 U168 ( .B1(n29), .B2(n97), .C1(n31), .C2(n98), .A(n159), .ZN(n81)
         );
  AOI22_X1 U169 ( .A1(A[20]), .A2(n94), .B1(A[21]), .B2(n95), .ZN(n159) );
  AOI221_X1 U170 ( .B1(n94), .B2(A[16]), .C1(n95), .C2(A[17]), .A(n35), .ZN(
        n141) );
  AOI22_X1 U171 ( .A1(A[15]), .A2(n58), .B1(A[14]), .B2(n59), .ZN(n160) );
  AOI221_X1 U172 ( .B1(n123), .B2(n112), .C1(n119), .C2(n114), .A(n14), .ZN(
        n110) );
  NAND2_X1 U173 ( .A1(\A[31] ), .A2(SH[3]), .ZN(n135) );
  OAI221_X1 U174 ( .B1(n56), .B2(n19), .C1(n57), .C2(n18), .A(n161), .ZN(n119)
         );
  AOI22_X1 U175 ( .A1(A[27]), .A2(n58), .B1(A[26]), .B2(n59), .ZN(n161) );
  MUX2_X1 U176 ( .A(A[30]), .B(\A[31] ), .S(n98), .Z(n123) );
  AOI221_X1 U177 ( .B1(n94), .B2(A[12]), .C1(n95), .C2(A[13]), .A(n162), .ZN(
        n104) );
  OAI22_X1 U178 ( .A1(n43), .A2(n97), .B1(n45), .B2(n98), .ZN(n162) );
  OAI221_X1 U179 ( .B1(n85), .B2(n88), .C1(n139), .C2(n7), .A(n163), .ZN(B[0])
         );
  AOI222_X1 U180 ( .A1(n66), .A2(n36), .B1(n55), .B2(n164), .C1(n64), .C2(n44), 
        .ZN(n163) );
  AOI221_X1 U181 ( .B1(n94), .B2(A[10]), .C1(n95), .C2(A[11]), .A(n165), .ZN(
        n68) );
  OAI22_X1 U182 ( .A1(n46), .A2(n97), .B1(n47), .B2(n98), .ZN(n165) );
  OAI221_X1 U183 ( .B1(n56), .B2(n53), .C1(n57), .C2(n52), .A(n167), .ZN(n164)
         );
  AOI22_X1 U184 ( .A1(A[1]), .A2(n58), .B1(A[0]), .B2(n59), .ZN(n167) );
  NAND2_X1 U185 ( .A1(n114), .A2(n7), .ZN(n61) );
  AOI221_X1 U186 ( .B1(n94), .B2(A[14]), .C1(n95), .C2(A[15]), .A(n40), .ZN(
        n149) );
  AOI22_X1 U187 ( .A1(A[13]), .A2(n58), .B1(A[12]), .B2(n59), .ZN(n168) );
  AND2_X1 U188 ( .A1(SH[2]), .A2(n166), .ZN(n66) );
  AND2_X1 U189 ( .A1(SH[3]), .A2(n7), .ZN(n166) );
  AOI221_X1 U190 ( .B1(n72), .B2(n112), .C1(n71), .C2(n114), .A(n8), .ZN(n139)
         );
  AOI22_X1 U191 ( .A1(n136), .A2(n115), .B1(n122), .B2(n116), .ZN(n169) );
  OAI221_X1 U192 ( .B1(n56), .B2(n21), .C1(n57), .C2(n20), .A(n170), .ZN(n116)
         );
  AOI22_X1 U193 ( .A1(A[25]), .A2(n58), .B1(A[24]), .B2(n59), .ZN(n170) );
  AND2_X1 U194 ( .A1(SH[3]), .A2(n3), .ZN(n122) );
  OAI221_X1 U195 ( .B1(n56), .B2(n17), .C1(n57), .C2(n12), .A(n171), .ZN(n115)
         );
  AOI22_X1 U196 ( .A1(A[29]), .A2(n58), .B1(A[28]), .B2(n59), .ZN(n171) );
  AND2_X1 U197 ( .A1(SH[2]), .A2(SH[3]), .ZN(n136) );
  OAI221_X1 U198 ( .B1(n56), .B2(n31), .C1(n29), .C2(n57), .A(n172), .ZN(n71)
         );
  AOI22_X1 U199 ( .A1(A[17]), .A2(n58), .B1(A[16]), .B2(n59), .ZN(n172) );
  OAI221_X1 U200 ( .B1(n97), .B2(n27), .C1(n28), .C2(n98), .A(n173), .ZN(n72)
         );
  AOI22_X1 U201 ( .A1(A[22]), .A2(n94), .B1(A[23]), .B2(n95), .ZN(n173) );
  NAND2_X1 U202 ( .A1(n112), .A2(n7), .ZN(n88) );
  NOR2_X1 U203 ( .A1(n3), .A2(SH[3]), .ZN(n112) );
  AOI221_X1 U204 ( .B1(n94), .B2(A[6]), .C1(n95), .C2(A[7]), .A(n174), .ZN(n85) );
  OAI22_X1 U205 ( .A1(n50), .A2(n97), .B1(n51), .B2(n98), .ZN(n174) );
  NAND2_X1 U206 ( .A1(SH[0]), .A2(n2), .ZN(n97) );
endmodule


module SHIFTER_GENERIC_N32_DW_lbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] ,
         \ML_int[5][31] , \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] ,
         \ML_int[5][15] , \ML_int[5][14] , \ML_int[5][13] , \ML_int[5][12] ,
         \ML_int[5][11] , \ML_int[5][10] , \ML_int[5][9] , \ML_int[5][8] ,
         \ML_int[5][7] , \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] ,
         \ML_int[5][3] , \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;
  assign B[31] = \ML_int[5][31] ;
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[8] = \ML_int[5][8] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n15), .Z(
        \ML_int[5][31] ) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n15), .Z(
        \ML_int[5][30] ) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n15), .Z(
        \ML_int[5][29] ) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n15), .Z(
        \ML_int[5][28] ) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n15), .Z(
        \ML_int[5][27] ) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n15), .Z(
        \ML_int[5][26] ) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n15), .Z(
        \ML_int[5][25] ) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n15), .Z(
        \ML_int[5][24] ) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n14), .Z(
        \ML_int[5][23] ) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n14), .Z(
        \ML_int[5][22] ) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n14), .Z(
        \ML_int[5][21] ) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n14), .Z(
        \ML_int[5][20] ) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n14), .Z(
        \ML_int[5][19] ) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n14), .Z(
        \ML_int[5][18] ) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n14), .Z(
        \ML_int[5][17] ) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n14), .Z(
        \ML_int[5][16] ) );
  MUX2_X1 M0_4_15 ( .A(\ML_int[4][15] ), .B(\ML_int[4][31] ), .S(n14), .Z(
        \ML_int[5][15] ) );
  MUX2_X1 M0_4_14 ( .A(\ML_int[4][14] ), .B(\ML_int[4][30] ), .S(n14), .Z(
        \ML_int[5][14] ) );
  MUX2_X1 M0_4_13 ( .A(\ML_int[4][13] ), .B(\ML_int[4][29] ), .S(n14), .Z(
        \ML_int[5][13] ) );
  MUX2_X1 M0_4_12 ( .A(\ML_int[4][12] ), .B(\ML_int[4][28] ), .S(n14), .Z(
        \ML_int[5][12] ) );
  MUX2_X1 M0_4_11 ( .A(\ML_int[4][11] ), .B(\ML_int[4][27] ), .S(n13), .Z(
        \ML_int[5][11] ) );
  MUX2_X1 M0_4_10 ( .A(\ML_int[4][10] ), .B(\ML_int[4][26] ), .S(n13), .Z(
        \ML_int[5][10] ) );
  MUX2_X1 M0_4_9 ( .A(\ML_int[4][9] ), .B(\ML_int[4][25] ), .S(n13), .Z(
        \ML_int[5][9] ) );
  MUX2_X1 M0_4_8 ( .A(\ML_int[4][8] ), .B(\ML_int[4][24] ), .S(n13), .Z(
        \ML_int[5][8] ) );
  MUX2_X1 M0_4_7 ( .A(\ML_int[4][7] ), .B(\ML_int[4][23] ), .S(n13), .Z(
        \ML_int[5][7] ) );
  MUX2_X1 M0_4_6 ( .A(\ML_int[4][6] ), .B(\ML_int[4][22] ), .S(n13), .Z(
        \ML_int[5][6] ) );
  MUX2_X1 M0_4_5 ( .A(\ML_int[4][5] ), .B(\ML_int[4][21] ), .S(n13), .Z(
        \ML_int[5][5] ) );
  MUX2_X1 M0_4_4 ( .A(\ML_int[4][4] ), .B(\ML_int[4][20] ), .S(n13), .Z(
        \ML_int[5][4] ) );
  MUX2_X1 M0_4_3 ( .A(\ML_int[4][3] ), .B(\ML_int[4][19] ), .S(n13), .Z(
        \ML_int[5][3] ) );
  MUX2_X1 M0_4_2 ( .A(\ML_int[4][2] ), .B(\ML_int[4][18] ), .S(n13), .Z(
        \ML_int[5][2] ) );
  MUX2_X1 M0_4_1 ( .A(\ML_int[4][1] ), .B(\ML_int[4][17] ), .S(n13), .Z(
        \ML_int[5][1] ) );
  MUX2_X1 M0_4_0 ( .A(\ML_int[4][0] ), .B(\ML_int[4][16] ), .S(n13), .Z(
        \ML_int[5][0] ) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n12), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n12), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n12), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n12), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n12), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n12), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n12), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n12), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n11), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n11), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n11), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n11), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n11), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n11), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n11), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n11), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n11), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n11), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n11), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n11), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n10), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n10), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n10), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n10), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M0_3_7 ( .A(\ML_int[3][7] ), .B(\ML_int[3][31] ), .S(n10), .Z(
        \ML_int[4][7] ) );
  MUX2_X1 M0_3_6 ( .A(\ML_int[3][6] ), .B(\ML_int[3][30] ), .S(n10), .Z(
        \ML_int[4][6] ) );
  MUX2_X1 M0_3_5 ( .A(\ML_int[3][5] ), .B(\ML_int[3][29] ), .S(n10), .Z(
        \ML_int[4][5] ) );
  MUX2_X1 M0_3_4 ( .A(\ML_int[3][4] ), .B(\ML_int[3][28] ), .S(n10), .Z(
        \ML_int[4][4] ) );
  MUX2_X1 M0_3_3 ( .A(\ML_int[3][3] ), .B(\ML_int[3][27] ), .S(n10), .Z(
        \ML_int[4][3] ) );
  MUX2_X1 M0_3_2 ( .A(\ML_int[3][2] ), .B(\ML_int[3][26] ), .S(n10), .Z(
        \ML_int[4][2] ) );
  MUX2_X1 M0_3_1 ( .A(\ML_int[3][1] ), .B(\ML_int[3][25] ), .S(n10), .Z(
        \ML_int[4][1] ) );
  MUX2_X1 M0_3_0 ( .A(\ML_int[3][0] ), .B(\ML_int[3][24] ), .S(n10), .Z(
        \ML_int[4][0] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n9), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n9), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n9), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n9), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n9), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n9), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n9), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n9), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n8), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n8), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n8), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n8), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n8), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n8), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n8), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n8), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n8), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n8), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n8), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n8), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n7), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n7), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n7), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n7), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n7), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n7), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n7), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n7), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M0_2_3 ( .A(\ML_int[2][3] ), .B(\ML_int[2][31] ), .S(n7), .Z(
        \ML_int[3][3] ) );
  MUX2_X1 M0_2_2 ( .A(\ML_int[2][2] ), .B(\ML_int[2][30] ), .S(n7), .Z(
        \ML_int[3][2] ) );
  MUX2_X1 M0_2_1 ( .A(\ML_int[2][1] ), .B(\ML_int[2][29] ), .S(n7), .Z(
        \ML_int[3][1] ) );
  MUX2_X1 M0_2_0 ( .A(\ML_int[2][0] ), .B(\ML_int[2][28] ), .S(n7), .Z(
        \ML_int[3][0] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n6), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n6), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n6), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n6), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n6), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n6), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n6), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n6), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n5), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n5), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n5), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n5), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n5), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n5), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n5), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n5), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n5), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n5), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n5), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n5), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n4), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n4), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n4), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n4), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n4), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n4), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n4), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n4), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n4), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n4), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M0_1_1 ( .A(\ML_int[1][1] ), .B(\ML_int[1][31] ), .S(n4), .Z(
        \ML_int[2][1] ) );
  MUX2_X1 M0_1_0 ( .A(\ML_int[1][0] ), .B(\ML_int[1][30] ), .S(n4), .Z(
        \ML_int[2][0] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n3), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n3), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n3), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n3), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n3), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n3), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n3), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n3), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n2), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n2), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n2), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n2), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n2), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n2), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n2), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n2), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n2), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n2), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n2), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n2), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n1), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n1), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n1), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n1), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n1), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n1), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n1), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n1), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n1), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n1), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n1), .Z(\ML_int[1][1] ) );
  MUX2_X1 M0_0_0 ( .A(A[0]), .B(A[31]), .S(n1), .Z(\ML_int[1][0] ) );
  BUF_X1 U2 ( .A(SH[4]), .Z(n14) );
  BUF_X1 U3 ( .A(SH[4]), .Z(n13) );
  BUF_X1 U4 ( .A(SH[4]), .Z(n15) );
  BUF_X1 U5 ( .A(SH[1]), .Z(n5) );
  BUF_X1 U6 ( .A(SH[1]), .Z(n4) );
  BUF_X1 U7 ( .A(SH[2]), .Z(n8) );
  BUF_X1 U8 ( .A(SH[2]), .Z(n7) );
  BUF_X1 U9 ( .A(SH[0]), .Z(n2) );
  BUF_X1 U10 ( .A(SH[0]), .Z(n1) );
  BUF_X1 U11 ( .A(SH[3]), .Z(n11) );
  BUF_X1 U12 ( .A(SH[3]), .Z(n10) );
  BUF_X1 U13 ( .A(SH[1]), .Z(n6) );
  BUF_X1 U14 ( .A(SH[2]), .Z(n9) );
  BUF_X1 U15 ( .A(SH[0]), .Z(n3) );
  BUF_X1 U16 ( .A(SH[3]), .Z(n12) );
endmodule


module SHIFTER_GENERIC_N32_DW_rbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \MR_int[1][31] , \MR_int[1][30] , \MR_int[1][29] , \MR_int[1][28] ,
         \MR_int[1][27] , \MR_int[1][26] , \MR_int[1][25] , \MR_int[1][24] ,
         \MR_int[1][23] , \MR_int[1][22] , \MR_int[1][21] , \MR_int[1][20] ,
         \MR_int[1][19] , \MR_int[1][18] , \MR_int[1][17] , \MR_int[1][16] ,
         \MR_int[1][15] , \MR_int[1][14] , \MR_int[1][13] , \MR_int[1][12] ,
         \MR_int[1][11] , \MR_int[1][10] , \MR_int[1][9] , \MR_int[1][8] ,
         \MR_int[1][7] , \MR_int[1][6] , \MR_int[1][5] , \MR_int[1][4] ,
         \MR_int[1][3] , \MR_int[1][2] , \MR_int[1][1] , \MR_int[1][0] ,
         \MR_int[2][31] , \MR_int[2][30] , \MR_int[2][29] , \MR_int[2][28] ,
         \MR_int[2][27] , \MR_int[2][26] , \MR_int[2][25] , \MR_int[2][24] ,
         \MR_int[2][23] , \MR_int[2][22] , \MR_int[2][21] , \MR_int[2][20] ,
         \MR_int[2][19] , \MR_int[2][18] , \MR_int[2][17] , \MR_int[2][16] ,
         \MR_int[2][15] , \MR_int[2][14] , \MR_int[2][13] , \MR_int[2][12] ,
         \MR_int[2][11] , \MR_int[2][10] , \MR_int[2][9] , \MR_int[2][8] ,
         \MR_int[2][7] , \MR_int[2][6] , \MR_int[2][5] , \MR_int[2][4] ,
         \MR_int[2][3] , \MR_int[2][2] , \MR_int[2][1] , \MR_int[2][0] ,
         \MR_int[3][31] , \MR_int[3][30] , \MR_int[3][29] , \MR_int[3][28] ,
         \MR_int[3][27] , \MR_int[3][26] , \MR_int[3][25] , \MR_int[3][24] ,
         \MR_int[3][23] , \MR_int[3][22] , \MR_int[3][21] , \MR_int[3][20] ,
         \MR_int[3][19] , \MR_int[3][18] , \MR_int[3][17] , \MR_int[3][16] ,
         \MR_int[3][15] , \MR_int[3][14] , \MR_int[3][13] , \MR_int[3][12] ,
         \MR_int[3][11] , \MR_int[3][10] , \MR_int[3][9] , \MR_int[3][8] ,
         \MR_int[3][7] , \MR_int[3][6] , \MR_int[3][5] , \MR_int[3][4] ,
         \MR_int[3][3] , \MR_int[3][2] , \MR_int[3][1] , \MR_int[3][0] ,
         \MR_int[4][31] , \MR_int[4][30] , \MR_int[4][29] , \MR_int[4][28] ,
         \MR_int[4][27] , \MR_int[4][26] , \MR_int[4][25] , \MR_int[4][24] ,
         \MR_int[4][23] , \MR_int[4][22] , \MR_int[4][21] , \MR_int[4][20] ,
         \MR_int[4][19] , \MR_int[4][18] , \MR_int[4][17] , \MR_int[4][16] ,
         \MR_int[4][15] , \MR_int[4][14] , \MR_int[4][13] , \MR_int[4][12] ,
         \MR_int[4][11] , \MR_int[4][10] , \MR_int[4][9] , \MR_int[4][8] ,
         \MR_int[4][7] , \MR_int[4][6] , \MR_int[4][5] , \MR_int[4][4] ,
         \MR_int[4][3] , \MR_int[4][2] , \MR_int[4][1] , \MR_int[4][0] ,
         \MR_int[5][31] , \MR_int[5][30] , \MR_int[5][29] , \MR_int[5][28] ,
         \MR_int[5][27] , \MR_int[5][26] , \MR_int[5][25] , \MR_int[5][24] ,
         \MR_int[5][23] , \MR_int[5][22] , \MR_int[5][21] , \MR_int[5][20] ,
         \MR_int[5][19] , \MR_int[5][18] , \MR_int[5][17] , \MR_int[5][16] ,
         \MR_int[5][15] , \MR_int[5][14] , \MR_int[5][13] , \MR_int[5][12] ,
         \MR_int[5][11] , \MR_int[5][10] , \MR_int[5][9] , \MR_int[5][8] ,
         \MR_int[5][7] , \MR_int[5][6] , \MR_int[5][5] , \MR_int[5][4] ,
         \MR_int[5][3] , \MR_int[5][2] , \MR_int[5][1] , \MR_int[5][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;
  assign B[31] = \MR_int[5][31] ;
  assign B[30] = \MR_int[5][30] ;
  assign B[29] = \MR_int[5][29] ;
  assign B[28] = \MR_int[5][28] ;
  assign B[27] = \MR_int[5][27] ;
  assign B[26] = \MR_int[5][26] ;
  assign B[25] = \MR_int[5][25] ;
  assign B[24] = \MR_int[5][24] ;
  assign B[23] = \MR_int[5][23] ;
  assign B[22] = \MR_int[5][22] ;
  assign B[21] = \MR_int[5][21] ;
  assign B[20] = \MR_int[5][20] ;
  assign B[19] = \MR_int[5][19] ;
  assign B[18] = \MR_int[5][18] ;
  assign B[17] = \MR_int[5][17] ;
  assign B[16] = \MR_int[5][16] ;
  assign B[15] = \MR_int[5][15] ;
  assign B[14] = \MR_int[5][14] ;
  assign B[13] = \MR_int[5][13] ;
  assign B[12] = \MR_int[5][12] ;
  assign B[11] = \MR_int[5][11] ;
  assign B[10] = \MR_int[5][10] ;
  assign B[9] = \MR_int[5][9] ;
  assign B[8] = \MR_int[5][8] ;
  assign B[7] = \MR_int[5][7] ;
  assign B[6] = \MR_int[5][6] ;
  assign B[5] = \MR_int[5][5] ;
  assign B[4] = \MR_int[5][4] ;
  assign B[3] = \MR_int[5][3] ;
  assign B[2] = \MR_int[5][2] ;
  assign B[1] = \MR_int[5][1] ;
  assign B[0] = \MR_int[5][0] ;

  MUX2_X1 M1_4_31 ( .A(\MR_int[4][31] ), .B(\MR_int[4][15] ), .S(n15), .Z(
        \MR_int[5][31] ) );
  MUX2_X1 M1_4_30 ( .A(\MR_int[4][30] ), .B(\MR_int[4][14] ), .S(n15), .Z(
        \MR_int[5][30] ) );
  MUX2_X1 M1_4_29 ( .A(\MR_int[4][29] ), .B(\MR_int[4][13] ), .S(n15), .Z(
        \MR_int[5][29] ) );
  MUX2_X1 M1_4_28 ( .A(\MR_int[4][28] ), .B(\MR_int[4][12] ), .S(n15), .Z(
        \MR_int[5][28] ) );
  MUX2_X1 M1_4_27 ( .A(\MR_int[4][27] ), .B(\MR_int[4][11] ), .S(n15), .Z(
        \MR_int[5][27] ) );
  MUX2_X1 M1_4_26 ( .A(\MR_int[4][26] ), .B(\MR_int[4][10] ), .S(n15), .Z(
        \MR_int[5][26] ) );
  MUX2_X1 M1_4_25 ( .A(\MR_int[4][25] ), .B(\MR_int[4][9] ), .S(n15), .Z(
        \MR_int[5][25] ) );
  MUX2_X1 M1_4_24 ( .A(\MR_int[4][24] ), .B(\MR_int[4][8] ), .S(n15), .Z(
        \MR_int[5][24] ) );
  MUX2_X1 M1_4_23 ( .A(\MR_int[4][23] ), .B(\MR_int[4][7] ), .S(n14), .Z(
        \MR_int[5][23] ) );
  MUX2_X1 M1_4_22 ( .A(\MR_int[4][22] ), .B(\MR_int[4][6] ), .S(n14), .Z(
        \MR_int[5][22] ) );
  MUX2_X1 M1_4_21 ( .A(\MR_int[4][21] ), .B(\MR_int[4][5] ), .S(n14), .Z(
        \MR_int[5][21] ) );
  MUX2_X1 M1_4_20 ( .A(\MR_int[4][20] ), .B(\MR_int[4][4] ), .S(n14), .Z(
        \MR_int[5][20] ) );
  MUX2_X1 M1_4_19 ( .A(\MR_int[4][19] ), .B(\MR_int[4][3] ), .S(n14), .Z(
        \MR_int[5][19] ) );
  MUX2_X1 M1_4_18 ( .A(\MR_int[4][18] ), .B(\MR_int[4][2] ), .S(n14), .Z(
        \MR_int[5][18] ) );
  MUX2_X1 M1_4_17 ( .A(\MR_int[4][17] ), .B(\MR_int[4][1] ), .S(n14), .Z(
        \MR_int[5][17] ) );
  MUX2_X1 M1_4_16 ( .A(\MR_int[4][16] ), .B(\MR_int[4][0] ), .S(n14), .Z(
        \MR_int[5][16] ) );
  MUX2_X1 M1_4_15 ( .A(\MR_int[4][15] ), .B(\MR_int[4][31] ), .S(n14), .Z(
        \MR_int[5][15] ) );
  MUX2_X1 M1_4_14 ( .A(\MR_int[4][14] ), .B(\MR_int[4][30] ), .S(n14), .Z(
        \MR_int[5][14] ) );
  MUX2_X1 M1_4_13 ( .A(\MR_int[4][13] ), .B(\MR_int[4][29] ), .S(n14), .Z(
        \MR_int[5][13] ) );
  MUX2_X1 M1_4_12 ( .A(\MR_int[4][12] ), .B(\MR_int[4][28] ), .S(n14), .Z(
        \MR_int[5][12] ) );
  MUX2_X1 M1_4_11 ( .A(\MR_int[4][11] ), .B(\MR_int[4][27] ), .S(n13), .Z(
        \MR_int[5][11] ) );
  MUX2_X1 M1_4_10 ( .A(\MR_int[4][10] ), .B(\MR_int[4][26] ), .S(n13), .Z(
        \MR_int[5][10] ) );
  MUX2_X1 M1_4_9 ( .A(\MR_int[4][9] ), .B(\MR_int[4][25] ), .S(n13), .Z(
        \MR_int[5][9] ) );
  MUX2_X1 M1_4_8 ( .A(\MR_int[4][8] ), .B(\MR_int[4][24] ), .S(n13), .Z(
        \MR_int[5][8] ) );
  MUX2_X1 M1_4_7 ( .A(\MR_int[4][7] ), .B(\MR_int[4][23] ), .S(n13), .Z(
        \MR_int[5][7] ) );
  MUX2_X1 M1_4_6 ( .A(\MR_int[4][6] ), .B(\MR_int[4][22] ), .S(n13), .Z(
        \MR_int[5][6] ) );
  MUX2_X1 M1_4_5 ( .A(\MR_int[4][5] ), .B(\MR_int[4][21] ), .S(n13), .Z(
        \MR_int[5][5] ) );
  MUX2_X1 M1_4_4 ( .A(\MR_int[4][4] ), .B(\MR_int[4][20] ), .S(n13), .Z(
        \MR_int[5][4] ) );
  MUX2_X1 M1_4_3 ( .A(\MR_int[4][3] ), .B(\MR_int[4][19] ), .S(n13), .Z(
        \MR_int[5][3] ) );
  MUX2_X1 M1_4_2 ( .A(\MR_int[4][2] ), .B(\MR_int[4][18] ), .S(n13), .Z(
        \MR_int[5][2] ) );
  MUX2_X1 M1_4_1 ( .A(\MR_int[4][1] ), .B(\MR_int[4][17] ), .S(n13), .Z(
        \MR_int[5][1] ) );
  MUX2_X1 M1_4_0 ( .A(\MR_int[4][0] ), .B(\MR_int[4][16] ), .S(n13), .Z(
        \MR_int[5][0] ) );
  MUX2_X1 M1_3_31_0 ( .A(\MR_int[3][31] ), .B(\MR_int[3][7] ), .S(n12), .Z(
        \MR_int[4][31] ) );
  MUX2_X1 M1_3_30_0 ( .A(\MR_int[3][30] ), .B(\MR_int[3][6] ), .S(n12), .Z(
        \MR_int[4][30] ) );
  MUX2_X1 M1_3_29_0 ( .A(\MR_int[3][29] ), .B(\MR_int[3][5] ), .S(n12), .Z(
        \MR_int[4][29] ) );
  MUX2_X1 M1_3_28_0 ( .A(\MR_int[3][28] ), .B(\MR_int[3][4] ), .S(n12), .Z(
        \MR_int[4][28] ) );
  MUX2_X1 M1_3_27_0 ( .A(\MR_int[3][27] ), .B(\MR_int[3][3] ), .S(n12), .Z(
        \MR_int[4][27] ) );
  MUX2_X1 M1_3_26_0 ( .A(\MR_int[3][26] ), .B(\MR_int[3][2] ), .S(n12), .Z(
        \MR_int[4][26] ) );
  MUX2_X1 M1_3_25_0 ( .A(\MR_int[3][25] ), .B(\MR_int[3][1] ), .S(n12), .Z(
        \MR_int[4][25] ) );
  MUX2_X1 M1_3_24_0 ( .A(\MR_int[3][24] ), .B(\MR_int[3][0] ), .S(n12), .Z(
        \MR_int[4][24] ) );
  MUX2_X1 M1_3_23_0 ( .A(\MR_int[3][23] ), .B(\MR_int[3][31] ), .S(n11), .Z(
        \MR_int[4][23] ) );
  MUX2_X1 M1_3_22_0 ( .A(\MR_int[3][22] ), .B(\MR_int[3][30] ), .S(n11), .Z(
        \MR_int[4][22] ) );
  MUX2_X1 M1_3_21_0 ( .A(\MR_int[3][21] ), .B(\MR_int[3][29] ), .S(n11), .Z(
        \MR_int[4][21] ) );
  MUX2_X1 M1_3_20_0 ( .A(\MR_int[3][20] ), .B(\MR_int[3][28] ), .S(n11), .Z(
        \MR_int[4][20] ) );
  MUX2_X1 M1_3_19_0 ( .A(\MR_int[3][19] ), .B(\MR_int[3][27] ), .S(n11), .Z(
        \MR_int[4][19] ) );
  MUX2_X1 M1_3_18_0 ( .A(\MR_int[3][18] ), .B(\MR_int[3][26] ), .S(n11), .Z(
        \MR_int[4][18] ) );
  MUX2_X1 M1_3_17_0 ( .A(\MR_int[3][17] ), .B(\MR_int[3][25] ), .S(n11), .Z(
        \MR_int[4][17] ) );
  MUX2_X1 M1_3_16_0 ( .A(\MR_int[3][16] ), .B(\MR_int[3][24] ), .S(n11), .Z(
        \MR_int[4][16] ) );
  MUX2_X1 M1_3_15_0 ( .A(\MR_int[3][15] ), .B(\MR_int[3][23] ), .S(n11), .Z(
        \MR_int[4][15] ) );
  MUX2_X1 M1_3_14_0 ( .A(\MR_int[3][14] ), .B(\MR_int[3][22] ), .S(n11), .Z(
        \MR_int[4][14] ) );
  MUX2_X1 M1_3_13_0 ( .A(\MR_int[3][13] ), .B(\MR_int[3][21] ), .S(n11), .Z(
        \MR_int[4][13] ) );
  MUX2_X1 M1_3_12_0 ( .A(\MR_int[3][12] ), .B(\MR_int[3][20] ), .S(n11), .Z(
        \MR_int[4][12] ) );
  MUX2_X1 M1_3_11_0 ( .A(\MR_int[3][11] ), .B(\MR_int[3][19] ), .S(n10), .Z(
        \MR_int[4][11] ) );
  MUX2_X1 M1_3_10_0 ( .A(\MR_int[3][10] ), .B(\MR_int[3][18] ), .S(n10), .Z(
        \MR_int[4][10] ) );
  MUX2_X1 M1_3_9_0 ( .A(\MR_int[3][9] ), .B(\MR_int[3][17] ), .S(n10), .Z(
        \MR_int[4][9] ) );
  MUX2_X1 M1_3_8_0 ( .A(\MR_int[3][8] ), .B(\MR_int[3][16] ), .S(n10), .Z(
        \MR_int[4][8] ) );
  MUX2_X1 M1_3_7 ( .A(\MR_int[3][7] ), .B(\MR_int[3][15] ), .S(n10), .Z(
        \MR_int[4][7] ) );
  MUX2_X1 M1_3_6 ( .A(\MR_int[3][6] ), .B(\MR_int[3][14] ), .S(n10), .Z(
        \MR_int[4][6] ) );
  MUX2_X1 M1_3_5 ( .A(\MR_int[3][5] ), .B(\MR_int[3][13] ), .S(n10), .Z(
        \MR_int[4][5] ) );
  MUX2_X1 M1_3_4 ( .A(\MR_int[3][4] ), .B(\MR_int[3][12] ), .S(n10), .Z(
        \MR_int[4][4] ) );
  MUX2_X1 M1_3_3 ( .A(\MR_int[3][3] ), .B(\MR_int[3][11] ), .S(n10), .Z(
        \MR_int[4][3] ) );
  MUX2_X1 M1_3_2 ( .A(\MR_int[3][2] ), .B(\MR_int[3][10] ), .S(n10), .Z(
        \MR_int[4][2] ) );
  MUX2_X1 M1_3_1 ( .A(\MR_int[3][1] ), .B(\MR_int[3][9] ), .S(n10), .Z(
        \MR_int[4][1] ) );
  MUX2_X1 M1_3_0 ( .A(\MR_int[3][0] ), .B(\MR_int[3][8] ), .S(n10), .Z(
        \MR_int[4][0] ) );
  MUX2_X1 M1_2_31_0 ( .A(\MR_int[2][31] ), .B(\MR_int[2][3] ), .S(n9), .Z(
        \MR_int[3][31] ) );
  MUX2_X1 M1_2_30_0 ( .A(\MR_int[2][30] ), .B(\MR_int[2][2] ), .S(n9), .Z(
        \MR_int[3][30] ) );
  MUX2_X1 M1_2_29_0 ( .A(\MR_int[2][29] ), .B(\MR_int[2][1] ), .S(n9), .Z(
        \MR_int[3][29] ) );
  MUX2_X1 M1_2_28_0 ( .A(\MR_int[2][28] ), .B(\MR_int[2][0] ), .S(n9), .Z(
        \MR_int[3][28] ) );
  MUX2_X1 M1_2_27_0 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n9), .Z(
        \MR_int[3][27] ) );
  MUX2_X1 M1_2_26_0 ( .A(\MR_int[2][26] ), .B(\MR_int[2][30] ), .S(n9), .Z(
        \MR_int[3][26] ) );
  MUX2_X1 M1_2_25_0 ( .A(\MR_int[2][25] ), .B(\MR_int[2][29] ), .S(n9), .Z(
        \MR_int[3][25] ) );
  MUX2_X1 M1_2_24_0 ( .A(\MR_int[2][24] ), .B(\MR_int[2][28] ), .S(n9), .Z(
        \MR_int[3][24] ) );
  MUX2_X1 M1_2_23_0 ( .A(\MR_int[2][23] ), .B(\MR_int[2][27] ), .S(n8), .Z(
        \MR_int[3][23] ) );
  MUX2_X1 M1_2_22_0 ( .A(\MR_int[2][22] ), .B(\MR_int[2][26] ), .S(n8), .Z(
        \MR_int[3][22] ) );
  MUX2_X1 M1_2_21_0 ( .A(\MR_int[2][21] ), .B(\MR_int[2][25] ), .S(n8), .Z(
        \MR_int[3][21] ) );
  MUX2_X1 M1_2_20_0 ( .A(\MR_int[2][20] ), .B(\MR_int[2][24] ), .S(n8), .Z(
        \MR_int[3][20] ) );
  MUX2_X1 M1_2_19_0 ( .A(\MR_int[2][19] ), .B(\MR_int[2][23] ), .S(n8), .Z(
        \MR_int[3][19] ) );
  MUX2_X1 M1_2_18_0 ( .A(\MR_int[2][18] ), .B(\MR_int[2][22] ), .S(n8), .Z(
        \MR_int[3][18] ) );
  MUX2_X1 M1_2_17_0 ( .A(\MR_int[2][17] ), .B(\MR_int[2][21] ), .S(n8), .Z(
        \MR_int[3][17] ) );
  MUX2_X1 M1_2_16_0 ( .A(\MR_int[2][16] ), .B(\MR_int[2][20] ), .S(n8), .Z(
        \MR_int[3][16] ) );
  MUX2_X1 M1_2_15_0 ( .A(\MR_int[2][15] ), .B(\MR_int[2][19] ), .S(n8), .Z(
        \MR_int[3][15] ) );
  MUX2_X1 M1_2_14_0 ( .A(\MR_int[2][14] ), .B(\MR_int[2][18] ), .S(n8), .Z(
        \MR_int[3][14] ) );
  MUX2_X1 M1_2_13_0 ( .A(\MR_int[2][13] ), .B(\MR_int[2][17] ), .S(n8), .Z(
        \MR_int[3][13] ) );
  MUX2_X1 M1_2_12_0 ( .A(\MR_int[2][12] ), .B(\MR_int[2][16] ), .S(n8), .Z(
        \MR_int[3][12] ) );
  MUX2_X1 M1_2_11_0 ( .A(\MR_int[2][11] ), .B(\MR_int[2][15] ), .S(n7), .Z(
        \MR_int[3][11] ) );
  MUX2_X1 M1_2_10_0 ( .A(\MR_int[2][10] ), .B(\MR_int[2][14] ), .S(n7), .Z(
        \MR_int[3][10] ) );
  MUX2_X1 M1_2_9_0 ( .A(\MR_int[2][9] ), .B(\MR_int[2][13] ), .S(n7), .Z(
        \MR_int[3][9] ) );
  MUX2_X1 M1_2_8_0 ( .A(\MR_int[2][8] ), .B(\MR_int[2][12] ), .S(n7), .Z(
        \MR_int[3][8] ) );
  MUX2_X1 M1_2_7_0 ( .A(\MR_int[2][7] ), .B(\MR_int[2][11] ), .S(n7), .Z(
        \MR_int[3][7] ) );
  MUX2_X1 M1_2_6_0 ( .A(\MR_int[2][6] ), .B(\MR_int[2][10] ), .S(n7), .Z(
        \MR_int[3][6] ) );
  MUX2_X1 M1_2_5_0 ( .A(\MR_int[2][5] ), .B(\MR_int[2][9] ), .S(n7), .Z(
        \MR_int[3][5] ) );
  MUX2_X1 M1_2_4_0 ( .A(\MR_int[2][4] ), .B(\MR_int[2][8] ), .S(n7), .Z(
        \MR_int[3][4] ) );
  MUX2_X1 M1_2_3 ( .A(\MR_int[2][3] ), .B(\MR_int[2][7] ), .S(n7), .Z(
        \MR_int[3][3] ) );
  MUX2_X1 M1_2_2 ( .A(\MR_int[2][2] ), .B(\MR_int[2][6] ), .S(n7), .Z(
        \MR_int[3][2] ) );
  MUX2_X1 M1_2_1 ( .A(\MR_int[2][1] ), .B(\MR_int[2][5] ), .S(n7), .Z(
        \MR_int[3][1] ) );
  MUX2_X1 M1_2_0 ( .A(\MR_int[2][0] ), .B(\MR_int[2][4] ), .S(n7), .Z(
        \MR_int[3][0] ) );
  MUX2_X1 M1_1_31_0 ( .A(\MR_int[1][31] ), .B(\MR_int[1][1] ), .S(n6), .Z(
        \MR_int[2][31] ) );
  MUX2_X1 M1_1_30_0 ( .A(\MR_int[1][30] ), .B(\MR_int[1][0] ), .S(n6), .Z(
        \MR_int[2][30] ) );
  MUX2_X1 M1_1_29_0 ( .A(\MR_int[1][29] ), .B(\MR_int[1][31] ), .S(n6), .Z(
        \MR_int[2][29] ) );
  MUX2_X1 M1_1_28_0 ( .A(\MR_int[1][28] ), .B(\MR_int[1][30] ), .S(n6), .Z(
        \MR_int[2][28] ) );
  MUX2_X1 M1_1_27_0 ( .A(\MR_int[1][27] ), .B(\MR_int[1][29] ), .S(n6), .Z(
        \MR_int[2][27] ) );
  MUX2_X1 M1_1_26_0 ( .A(\MR_int[1][26] ), .B(\MR_int[1][28] ), .S(n6), .Z(
        \MR_int[2][26] ) );
  MUX2_X1 M1_1_25_0 ( .A(\MR_int[1][25] ), .B(\MR_int[1][27] ), .S(n6), .Z(
        \MR_int[2][25] ) );
  MUX2_X1 M1_1_24_0 ( .A(\MR_int[1][24] ), .B(\MR_int[1][26] ), .S(n6), .Z(
        \MR_int[2][24] ) );
  MUX2_X1 M1_1_23_0 ( .A(\MR_int[1][23] ), .B(\MR_int[1][25] ), .S(n5), .Z(
        \MR_int[2][23] ) );
  MUX2_X1 M1_1_22_0 ( .A(\MR_int[1][22] ), .B(\MR_int[1][24] ), .S(n5), .Z(
        \MR_int[2][22] ) );
  MUX2_X1 M1_1_21_0 ( .A(\MR_int[1][21] ), .B(\MR_int[1][23] ), .S(n5), .Z(
        \MR_int[2][21] ) );
  MUX2_X1 M1_1_20_0 ( .A(\MR_int[1][20] ), .B(\MR_int[1][22] ), .S(n5), .Z(
        \MR_int[2][20] ) );
  MUX2_X1 M1_1_19_0 ( .A(\MR_int[1][19] ), .B(\MR_int[1][21] ), .S(n5), .Z(
        \MR_int[2][19] ) );
  MUX2_X1 M1_1_18_0 ( .A(\MR_int[1][18] ), .B(\MR_int[1][20] ), .S(n5), .Z(
        \MR_int[2][18] ) );
  MUX2_X1 M1_1_17_0 ( .A(\MR_int[1][17] ), .B(\MR_int[1][19] ), .S(n5), .Z(
        \MR_int[2][17] ) );
  MUX2_X1 M1_1_16_0 ( .A(\MR_int[1][16] ), .B(\MR_int[1][18] ), .S(n5), .Z(
        \MR_int[2][16] ) );
  MUX2_X1 M1_1_15_0 ( .A(\MR_int[1][15] ), .B(\MR_int[1][17] ), .S(n5), .Z(
        \MR_int[2][15] ) );
  MUX2_X1 M1_1_14_0 ( .A(\MR_int[1][14] ), .B(\MR_int[1][16] ), .S(n5), .Z(
        \MR_int[2][14] ) );
  MUX2_X1 M1_1_13_0 ( .A(\MR_int[1][13] ), .B(\MR_int[1][15] ), .S(n5), .Z(
        \MR_int[2][13] ) );
  MUX2_X1 M1_1_12_0 ( .A(\MR_int[1][12] ), .B(\MR_int[1][14] ), .S(n5), .Z(
        \MR_int[2][12] ) );
  MUX2_X1 M1_1_11_0 ( .A(\MR_int[1][11] ), .B(\MR_int[1][13] ), .S(n4), .Z(
        \MR_int[2][11] ) );
  MUX2_X1 M1_1_10_0 ( .A(\MR_int[1][10] ), .B(\MR_int[1][12] ), .S(n4), .Z(
        \MR_int[2][10] ) );
  MUX2_X1 M1_1_9_0 ( .A(\MR_int[1][9] ), .B(\MR_int[1][11] ), .S(n4), .Z(
        \MR_int[2][9] ) );
  MUX2_X1 M1_1_8_0 ( .A(\MR_int[1][8] ), .B(\MR_int[1][10] ), .S(n4), .Z(
        \MR_int[2][8] ) );
  MUX2_X1 M1_1_7_0 ( .A(\MR_int[1][7] ), .B(\MR_int[1][9] ), .S(n4), .Z(
        \MR_int[2][7] ) );
  MUX2_X1 M1_1_6_0 ( .A(\MR_int[1][6] ), .B(\MR_int[1][8] ), .S(n4), .Z(
        \MR_int[2][6] ) );
  MUX2_X1 M1_1_5_0 ( .A(\MR_int[1][5] ), .B(\MR_int[1][7] ), .S(n4), .Z(
        \MR_int[2][5] ) );
  MUX2_X1 M1_1_4_0 ( .A(\MR_int[1][4] ), .B(\MR_int[1][6] ), .S(n4), .Z(
        \MR_int[2][4] ) );
  MUX2_X1 M1_1_3_0 ( .A(\MR_int[1][3] ), .B(\MR_int[1][5] ), .S(n4), .Z(
        \MR_int[2][3] ) );
  MUX2_X1 M1_1_2_0 ( .A(\MR_int[1][2] ), .B(\MR_int[1][4] ), .S(n4), .Z(
        \MR_int[2][2] ) );
  MUX2_X1 M1_1_1 ( .A(\MR_int[1][1] ), .B(\MR_int[1][3] ), .S(n4), .Z(
        \MR_int[2][1] ) );
  MUX2_X1 M1_1_0 ( .A(\MR_int[1][0] ), .B(\MR_int[1][2] ), .S(n4), .Z(
        \MR_int[2][0] ) );
  MUX2_X1 M1_0_31_0 ( .A(A[31]), .B(A[0]), .S(n3), .Z(\MR_int[1][31] ) );
  MUX2_X1 M1_0_30_0 ( .A(A[30]), .B(A[31]), .S(n3), .Z(\MR_int[1][30] ) );
  MUX2_X1 M1_0_29_0 ( .A(A[29]), .B(A[30]), .S(n3), .Z(\MR_int[1][29] ) );
  MUX2_X1 M1_0_28_0 ( .A(A[28]), .B(A[29]), .S(n3), .Z(\MR_int[1][28] ) );
  MUX2_X1 M1_0_27_0 ( .A(A[27]), .B(A[28]), .S(n3), .Z(\MR_int[1][27] ) );
  MUX2_X1 M1_0_26_0 ( .A(A[26]), .B(A[27]), .S(n3), .Z(\MR_int[1][26] ) );
  MUX2_X1 M1_0_25_0 ( .A(A[25]), .B(A[26]), .S(n3), .Z(\MR_int[1][25] ) );
  MUX2_X1 M1_0_24_0 ( .A(A[24]), .B(A[25]), .S(n3), .Z(\MR_int[1][24] ) );
  MUX2_X1 M1_0_23_0 ( .A(A[23]), .B(A[24]), .S(n2), .Z(\MR_int[1][23] ) );
  MUX2_X1 M1_0_22_0 ( .A(A[22]), .B(A[23]), .S(n2), .Z(\MR_int[1][22] ) );
  MUX2_X1 M1_0_21_0 ( .A(A[21]), .B(A[22]), .S(n2), .Z(\MR_int[1][21] ) );
  MUX2_X1 M1_0_20_0 ( .A(A[20]), .B(A[21]), .S(n2), .Z(\MR_int[1][20] ) );
  MUX2_X1 M1_0_19_0 ( .A(A[19]), .B(A[20]), .S(n2), .Z(\MR_int[1][19] ) );
  MUX2_X1 M1_0_18_0 ( .A(A[18]), .B(A[19]), .S(n2), .Z(\MR_int[1][18] ) );
  MUX2_X1 M1_0_17_0 ( .A(A[17]), .B(A[18]), .S(n2), .Z(\MR_int[1][17] ) );
  MUX2_X1 M1_0_16_0 ( .A(A[16]), .B(A[17]), .S(n2), .Z(\MR_int[1][16] ) );
  MUX2_X1 M1_0_15_0 ( .A(A[15]), .B(A[16]), .S(n2), .Z(\MR_int[1][15] ) );
  MUX2_X1 M1_0_14_0 ( .A(A[14]), .B(A[15]), .S(n2), .Z(\MR_int[1][14] ) );
  MUX2_X1 M1_0_13_0 ( .A(A[13]), .B(A[14]), .S(n2), .Z(\MR_int[1][13] ) );
  MUX2_X1 M1_0_12_0 ( .A(A[12]), .B(A[13]), .S(n2), .Z(\MR_int[1][12] ) );
  MUX2_X1 M1_0_11_0 ( .A(A[11]), .B(A[12]), .S(n1), .Z(\MR_int[1][11] ) );
  MUX2_X1 M1_0_10_0 ( .A(A[10]), .B(A[11]), .S(n1), .Z(\MR_int[1][10] ) );
  MUX2_X1 M1_0_9_0 ( .A(A[9]), .B(A[10]), .S(n1), .Z(\MR_int[1][9] ) );
  MUX2_X1 M1_0_8_0 ( .A(A[8]), .B(A[9]), .S(n1), .Z(\MR_int[1][8] ) );
  MUX2_X1 M1_0_7_0 ( .A(A[7]), .B(A[8]), .S(n1), .Z(\MR_int[1][7] ) );
  MUX2_X1 M1_0_6_0 ( .A(A[6]), .B(A[7]), .S(n1), .Z(\MR_int[1][6] ) );
  MUX2_X1 M1_0_5_0 ( .A(A[5]), .B(A[6]), .S(n1), .Z(\MR_int[1][5] ) );
  MUX2_X1 M1_0_4_0 ( .A(A[4]), .B(A[5]), .S(n1), .Z(\MR_int[1][4] ) );
  MUX2_X1 M1_0_3_0 ( .A(A[3]), .B(A[4]), .S(n1), .Z(\MR_int[1][3] ) );
  MUX2_X1 M1_0_2_0 ( .A(A[2]), .B(A[3]), .S(n1), .Z(\MR_int[1][2] ) );
  MUX2_X1 M1_0_1_0 ( .A(A[1]), .B(A[2]), .S(n1), .Z(\MR_int[1][1] ) );
  MUX2_X1 M1_0_0 ( .A(A[0]), .B(A[1]), .S(n1), .Z(\MR_int[1][0] ) );
  BUF_X1 U2 ( .A(SH[4]), .Z(n14) );
  BUF_X1 U3 ( .A(SH[4]), .Z(n13) );
  BUF_X1 U4 ( .A(SH[4]), .Z(n15) );
  BUF_X1 U5 ( .A(SH[1]), .Z(n5) );
  BUF_X1 U6 ( .A(SH[1]), .Z(n4) );
  BUF_X1 U7 ( .A(SH[2]), .Z(n8) );
  BUF_X1 U8 ( .A(SH[2]), .Z(n7) );
  BUF_X1 U9 ( .A(SH[0]), .Z(n2) );
  BUF_X1 U10 ( .A(SH[0]), .Z(n1) );
  BUF_X1 U11 ( .A(SH[3]), .Z(n11) );
  BUF_X1 U12 ( .A(SH[3]), .Z(n10) );
  BUF_X1 U13 ( .A(SH[1]), .Z(n6) );
  BUF_X1 U14 ( .A(SH[2]), .Z(n9) );
  BUF_X1 U15 ( .A(SH[0]), .Z(n3) );
  BUF_X1 U16 ( .A(SH[3]), .Z(n12) );
endmodule


module SHIFTER_GENERIC_N32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE, 
        OUTPUT );
  input [31:0] A;
  input [4:0] B;
  output [31:0] OUTPUT;
  input LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n19, n20, n93, n94, n95, n96, n97, n98, n99;

  SHIFTER_GENERIC_N32_DW01_ash_0 sll_49 ( .A(A), .DATA_TC(1'b0), .SH({n97, 
        B[3:0]}), .SH_TC(1'b0), .B({N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234}) );
  SHIFTER_GENERIC_N32_DW_sla_0 sla_47 ( .A(A), .SH({n97, B[3:0]}), .SH_TC(1'b0), .B({N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, 
        N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, 
        N209, N208, N207, N206, N205, N204, N203, N202}) );
  SHIFTER_GENERIC_N32_DW_rash_0 srl_42 ( .A(A), .DATA_TC(1'b0), .SH({n97, 
        B[3:0]}), .SH_TC(1'b0), .B({N168, N167, N166, N165, N164, N163, N162, 
        N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, 
        N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, 
        N137}) );
  SHIFTER_GENERIC_N32_DW_sra_0 sra_40 ( .A(A), .SH({n97, B[3:0]}), .SH_TC(1'b0), .B({N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, 
        N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, 
        N112, N111, N110, N109, N108, N107, N106, N105}) );
  SHIFTER_GENERIC_N32_DW_lbsh_0 rol_33 ( .A(A), .SH({n97, B[3:0]}), .SH_TC(
        1'b0), .B({N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, 
        N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, 
        N44, N43, N42, N41, N40, N39}) );
  SHIFTER_GENERIC_N32_DW_rbsh_0 ror_31 ( .A(A), .SH({n97, B[3:0]}), .SH_TC(
        1'b0), .B({N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7}) );
  AOI222_X1 U5 ( .A1(N211), .A2(n96), .B1(N114), .B2(n93), .C1(N146), .C2(n12), 
        .ZN(n22) );
  AOI222_X1 U6 ( .A1(N210), .A2(n96), .B1(N113), .B2(n93), .C1(N145), .C2(n12), 
        .ZN(n30) );
  AOI222_X1 U7 ( .A1(N209), .A2(n96), .B1(N112), .B2(n93), .C1(N144), .C2(n12), 
        .ZN(n32) );
  AOI222_X1 U8 ( .A1(N208), .A2(n96), .B1(N111), .B2(n93), .C1(N143), .C2(n12), 
        .ZN(n34) );
  AOI222_X1 U9 ( .A1(N207), .A2(n96), .B1(N110), .B2(n93), .C1(N142), .C2(n12), 
        .ZN(n36) );
  AOI222_X1 U10 ( .A1(N206), .A2(n96), .B1(N109), .B2(n93), .C1(N141), .C2(n12), .ZN(n38) );
  AOI222_X1 U13 ( .A1(N205), .A2(n96), .B1(N108), .B2(n93), .C1(N140), .C2(n12), .ZN(n40) );
  AOI222_X1 U14 ( .A1(N232), .A2(n95), .B1(N135), .B2(n20), .C1(N167), .C2(n11), .ZN(n44) );
  AOI222_X1 U15 ( .A1(N231), .A2(n95), .B1(N134), .B2(n20), .C1(N166), .C2(n11), .ZN(n48) );
  AOI222_X1 U16 ( .A1(N230), .A2(n95), .B1(N133), .B2(n20), .C1(N165), .C2(n11), .ZN(n50) );
  AOI222_X1 U17 ( .A1(N229), .A2(n95), .B1(N132), .B2(n20), .C1(N164), .C2(n11), .ZN(n52) );
  AOI222_X1 U18 ( .A1(N228), .A2(n95), .B1(N131), .B2(n20), .C1(N163), .C2(n11), .ZN(n54) );
  AOI222_X1 U19 ( .A1(N227), .A2(n95), .B1(N130), .B2(n20), .C1(N162), .C2(n11), .ZN(n56) );
  AOI222_X1 U20 ( .A1(N226), .A2(n95), .B1(N129), .B2(n20), .C1(N161), .C2(n11), .ZN(n58) );
  AOI222_X1 U21 ( .A1(N225), .A2(n95), .B1(N128), .B2(n20), .C1(N160), .C2(n11), .ZN(n60) );
  AOI222_X1 U22 ( .A1(N224), .A2(n95), .B1(N127), .B2(n20), .C1(N159), .C2(n11), .ZN(n62) );
  AOI222_X1 U23 ( .A1(N223), .A2(n95), .B1(N126), .B2(n20), .C1(N158), .C2(n11), .ZN(n64) );
  AOI222_X1 U24 ( .A1(N222), .A2(n95), .B1(N125), .B2(n20), .C1(N157), .C2(n11), .ZN(n66) );
  AOI222_X1 U25 ( .A1(N221), .A2(n94), .B1(N124), .B2(n19), .C1(N156), .C2(n10), .ZN(n70) );
  AOI222_X1 U26 ( .A1(N220), .A2(n94), .B1(N123), .B2(n19), .C1(N155), .C2(n10), .ZN(n72) );
  AOI222_X1 U27 ( .A1(N219), .A2(n94), .B1(N122), .B2(n19), .C1(N154), .C2(n10), .ZN(n74) );
  AOI222_X1 U28 ( .A1(N218), .A2(n94), .B1(N121), .B2(n19), .C1(N153), .C2(n10), .ZN(n76) );
  AOI222_X1 U29 ( .A1(N217), .A2(n94), .B1(N120), .B2(n19), .C1(N152), .C2(n10), .ZN(n78) );
  AOI222_X1 U30 ( .A1(N216), .A2(n94), .B1(N119), .B2(n19), .C1(N151), .C2(n10), .ZN(n80) );
  AOI222_X1 U31 ( .A1(N215), .A2(n94), .B1(N118), .B2(n19), .C1(N150), .C2(n10), .ZN(n82) );
  AOI222_X1 U32 ( .A1(N214), .A2(n94), .B1(N117), .B2(n19), .C1(N149), .C2(n10), .ZN(n84) );
  AOI222_X1 U33 ( .A1(N213), .A2(n94), .B1(N116), .B2(n19), .C1(N148), .C2(n10), .ZN(n86) );
  AOI222_X1 U34 ( .A1(N212), .A2(n94), .B1(N115), .B2(n19), .C1(N147), .C2(n10), .ZN(n88) );
  AOI222_X1 U35 ( .A1(N204), .A2(n95), .B1(N107), .B2(n20), .C1(N139), .C2(n11), .ZN(n46) );
  AOI222_X1 U36 ( .A1(N203), .A2(n94), .B1(N106), .B2(n19), .C1(N138), .C2(n10), .ZN(n68) );
  AOI222_X1 U37 ( .A1(N70), .A2(n9), .B1(N265), .B2(n6), .C1(N38), .C2(n3), 
        .ZN(n41) );
  AOI222_X1 U38 ( .A1(N48), .A2(n9), .B1(N243), .B2(n6), .C1(N16), .C2(n3), 
        .ZN(n21) );
  AOI222_X1 U39 ( .A1(N47), .A2(n9), .B1(N242), .B2(n6), .C1(N15), .C2(n3), 
        .ZN(n29) );
  AOI222_X1 U40 ( .A1(N46), .A2(n9), .B1(N241), .B2(n6), .C1(N14), .C2(n3), 
        .ZN(n31) );
  AOI222_X1 U41 ( .A1(N45), .A2(n9), .B1(N240), .B2(n6), .C1(N13), .C2(n3), 
        .ZN(n33) );
  AOI222_X1 U42 ( .A1(N44), .A2(n9), .B1(N239), .B2(n6), .C1(N12), .C2(n3), 
        .ZN(n35) );
  AOI222_X1 U43 ( .A1(N43), .A2(n9), .B1(N238), .B2(n6), .C1(N11), .C2(n3), 
        .ZN(n37) );
  AOI222_X1 U44 ( .A1(N42), .A2(n9), .B1(N237), .B2(n6), .C1(N10), .C2(n3), 
        .ZN(n39) );
  AOI222_X1 U45 ( .A1(N69), .A2(n8), .B1(N264), .B2(n5), .C1(N37), .C2(n2), 
        .ZN(n43) );
  AOI222_X1 U46 ( .A1(N68), .A2(n8), .B1(N263), .B2(n5), .C1(N36), .C2(n2), 
        .ZN(n47) );
  AOI222_X1 U47 ( .A1(N67), .A2(n8), .B1(N262), .B2(n5), .C1(N35), .C2(n2), 
        .ZN(n49) );
  AOI222_X1 U48 ( .A1(N66), .A2(n8), .B1(N261), .B2(n5), .C1(N34), .C2(n2), 
        .ZN(n51) );
  AOI222_X1 U49 ( .A1(N65), .A2(n8), .B1(N260), .B2(n5), .C1(N33), .C2(n2), 
        .ZN(n53) );
  AOI222_X1 U50 ( .A1(N64), .A2(n8), .B1(N259), .B2(n5), .C1(N32), .C2(n2), 
        .ZN(n55) );
  AOI222_X1 U51 ( .A1(N63), .A2(n8), .B1(N258), .B2(n5), .C1(N31), .C2(n2), 
        .ZN(n57) );
  AOI222_X1 U52 ( .A1(N62), .A2(n8), .B1(N257), .B2(n5), .C1(N30), .C2(n2), 
        .ZN(n59) );
  AOI222_X1 U53 ( .A1(N61), .A2(n8), .B1(N256), .B2(n5), .C1(N29), .C2(n2), 
        .ZN(n61) );
  AOI222_X1 U54 ( .A1(N60), .A2(n8), .B1(N255), .B2(n5), .C1(N28), .C2(n2), 
        .ZN(n63) );
  AOI222_X1 U55 ( .A1(N59), .A2(n8), .B1(N254), .B2(n5), .C1(N27), .C2(n2), 
        .ZN(n65) );
  AOI222_X1 U56 ( .A1(N58), .A2(n7), .B1(N253), .B2(n4), .C1(N26), .C2(n1), 
        .ZN(n69) );
  AOI222_X1 U57 ( .A1(N57), .A2(n7), .B1(N252), .B2(n4), .C1(N25), .C2(n1), 
        .ZN(n71) );
  AOI222_X1 U58 ( .A1(N56), .A2(n7), .B1(N251), .B2(n4), .C1(N24), .C2(n1), 
        .ZN(n73) );
  AOI222_X1 U59 ( .A1(N55), .A2(n7), .B1(N250), .B2(n4), .C1(N23), .C2(n1), 
        .ZN(n75) );
  AOI222_X1 U60 ( .A1(N54), .A2(n7), .B1(N249), .B2(n4), .C1(N22), .C2(n1), 
        .ZN(n77) );
  AOI222_X1 U61 ( .A1(N53), .A2(n7), .B1(N248), .B2(n4), .C1(N21), .C2(n1), 
        .ZN(n79) );
  AOI222_X1 U62 ( .A1(N52), .A2(n7), .B1(N247), .B2(n4), .C1(N20), .C2(n1), 
        .ZN(n81) );
  AOI222_X1 U63 ( .A1(N51), .A2(n7), .B1(N246), .B2(n4), .C1(N19), .C2(n1), 
        .ZN(n83) );
  AOI222_X1 U64 ( .A1(N50), .A2(n7), .B1(N245), .B2(n4), .C1(N18), .C2(n1), 
        .ZN(n85) );
  AOI222_X1 U65 ( .A1(N49), .A2(n7), .B1(N244), .B2(n4), .C1(N17), .C2(n1), 
        .ZN(n87) );
  AOI222_X1 U66 ( .A1(N41), .A2(n8), .B1(N236), .B2(n5), .C1(N9), .C2(n2), 
        .ZN(n45) );
  AOI222_X1 U67 ( .A1(N40), .A2(n7), .B1(N235), .B2(n4), .C1(N8), .C2(n1), 
        .ZN(n67) );
  AOI222_X1 U68 ( .A1(N39), .A2(n7), .B1(N234), .B2(n4), .C1(N7), .C2(n1), 
        .ZN(n89) );
  BUF_X1 U69 ( .A(n24), .Z(n20) );
  BUF_X1 U70 ( .A(n24), .Z(n19) );
  BUF_X1 U71 ( .A(n25), .Z(n11) );
  BUF_X1 U72 ( .A(n25), .Z(n10) );
  BUF_X1 U73 ( .A(n24), .Z(n93) );
  BUF_X1 U74 ( .A(n25), .Z(n12) );
  BUF_X1 U75 ( .A(B[4]), .Z(n97) );
  NAND2_X1 U76 ( .A1(n41), .A2(n42), .ZN(OUTPUT[31]) );
  NAND2_X1 U77 ( .A1(n43), .A2(n44), .ZN(OUTPUT[30]) );
  NAND2_X1 U78 ( .A1(n47), .A2(n48), .ZN(OUTPUT[29]) );
  NAND2_X1 U79 ( .A1(n49), .A2(n50), .ZN(OUTPUT[28]) );
  NAND2_X1 U80 ( .A1(n51), .A2(n52), .ZN(OUTPUT[27]) );
  NAND2_X1 U81 ( .A1(n53), .A2(n54), .ZN(OUTPUT[26]) );
  NAND2_X1 U82 ( .A1(n55), .A2(n56), .ZN(OUTPUT[25]) );
  NAND2_X1 U83 ( .A1(n57), .A2(n58), .ZN(OUTPUT[24]) );
  NAND2_X1 U84 ( .A1(n59), .A2(n60), .ZN(OUTPUT[23]) );
  NAND2_X1 U85 ( .A1(n61), .A2(n62), .ZN(OUTPUT[22]) );
  NAND2_X1 U86 ( .A1(n63), .A2(n64), .ZN(OUTPUT[21]) );
  NAND2_X1 U87 ( .A1(n65), .A2(n66), .ZN(OUTPUT[20]) );
  NAND2_X1 U88 ( .A1(n69), .A2(n70), .ZN(OUTPUT[19]) );
  NAND2_X1 U89 ( .A1(n71), .A2(n72), .ZN(OUTPUT[18]) );
  NAND2_X1 U90 ( .A1(n73), .A2(n74), .ZN(OUTPUT[17]) );
  NAND2_X1 U91 ( .A1(n75), .A2(n76), .ZN(OUTPUT[16]) );
  NAND2_X1 U92 ( .A1(n77), .A2(n78), .ZN(OUTPUT[15]) );
  NAND2_X1 U93 ( .A1(n79), .A2(n80), .ZN(OUTPUT[14]) );
  NAND2_X1 U94 ( .A1(n81), .A2(n82), .ZN(OUTPUT[13]) );
  NAND2_X1 U95 ( .A1(n83), .A2(n84), .ZN(OUTPUT[12]) );
  NAND2_X1 U96 ( .A1(n85), .A2(n86), .ZN(OUTPUT[11]) );
  NAND2_X1 U97 ( .A1(n87), .A2(n88), .ZN(OUTPUT[10]) );
  NAND2_X1 U98 ( .A1(n21), .A2(n22), .ZN(OUTPUT[9]) );
  NAND2_X1 U99 ( .A1(n29), .A2(n30), .ZN(OUTPUT[8]) );
  NAND2_X1 U100 ( .A1(n31), .A2(n32), .ZN(OUTPUT[7]) );
  NAND2_X1 U101 ( .A1(n33), .A2(n34), .ZN(OUTPUT[6]) );
  NAND2_X1 U102 ( .A1(n35), .A2(n36), .ZN(OUTPUT[5]) );
  NAND2_X1 U103 ( .A1(n37), .A2(n38), .ZN(OUTPUT[4]) );
  AOI222_X1 U104 ( .A1(N233), .A2(n96), .B1(N136), .B2(n93), .C1(N168), .C2(
        n12), .ZN(n42) );
  AOI222_X1 U105 ( .A1(N202), .A2(n94), .B1(N105), .B2(n19), .C1(N137), .C2(
        n10), .ZN(n90) );
  BUF_X1 U106 ( .A(n27), .Z(n5) );
  BUF_X1 U107 ( .A(n27), .Z(n4) );
  BUF_X1 U108 ( .A(n28), .Z(n2) );
  BUF_X1 U109 ( .A(n28), .Z(n1) );
  BUF_X1 U110 ( .A(n26), .Z(n8) );
  BUF_X1 U111 ( .A(n26), .Z(n7) );
  BUF_X1 U112 ( .A(n23), .Z(n95) );
  BUF_X1 U113 ( .A(n23), .Z(n94) );
  BUF_X1 U114 ( .A(n27), .Z(n6) );
  BUF_X1 U115 ( .A(n28), .Z(n3) );
  BUF_X1 U116 ( .A(n26), .Z(n9) );
  BUF_X1 U117 ( .A(n23), .Z(n96) );
  AND2_X1 U118 ( .A1(n92), .A2(n98), .ZN(n24) );
  AND2_X1 U119 ( .A1(n91), .A2(n98), .ZN(n25) );
  NAND2_X1 U120 ( .A1(n39), .A2(n40), .ZN(OUTPUT[3]) );
  NAND2_X1 U121 ( .A1(n45), .A2(n46), .ZN(OUTPUT[2]) );
  NAND2_X1 U122 ( .A1(n67), .A2(n68), .ZN(OUTPUT[1]) );
  NOR2_X1 U123 ( .A1(LEFT_RIGHT), .A2(SHIFT_ROTATE), .ZN(n28) );
  NOR2_X1 U124 ( .A1(n98), .A2(SHIFT_ROTATE), .ZN(n26) );
  NOR2_X1 U125 ( .A1(n99), .A2(LOGIC_ARITH), .ZN(n92) );
  INV_X1 U126 ( .A(SHIFT_ROTATE), .ZN(n99) );
  AND2_X1 U127 ( .A1(LEFT_RIGHT), .A2(n92), .ZN(n23) );
  AND2_X1 U128 ( .A1(LEFT_RIGHT), .A2(n91), .ZN(n27) );
  INV_X1 U129 ( .A(LEFT_RIGHT), .ZN(n98) );
  AND2_X1 U130 ( .A1(LOGIC_ARITH), .A2(SHIFT_ROTATE), .ZN(n91) );
  NAND2_X1 U131 ( .A1(n89), .A2(n90), .ZN(OUTPUT[0]) );
endmodule


module G_0 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_43 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_0 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_0 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_43 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_0 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_52 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module G_42 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_42 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_42 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_42 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_42 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_41 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_41 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_41 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_41 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_41 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_40 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_40 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_40 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_40 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_40 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_39 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_39 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_39 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_39 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_39 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_38 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_38 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_38 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_38 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_38 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_37 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_37 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_37 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_37 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_37 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_36 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_36 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_36 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_36 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_36 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_35 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_35 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_35 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_35 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_35 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_34 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_34 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_34 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_34 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_34 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_33 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_33 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_33 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_33 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_33 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_32 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_32 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_32 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_32 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_32 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_31 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_31 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_31 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_31 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_31 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_30 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_30 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_30 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_30 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_30 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_29 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_29 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_29 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_29 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_29 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_28 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_28 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_28 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_28 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_28 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_27 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_27 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_27 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_27 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_27 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_26 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_26 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_26 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_26 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_26 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_25 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_25 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_25 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_25 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_25 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_24 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_24 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_24 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_24 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_24 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_23 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_23 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_23 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_23 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_23 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_22 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_22 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_22 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_22 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_22 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_21 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_21 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_21 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_21 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_21 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_20 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_20 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_20 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_20 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_20 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_19 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_19 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_19 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_19 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_19 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_18 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_18 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_18 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_18 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_18 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_17 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_17 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_17 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_17 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_17 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_16 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_16 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_16 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_16 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_16 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_15 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_15 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_15 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_15 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_15 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_14 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_14 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_14 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_14 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_14 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_13 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_13 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_13 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_13 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_13 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_51 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module G_12 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_12 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_12 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_12 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_12 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_11 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_11 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_11 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_11 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_11 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_10 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_10 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_10 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_10 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_10 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_9 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_9 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_9 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_9 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_9 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_8 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_8 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_8 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_8 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_8 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_7 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_7 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_7 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_7 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_7 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_6 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_6 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_6 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_6 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_6 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_50 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module G_5 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_5 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_5 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_5 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_5 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_4 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_4 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_4 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_4 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_4 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_3 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_3 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_3 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_3 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_3 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_49 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module G_48 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module G_2 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_2 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_2 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_2 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_2 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_1 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module P_1 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_1 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_1 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_1 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_47 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module G_46 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module G_45 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module G_44 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n3) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   \gi[32][4] , \gi[32][3] , \gi[32][2] , \gi[32][1] , \gi[32][0] ,
         \gi[31][0] , \gi[30][0] , \gi[29][0] , \gi[28][4] , \gi[28][2] ,
         \gi[28][1] , \gi[28][0] , \gi[27][0] , \gi[26][0] , \gi[25][0] ,
         \gi[24][3] , \gi[24][2] , \gi[24][1] , \gi[24][0] , \gi[23][0] ,
         \gi[22][0] , \gi[21][0] , \gi[20][2] , \gi[20][1] , \gi[20][0] ,
         \gi[19][0] , \gi[18][0] , \gi[17][0] , \gi[16][3] , \gi[16][2] ,
         \gi[16][1] , \gi[16][0] , \gi[15][0] , \gi[14][0] , \gi[13][0] ,
         \gi[12][2] , \gi[12][1] , \gi[12][0] , \gi[11][0] , \gi[10][0] ,
         \gi[9][0] , \gi[8][2] , \gi[8][1] , \gi[8][0] , \gi[7][0] ,
         \gi[6][0] , \gi[5][0] , \gi[4][1] , \gi[4][0] , \gi[3][0] ,
         \gi[2][1] , \gi[2][0] , \gi[1][0] , \gi[0][0] , \pi[32][4] ,
         \pi[32][3] , \pi[32][2] , \pi[32][1] , \pi[32][0] , \pi[31][0] ,
         \pi[30][0] , \pi[29][0] , \pi[28][4] , \pi[28][2] , \pi[28][1] ,
         \pi[28][0] , \pi[27][0] , \pi[26][0] , \pi[25][0] , \pi[24][3] ,
         \pi[24][2] , \pi[24][1] , \pi[24][0] , \pi[23][0] , \pi[22][0] ,
         \pi[21][0] , \pi[20][2] , \pi[20][1] , \pi[20][0] , \pi[19][0] ,
         \pi[18][0] , \pi[17][0] , \pi[16][3] , \pi[16][2] , \pi[16][1] ,
         \pi[16][0] , \pi[15][0] , \pi[14][0] , \pi[13][0] , \pi[12][2] ,
         \pi[12][1] , \pi[12][0] , \pi[11][0] , \pi[10][0] , \pi[9][0] ,
         \pi[8][2] , \pi[8][1] , \pi[8][0] , \pi[7][0] , \pi[6][0] ,
         \pi[5][0] , \pi[4][1] , \pi[4][0] , \pi[3][0] , \pi[2][0] ,
         \pi[0][0] ;

  XOR2_X1 U34 ( .A(B[8]), .B(A[8]), .Z(\pi[9][0] ) );
  XOR2_X1 U35 ( .A(B[7]), .B(A[7]), .Z(\pi[8][0] ) );
  XOR2_X1 U36 ( .A(B[6]), .B(A[6]), .Z(\pi[7][0] ) );
  XOR2_X1 U37 ( .A(B[5]), .B(A[5]), .Z(\pi[6][0] ) );
  XOR2_X1 U38 ( .A(B[4]), .B(A[4]), .Z(\pi[5][0] ) );
  XOR2_X1 U39 ( .A(B[3]), .B(A[3]), .Z(\pi[4][0] ) );
  XOR2_X1 U40 ( .A(B[2]), .B(A[2]), .Z(\pi[3][0] ) );
  XOR2_X1 U41 ( .A(B[31]), .B(A[31]), .Z(\pi[32][0] ) );
  XOR2_X1 U42 ( .A(B[30]), .B(A[30]), .Z(\pi[31][0] ) );
  XOR2_X1 U43 ( .A(B[29]), .B(A[29]), .Z(\pi[30][0] ) );
  XOR2_X1 U44 ( .A(B[1]), .B(A[1]), .Z(\pi[2][0] ) );
  XOR2_X1 U45 ( .A(B[28]), .B(A[28]), .Z(\pi[29][0] ) );
  XOR2_X1 U46 ( .A(B[27]), .B(A[27]), .Z(\pi[28][0] ) );
  XOR2_X1 U47 ( .A(B[26]), .B(A[26]), .Z(\pi[27][0] ) );
  XOR2_X1 U48 ( .A(B[25]), .B(A[25]), .Z(\pi[26][0] ) );
  XOR2_X1 U49 ( .A(B[24]), .B(A[24]), .Z(\pi[25][0] ) );
  XOR2_X1 U50 ( .A(B[23]), .B(A[23]), .Z(\pi[24][0] ) );
  XOR2_X1 U51 ( .A(B[22]), .B(A[22]), .Z(\pi[23][0] ) );
  XOR2_X1 U52 ( .A(B[21]), .B(A[21]), .Z(\pi[22][0] ) );
  XOR2_X1 U53 ( .A(B[20]), .B(A[20]), .Z(\pi[21][0] ) );
  XOR2_X1 U54 ( .A(B[19]), .B(A[19]), .Z(\pi[20][0] ) );
  XOR2_X1 U55 ( .A(B[18]), .B(A[18]), .Z(\pi[19][0] ) );
  XOR2_X1 U56 ( .A(B[17]), .B(A[17]), .Z(\pi[18][0] ) );
  XOR2_X1 U57 ( .A(B[16]), .B(A[16]), .Z(\pi[17][0] ) );
  XOR2_X1 U58 ( .A(B[15]), .B(A[15]), .Z(\pi[16][0] ) );
  XOR2_X1 U59 ( .A(B[14]), .B(A[14]), .Z(\pi[15][0] ) );
  XOR2_X1 U60 ( .A(B[13]), .B(A[13]), .Z(\pi[14][0] ) );
  XOR2_X1 U61 ( .A(B[12]), .B(A[12]), .Z(\pi[13][0] ) );
  XOR2_X1 U62 ( .A(B[11]), .B(A[11]), .Z(\pi[12][0] ) );
  XOR2_X1 U63 ( .A(B[10]), .B(A[10]), .Z(\pi[11][0] ) );
  XOR2_X1 U64 ( .A(B[9]), .B(A[9]), .Z(\pi[10][0] ) );
  XOR2_X1 U65 ( .A(B[0]), .B(A[0]), .Z(\pi[0][0] ) );
  G_0 g_port0_0_1 ( .G1(\gi[0][0] ), .P(\pi[0][0] ), .G2(Cin), .Co(\gi[1][0] )
         );
  PG_0 pg_port2_1_1 ( .G1(\gi[1][0] ), .P1(1'b0), .G2(\gi[0][0] ), .P2(
        \pi[0][0] ) );
  G_52 g_port1_1_2 ( .G1(\gi[2][0] ), .P(\pi[2][0] ), .G2(\gi[1][0] ), .Co(
        \gi[2][1] ) );
  PG_42 pg_port2_1_3 ( .G1(\gi[3][0] ), .P1(\pi[3][0] ), .G2(\gi[2][0] ), .P2(
        \pi[2][0] ) );
  PG_41 pg_port2_1_4 ( .G1(\gi[4][0] ), .P1(\pi[4][0] ), .G2(\gi[3][0] ), .P2(
        \pi[3][0] ), .gout(\gi[4][1] ), .pout(\pi[4][1] ) );
  PG_40 pg_port2_1_5 ( .G1(\gi[5][0] ), .P1(\pi[5][0] ), .G2(\gi[4][0] ), .P2(
        \pi[4][0] ) );
  PG_39 pg_port2_1_6 ( .G1(\gi[6][0] ), .P1(\pi[6][0] ), .G2(\gi[5][0] ), .P2(
        \pi[5][0] ) );
  PG_38 pg_port2_1_7 ( .G1(\gi[7][0] ), .P1(\pi[7][0] ), .G2(\gi[6][0] ), .P2(
        \pi[6][0] ) );
  PG_37 pg_port2_1_8 ( .G1(\gi[8][0] ), .P1(\pi[8][0] ), .G2(\gi[7][0] ), .P2(
        \pi[7][0] ), .gout(\gi[8][1] ), .pout(\pi[8][1] ) );
  PG_36 pg_port2_1_9 ( .G1(\gi[9][0] ), .P1(\pi[9][0] ), .G2(\gi[8][0] ), .P2(
        \pi[8][0] ) );
  PG_35 pg_port2_1_10 ( .G1(\gi[10][0] ), .P1(\pi[10][0] ), .G2(\gi[9][0] ), 
        .P2(\pi[9][0] ) );
  PG_34 pg_port2_1_11 ( .G1(\gi[11][0] ), .P1(\pi[11][0] ), .G2(\gi[10][0] ), 
        .P2(\pi[10][0] ) );
  PG_33 pg_port2_1_12 ( .G1(\gi[12][0] ), .P1(\pi[12][0] ), .G2(\gi[11][0] ), 
        .P2(\pi[11][0] ), .gout(\gi[12][1] ), .pout(\pi[12][1] ) );
  PG_32 pg_port2_1_13 ( .G1(\gi[13][0] ), .P1(\pi[13][0] ), .G2(\gi[12][0] ), 
        .P2(\pi[12][0] ) );
  PG_31 pg_port2_1_14 ( .G1(\gi[14][0] ), .P1(\pi[14][0] ), .G2(\gi[13][0] ), 
        .P2(\pi[13][0] ) );
  PG_30 pg_port2_1_15 ( .G1(\gi[15][0] ), .P1(\pi[15][0] ), .G2(\gi[14][0] ), 
        .P2(\pi[14][0] ) );
  PG_29 pg_port2_1_16 ( .G1(\gi[16][0] ), .P1(\pi[16][0] ), .G2(\gi[15][0] ), 
        .P2(\pi[15][0] ), .gout(\gi[16][1] ), .pout(\pi[16][1] ) );
  PG_28 pg_port2_1_17 ( .G1(\gi[17][0] ), .P1(\pi[17][0] ), .G2(\gi[16][0] ), 
        .P2(\pi[16][0] ) );
  PG_27 pg_port2_1_18 ( .G1(\gi[18][0] ), .P1(\pi[18][0] ), .G2(\gi[17][0] ), 
        .P2(\pi[17][0] ) );
  PG_26 pg_port2_1_19 ( .G1(\gi[19][0] ), .P1(\pi[19][0] ), .G2(\gi[18][0] ), 
        .P2(\pi[18][0] ) );
  PG_25 pg_port2_1_20 ( .G1(\gi[20][0] ), .P1(\pi[20][0] ), .G2(\gi[19][0] ), 
        .P2(\pi[19][0] ), .gout(\gi[20][1] ), .pout(\pi[20][1] ) );
  PG_24 pg_port2_1_21 ( .G1(\gi[21][0] ), .P1(\pi[21][0] ), .G2(\gi[20][0] ), 
        .P2(\pi[20][0] ) );
  PG_23 pg_port2_1_22 ( .G1(\gi[22][0] ), .P1(\pi[22][0] ), .G2(\gi[21][0] ), 
        .P2(\pi[21][0] ) );
  PG_22 pg_port2_1_23 ( .G1(\gi[23][0] ), .P1(\pi[23][0] ), .G2(\gi[22][0] ), 
        .P2(\pi[22][0] ) );
  PG_21 pg_port2_1_24 ( .G1(\gi[24][0] ), .P1(\pi[24][0] ), .G2(\gi[23][0] ), 
        .P2(\pi[23][0] ), .gout(\gi[24][1] ), .pout(\pi[24][1] ) );
  PG_20 pg_port2_1_25 ( .G1(\gi[25][0] ), .P1(\pi[25][0] ), .G2(\gi[24][0] ), 
        .P2(\pi[24][0] ) );
  PG_19 pg_port2_1_26 ( .G1(\gi[26][0] ), .P1(\pi[26][0] ), .G2(\gi[25][0] ), 
        .P2(\pi[25][0] ) );
  PG_18 pg_port2_1_27 ( .G1(\gi[27][0] ), .P1(\pi[27][0] ), .G2(\gi[26][0] ), 
        .P2(\pi[26][0] ) );
  PG_17 pg_port2_1_28 ( .G1(\gi[28][0] ), .P1(\pi[28][0] ), .G2(\gi[27][0] ), 
        .P2(\pi[27][0] ), .gout(\gi[28][1] ), .pout(\pi[28][1] ) );
  PG_16 pg_port2_1_29 ( .G1(\gi[29][0] ), .P1(\pi[29][0] ), .G2(\gi[28][0] ), 
        .P2(\pi[28][0] ) );
  PG_15 pg_port2_1_30 ( .G1(\gi[30][0] ), .P1(\pi[30][0] ), .G2(\gi[29][0] ), 
        .P2(\pi[29][0] ) );
  PG_14 pg_port2_1_31 ( .G1(\gi[31][0] ), .P1(\pi[31][0] ), .G2(\gi[30][0] ), 
        .P2(\pi[30][0] ) );
  PG_13 pg_port2_1_32 ( .G1(\gi[32][0] ), .P1(\pi[32][0] ), .G2(\gi[31][0] ), 
        .P2(\pi[31][0] ), .gout(\gi[32][1] ), .pout(\pi[32][1] ) );
  G_51 g_port_0 ( .G1(\gi[4][1] ), .P(\pi[4][1] ), .G2(\gi[2][1] ), .Co(Co[0])
         );
  PG_12 pg_port2_0_1_2 ( .G1(\gi[8][1] ), .P1(\pi[8][1] ), .G2(\gi[4][1] ), 
        .P2(\pi[4][1] ), .gout(\gi[8][2] ), .pout(\pi[8][2] ) );
  PG_11 pg_port2_0_2_3 ( .G1(\gi[12][1] ), .P1(\pi[12][1] ), .G2(\gi[8][1] ), 
        .P2(\pi[8][1] ), .gout(\gi[12][2] ), .pout(\pi[12][2] ) );
  PG_10 pg_port2_0_3_4 ( .G1(\gi[16][1] ), .P1(\pi[16][1] ), .G2(\gi[12][1] ), 
        .P2(\pi[12][1] ), .gout(\gi[16][2] ), .pout(\pi[16][2] ) );
  PG_9 pg_port2_0_4_5 ( .G1(\gi[20][1] ), .P1(\pi[20][1] ), .G2(\gi[16][1] ), 
        .P2(\pi[16][1] ), .gout(\gi[20][2] ), .pout(\pi[20][2] ) );
  PG_8 pg_port2_0_5_6 ( .G1(\gi[24][1] ), .P1(\pi[24][1] ), .G2(\gi[20][1] ), 
        .P2(\pi[20][1] ), .gout(\gi[24][2] ), .pout(\pi[24][2] ) );
  PG_7 pg_port2_0_6_7 ( .G1(\gi[28][1] ), .P1(\pi[28][1] ), .G2(\gi[24][1] ), 
        .P2(\pi[24][1] ), .gout(\gi[28][2] ), .pout(\pi[28][2] ) );
  PG_6 pg_port2_0_7_8 ( .G1(\gi[32][1] ), .P1(\pi[32][1] ), .G2(\gi[28][1] ), 
        .P2(\pi[28][1] ), .gout(\gi[32][2] ), .pout(\pi[32][2] ) );
  G_50 g_port_1_2 ( .G1(\gi[8][2] ), .P(\pi[8][2] ), .G2(Co[0]), .Co(Co[1]) );
  PG_5 pg_port2_1_1_4 ( .G1(\gi[16][2] ), .P1(\pi[16][2] ), .G2(\gi[12][2] ), 
        .P2(\pi[12][2] ), .gout(\gi[16][3] ), .pout(\pi[16][3] ) );
  PG_4 pg_port2_1_2_6 ( .G1(\gi[24][2] ), .P1(\pi[24][2] ), .G2(\gi[20][2] ), 
        .P2(\pi[20][2] ), .gout(\gi[24][3] ), .pout(\pi[24][3] ) );
  PG_3 pg_port2_1_3_8 ( .G1(\gi[32][2] ), .P1(\pi[32][2] ), .G2(\gi[28][2] ), 
        .P2(\pi[28][2] ), .gout(\gi[32][3] ), .pout(\pi[32][3] ) );
  G_49 g_port_2_3 ( .G1(\gi[12][2] ), .P(\pi[12][2] ), .G2(Co[1]), .Co(Co[2])
         );
  G_48 g_port_2_4 ( .G1(\gi[16][3] ), .P(\pi[16][3] ), .G2(Co[1]), .Co(Co[3])
         );
  PG_2 pg_port2_2_1_7 ( .G1(\gi[28][2] ), .P1(\pi[28][2] ), .G2(\gi[24][3] ), 
        .P2(\pi[24][3] ), .gout(\gi[28][4] ), .pout(\pi[28][4] ) );
  PG_1 pg_port2_2_1_8 ( .G1(\gi[32][3] ), .P1(\pi[32][3] ), .G2(\gi[24][3] ), 
        .P2(\pi[24][3] ), .gout(\gi[32][4] ), .pout(\pi[32][4] ) );
  G_47 g_port_3_5 ( .G1(\gi[20][2] ), .P(\pi[20][2] ), .G2(Co[3]), .Co(Co[4])
         );
  G_46 g_port_3_6 ( .G1(\gi[24][3] ), .P(\pi[24][3] ), .G2(Co[3]), .Co(Co[5])
         );
  G_45 g_port_3_7 ( .G1(\gi[28][4] ), .P(\pi[28][4] ), .G2(Co[3]), .Co(Co[6])
         );
  G_44 g_port_3_8 ( .G1(\gi[32][4] ), .P(\pi[32][4] ), .G2(Co[3]), .Co(Co[7])
         );
  AND2_X1 U2 ( .A1(B[31]), .A2(A[31]), .ZN(\gi[32][0] ) );
  AND2_X1 U3 ( .A1(B[15]), .A2(A[15]), .ZN(\gi[16][0] ) );
  AND2_X1 U4 ( .A1(B[14]), .A2(A[14]), .ZN(\gi[15][0] ) );
  AND2_X1 U5 ( .A1(B[19]), .A2(A[19]), .ZN(\gi[20][0] ) );
  AND2_X1 U6 ( .A1(B[18]), .A2(A[18]), .ZN(\gi[19][0] ) );
  AND2_X1 U7 ( .A1(B[23]), .A2(A[23]), .ZN(\gi[24][0] ) );
  AND2_X1 U8 ( .A1(B[22]), .A2(A[22]), .ZN(\gi[23][0] ) );
  AND2_X1 U9 ( .A1(B[27]), .A2(A[27]), .ZN(\gi[28][0] ) );
  AND2_X1 U10 ( .A1(B[26]), .A2(A[26]), .ZN(\gi[27][0] ) );
  AND2_X1 U11 ( .A1(B[30]), .A2(A[30]), .ZN(\gi[31][0] ) );
  AND2_X1 U12 ( .A1(B[7]), .A2(A[7]), .ZN(\gi[8][0] ) );
  AND2_X1 U13 ( .A1(B[6]), .A2(A[6]), .ZN(\gi[7][0] ) );
  AND2_X1 U14 ( .A1(B[11]), .A2(A[11]), .ZN(\gi[12][0] ) );
  AND2_X1 U15 ( .A1(B[10]), .A2(A[10]), .ZN(\gi[11][0] ) );
  AND2_X1 U16 ( .A1(B[3]), .A2(A[3]), .ZN(\gi[4][0] ) );
  AND2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(\gi[3][0] ) );
  AND2_X1 U18 ( .A1(B[0]), .A2(A[0]), .ZN(\gi[0][0] ) );
  AND2_X1 U19 ( .A1(B[1]), .A2(A[1]), .ZN(\gi[2][0] ) );
  AND2_X1 U20 ( .A1(B[4]), .A2(A[4]), .ZN(\gi[5][0] ) );
  AND2_X1 U21 ( .A1(B[5]), .A2(A[5]), .ZN(\gi[6][0] ) );
  AND2_X1 U22 ( .A1(B[8]), .A2(A[8]), .ZN(\gi[9][0] ) );
  AND2_X1 U23 ( .A1(B[9]), .A2(A[9]), .ZN(\gi[10][0] ) );
  AND2_X1 U24 ( .A1(B[12]), .A2(A[12]), .ZN(\gi[13][0] ) );
  AND2_X1 U25 ( .A1(B[13]), .A2(A[13]), .ZN(\gi[14][0] ) );
  AND2_X1 U26 ( .A1(B[16]), .A2(A[16]), .ZN(\gi[17][0] ) );
  AND2_X1 U27 ( .A1(B[17]), .A2(A[17]), .ZN(\gi[18][0] ) );
  AND2_X1 U28 ( .A1(B[20]), .A2(A[20]), .ZN(\gi[21][0] ) );
  AND2_X1 U29 ( .A1(B[21]), .A2(A[21]), .ZN(\gi[22][0] ) );
  AND2_X1 U30 ( .A1(B[24]), .A2(A[24]), .ZN(\gi[25][0] ) );
  AND2_X1 U31 ( .A1(B[25]), .A2(A[25]), .ZN(\gi[26][0] ) );
  AND2_X1 U32 ( .A1(B[28]), .A2(A[28]), .ZN(\gi[29][0] ) );
  AND2_X1 U33 ( .A1(B[29]), .A2(A[29]), .ZN(\gi[30][0] ) );
endmodule


module RCA_NBIT4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_32 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_32 UIV ( .A(S), .Y(SB) );
  ND2_96 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_95 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_94 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31 UIV ( .A(S), .Y(SB) );
  ND2_93 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_92 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_91 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30 UIV ( .A(S), .Y(SB) );
  ND2_90 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_89 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_88 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_29 UIV ( .A(S), .Y(SB) );
  ND2_87 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_86 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_85 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_32 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_29 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_0 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_28 UIV ( .A(S), .Y(SB) );
  ND2_84 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_83 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_82 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_27 UIV ( .A(S), .Y(SB) );
  ND2_81 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_80 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_79 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_26 UIV ( .A(S), .Y(SB) );
  ND2_78 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_77 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_76 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_25 UIV ( .A(S), .Y(SB) );
  ND2_75 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_74 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_73 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_28 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_27 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_26 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_25 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_7 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_24 UIV ( .A(S), .Y(SB) );
  ND2_72 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_71 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_70 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_23 UIV ( .A(S), .Y(SB) );
  ND2_69 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_68 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_67 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_22 UIV ( .A(S), .Y(SB) );
  ND2_66 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_65 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_64 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_21 UIV ( .A(S), .Y(SB) );
  ND2_63 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_62 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_61 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_24 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_23 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_22 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_21 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_6 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_20 UIV ( .A(S), .Y(SB) );
  ND2_60 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_59 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_58 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_19 UIV ( .A(S), .Y(SB) );
  ND2_57 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_56 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_55 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_18 UIV ( .A(S), .Y(SB) );
  ND2_54 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_53 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_52 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_17 UIV ( .A(S), .Y(SB) );
  ND2_51 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_50 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_49 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_20 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_19 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_18 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_17 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_5 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_16 UIV ( .A(S), .Y(SB) );
  ND2_48 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_47 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_46 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_15 UIV ( .A(S), .Y(SB) );
  ND2_45 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_44 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_43 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_14 UIV ( .A(S), .Y(SB) );
  ND2_42 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_41 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_40 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_13 UIV ( .A(S), .Y(SB) );
  ND2_39 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_38 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_37 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_16 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_15 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_14 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_13 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_4 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_12 UIV ( .A(S), .Y(SB) );
  ND2_36 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_35 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_34 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_11 UIV ( .A(S), .Y(SB) );
  ND2_33 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_32 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_31 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_10 UIV ( .A(S), .Y(SB) );
  ND2_30 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_29 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_28 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_9 UIV ( .A(S), .Y(SB) );
  ND2_27 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_26 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_25 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_12 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_11 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_10 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_9 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_3 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_8 UIV ( .A(S), .Y(SB) );
  ND2_24 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_23 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_22 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_7 UIV ( .A(S), .Y(SB) );
  ND2_21 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_20 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_19 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_6 UIV ( .A(S), .Y(SB) );
  ND2_18 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_17 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_16 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_5 UIV ( .A(S), .Y(SB) );
  ND2_15 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_14 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_13 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_8 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_7 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_6 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_5 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_2 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_4 UIV ( .A(S), .Y(SB) );
  ND2_12 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_11 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_10 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_3 UIV ( .A(S), .Y(SB) );
  ND2_9 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_8 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_7 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_2 UIV ( .A(S), .Y(SB) );
  ND2_6 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_5 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_4 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_1 UIV ( .A(S), .Y(SB) );
  ND2_3 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_2 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_1 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_4 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_3 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_2 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_1 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_1 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSB_NBIT4_0 CSBI_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSB_NBIT4_7 CSBI_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSB_NBIT4_6 CSBI_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  CSB_NBIT4_5 CSBI_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(S[15:12]) );
  CSB_NBIT4_4 CSBI_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(S[19:16]) );
  CSB_NBIT4_3 CSBI_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(S[23:20]) );
  CSB_NBIT4_2 CSBI_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(S[27:24]) );
  CSB_NBIT4_1 CSBI_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28]) );
endmodule


module P4_ADDER_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [6:0] Cout_gen;

  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 carry_logic ( .A(A), .B(B), .Cin(Cin), 
        .Co({Cout, Cout_gen}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 sum_logic ( .A(A), .B(B), .Ci({
        Cout_gen, Cin}), .S(S) );
endmodule


module ALU_N32 ( CLK, .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , 
        \FUNC[1] , \FUNC[0] }), DATA1, DATA2, OUT_ALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUT_ALU;
  input CLK, \FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   Cout_i, \OUTPUT3[0] , LOGIC_ARITH_i, LEFT_RIGHT_i, Cin_i, N139, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163,
         N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174,
         N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185,
         N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, n48, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n49, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174;
  wire   [5:0] FUNC;
  wire   [31:0] OUTPUT_alu_i;
  wire   [31:0] OUTPUT4;
  wire   [31:0] OUTPUT2;
  wire   [31:0] OUTPUT1;
  wire   [31:0] data1i;
  wire   [31:0] data2i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  DLH_X1 Cin_i_reg ( .G(n19), .D(n1), .Q(Cin_i) );
  DLH_X1 \data2i_reg[31]  ( .G(n19), .D(N205), .Q(data2i[31]) );
  DLH_X1 \data2i_reg[30]  ( .G(n19), .D(N204), .Q(data2i[30]) );
  DLH_X1 \data2i_reg[29]  ( .G(n19), .D(N203), .Q(data2i[29]) );
  DLH_X1 \data2i_reg[28]  ( .G(n19), .D(N202), .Q(data2i[28]) );
  DLH_X1 \data2i_reg[27]  ( .G(n19), .D(N201), .Q(data2i[27]) );
  DLH_X1 \data2i_reg[26]  ( .G(n19), .D(N200), .Q(data2i[26]) );
  DLH_X1 \data2i_reg[25]  ( .G(n19), .D(N199), .Q(data2i[25]) );
  DLH_X1 \data2i_reg[24]  ( .G(n19), .D(N198), .Q(data2i[24]) );
  DLH_X1 \data2i_reg[23]  ( .G(n19), .D(N197), .Q(data2i[23]) );
  DLH_X1 \data2i_reg[22]  ( .G(n19), .D(N196), .Q(data2i[22]) );
  DLH_X1 \data2i_reg[21]  ( .G(n19), .D(N195), .Q(data2i[21]) );
  DLH_X1 \data2i_reg[20]  ( .G(n19), .D(N194), .Q(data2i[20]) );
  DLH_X1 \data2i_reg[19]  ( .G(n19), .D(N193), .Q(data2i[19]) );
  DLH_X1 \data2i_reg[18]  ( .G(n19), .D(N192), .Q(data2i[18]) );
  DLH_X1 \data2i_reg[17]  ( .G(n19), .D(N191), .Q(data2i[17]) );
  DLH_X1 \data2i_reg[16]  ( .G(n19), .D(N190), .Q(data2i[16]) );
  DLH_X1 \data2i_reg[15]  ( .G(n19), .D(N189), .Q(data2i[15]) );
  DLH_X1 \data2i_reg[14]  ( .G(n19), .D(N188), .Q(data2i[14]) );
  DLH_X1 \data2i_reg[13]  ( .G(n19), .D(N187), .Q(data2i[13]) );
  DLH_X1 \data2i_reg[12]  ( .G(n19), .D(N186), .Q(data2i[12]) );
  DLH_X1 \data2i_reg[11]  ( .G(n19), .D(N185), .Q(data2i[11]) );
  DLH_X1 \data2i_reg[10]  ( .G(n19), .D(N184), .Q(data2i[10]) );
  DLH_X1 \data2i_reg[9]  ( .G(n19), .D(N183), .Q(data2i[9]) );
  DLH_X1 \data2i_reg[8]  ( .G(n20), .D(N182), .Q(data2i[8]) );
  DLH_X1 \data2i_reg[7]  ( .G(n20), .D(N181), .Q(data2i[7]) );
  DLH_X1 \data2i_reg[6]  ( .G(n20), .D(N180), .Q(data2i[6]) );
  DLH_X1 \data2i_reg[5]  ( .G(n20), .D(N179), .Q(data2i[5]) );
  DLH_X1 \data2i_reg[4]  ( .G(n20), .D(N178), .Q(data2i[4]) );
  DLH_X1 \data2i_reg[3]  ( .G(n20), .D(N177), .Q(data2i[3]) );
  DLH_X1 \data2i_reg[2]  ( .G(n20), .D(N176), .Q(data2i[2]) );
  DLH_X1 \data2i_reg[1]  ( .G(n20), .D(N175), .Q(data2i[1]) );
  DLH_X1 \data2i_reg[0]  ( .G(n20), .D(N174), .Q(data2i[0]) );
  DLH_X1 \data1i_reg[31]  ( .G(n20), .D(DATA1[31]), .Q(data1i[31]) );
  DLH_X1 \data1i_reg[30]  ( .G(n20), .D(DATA1[30]), .Q(data1i[30]) );
  DLH_X1 \data1i_reg[29]  ( .G(n20), .D(DATA1[29]), .Q(data1i[29]) );
  DLH_X1 \data1i_reg[28]  ( .G(n20), .D(DATA1[28]), .Q(data1i[28]) );
  DLH_X1 \data1i_reg[27]  ( .G(n20), .D(DATA1[27]), .Q(data1i[27]) );
  DLH_X1 \data1i_reg[26]  ( .G(n20), .D(DATA1[26]), .Q(data1i[26]) );
  DLH_X1 \data1i_reg[25]  ( .G(n20), .D(DATA1[25]), .Q(data1i[25]) );
  DLH_X1 \data1i_reg[24]  ( .G(n20), .D(DATA1[24]), .Q(data1i[24]) );
  DLH_X1 \data1i_reg[23]  ( .G(n20), .D(DATA1[23]), .Q(data1i[23]) );
  DLH_X1 \data1i_reg[22]  ( .G(n20), .D(DATA1[22]), .Q(data1i[22]) );
  DLH_X1 \data1i_reg[21]  ( .G(n20), .D(DATA1[21]), .Q(data1i[21]) );
  DLH_X1 \data1i_reg[20]  ( .G(n20), .D(DATA1[20]), .Q(data1i[20]) );
  DLH_X1 \data1i_reg[19]  ( .G(n20), .D(DATA1[19]), .Q(data1i[19]) );
  DLH_X1 \data1i_reg[18]  ( .G(n20), .D(DATA1[18]), .Q(data1i[18]) );
  DLH_X1 \data1i_reg[17]  ( .G(n20), .D(DATA1[17]), .Q(data1i[17]) );
  DLH_X1 \data1i_reg[16]  ( .G(n20), .D(DATA1[16]), .Q(data1i[16]) );
  DLH_X1 \data1i_reg[15]  ( .G(n20), .D(DATA1[15]), .Q(data1i[15]) );
  DLH_X1 \data1i_reg[14]  ( .G(n20), .D(DATA1[14]), .Q(data1i[14]) );
  DLH_X1 \data1i_reg[13]  ( .G(n21), .D(DATA1[13]), .Q(data1i[13]) );
  DLH_X1 \data1i_reg[12]  ( .G(n21), .D(DATA1[12]), .Q(data1i[12]) );
  DLH_X1 \data1i_reg[11]  ( .G(n21), .D(DATA1[11]), .Q(data1i[11]) );
  DLH_X1 \data1i_reg[10]  ( .G(n21), .D(DATA1[10]), .Q(data1i[10]) );
  DLH_X1 \data1i_reg[9]  ( .G(n21), .D(DATA1[9]), .Q(data1i[9]) );
  DLH_X1 \data1i_reg[8]  ( .G(n21), .D(DATA1[8]), .Q(data1i[8]) );
  DLH_X1 \data1i_reg[7]  ( .G(n21), .D(DATA1[7]), .Q(data1i[7]) );
  DLH_X1 \data1i_reg[6]  ( .G(n21), .D(DATA1[6]), .Q(data1i[6]) );
  DLH_X1 \data1i_reg[5]  ( .G(n21), .D(DATA1[5]), .Q(data1i[5]) );
  DLH_X1 \data1i_reg[4]  ( .G(n21), .D(DATA1[4]), .Q(data1i[4]) );
  DLH_X1 \data1i_reg[3]  ( .G(n21), .D(DATA1[3]), .Q(data1i[3]) );
  DLH_X1 \data1i_reg[2]  ( .G(n21), .D(DATA1[2]), .Q(data1i[2]) );
  DLH_X1 \data1i_reg[1]  ( .G(n21), .D(DATA1[1]), .Q(data1i[1]) );
  DLH_X1 \data1i_reg[0]  ( .G(n21), .D(DATA1[0]), .Q(data1i[0]) );
  DLH_X1 LOGIC_ARITH_i_reg ( .G(n15), .D(n164), .Q(LOGIC_ARITH_i) );
  DLH_X1 LEFT_RIGHT_i_reg ( .G(n15), .D(n164), .Q(LEFT_RIGHT_i) );
  DLH_X1 \OUTPUT_alu_i_reg[0]  ( .G(n16), .D(N142), .Q(OUTPUT_alu_i[0]) );
  DFF_X1 \OUT_ALU_reg[0]  ( .D(OUTPUT_alu_i[0]), .CK(CLK), .Q(OUT_ALU[0]) );
  DLH_X1 \OUTPUT_alu_i_reg[1]  ( .G(n16), .D(N143), .Q(OUTPUT_alu_i[1]) );
  DFF_X1 \OUT_ALU_reg[1]  ( .D(OUTPUT_alu_i[1]), .CK(CLK), .Q(OUT_ALU[1]) );
  DLH_X1 \OUTPUT_alu_i_reg[2]  ( .G(n16), .D(N144), .Q(OUTPUT_alu_i[2]) );
  DFF_X1 \OUT_ALU_reg[2]  ( .D(OUTPUT_alu_i[2]), .CK(CLK), .Q(OUT_ALU[2]) );
  DLH_X1 \OUTPUT_alu_i_reg[3]  ( .G(n16), .D(N145), .Q(OUTPUT_alu_i[3]) );
  DFF_X1 \OUT_ALU_reg[3]  ( .D(OUTPUT_alu_i[3]), .CK(CLK), .Q(OUT_ALU[3]) );
  DLH_X1 \OUTPUT_alu_i_reg[4]  ( .G(n16), .D(N146), .Q(OUTPUT_alu_i[4]) );
  DFF_X1 \OUT_ALU_reg[4]  ( .D(OUTPUT_alu_i[4]), .CK(CLK), .Q(OUT_ALU[4]) );
  DLH_X1 \OUTPUT_alu_i_reg[5]  ( .G(n16), .D(N147), .Q(OUTPUT_alu_i[5]) );
  DFF_X1 \OUT_ALU_reg[5]  ( .D(OUTPUT_alu_i[5]), .CK(CLK), .Q(OUT_ALU[5]) );
  DLH_X1 \OUTPUT_alu_i_reg[6]  ( .G(n16), .D(N148), .Q(OUTPUT_alu_i[6]) );
  DFF_X1 \OUT_ALU_reg[6]  ( .D(OUTPUT_alu_i[6]), .CK(CLK), .Q(OUT_ALU[6]) );
  DLH_X1 \OUTPUT_alu_i_reg[7]  ( .G(n16), .D(N149), .Q(OUTPUT_alu_i[7]) );
  DFF_X1 \OUT_ALU_reg[7]  ( .D(OUTPUT_alu_i[7]), .CK(CLK), .Q(OUT_ALU[7]) );
  DLH_X1 \OUTPUT_alu_i_reg[8]  ( .G(n16), .D(N150), .Q(OUTPUT_alu_i[8]) );
  DFF_X1 \OUT_ALU_reg[8]  ( .D(OUTPUT_alu_i[8]), .CK(CLK), .Q(OUT_ALU[8]) );
  DLH_X1 \OUTPUT_alu_i_reg[9]  ( .G(n16), .D(N151), .Q(OUTPUT_alu_i[9]) );
  DFF_X1 \OUT_ALU_reg[9]  ( .D(OUTPUT_alu_i[9]), .CK(CLK), .Q(OUT_ALU[9]) );
  DLH_X1 \OUTPUT_alu_i_reg[10]  ( .G(n16), .D(N152), .Q(OUTPUT_alu_i[10]) );
  DFF_X1 \OUT_ALU_reg[10]  ( .D(OUTPUT_alu_i[10]), .CK(CLK), .Q(OUT_ALU[10])
         );
  DLH_X1 \OUTPUT_alu_i_reg[11]  ( .G(n17), .D(N153), .Q(OUTPUT_alu_i[11]) );
  DFF_X1 \OUT_ALU_reg[11]  ( .D(OUTPUT_alu_i[11]), .CK(CLK), .Q(OUT_ALU[11])
         );
  DLH_X1 \OUTPUT_alu_i_reg[12]  ( .G(n17), .D(N154), .Q(OUTPUT_alu_i[12]) );
  DFF_X1 \OUT_ALU_reg[12]  ( .D(OUTPUT_alu_i[12]), .CK(CLK), .Q(OUT_ALU[12])
         );
  DLH_X1 \OUTPUT_alu_i_reg[13]  ( .G(n17), .D(N155), .Q(OUTPUT_alu_i[13]) );
  DFF_X1 \OUT_ALU_reg[13]  ( .D(OUTPUT_alu_i[13]), .CK(CLK), .Q(OUT_ALU[13])
         );
  DLH_X1 \OUTPUT_alu_i_reg[14]  ( .G(n17), .D(N156), .Q(OUTPUT_alu_i[14]) );
  DFF_X1 \OUT_ALU_reg[14]  ( .D(OUTPUT_alu_i[14]), .CK(CLK), .Q(OUT_ALU[14])
         );
  DLH_X1 \OUTPUT_alu_i_reg[15]  ( .G(n17), .D(N157), .Q(OUTPUT_alu_i[15]) );
  DFF_X1 \OUT_ALU_reg[15]  ( .D(OUTPUT_alu_i[15]), .CK(CLK), .Q(OUT_ALU[15])
         );
  DLH_X1 \OUTPUT_alu_i_reg[16]  ( .G(n17), .D(N158), .Q(OUTPUT_alu_i[16]) );
  DFF_X1 \OUT_ALU_reg[16]  ( .D(OUTPUT_alu_i[16]), .CK(CLK), .Q(OUT_ALU[16])
         );
  DLH_X1 \OUTPUT_alu_i_reg[17]  ( .G(n17), .D(N159), .Q(OUTPUT_alu_i[17]) );
  DFF_X1 \OUT_ALU_reg[17]  ( .D(OUTPUT_alu_i[17]), .CK(CLK), .Q(OUT_ALU[17])
         );
  DLH_X1 \OUTPUT_alu_i_reg[18]  ( .G(n17), .D(N160), .Q(OUTPUT_alu_i[18]) );
  DFF_X1 \OUT_ALU_reg[18]  ( .D(OUTPUT_alu_i[18]), .CK(CLK), .Q(OUT_ALU[18])
         );
  DLH_X1 \OUTPUT_alu_i_reg[19]  ( .G(n17), .D(N161), .Q(OUTPUT_alu_i[19]) );
  DFF_X1 \OUT_ALU_reg[19]  ( .D(OUTPUT_alu_i[19]), .CK(CLK), .Q(OUT_ALU[19])
         );
  DLH_X1 \OUTPUT_alu_i_reg[20]  ( .G(n17), .D(N162), .Q(OUTPUT_alu_i[20]) );
  DFF_X1 \OUT_ALU_reg[20]  ( .D(OUTPUT_alu_i[20]), .CK(CLK), .Q(OUT_ALU[20])
         );
  DLH_X1 \OUTPUT_alu_i_reg[21]  ( .G(n17), .D(N163), .Q(OUTPUT_alu_i[21]) );
  DFF_X1 \OUT_ALU_reg[21]  ( .D(OUTPUT_alu_i[21]), .CK(CLK), .Q(OUT_ALU[21])
         );
  DLH_X1 \OUTPUT_alu_i_reg[22]  ( .G(n18), .D(N164), .Q(OUTPUT_alu_i[22]) );
  DFF_X1 \OUT_ALU_reg[22]  ( .D(OUTPUT_alu_i[22]), .CK(CLK), .Q(OUT_ALU[22])
         );
  DLH_X1 \OUTPUT_alu_i_reg[23]  ( .G(n18), .D(N165), .Q(OUTPUT_alu_i[23]) );
  DFF_X1 \OUT_ALU_reg[23]  ( .D(OUTPUT_alu_i[23]), .CK(CLK), .Q(OUT_ALU[23])
         );
  DLH_X1 \OUTPUT_alu_i_reg[24]  ( .G(n18), .D(N166), .Q(OUTPUT_alu_i[24]) );
  DFF_X1 \OUT_ALU_reg[24]  ( .D(OUTPUT_alu_i[24]), .CK(CLK), .Q(OUT_ALU[24])
         );
  DLH_X1 \OUTPUT_alu_i_reg[25]  ( .G(n18), .D(N167), .Q(OUTPUT_alu_i[25]) );
  DFF_X1 \OUT_ALU_reg[25]  ( .D(OUTPUT_alu_i[25]), .CK(CLK), .Q(OUT_ALU[25])
         );
  DLH_X1 \OUTPUT_alu_i_reg[26]  ( .G(n18), .D(N168), .Q(OUTPUT_alu_i[26]) );
  DFF_X1 \OUT_ALU_reg[26]  ( .D(OUTPUT_alu_i[26]), .CK(CLK), .Q(OUT_ALU[26])
         );
  DLH_X1 \OUTPUT_alu_i_reg[27]  ( .G(n18), .D(N169), .Q(OUTPUT_alu_i[27]) );
  DFF_X1 \OUT_ALU_reg[27]  ( .D(OUTPUT_alu_i[27]), .CK(CLK), .Q(OUT_ALU[27])
         );
  DLH_X1 \OUTPUT_alu_i_reg[28]  ( .G(n18), .D(N170), .Q(OUTPUT_alu_i[28]) );
  DFF_X1 \OUT_ALU_reg[28]  ( .D(OUTPUT_alu_i[28]), .CK(CLK), .Q(OUT_ALU[28])
         );
  DLH_X1 \OUTPUT_alu_i_reg[29]  ( .G(n18), .D(N171), .Q(OUTPUT_alu_i[29]) );
  DFF_X1 \OUT_ALU_reg[29]  ( .D(OUTPUT_alu_i[29]), .CK(CLK), .Q(OUT_ALU[29])
         );
  DLH_X1 \OUTPUT_alu_i_reg[30]  ( .G(n18), .D(N172), .Q(OUTPUT_alu_i[30]) );
  DFF_X1 \OUT_ALU_reg[30]  ( .D(OUTPUT_alu_i[30]), .CK(CLK), .Q(OUT_ALU[30])
         );
  DLH_X1 \OUTPUT_alu_i_reg[31]  ( .G(n18), .D(N173), .Q(OUTPUT_alu_i[31]) );
  DFF_X1 \OUT_ALU_reg[31]  ( .D(OUTPUT_alu_i[31]), .CK(CLK), .Q(OUT_ALU[31])
         );
  NAND3_X1 U221 ( .A1(n144), .A2(n143), .A3(n152), .ZN(n149) );
  NAND3_X1 U222 ( .A1(n133), .A2(n168), .A3(FUNC[2]), .ZN(n143) );
  NAND3_X1 U223 ( .A1(n147), .A2(n168), .A3(FUNC[2]), .ZN(n122) );
  logic_N32 log ( .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , 
        \FUNC[0] }), .DATA1(DATA1), .DATA2({DATA2[31:4], n26, n24, DATA2[1:0]}), .OUT_ALU(OUTPUT4) );
  comparator comp ( .DATA1(OUTPUT2), .DATA2i(Cout_i), .tipo({\FUNC[5] , 
        \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }), .OUTALU({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, \OUTPUT3[0] }) );
  SHIFTER_GENERIC_N32 shifter ( .A(DATA1), .B({DATA2[4], n26, n24, DATA2[1:0]}), .LOGIC_ARITH(LOGIC_ARITH_i), .LEFT_RIGHT(LEFT_RIGHT_i), .SHIFT_ROTATE(1'b1), 
        .OUTPUT(OUTPUT1) );
  P4_ADDER_NBIT32 adder ( .A(data1i), .B(data2i), .Cin(Cin_i), .S(OUTPUT2), 
        .Cout(Cout_i) );
  BUF_X1 U4 ( .A(N139), .Z(n20) );
  BUF_X1 U5 ( .A(n53), .Z(n8) );
  BUF_X1 U6 ( .A(n53), .Z(n9) );
  INV_X1 U7 ( .A(n1), .ZN(n11) );
  INV_X1 U8 ( .A(n1), .ZN(n12) );
  BUF_X1 U9 ( .A(N139), .Z(n19) );
  BUF_X1 U10 ( .A(n162), .Z(n2) );
  BUF_X1 U11 ( .A(n162), .Z(n3) );
  BUF_X1 U12 ( .A(n162), .Z(n4) );
  BUF_X1 U13 ( .A(n53), .Z(n10) );
  BUF_X1 U14 ( .A(N139), .Z(n21) );
  BUF_X1 U15 ( .A(N141), .Z(n17) );
  BUF_X1 U16 ( .A(N141), .Z(n16) );
  BUF_X1 U17 ( .A(N141), .Z(n18) );
  AOI21_X1 U18 ( .B1(n152), .B2(n120), .A(n171), .ZN(n134) );
  BUF_X1 U19 ( .A(n54), .Z(n5) );
  BUF_X1 U20 ( .A(n54), .Z(n6) );
  BUF_X1 U21 ( .A(n54), .Z(n7) );
  OR3_X1 U22 ( .A1(n134), .A2(n135), .A3(n55), .ZN(n1) );
  INV_X1 U23 ( .A(n50), .ZN(n162) );
  NAND2_X1 U24 ( .A1(n132), .A2(n123), .ZN(n130) );
  NAND2_X1 U25 ( .A1(n124), .A2(n171), .ZN(n140) );
  OR3_X1 U26 ( .A1(n134), .A2(n135), .A3(n50), .ZN(n53) );
  OR2_X1 U27 ( .A1(n10), .A2(n55), .ZN(N139) );
  OR3_X1 U28 ( .A1(n19), .A2(n15), .A3(n7), .ZN(N141) );
  INV_X1 U29 ( .A(n142), .ZN(n167) );
  NAND2_X1 U30 ( .A1(n51), .A2(n52), .ZN(N173) );
  NAND2_X1 U31 ( .A1(OUTPUT1[31]), .A2(n13), .ZN(n51) );
  AOI22_X1 U32 ( .A1(OUTPUT2[31]), .A2(n8), .B1(OUTPUT4[31]), .B2(n5), .ZN(n52) );
  NAND2_X1 U33 ( .A1(n56), .A2(n57), .ZN(N172) );
  NAND2_X1 U34 ( .A1(OUTPUT1[30]), .A2(n15), .ZN(n56) );
  AOI22_X1 U35 ( .A1(OUTPUT2[30]), .A2(n8), .B1(OUTPUT4[30]), .B2(n5), .ZN(n57) );
  NAND2_X1 U36 ( .A1(n58), .A2(n59), .ZN(N171) );
  NAND2_X1 U37 ( .A1(OUTPUT1[29]), .A2(n15), .ZN(n58) );
  AOI22_X1 U38 ( .A1(OUTPUT2[29]), .A2(n8), .B1(OUTPUT4[29]), .B2(n5), .ZN(n59) );
  NAND2_X1 U39 ( .A1(n60), .A2(n61), .ZN(N170) );
  NAND2_X1 U40 ( .A1(OUTPUT1[28]), .A2(n15), .ZN(n60) );
  AOI22_X1 U41 ( .A1(OUTPUT2[28]), .A2(n8), .B1(OUTPUT4[28]), .B2(n5), .ZN(n61) );
  NAND2_X1 U42 ( .A1(n62), .A2(n63), .ZN(N169) );
  NAND2_X1 U43 ( .A1(OUTPUT1[27]), .A2(n15), .ZN(n62) );
  AOI22_X1 U44 ( .A1(OUTPUT2[27]), .A2(n8), .B1(OUTPUT4[27]), .B2(n5), .ZN(n63) );
  NAND2_X1 U45 ( .A1(n64), .A2(n65), .ZN(N168) );
  NAND2_X1 U46 ( .A1(OUTPUT1[26]), .A2(n15), .ZN(n64) );
  AOI22_X1 U47 ( .A1(OUTPUT2[26]), .A2(n8), .B1(OUTPUT4[26]), .B2(n5), .ZN(n65) );
  NAND2_X1 U48 ( .A1(n66), .A2(n67), .ZN(N167) );
  NAND2_X1 U49 ( .A1(OUTPUT1[25]), .A2(n15), .ZN(n66) );
  AOI22_X1 U50 ( .A1(OUTPUT2[25]), .A2(n8), .B1(OUTPUT4[25]), .B2(n5), .ZN(n67) );
  NAND2_X1 U51 ( .A1(n68), .A2(n69), .ZN(N166) );
  NAND2_X1 U52 ( .A1(OUTPUT1[24]), .A2(n15), .ZN(n68) );
  AOI22_X1 U53 ( .A1(OUTPUT2[24]), .A2(n8), .B1(OUTPUT4[24]), .B2(n5), .ZN(n69) );
  NAND2_X1 U54 ( .A1(n70), .A2(n71), .ZN(N165) );
  NAND2_X1 U55 ( .A1(OUTPUT1[23]), .A2(n14), .ZN(n70) );
  AOI22_X1 U56 ( .A1(OUTPUT2[23]), .A2(n8), .B1(OUTPUT4[23]), .B2(n5), .ZN(n71) );
  NAND2_X1 U57 ( .A1(n72), .A2(n73), .ZN(N164) );
  NAND2_X1 U58 ( .A1(OUTPUT1[22]), .A2(n14), .ZN(n72) );
  AOI22_X1 U59 ( .A1(OUTPUT2[22]), .A2(n8), .B1(OUTPUT4[22]), .B2(n5), .ZN(n73) );
  NAND2_X1 U60 ( .A1(n74), .A2(n75), .ZN(N163) );
  NAND2_X1 U61 ( .A1(OUTPUT1[21]), .A2(n14), .ZN(n74) );
  AOI22_X1 U62 ( .A1(OUTPUT2[21]), .A2(n8), .B1(OUTPUT4[21]), .B2(n5), .ZN(n75) );
  NAND2_X1 U63 ( .A1(n76), .A2(n77), .ZN(N162) );
  NAND2_X1 U64 ( .A1(OUTPUT1[20]), .A2(n14), .ZN(n76) );
  AOI22_X1 U65 ( .A1(OUTPUT2[20]), .A2(n8), .B1(OUTPUT4[20]), .B2(n5), .ZN(n77) );
  NAND2_X1 U66 ( .A1(n78), .A2(n79), .ZN(N161) );
  NAND2_X1 U67 ( .A1(OUTPUT1[19]), .A2(n14), .ZN(n78) );
  AOI22_X1 U68 ( .A1(OUTPUT2[19]), .A2(n9), .B1(OUTPUT4[19]), .B2(n6), .ZN(n79) );
  NAND2_X1 U69 ( .A1(n80), .A2(n81), .ZN(N160) );
  NAND2_X1 U70 ( .A1(OUTPUT1[18]), .A2(n14), .ZN(n80) );
  AOI22_X1 U71 ( .A1(OUTPUT2[18]), .A2(n9), .B1(OUTPUT4[18]), .B2(n6), .ZN(n81) );
  NAND2_X1 U72 ( .A1(n82), .A2(n83), .ZN(N159) );
  NAND2_X1 U73 ( .A1(OUTPUT1[17]), .A2(n14), .ZN(n82) );
  AOI22_X1 U74 ( .A1(OUTPUT2[17]), .A2(n9), .B1(OUTPUT4[17]), .B2(n6), .ZN(n83) );
  NAND2_X1 U75 ( .A1(n84), .A2(n85), .ZN(N158) );
  NAND2_X1 U76 ( .A1(OUTPUT1[16]), .A2(n14), .ZN(n84) );
  AOI22_X1 U77 ( .A1(OUTPUT2[16]), .A2(n9), .B1(OUTPUT4[16]), .B2(n6), .ZN(n85) );
  NAND2_X1 U78 ( .A1(n86), .A2(n87), .ZN(N157) );
  NAND2_X1 U79 ( .A1(OUTPUT1[15]), .A2(n14), .ZN(n86) );
  AOI22_X1 U80 ( .A1(OUTPUT2[15]), .A2(n9), .B1(OUTPUT4[15]), .B2(n6), .ZN(n87) );
  NAND2_X1 U81 ( .A1(n88), .A2(n89), .ZN(N156) );
  NAND2_X1 U82 ( .A1(OUTPUT1[14]), .A2(n14), .ZN(n88) );
  AOI22_X1 U83 ( .A1(OUTPUT2[14]), .A2(n9), .B1(OUTPUT4[14]), .B2(n6), .ZN(n89) );
  NAND2_X1 U84 ( .A1(n90), .A2(n91), .ZN(N155) );
  NAND2_X1 U85 ( .A1(OUTPUT1[13]), .A2(n14), .ZN(n90) );
  AOI22_X1 U86 ( .A1(OUTPUT2[13]), .A2(n9), .B1(OUTPUT4[13]), .B2(n6), .ZN(n91) );
  NAND2_X1 U87 ( .A1(n92), .A2(n93), .ZN(N154) );
  NAND2_X1 U88 ( .A1(OUTPUT1[12]), .A2(n13), .ZN(n92) );
  AOI22_X1 U89 ( .A1(OUTPUT2[12]), .A2(n9), .B1(OUTPUT4[12]), .B2(n6), .ZN(n93) );
  NAND2_X1 U90 ( .A1(n94), .A2(n95), .ZN(N153) );
  NAND2_X1 U91 ( .A1(OUTPUT1[11]), .A2(n13), .ZN(n94) );
  AOI22_X1 U92 ( .A1(OUTPUT2[11]), .A2(n9), .B1(OUTPUT4[11]), .B2(n6), .ZN(n95) );
  NAND2_X1 U93 ( .A1(n96), .A2(n97), .ZN(N152) );
  NAND2_X1 U94 ( .A1(OUTPUT1[10]), .A2(n13), .ZN(n96) );
  AOI22_X1 U95 ( .A1(OUTPUT2[10]), .A2(n9), .B1(OUTPUT4[10]), .B2(n6), .ZN(n97) );
  NAND2_X1 U96 ( .A1(n98), .A2(n99), .ZN(N151) );
  NAND2_X1 U97 ( .A1(OUTPUT1[9]), .A2(n13), .ZN(n98) );
  AOI22_X1 U98 ( .A1(OUTPUT2[9]), .A2(n9), .B1(OUTPUT4[9]), .B2(n6), .ZN(n99)
         );
  NAND2_X1 U99 ( .A1(n100), .A2(n101), .ZN(N150) );
  NAND2_X1 U100 ( .A1(OUTPUT1[8]), .A2(n13), .ZN(n100) );
  AOI22_X1 U101 ( .A1(OUTPUT2[8]), .A2(n9), .B1(OUTPUT4[8]), .B2(n6), .ZN(n101) );
  NAND2_X1 U102 ( .A1(n102), .A2(n103), .ZN(N149) );
  NAND2_X1 U103 ( .A1(OUTPUT1[7]), .A2(n13), .ZN(n102) );
  AOI22_X1 U104 ( .A1(OUTPUT2[7]), .A2(n10), .B1(OUTPUT4[7]), .B2(n7), .ZN(
        n103) );
  NAND2_X1 U105 ( .A1(n104), .A2(n105), .ZN(N148) );
  NAND2_X1 U106 ( .A1(OUTPUT1[6]), .A2(n13), .ZN(n104) );
  AOI22_X1 U107 ( .A1(OUTPUT2[6]), .A2(n10), .B1(OUTPUT4[6]), .B2(n7), .ZN(
        n105) );
  NAND2_X1 U108 ( .A1(n106), .A2(n107), .ZN(N147) );
  NAND2_X1 U109 ( .A1(OUTPUT1[5]), .A2(n14), .ZN(n106) );
  AOI22_X1 U110 ( .A1(OUTPUT2[5]), .A2(n10), .B1(OUTPUT4[5]), .B2(n7), .ZN(
        n107) );
  NAND2_X1 U111 ( .A1(n108), .A2(n109), .ZN(N146) );
  NAND2_X1 U112 ( .A1(OUTPUT1[4]), .A2(n13), .ZN(n108) );
  AOI22_X1 U113 ( .A1(OUTPUT2[4]), .A2(n10), .B1(OUTPUT4[4]), .B2(n7), .ZN(
        n109) );
  INV_X1 U114 ( .A(n48), .ZN(n164) );
  INV_X1 U115 ( .A(n27), .ZN(n26) );
  OAI221_X1 U116 ( .B1(n173), .B2(n118), .C1(n119), .C2(n120), .A(n165), .ZN(
        n54) );
  INV_X1 U117 ( .A(n121), .ZN(n165) );
  OAI22_X1 U118 ( .A1(n122), .A2(n170), .B1(n123), .B2(n124), .ZN(n121) );
  INV_X1 U119 ( .A(n125), .ZN(n170) );
  OAI221_X1 U120 ( .B1(n127), .B2(n118), .C1(n119), .C2(n136), .A(n137), .ZN(
        n55) );
  AOI221_X1 U121 ( .B1(n138), .B2(n125), .C1(n139), .C2(n140), .A(n141), .ZN(
        n137) );
  NAND2_X1 U122 ( .A1(n143), .A2(n144), .ZN(n139) );
  OAI211_X1 U123 ( .C1(n142), .C2(n161), .A(n118), .B(n126), .ZN(n138) );
  OAI221_X1 U124 ( .B1(n124), .B2(n120), .C1(n127), .C2(n132), .A(n148), .ZN(
        n50) );
  AOI222_X1 U125 ( .A1(n163), .A2(n140), .B1(n174), .B2(n149), .C1(n150), .C2(
        n151), .ZN(n148) );
  INV_X1 U126 ( .A(n136), .ZN(n163) );
  NOR2_X1 U127 ( .A1(n168), .A2(n169), .ZN(n153) );
  BUF_X1 U128 ( .A(N206), .Z(n15) );
  AOI21_X1 U129 ( .B1(n122), .B2(n152), .A(n127), .ZN(n135) );
  BUF_X1 U130 ( .A(N206), .Z(n14) );
  BUF_X1 U131 ( .A(N206), .Z(n13) );
  NOR3_X1 U132 ( .A1(n166), .A2(n124), .A3(n142), .ZN(n141) );
  OAI22_X1 U133 ( .A1(DATA2[1]), .A2(n11), .B1(n2), .B2(n23), .ZN(N175) );
  OAI22_X1 U134 ( .A1(n24), .A2(n11), .B1(n2), .B2(n25), .ZN(N176) );
  OAI22_X1 U135 ( .A1(DATA2[0]), .A2(n11), .B1(n2), .B2(n22), .ZN(N174) );
  OAI22_X1 U136 ( .A1(DATA2[24]), .A2(n11), .B1(n4), .B2(n36), .ZN(N198) );
  INV_X1 U137 ( .A(DATA2[24]), .ZN(n36) );
  OAI22_X1 U138 ( .A1(DATA2[25]), .A2(n12), .B1(n4), .B2(n35), .ZN(N199) );
  INV_X1 U139 ( .A(DATA2[25]), .ZN(n35) );
  OAI22_X1 U140 ( .A1(DATA2[26]), .A2(n11), .B1(n4), .B2(n34), .ZN(N200) );
  INV_X1 U141 ( .A(DATA2[26]), .ZN(n34) );
  OAI22_X1 U142 ( .A1(DATA2[27]), .A2(n12), .B1(n4), .B2(n33), .ZN(N201) );
  INV_X1 U143 ( .A(DATA2[27]), .ZN(n33) );
  OAI22_X1 U144 ( .A1(DATA2[28]), .A2(n11), .B1(n4), .B2(n32), .ZN(N202) );
  INV_X1 U145 ( .A(DATA2[28]), .ZN(n32) );
  OAI22_X1 U146 ( .A1(DATA2[29]), .A2(n12), .B1(n4), .B2(n31), .ZN(N203) );
  INV_X1 U147 ( .A(DATA2[29]), .ZN(n31) );
  OAI22_X1 U148 ( .A1(DATA2[30]), .A2(n11), .B1(n4), .B2(n30), .ZN(N204) );
  INV_X1 U149 ( .A(DATA2[30]), .ZN(n30) );
  OAI22_X1 U150 ( .A1(DATA2[31]), .A2(n12), .B1(n4), .B2(n29), .ZN(N205) );
  INV_X1 U151 ( .A(DATA2[31]), .ZN(n29) );
  OAI22_X1 U152 ( .A1(n26), .A2(n11), .B1(n2), .B2(n27), .ZN(N177) );
  OAI22_X1 U153 ( .A1(DATA2[4]), .A2(n11), .B1(n2), .B2(n28), .ZN(N178) );
  OAI22_X1 U154 ( .A1(DATA2[5]), .A2(n11), .B1(n2), .B2(n160), .ZN(N179) );
  INV_X1 U155 ( .A(DATA2[5]), .ZN(n160) );
  OAI22_X1 U156 ( .A1(DATA2[6]), .A2(n11), .B1(n2), .B2(n159), .ZN(N180) );
  INV_X1 U157 ( .A(DATA2[6]), .ZN(n159) );
  OAI22_X1 U158 ( .A1(DATA2[7]), .A2(n11), .B1(n2), .B2(n158), .ZN(N181) );
  INV_X1 U159 ( .A(DATA2[7]), .ZN(n158) );
  OAI22_X1 U160 ( .A1(DATA2[8]), .A2(n11), .B1(n2), .B2(n157), .ZN(N182) );
  INV_X1 U161 ( .A(DATA2[8]), .ZN(n157) );
  OAI22_X1 U162 ( .A1(DATA2[9]), .A2(n11), .B1(n2), .B2(n156), .ZN(N183) );
  INV_X1 U163 ( .A(DATA2[9]), .ZN(n156) );
  OAI22_X1 U164 ( .A1(DATA2[10]), .A2(n11), .B1(n2), .B2(n155), .ZN(N184) );
  INV_X1 U165 ( .A(DATA2[10]), .ZN(n155) );
  OAI22_X1 U166 ( .A1(DATA2[11]), .A2(n11), .B1(n2), .B2(n154), .ZN(N185) );
  INV_X1 U167 ( .A(DATA2[11]), .ZN(n154) );
  OAI22_X1 U168 ( .A1(DATA2[12]), .A2(n12), .B1(n3), .B2(n49), .ZN(N186) );
  INV_X1 U169 ( .A(DATA2[12]), .ZN(n49) );
  OAI22_X1 U170 ( .A1(DATA2[13]), .A2(n12), .B1(n3), .B2(n47), .ZN(N187) );
  INV_X1 U171 ( .A(DATA2[13]), .ZN(n47) );
  OAI22_X1 U172 ( .A1(DATA2[14]), .A2(n12), .B1(n3), .B2(n46), .ZN(N188) );
  INV_X1 U173 ( .A(DATA2[14]), .ZN(n46) );
  OAI22_X1 U174 ( .A1(DATA2[15]), .A2(n12), .B1(n3), .B2(n45), .ZN(N189) );
  INV_X1 U175 ( .A(DATA2[15]), .ZN(n45) );
  OAI22_X1 U176 ( .A1(DATA2[16]), .A2(n12), .B1(n3), .B2(n44), .ZN(N190) );
  INV_X1 U177 ( .A(DATA2[16]), .ZN(n44) );
  OAI22_X1 U178 ( .A1(DATA2[17]), .A2(n12), .B1(n3), .B2(n43), .ZN(N191) );
  INV_X1 U179 ( .A(DATA2[17]), .ZN(n43) );
  OAI22_X1 U180 ( .A1(DATA2[18]), .A2(n12), .B1(n3), .B2(n42), .ZN(N192) );
  INV_X1 U181 ( .A(DATA2[18]), .ZN(n42) );
  OAI22_X1 U182 ( .A1(DATA2[19]), .A2(n12), .B1(n3), .B2(n41), .ZN(N193) );
  INV_X1 U183 ( .A(DATA2[19]), .ZN(n41) );
  OAI22_X1 U184 ( .A1(DATA2[20]), .A2(n12), .B1(n3), .B2(n40), .ZN(N194) );
  INV_X1 U185 ( .A(DATA2[20]), .ZN(n40) );
  OAI22_X1 U186 ( .A1(DATA2[21]), .A2(n12), .B1(n3), .B2(n39), .ZN(N195) );
  INV_X1 U187 ( .A(DATA2[21]), .ZN(n39) );
  OAI22_X1 U188 ( .A1(DATA2[22]), .A2(n12), .B1(n3), .B2(n38), .ZN(N196) );
  INV_X1 U189 ( .A(DATA2[22]), .ZN(n38) );
  OAI22_X1 U190 ( .A1(DATA2[23]), .A2(n12), .B1(n3), .B2(n37), .ZN(N197) );
  INV_X1 U191 ( .A(DATA2[23]), .ZN(n37) );
  NAND2_X1 U192 ( .A1(n146), .A2(n133), .ZN(n152) );
  AND2_X1 U193 ( .A1(n127), .A2(n173), .ZN(n124) );
  NAND4_X1 U194 ( .A1(n122), .A2(n152), .A3(n126), .A4(n132), .ZN(n151) );
  NAND2_X1 U195 ( .A1(n153), .A2(n147), .ZN(n120) );
  NAND2_X1 U196 ( .A1(n168), .A2(n169), .ZN(n142) );
  NAND2_X1 U197 ( .A1(n146), .A2(n147), .ZN(n118) );
  NAND2_X1 U198 ( .A1(n147), .A2(n167), .ZN(n132) );
  NAND2_X1 U199 ( .A1(n153), .A2(n133), .ZN(n126) );
  INV_X1 U200 ( .A(n129), .ZN(n171) );
  NAND2_X1 U201 ( .A1(n119), .A2(n171), .ZN(n125) );
  NAND2_X1 U202 ( .A1(n153), .A2(n145), .ZN(n136) );
  INV_X1 U203 ( .A(n119), .ZN(n174) );
  NAND2_X1 U204 ( .A1(n146), .A2(n145), .ZN(n144) );
  INV_X1 U205 ( .A(n145), .ZN(n161) );
  NAND2_X1 U206 ( .A1(n129), .A2(n130), .ZN(n48) );
  NAND2_X1 U207 ( .A1(n167), .A2(n133), .ZN(n123) );
  INV_X1 U208 ( .A(n150), .ZN(n173) );
  NAND2_X1 U209 ( .A1(n110), .A2(n111), .ZN(N145) );
  NAND2_X1 U210 ( .A1(OUTPUT1[3]), .A2(n13), .ZN(n110) );
  AOI22_X1 U211 ( .A1(OUTPUT2[3]), .A2(n10), .B1(OUTPUT4[3]), .B2(n7), .ZN(
        n111) );
  NAND2_X1 U212 ( .A1(n112), .A2(n113), .ZN(N144) );
  NAND2_X1 U213 ( .A1(OUTPUT1[2]), .A2(n13), .ZN(n112) );
  AOI22_X1 U214 ( .A1(OUTPUT2[2]), .A2(n10), .B1(OUTPUT4[2]), .B2(n7), .ZN(
        n113) );
  NAND2_X1 U215 ( .A1(n114), .A2(n115), .ZN(N143) );
  NAND2_X1 U216 ( .A1(OUTPUT1[1]), .A2(n13), .ZN(n114) );
  AOI22_X1 U217 ( .A1(OUTPUT2[1]), .A2(n10), .B1(OUTPUT4[1]), .B2(n7), .ZN(
        n115) );
  NOR2_X1 U218 ( .A1(FUNC[5]), .A2(FUNC[4]), .ZN(n147) );
  OAI211_X1 U219 ( .C1(n126), .C2(n127), .A(n128), .B(n48), .ZN(N206) );
  OAI21_X1 U220 ( .B1(n131), .B2(n130), .A(n174), .ZN(n128) );
  NOR3_X1 U224 ( .A1(n169), .A2(FUNC[3]), .A3(n161), .ZN(n131) );
  NOR2_X1 U225 ( .A1(n166), .A2(FUNC[4]), .ZN(n145) );
  NOR2_X1 U226 ( .A1(n168), .A2(FUNC[2]), .ZN(n146) );
  NAND2_X1 U227 ( .A1(FUNC[0]), .A2(n172), .ZN(n127) );
  NAND2_X1 U228 ( .A1(FUNC[0]), .A2(FUNC[1]), .ZN(n119) );
  INV_X1 U229 ( .A(FUNC[2]), .ZN(n169) );
  INV_X1 U230 ( .A(FUNC[3]), .ZN(n168) );
  NOR2_X1 U231 ( .A1(FUNC[1]), .A2(FUNC[0]), .ZN(n150) );
  NOR2_X1 U232 ( .A1(n172), .A2(FUNC[0]), .ZN(n129) );
  INV_X1 U233 ( .A(FUNC[5]), .ZN(n166) );
  INV_X1 U234 ( .A(FUNC[1]), .ZN(n172) );
  AND2_X1 U235 ( .A1(FUNC[4]), .A2(n166), .ZN(n133) );
  INV_X1 U236 ( .A(DATA2[3]), .ZN(n27) );
  NAND2_X1 U237 ( .A1(n116), .A2(n117), .ZN(N142) );
  AOI22_X1 U238 ( .A1(\OUTPUT3[0] ), .A2(n55), .B1(OUTPUT1[0]), .B2(n15), .ZN(
        n116) );
  AOI22_X1 U239 ( .A1(OUTPUT2[0]), .A2(n10), .B1(OUTPUT4[0]), .B2(n7), .ZN(
        n117) );
  INV_X1 U240 ( .A(DATA2[0]), .ZN(n22) );
  INV_X1 U241 ( .A(DATA2[1]), .ZN(n23) );
  INV_X1 U242 ( .A(n25), .ZN(n24) );
  INV_X1 U243 ( .A(DATA2[2]), .ZN(n25) );
  INV_X1 U244 ( .A(DATA2[4]), .ZN(n28) );
endmodule


module zero_eval_NBIT32 ( \input , res );
  input [31:0] \input ;
  output res;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(\input [23]), .A2(\input [22]), .A3(\input [21]), .A4(
        \input [20]), .ZN(n6) );
  NOR4_X1 U2 ( .A1(\input [9]), .A2(\input [8]), .A3(\input [7]), .A4(
        \input [6]), .ZN(n10) );
  NOR4_X1 U3 ( .A1(\input [5]), .A2(\input [4]), .A3(\input [3]), .A4(
        \input [31]), .ZN(n9) );
  NOR4_X1 U4 ( .A1(\input [30]), .A2(\input [2]), .A3(\input [29]), .A4(
        \input [28]), .ZN(n8) );
  NOR4_X1 U5 ( .A1(\input [27]), .A2(\input [26]), .A3(\input [25]), .A4(
        \input [24]), .ZN(n7) );
  NAND4_X1 U6 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NOR4_X1 U7 ( .A1(\input [12]), .A2(\input [11]), .A3(\input [10]), .A4(
        \input [0]), .ZN(n3) );
  NOR4_X1 U8 ( .A1(\input [16]), .A2(\input [15]), .A3(\input [14]), .A4(
        \input [13]), .ZN(n4) );
  NOR4_X1 U9 ( .A1(\input [1]), .A2(\input [19]), .A3(\input [18]), .A4(
        \input [17]), .ZN(n5) );
  NOR2_X1 U10 ( .A1(n1), .A2(n2), .ZN(res) );
  NAND4_X1 U11 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
endmodule


module COND_BT_NBIT32 ( ZERO_BIT, OPCODE_0, branch_op, con_sign );
  input ZERO_BIT, OPCODE_0, branch_op;
  output con_sign;
  wire   n1;

  XOR2_X1 U3 ( .A(ZERO_BIT), .B(OPCODE_0), .Z(n1) );
  AND2_X1 U2 ( .A1(branch_op), .A2(n1), .ZN(con_sign) );
endmodule


module IV_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_160 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_160 UIV ( .A(S), .Y(SB) );
  ND2_480 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_479 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_478 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_159 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_159 UIV ( .A(S), .Y(SB) );
  ND2_477 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_476 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_475 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_158 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_158 UIV ( .A(S), .Y(SB) );
  ND2_474 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_473 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_472 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_157 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_157 UIV ( .A(S), .Y(SB) );
  ND2_471 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_470 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_469 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_156 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_156 UIV ( .A(S), .Y(SB) );
  ND2_468 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_467 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_466 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_155 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_155 UIV ( .A(S), .Y(SB) );
  ND2_465 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_464 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_463 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_154 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_154 UIV ( .A(S), .Y(SB) );
  ND2_462 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_461 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_460 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_153 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_153 UIV ( .A(S), .Y(SB) );
  ND2_459 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_458 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_457 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_152 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_152 UIV ( .A(S), .Y(SB) );
  ND2_456 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_455 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_454 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_151 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_151 UIV ( .A(S), .Y(SB) );
  ND2_453 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_452 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_451 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_150 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_150 UIV ( .A(S), .Y(SB) );
  ND2_450 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_449 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_448 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_149 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_149 UIV ( .A(S), .Y(SB) );
  ND2_447 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_446 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_445 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_148 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_148 UIV ( .A(S), .Y(SB) );
  ND2_444 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_443 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_442 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_147 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_147 UIV ( .A(S), .Y(SB) );
  ND2_441 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_440 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_439 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_146 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_146 UIV ( .A(S), .Y(SB) );
  ND2_438 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_437 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_436 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_145 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_145 UIV ( .A(S), .Y(SB) );
  ND2_435 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_434 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_433 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_144 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_144 UIV ( .A(S), .Y(SB) );
  ND2_432 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_431 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_430 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_143 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_143 UIV ( .A(S), .Y(SB) );
  ND2_429 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_428 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_427 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_142 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_142 UIV ( .A(S), .Y(SB) );
  ND2_426 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_425 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_424 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_141 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_141 UIV ( .A(S), .Y(SB) );
  ND2_423 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_422 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_421 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_140 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_140 UIV ( .A(S), .Y(SB) );
  ND2_420 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_419 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_418 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_139 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_139 UIV ( .A(S), .Y(SB) );
  ND2_417 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_416 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_415 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_138 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_138 UIV ( .A(S), .Y(SB) );
  ND2_414 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_413 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_412 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_137 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_137 UIV ( .A(S), .Y(SB) );
  ND2_411 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_410 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_409 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_136 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_136 UIV ( .A(S), .Y(SB) );
  ND2_408 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_407 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_406 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_135 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_135 UIV ( .A(S), .Y(SB) );
  ND2_405 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_404 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_403 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_134 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_134 UIV ( .A(S), .Y(SB) );
  ND2_402 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_401 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_400 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_133 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_133 UIV ( .A(S), .Y(SB) );
  ND2_399 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_398 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_397 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_132 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_132 UIV ( .A(S), .Y(SB) );
  ND2_396 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_395 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_394 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_131 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_131 UIV ( .A(S), .Y(SB) );
  ND2_393 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_392 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_391 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_130 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_130 UIV ( .A(S), .Y(SB) );
  ND2_390 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_389 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_388 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_129 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_129 UIV ( .A(S), .Y(SB) );
  ND2_387 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_386 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_385 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_160 gen1_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_159 gen1_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_158 gen1_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_157 gen1_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_156 gen1_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_155 gen1_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_154 gen1_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_153 gen1_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_152 gen1_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_151 gen1_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_150 gen1_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_149 gen1_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_148 gen1_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_147 gen1_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_146 gen1_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_145 gen1_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_144 gen1_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_143 gen1_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_142 gen1_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_141 gen1_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_140 gen1_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_139 gen1_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_138 gen1_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_137 gen1_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_136 gen1_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_135 gen1_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_134 gen1_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_133 gen1_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_132 gen1_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_131 gen1_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_130 gen1_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_129 gen1_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module FF_6 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n1, n2, n5, n6;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n1), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n2), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n2) );
  INV_X1 U6 ( .A(RESET), .ZN(n1) );
endmodule


module regFFD_NBIT32_5 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module FF_5 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n1, n2, n5, n6;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n1), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n2), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n2) );
  INV_X1 U6 ( .A(RESET), .ZN(n1) );
endmodule


module regFFD_NBIT32_4 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT5_2 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \Q_reg[4]  ( .D(n16), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n21) );
  DFFR_X1 \Q_reg[3]  ( .D(n17), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n22) );
  DFFR_X1 \Q_reg[2]  ( .D(n18), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n23) );
  DFFR_X1 \Q_reg[1]  ( .D(n19), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n24) );
  DFFR_X1 \Q_reg[0]  ( .D(n20), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n25) );
  OAI21_X1 U2 ( .B1(n25), .B2(ENABLE), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(ENABLE), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(ENABLE), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(ENABLE), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(ENABLE), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n26) );
endmodule


module FF_4 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n2, n4;

  SDFF_X1 Q_reg ( .D(RESET), .SI(1'b0), .SE(n4), .CK(CLK), .Q(Q) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n2), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n2) );
endmodule


module regFFD_NBIT6_1 ( CK, RESET, ENABLE, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET, ENABLE;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36;

  DFFR_X1 \Q_reg[5]  ( .D(n19), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n25) );
  DFFR_X1 \Q_reg[4]  ( .D(n20), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n26) );
  DFFR_X1 \Q_reg[3]  ( .D(n21), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n27) );
  DFFR_X1 \Q_reg[2]  ( .D(n22), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n28) );
  DFFR_X1 \Q_reg[1]  ( .D(n23), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n29) );
  DFFR_X1 \Q_reg[0]  ( .D(n24), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n30) );
  OAI21_X1 U2 ( .B1(n30), .B2(ENABLE), .A(n36), .ZN(n24) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n36) );
  OAI21_X1 U4 ( .B1(n29), .B2(ENABLE), .A(n35), .ZN(n23) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n35) );
  OAI21_X1 U6 ( .B1(n28), .B2(ENABLE), .A(n34), .ZN(n22) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n34) );
  OAI21_X1 U8 ( .B1(n27), .B2(ENABLE), .A(n33), .ZN(n21) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n33) );
  OAI21_X1 U10 ( .B1(n26), .B2(ENABLE), .A(n32), .ZN(n20) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n32) );
  OAI21_X1 U12 ( .B1(n25), .B2(ENABLE), .A(n31), .ZN(n19) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n31) );
endmodule


module IV_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_128 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_128 UIV ( .A(S), .Y(SB) );
  ND2_384 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_383 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_382 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_127 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_127 UIV ( .A(S), .Y(SB) );
  ND2_381 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_380 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_379 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_126 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_126 UIV ( .A(S), .Y(SB) );
  ND2_378 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_377 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_376 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_125 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_125 UIV ( .A(S), .Y(SB) );
  ND2_375 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_374 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_373 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_124 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_124 UIV ( .A(S), .Y(SB) );
  ND2_372 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_371 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_370 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_123 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_123 UIV ( .A(S), .Y(SB) );
  ND2_369 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_368 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_367 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_122 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_122 UIV ( .A(S), .Y(SB) );
  ND2_366 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_365 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_364 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_121 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_121 UIV ( .A(S), .Y(SB) );
  ND2_363 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_362 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_361 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_120 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_120 UIV ( .A(S), .Y(SB) );
  ND2_360 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_359 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_358 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_119 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_119 UIV ( .A(S), .Y(SB) );
  ND2_357 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_356 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_355 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_118 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_118 UIV ( .A(S), .Y(SB) );
  ND2_354 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_353 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_352 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_117 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_117 UIV ( .A(S), .Y(SB) );
  ND2_351 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_350 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_349 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_116 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_116 UIV ( .A(S), .Y(SB) );
  ND2_348 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_347 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_346 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_115 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_115 UIV ( .A(S), .Y(SB) );
  ND2_345 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_344 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_343 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_114 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_114 UIV ( .A(S), .Y(SB) );
  ND2_342 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_341 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_340 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_113 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_113 UIV ( .A(S), .Y(SB) );
  ND2_339 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_338 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_337 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_112 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_112 UIV ( .A(S), .Y(SB) );
  ND2_336 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_335 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_334 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_111 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_111 UIV ( .A(S), .Y(SB) );
  ND2_333 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_332 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_331 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_110 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_110 UIV ( .A(S), .Y(SB) );
  ND2_330 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_329 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_328 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_109 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_109 UIV ( .A(S), .Y(SB) );
  ND2_327 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_326 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_325 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_108 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_108 UIV ( .A(S), .Y(SB) );
  ND2_324 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_323 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_322 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_107 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_107 UIV ( .A(S), .Y(SB) );
  ND2_321 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_320 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_319 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_106 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_106 UIV ( .A(S), .Y(SB) );
  ND2_318 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_317 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_316 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_105 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_105 UIV ( .A(S), .Y(SB) );
  ND2_315 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_314 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_313 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_104 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_104 UIV ( .A(S), .Y(SB) );
  ND2_312 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_311 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_310 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_103 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_103 UIV ( .A(S), .Y(SB) );
  ND2_309 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_308 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_307 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_102 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_102 UIV ( .A(S), .Y(SB) );
  ND2_306 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_305 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_304 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_101 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_101 UIV ( .A(S), .Y(SB) );
  ND2_303 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_302 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_301 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_100 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_100 UIV ( .A(S), .Y(SB) );
  ND2_300 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_299 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_298 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_99 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_99 UIV ( .A(S), .Y(SB) );
  ND2_297 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_296 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_295 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_98 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_98 UIV ( .A(S), .Y(SB) );
  ND2_294 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_293 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_292 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_97 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_97 UIV ( .A(S), .Y(SB) );
  ND2_291 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_290 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_289 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_128 gen1_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_127 gen1_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_126 gen1_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_125 gen1_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_124 gen1_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_123 gen1_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_122 gen1_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_121 gen1_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_120 gen1_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_119 gen1_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_118 gen1_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_117 gen1_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_116 gen1_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_115 gen1_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_114 gen1_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_113 gen1_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_112 gen1_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_111 gen1_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_110 gen1_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_109 gen1_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_108 gen1_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_107 gen1_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_106 gen1_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_105 gen1_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_104 gen1_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_103 gen1_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_102 gen1_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_101 gen1_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_100 gen1_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_99 gen1_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_98 gen1_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_97 gen1_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module load_data ( data_in, signed_val, load_op, load_type, data_out );
  input [31:0] data_in;
  input [1:0] load_type;
  output [31:0] data_out;
  input signed_val, load_op;
  wire   N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n1, n2, n3, n31, n32;

  DLH_X1 \data_out_reg[31]  ( .G(load_op), .D(N67), .Q(data_out[31]) );
  DLH_X1 \data_out_reg[30]  ( .G(load_op), .D(N66), .Q(data_out[30]) );
  DLH_X1 \data_out_reg[29]  ( .G(load_op), .D(N65), .Q(data_out[29]) );
  DLH_X1 \data_out_reg[28]  ( .G(load_op), .D(N64), .Q(data_out[28]) );
  DLH_X1 \data_out_reg[27]  ( .G(load_op), .D(N63), .Q(data_out[27]) );
  DLH_X1 \data_out_reg[26]  ( .G(load_op), .D(N62), .Q(data_out[26]) );
  DLH_X1 \data_out_reg[25]  ( .G(load_op), .D(N61), .Q(data_out[25]) );
  DLH_X1 \data_out_reg[24]  ( .G(load_op), .D(N60), .Q(data_out[24]) );
  DLH_X1 \data_out_reg[23]  ( .G(load_op), .D(N59), .Q(data_out[23]) );
  DLH_X1 \data_out_reg[22]  ( .G(load_op), .D(N58), .Q(data_out[22]) );
  DLH_X1 \data_out_reg[21]  ( .G(load_op), .D(N57), .Q(data_out[21]) );
  DLH_X1 \data_out_reg[20]  ( .G(load_op), .D(N56), .Q(data_out[20]) );
  DLH_X1 \data_out_reg[19]  ( .G(load_op), .D(N55), .Q(data_out[19]) );
  DLH_X1 \data_out_reg[18]  ( .G(load_op), .D(N54), .Q(data_out[18]) );
  DLH_X1 \data_out_reg[17]  ( .G(load_op), .D(N53), .Q(data_out[17]) );
  DLH_X1 \data_out_reg[16]  ( .G(load_op), .D(N52), .Q(data_out[16]) );
  DLH_X1 \data_out_reg[15]  ( .G(load_op), .D(N51), .Q(data_out[15]) );
  DLH_X1 \data_out_reg[14]  ( .G(load_op), .D(N50), .Q(data_out[14]) );
  DLH_X1 \data_out_reg[13]  ( .G(load_op), .D(N49), .Q(data_out[13]) );
  DLH_X1 \data_out_reg[12]  ( .G(load_op), .D(N48), .Q(data_out[12]) );
  DLH_X1 \data_out_reg[11]  ( .G(load_op), .D(N47), .Q(data_out[11]) );
  DLH_X1 \data_out_reg[10]  ( .G(load_op), .D(N46), .Q(data_out[10]) );
  DLH_X1 \data_out_reg[9]  ( .G(load_op), .D(N45), .Q(data_out[9]) );
  DLH_X1 \data_out_reg[8]  ( .G(load_op), .D(N44), .Q(data_out[8]) );
  DLH_X1 \data_out_reg[7]  ( .G(load_op), .D(N43), .Q(data_out[7]) );
  DLH_X1 \data_out_reg[6]  ( .G(load_op), .D(N42), .Q(data_out[6]) );
  DLH_X1 \data_out_reg[5]  ( .G(load_op), .D(N41), .Q(data_out[5]) );
  DLH_X1 \data_out_reg[4]  ( .G(load_op), .D(N40), .Q(data_out[4]) );
  DLH_X1 \data_out_reg[3]  ( .G(load_op), .D(N39), .Q(data_out[3]) );
  DLH_X1 \data_out_reg[2]  ( .G(load_op), .D(N38), .Q(data_out[2]) );
  DLH_X1 \data_out_reg[1]  ( .G(load_op), .D(N37), .Q(data_out[1]) );
  DLH_X1 \data_out_reg[0]  ( .G(load_op), .D(N36), .Q(data_out[0]) );
  INV_X1 U2 ( .A(n4), .ZN(n3) );
  BUF_X1 U3 ( .A(n5), .Z(n1) );
  BUF_X1 U4 ( .A(n5), .Z(n2) );
  OAI21_X1 U5 ( .B1(n4), .B2(n32), .A(n1), .ZN(N67) );
  NAND2_X1 U6 ( .A1(load_type[1]), .A2(load_type[0]), .ZN(n4) );
  NAND2_X1 U7 ( .A1(n31), .A2(n29), .ZN(n30) );
  INV_X1 U8 ( .A(load_type[0]), .ZN(n31) );
  OR2_X1 U9 ( .A1(load_type[1]), .A2(load_type[0]), .ZN(n29) );
  OR3_X1 U10 ( .A1(signed_val), .A2(n32), .A3(n29), .ZN(n5) );
  INV_X1 U11 ( .A(data_in[31]), .ZN(n32) );
  NAND2_X1 U12 ( .A1(n2), .A2(n28), .ZN(N44) );
  NAND2_X1 U13 ( .A1(data_in[8]), .A2(load_type[0]), .ZN(n28) );
  NAND2_X1 U14 ( .A1(n2), .A2(n27), .ZN(N45) );
  NAND2_X1 U15 ( .A1(data_in[9]), .A2(load_type[0]), .ZN(n27) );
  NAND2_X1 U16 ( .A1(n2), .A2(n26), .ZN(N46) );
  NAND2_X1 U17 ( .A1(data_in[10]), .A2(load_type[0]), .ZN(n26) );
  NAND2_X1 U18 ( .A1(n2), .A2(n25), .ZN(N47) );
  NAND2_X1 U19 ( .A1(data_in[11]), .A2(load_type[0]), .ZN(n25) );
  NAND2_X1 U20 ( .A1(n2), .A2(n24), .ZN(N48) );
  NAND2_X1 U21 ( .A1(data_in[12]), .A2(load_type[0]), .ZN(n24) );
  NAND2_X1 U22 ( .A1(n2), .A2(n23), .ZN(N49) );
  NAND2_X1 U23 ( .A1(data_in[13]), .A2(load_type[0]), .ZN(n23) );
  NAND2_X1 U24 ( .A1(n2), .A2(n22), .ZN(N50) );
  NAND2_X1 U25 ( .A1(data_in[14]), .A2(load_type[0]), .ZN(n22) );
  NAND2_X1 U26 ( .A1(n2), .A2(n21), .ZN(N51) );
  NAND2_X1 U27 ( .A1(data_in[15]), .A2(load_type[0]), .ZN(n21) );
  NAND2_X1 U28 ( .A1(n1), .A2(n16), .ZN(N56) );
  NAND2_X1 U29 ( .A1(data_in[20]), .A2(n3), .ZN(n16) );
  NAND2_X1 U30 ( .A1(n1), .A2(n15), .ZN(N57) );
  NAND2_X1 U31 ( .A1(data_in[21]), .A2(n3), .ZN(n15) );
  NAND2_X1 U32 ( .A1(n1), .A2(n14), .ZN(N58) );
  NAND2_X1 U33 ( .A1(data_in[22]), .A2(n3), .ZN(n14) );
  NAND2_X1 U34 ( .A1(n1), .A2(n13), .ZN(N59) );
  NAND2_X1 U35 ( .A1(data_in[23]), .A2(n3), .ZN(n13) );
  NAND2_X1 U36 ( .A1(n1), .A2(n12), .ZN(N60) );
  NAND2_X1 U37 ( .A1(data_in[24]), .A2(n3), .ZN(n12) );
  NAND2_X1 U38 ( .A1(n1), .A2(n11), .ZN(N61) );
  NAND2_X1 U39 ( .A1(data_in[25]), .A2(n3), .ZN(n11) );
  NAND2_X1 U40 ( .A1(n1), .A2(n10), .ZN(N62) );
  NAND2_X1 U41 ( .A1(data_in[26]), .A2(n3), .ZN(n10) );
  NAND2_X1 U42 ( .A1(n1), .A2(n9), .ZN(N63) );
  NAND2_X1 U43 ( .A1(data_in[27]), .A2(n3), .ZN(n9) );
  NAND2_X1 U44 ( .A1(n1), .A2(n8), .ZN(N64) );
  NAND2_X1 U45 ( .A1(data_in[28]), .A2(n3), .ZN(n8) );
  NAND2_X1 U46 ( .A1(n1), .A2(n7), .ZN(N65) );
  NAND2_X1 U47 ( .A1(data_in[29]), .A2(n3), .ZN(n7) );
  NAND2_X1 U48 ( .A1(n1), .A2(n6), .ZN(N66) );
  NAND2_X1 U49 ( .A1(data_in[30]), .A2(n3), .ZN(n6) );
  NAND2_X1 U50 ( .A1(n2), .A2(n20), .ZN(N52) );
  NAND2_X1 U51 ( .A1(data_in[16]), .A2(n3), .ZN(n20) );
  NAND2_X1 U52 ( .A1(n2), .A2(n19), .ZN(N53) );
  NAND2_X1 U53 ( .A1(data_in[17]), .A2(n3), .ZN(n19) );
  NAND2_X1 U54 ( .A1(n2), .A2(n18), .ZN(N54) );
  NAND2_X1 U55 ( .A1(data_in[18]), .A2(n3), .ZN(n18) );
  NAND2_X1 U56 ( .A1(n2), .A2(n17), .ZN(N55) );
  NAND2_X1 U57 ( .A1(data_in[19]), .A2(n3), .ZN(n17) );
  AND2_X1 U58 ( .A1(data_in[0]), .A2(n30), .ZN(N36) );
  AND2_X1 U59 ( .A1(data_in[1]), .A2(n30), .ZN(N37) );
  AND2_X1 U60 ( .A1(data_in[2]), .A2(n30), .ZN(N38) );
  AND2_X1 U61 ( .A1(data_in[3]), .A2(n30), .ZN(N39) );
  AND2_X1 U62 ( .A1(data_in[4]), .A2(n30), .ZN(N40) );
  AND2_X1 U63 ( .A1(data_in[5]), .A2(n30), .ZN(N41) );
  AND2_X1 U64 ( .A1(data_in[6]), .A2(n30), .ZN(N42) );
  AND2_X1 U65 ( .A1(data_in[7]), .A2(n30), .ZN(N43) );
endmodule


module regFFD_NBIT32_3 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT32_2 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module regFFD_NBIT5_1 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30;

  DFFR_X1 \Q_reg[4]  ( .D(n16), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n21) );
  DFFR_X1 \Q_reg[3]  ( .D(n17), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n22) );
  DFFR_X1 \Q_reg[2]  ( .D(n18), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n23) );
  DFFR_X1 \Q_reg[1]  ( .D(n19), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n24) );
  DFFR_X1 \Q_reg[0]  ( .D(n20), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n25) );
  OAI21_X1 U2 ( .B1(n25), .B2(ENABLE), .A(n30), .ZN(n20) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n24), .B2(ENABLE), .A(n29), .ZN(n19) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n23), .B2(ENABLE), .A(n28), .ZN(n18) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(ENABLE), .A(n27), .ZN(n17) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n21), .B2(ENABLE), .A(n26), .ZN(n16) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n26) );
endmodule


module FF_3 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n1, n2, n5, n6;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n1), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n2), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n2) );
  INV_X1 U6 ( .A(RESET), .ZN(n1) );
endmodule


module FF_2 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n1, n2, n5, n6;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n1), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n2), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n2) );
  INV_X1 U6 ( .A(RESET), .ZN(n1) );
endmodule


module FF_1 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n1, n2, n5, n6;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n1), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(Q), .B2(n2), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n2) );
  INV_X1 U6 ( .A(RESET), .ZN(n1) );
endmodule


module regFFD_NBIT32_1 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195;

  DFFR_X1 \Q_reg[31]  ( .D(n100), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n132) );
  DFFR_X1 \Q_reg[30]  ( .D(n101), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n133) );
  DFFR_X1 \Q_reg[29]  ( .D(n102), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n134) );
  DFFR_X1 \Q_reg[28]  ( .D(n103), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n135) );
  DFFR_X1 \Q_reg[27]  ( .D(n104), .CK(CK), .RN(n99), .Q(Q[27]), .QN(n136) );
  DFFR_X1 \Q_reg[26]  ( .D(n105), .CK(CK), .RN(n99), .Q(Q[26]), .QN(n137) );
  DFFR_X1 \Q_reg[25]  ( .D(n106), .CK(CK), .RN(n99), .Q(Q[25]), .QN(n138) );
  DFFR_X1 \Q_reg[24]  ( .D(n107), .CK(CK), .RN(n99), .Q(Q[24]), .QN(n139) );
  DFFR_X1 \Q_reg[23]  ( .D(n108), .CK(CK), .RN(n98), .Q(Q[23]), .QN(n140) );
  DFFR_X1 \Q_reg[22]  ( .D(n109), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n141) );
  DFFR_X1 \Q_reg[21]  ( .D(n110), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n142) );
  DFFR_X1 \Q_reg[20]  ( .D(n111), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n143) );
  DFFR_X1 \Q_reg[19]  ( .D(n112), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n144) );
  DFFR_X1 \Q_reg[18]  ( .D(n113), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n145) );
  DFFR_X1 \Q_reg[17]  ( .D(n114), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n146) );
  DFFR_X1 \Q_reg[16]  ( .D(n115), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n147) );
  DFFR_X1 \Q_reg[15]  ( .D(n116), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n148) );
  DFFR_X1 \Q_reg[14]  ( .D(n117), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n149) );
  DFFR_X1 \Q_reg[13]  ( .D(n118), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n150) );
  DFFR_X1 \Q_reg[12]  ( .D(n119), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n151) );
  DFFR_X1 \Q_reg[11]  ( .D(n120), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n152) );
  DFFR_X1 \Q_reg[10]  ( .D(n121), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n153) );
  DFFR_X1 \Q_reg[9]  ( .D(n122), .CK(CK), .RN(n97), .Q(Q[9]), .QN(n154) );
  DFFR_X1 \Q_reg[8]  ( .D(n123), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n155) );
  DFFR_X1 \Q_reg[7]  ( .D(n124), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n156) );
  DFFR_X1 \Q_reg[6]  ( .D(n125), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n157) );
  DFFR_X1 \Q_reg[5]  ( .D(n126), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n158) );
  DFFR_X1 \Q_reg[4]  ( .D(n127), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n159) );
  DFFR_X1 \Q_reg[3]  ( .D(n128), .CK(CK), .RN(n97), .Q(Q[3]), .QN(n160) );
  DFFR_X1 \Q_reg[2]  ( .D(n129), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n161) );
  DFFR_X1 \Q_reg[1]  ( .D(n130), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n162) );
  DFFR_X1 \Q_reg[0]  ( .D(n131), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n163) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n163), .B2(ENABLE), .A(n195), .ZN(n131) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[0]), .ZN(n195) );
  OAI21_X1 U7 ( .B1(n162), .B2(ENABLE), .A(n194), .ZN(n130) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n194) );
  OAI21_X1 U9 ( .B1(n161), .B2(ENABLE), .A(n193), .ZN(n129) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n193) );
  OAI21_X1 U11 ( .B1(n160), .B2(ENABLE), .A(n192), .ZN(n128) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n192) );
  OAI21_X1 U13 ( .B1(n159), .B2(ENABLE), .A(n191), .ZN(n127) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n191) );
  OAI21_X1 U15 ( .B1(n158), .B2(ENABLE), .A(n190), .ZN(n126) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n190) );
  OAI21_X1 U17 ( .B1(n157), .B2(ENABLE), .A(n189), .ZN(n125) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n189) );
  OAI21_X1 U19 ( .B1(n156), .B2(ENABLE), .A(n188), .ZN(n124) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n188) );
  OAI21_X1 U21 ( .B1(n155), .B2(ENABLE), .A(n187), .ZN(n123) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n187) );
  OAI21_X1 U23 ( .B1(n154), .B2(ENABLE), .A(n186), .ZN(n122) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n186) );
  OAI21_X1 U25 ( .B1(n153), .B2(ENABLE), .A(n185), .ZN(n121) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n185) );
  OAI21_X1 U27 ( .B1(n152), .B2(ENABLE), .A(n184), .ZN(n120) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n184) );
  OAI21_X1 U29 ( .B1(n151), .B2(ENABLE), .A(n183), .ZN(n119) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n183) );
  OAI21_X1 U31 ( .B1(n150), .B2(ENABLE), .A(n182), .ZN(n118) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n182) );
  OAI21_X1 U33 ( .B1(n149), .B2(ENABLE), .A(n181), .ZN(n117) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n181) );
  OAI21_X1 U35 ( .B1(n148), .B2(ENABLE), .A(n180), .ZN(n116) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n180) );
  OAI21_X1 U37 ( .B1(n147), .B2(ENABLE), .A(n179), .ZN(n115) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n179) );
  OAI21_X1 U39 ( .B1(n146), .B2(ENABLE), .A(n178), .ZN(n114) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n178) );
  OAI21_X1 U41 ( .B1(n145), .B2(ENABLE), .A(n177), .ZN(n113) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n177) );
  OAI21_X1 U43 ( .B1(n144), .B2(ENABLE), .A(n176), .ZN(n112) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n176) );
  OAI21_X1 U45 ( .B1(n143), .B2(ENABLE), .A(n175), .ZN(n111) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n175) );
  OAI21_X1 U47 ( .B1(n142), .B2(ENABLE), .A(n174), .ZN(n110) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n174) );
  OAI21_X1 U49 ( .B1(n141), .B2(ENABLE), .A(n173), .ZN(n109) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n173) );
  OAI21_X1 U51 ( .B1(n140), .B2(ENABLE), .A(n172), .ZN(n108) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(ENABLE), .ZN(n172) );
  OAI21_X1 U53 ( .B1(n139), .B2(ENABLE), .A(n171), .ZN(n107) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n171) );
  OAI21_X1 U55 ( .B1(n138), .B2(ENABLE), .A(n170), .ZN(n106) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n170) );
  OAI21_X1 U57 ( .B1(n137), .B2(ENABLE), .A(n169), .ZN(n105) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n169) );
  OAI21_X1 U59 ( .B1(n136), .B2(ENABLE), .A(n168), .ZN(n104) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n168) );
  OAI21_X1 U61 ( .B1(n135), .B2(ENABLE), .A(n167), .ZN(n103) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n167) );
  OAI21_X1 U63 ( .B1(n134), .B2(ENABLE), .A(n166), .ZN(n102) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n166) );
  OAI21_X1 U65 ( .B1(n133), .B2(ENABLE), .A(n165), .ZN(n101) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n132), .B2(ENABLE), .A(n164), .ZN(n100) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n164) );
endmodule


module IV_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_96 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_96 UIV ( .A(S), .Y(SB) );
  ND2_288 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_287 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_286 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_95 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_95 UIV ( .A(S), .Y(SB) );
  ND2_285 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_284 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_283 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_94 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_94 UIV ( .A(S), .Y(SB) );
  ND2_282 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_281 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_280 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_93 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_93 UIV ( .A(S), .Y(SB) );
  ND2_279 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_278 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_277 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_92 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_92 UIV ( .A(S), .Y(SB) );
  ND2_276 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_275 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_274 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_91 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_91 UIV ( .A(S), .Y(SB) );
  ND2_273 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_272 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_271 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_90 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_90 UIV ( .A(S), .Y(SB) );
  ND2_270 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_269 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_268 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_89 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_89 UIV ( .A(S), .Y(SB) );
  ND2_267 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_266 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_265 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_88 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_88 UIV ( .A(S), .Y(SB) );
  ND2_264 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_263 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_262 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_87 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_87 UIV ( .A(S), .Y(SB) );
  ND2_261 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_260 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_259 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_86 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_86 UIV ( .A(S), .Y(SB) );
  ND2_258 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_257 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_256 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_85 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_85 UIV ( .A(S), .Y(SB) );
  ND2_255 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_254 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_253 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_84 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_84 UIV ( .A(S), .Y(SB) );
  ND2_252 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_251 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_250 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_83 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_83 UIV ( .A(S), .Y(SB) );
  ND2_249 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_248 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_247 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_82 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_82 UIV ( .A(S), .Y(SB) );
  ND2_246 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_245 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_244 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_81 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_81 UIV ( .A(S), .Y(SB) );
  ND2_243 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_242 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_241 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_80 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_80 UIV ( .A(S), .Y(SB) );
  ND2_240 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_239 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_238 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_79 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_79 UIV ( .A(S), .Y(SB) );
  ND2_237 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_236 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_235 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_78 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_78 UIV ( .A(S), .Y(SB) );
  ND2_234 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_233 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_232 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_77 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_77 UIV ( .A(S), .Y(SB) );
  ND2_231 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_230 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_229 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_76 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_76 UIV ( .A(S), .Y(SB) );
  ND2_228 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_227 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_226 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_75 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_75 UIV ( .A(S), .Y(SB) );
  ND2_225 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_224 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_223 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_74 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_74 UIV ( .A(S), .Y(SB) );
  ND2_222 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_221 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_220 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_73 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_73 UIV ( .A(S), .Y(SB) );
  ND2_219 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_218 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_217 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_72 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_72 UIV ( .A(S), .Y(SB) );
  ND2_216 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_215 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_214 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_71 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_71 UIV ( .A(S), .Y(SB) );
  ND2_213 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_212 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_211 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_70 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_70 UIV ( .A(S), .Y(SB) );
  ND2_210 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_209 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_208 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_69 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_69 UIV ( .A(S), .Y(SB) );
  ND2_207 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_206 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_205 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_68 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_68 UIV ( .A(S), .Y(SB) );
  ND2_204 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_203 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_202 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_67 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_67 UIV ( .A(S), .Y(SB) );
  ND2_201 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_200 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_199 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_66 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_66 UIV ( .A(S), .Y(SB) );
  ND2_198 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_197 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_196 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_65 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_65 UIV ( .A(S), .Y(SB) );
  ND2_195 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_194 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_193 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_96 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_95 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_94 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_93 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_92 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_91 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_90 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_89 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_88 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_87 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_86 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_85 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_84 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_83 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_82 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_81 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_80 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_79 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_78 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_77 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_76 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_75 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_74 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_73 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_72 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_71 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_70 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_69 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_68 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_67 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_66 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_65 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_64 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_64 UIV ( .A(S), .Y(SB) );
  ND2_192 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_191 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_190 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_63 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_63 UIV ( .A(S), .Y(SB) );
  ND2_189 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_188 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_187 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_62 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_62 UIV ( .A(S), .Y(SB) );
  ND2_186 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_185 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_184 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_61 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_61 UIV ( .A(S), .Y(SB) );
  ND2_183 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_182 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_181 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_60 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_60 UIV ( .A(S), .Y(SB) );
  ND2_180 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_179 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_178 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_59 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_59 UIV ( .A(S), .Y(SB) );
  ND2_177 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_176 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_175 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_58 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_58 UIV ( .A(S), .Y(SB) );
  ND2_174 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_173 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_172 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_57 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_57 UIV ( .A(S), .Y(SB) );
  ND2_171 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_170 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_169 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_56 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_56 UIV ( .A(S), .Y(SB) );
  ND2_168 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_167 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_166 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_55 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_55 UIV ( .A(S), .Y(SB) );
  ND2_165 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_164 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_163 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_54 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_54 UIV ( .A(S), .Y(SB) );
  ND2_162 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_161 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_160 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_53 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_53 UIV ( .A(S), .Y(SB) );
  ND2_159 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_158 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_157 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_52 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_52 UIV ( .A(S), .Y(SB) );
  ND2_156 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_155 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_154 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_51 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_51 UIV ( .A(S), .Y(SB) );
  ND2_153 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_152 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_151 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_50 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_50 UIV ( .A(S), .Y(SB) );
  ND2_150 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_149 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_148 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_49 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_49 UIV ( .A(S), .Y(SB) );
  ND2_147 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_146 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_145 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_48 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_48 UIV ( .A(S), .Y(SB) );
  ND2_144 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_143 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_142 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_47 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_47 UIV ( .A(S), .Y(SB) );
  ND2_141 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_140 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_139 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_46 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_46 UIV ( .A(S), .Y(SB) );
  ND2_138 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_137 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_136 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_45 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_45 UIV ( .A(S), .Y(SB) );
  ND2_135 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_134 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_133 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_44 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_44 UIV ( .A(S), .Y(SB) );
  ND2_132 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_131 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_130 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_43 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_43 UIV ( .A(S), .Y(SB) );
  ND2_129 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_128 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_127 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_42 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_42 UIV ( .A(S), .Y(SB) );
  ND2_126 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_125 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_124 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_41 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_41 UIV ( .A(S), .Y(SB) );
  ND2_123 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_122 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_121 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_40 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_40 UIV ( .A(S), .Y(SB) );
  ND2_120 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_119 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_118 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_39 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_39 UIV ( .A(S), .Y(SB) );
  ND2_117 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_116 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_115 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_38 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_38 UIV ( .A(S), .Y(SB) );
  ND2_114 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_113 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_112 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_37 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_37 UIV ( .A(S), .Y(SB) );
  ND2_111 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_110 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_109 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_36 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_36 UIV ( .A(S), .Y(SB) );
  ND2_108 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_107 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_106 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_35 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_35 UIV ( .A(S), .Y(SB) );
  ND2_105 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_104 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_103 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_34 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_34 UIV ( .A(S), .Y(SB) );
  ND2_102 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_101 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_100 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_33 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_33 UIV ( .A(S), .Y(SB) );
  ND2_99 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_98 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_97 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_64 gen1_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_63 gen1_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_62 gen1_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_61 gen1_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_60 gen1_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_59 gen1_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_58 gen1_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_57 gen1_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_56 gen1_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_55 gen1_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_54 gen1_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_53 gen1_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_52 gen1_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_51 gen1_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_50 gen1_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_49 gen1_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_48 gen1_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_47 gen1_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_46 gen1_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_45 gen1_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_44 gen1_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_43 gen1_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_42 gen1_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_41 gen1_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_40 gen1_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_39 gen1_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_38 gen1_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_37 gen1_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_36 gen1_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_35 gen1_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_34 gen1_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_33 gen1_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[31]), .B(A[31]), .Z(SUM[31]) );
endmodule


module DATAPTH_NBIT32_REG_BIT5 ( CLK, RST, PC, IR, PC_OUT, NPC_LATCH_EN, 
        ir_LATCH_EN, signed_op, trap_cs, ret_cs, RF1, RF2, WF1, 
        regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond, sb_op, RM, 
        WM, EN3, S3, .instruction_alu({\instruction_alu[5] , 
        \instruction_alu[4] , \instruction_alu[3] , \instruction_alu[2] , 
        \instruction_alu[1] , \instruction_alu[0] }), DATA_MEM_ADDR, 
        DATA_MEM_IN, DATA_MEM_OUT, DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM
 );
  input [31:0] PC;
  input [31:0] IR;
  output [31:0] PC_OUT;
  output [31:0] DATA_MEM_ADDR;
  output [31:0] DATA_MEM_IN;
  input [31:0] DATA_MEM_OUT;
  input CLK, RST, NPC_LATCH_EN, ir_LATCH_EN, signed_op, trap_cs, ret_cs, RF1,
         RF2, WF1, regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond,
         sb_op, RM, WM, EN3, S3, \instruction_alu[5] , \instruction_alu[4] ,
         \instruction_alu[3] , \instruction_alu[2] , \instruction_alu[1] ,
         \instruction_alu[0] ;
  output DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM;
  wire   RM, WM, sel_npc, wr_signal_wb, signed_op_ex, wr_signal_exe, is_zero,
         cond, signed_op_mem, cond_mem, wr_signal_mem, sel_saved_reg, N13,
         wr_signal_mem1, sel_saved_reg_wb, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n57, n58, n59,
         n60, n61;
  wire   [5:0] instruction_alu;
  wire   [31:0] PC_fetch0;
  wire   [31:0] NPC;
  wire   [31:0] NPC_fetch1;
  wire   [31:0] PC_fetch1;
  wire   [31:0] PC_OUT_i;
  wire   [31:0] NPC_fetch;
  wire   [31:0] PC_fetch;
  wire   [31:0] ir_fetch;
  wire   [31:0] NPC_Dec;
  wire   [31:0] IR_Dec;
  wire   [4:0] RS1;
  wire   [4:0] RS2;
  wire   [4:0] RD;
  wire   [31:0] Imm;
  wire   [4:0] RD_wb;
  wire   [31:0] OUT_wb;
  wire   [31:0] regA;
  wire   [31:0] regB;
  wire   [31:0] NPC_ex;
  wire   [31:0] regA_ex;
  wire   [31:0] regB_ex;
  wire   [31:0] Imm_ex;
  wire   [4:0] RD_ex;
  wire   [5:0] IR_26_ex;
  wire   [31:0] LHI_ex;
  wire   [31:0] input1_ALU;
  wire   [31:0] input2_ALU;
  wire   [31:0] ALU_out;
  wire   [31:0] ALU_ex;
  wire   [31:0] NPC_mem;
  wire   [31:0] regB_mem;
  wire   [4:0] RD_mem;
  wire   [5:0] IR_26_mem;
  wire   [31:0] LMD_out;
  wire   [31:0] ALU_wb;
  wire   [31:0] LMD_wb;
  wire   [31:0] NPC_wb;
  wire   [31:0] OUT_data;
  assign DATA_MEM_RM = RM;
  assign DATA_MEM_WM = WM;

  DLH_X1 \DATA_MEM_ADDR_reg[31]  ( .G(n5), .D(ALU_ex[31]), .Q(
        DATA_MEM_ADDR[31]) );
  DLH_X1 \DATA_MEM_ADDR_reg[30]  ( .G(n5), .D(ALU_ex[30]), .Q(
        DATA_MEM_ADDR[30]) );
  DLH_X1 \DATA_MEM_ADDR_reg[29]  ( .G(n5), .D(ALU_ex[29]), .Q(
        DATA_MEM_ADDR[29]) );
  DLH_X1 \DATA_MEM_ADDR_reg[28]  ( .G(n5), .D(ALU_ex[28]), .Q(
        DATA_MEM_ADDR[28]) );
  DLH_X1 \DATA_MEM_ADDR_reg[27]  ( .G(n5), .D(ALU_ex[27]), .Q(
        DATA_MEM_ADDR[27]) );
  DLH_X1 \DATA_MEM_ADDR_reg[26]  ( .G(n5), .D(ALU_ex[26]), .Q(
        DATA_MEM_ADDR[26]) );
  DLH_X1 \DATA_MEM_ADDR_reg[25]  ( .G(n5), .D(ALU_ex[25]), .Q(
        DATA_MEM_ADDR[25]) );
  DLH_X1 \DATA_MEM_ADDR_reg[24]  ( .G(n5), .D(ALU_ex[24]), .Q(
        DATA_MEM_ADDR[24]) );
  DLH_X1 \DATA_MEM_ADDR_reg[23]  ( .G(n5), .D(ALU_ex[23]), .Q(
        DATA_MEM_ADDR[23]) );
  DLH_X1 \DATA_MEM_ADDR_reg[22]  ( .G(n5), .D(ALU_ex[22]), .Q(
        DATA_MEM_ADDR[22]) );
  DLH_X1 \DATA_MEM_ADDR_reg[21]  ( .G(n5), .D(ALU_ex[21]), .Q(
        DATA_MEM_ADDR[21]) );
  DLH_X1 \DATA_MEM_ADDR_reg[20]  ( .G(n6), .D(ALU_ex[20]), .Q(
        DATA_MEM_ADDR[20]) );
  DLH_X1 \DATA_MEM_ADDR_reg[19]  ( .G(n6), .D(ALU_ex[19]), .Q(
        DATA_MEM_ADDR[19]) );
  DLH_X1 \DATA_MEM_ADDR_reg[18]  ( .G(n6), .D(ALU_ex[18]), .Q(
        DATA_MEM_ADDR[18]) );
  DLH_X1 \DATA_MEM_ADDR_reg[17]  ( .G(n6), .D(ALU_ex[17]), .Q(
        DATA_MEM_ADDR[17]) );
  DLH_X1 \DATA_MEM_ADDR_reg[16]  ( .G(n6), .D(ALU_ex[16]), .Q(
        DATA_MEM_ADDR[16]) );
  DLH_X1 \DATA_MEM_ADDR_reg[15]  ( .G(n6), .D(ALU_ex[15]), .Q(
        DATA_MEM_ADDR[15]) );
  DLH_X1 \DATA_MEM_ADDR_reg[14]  ( .G(n6), .D(ALU_ex[14]), .Q(
        DATA_MEM_ADDR[14]) );
  DLH_X1 \DATA_MEM_ADDR_reg[13]  ( .G(n6), .D(ALU_ex[13]), .Q(
        DATA_MEM_ADDR[13]) );
  DLH_X1 \DATA_MEM_ADDR_reg[12]  ( .G(n6), .D(ALU_ex[12]), .Q(
        DATA_MEM_ADDR[12]) );
  DLH_X1 \DATA_MEM_ADDR_reg[11]  ( .G(n6), .D(ALU_ex[11]), .Q(
        DATA_MEM_ADDR[11]) );
  DLH_X1 \DATA_MEM_ADDR_reg[10]  ( .G(n6), .D(ALU_ex[10]), .Q(
        DATA_MEM_ADDR[10]) );
  DLH_X1 \DATA_MEM_ADDR_reg[9]  ( .G(n7), .D(ALU_ex[9]), .Q(DATA_MEM_ADDR[9])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[8]  ( .G(n7), .D(ALU_ex[8]), .Q(DATA_MEM_ADDR[8])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[7]  ( .G(n7), .D(ALU_ex[7]), .Q(DATA_MEM_ADDR[7])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[6]  ( .G(n7), .D(ALU_ex[6]), .Q(DATA_MEM_ADDR[6])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[5]  ( .G(n7), .D(ALU_ex[5]), .Q(DATA_MEM_ADDR[5])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[4]  ( .G(n7), .D(ALU_ex[4]), .Q(DATA_MEM_ADDR[4])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[3]  ( .G(n7), .D(ALU_ex[3]), .Q(DATA_MEM_ADDR[3])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[2]  ( .G(n7), .D(ALU_ex[2]), .Q(DATA_MEM_ADDR[2])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[1]  ( .G(n7), .D(ALU_ex[1]), .Q(DATA_MEM_ADDR[1])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[0]  ( .G(n7), .D(ALU_ex[0]), .Q(DATA_MEM_ADDR[0])
         );
  OAI33_X1 U80 ( .A1(n15), .A2(IR_Dec[31]), .A3(n2), .B1(n24), .B2(n13), .B3(
        n25), .ZN(n23) );
  XOR2_X1 U81 ( .A(IR_Dec[27]), .B(IR_Dec[26]), .Z(n25) );
  NAND3_X1 U82 ( .A1(n16), .A2(n14), .A3(n2), .ZN(n24) );
  NAND3_X1 U83 ( .A1(instruction_alu[2]), .A2(instruction_alu[1]), .A3(
        instruction_alu[4]), .ZN(n52) );
  regFFD_NBIT32_0 pipeline_PCING ( .CK(CLK), .RESET(n9), .ENABLE(1'b1), .D(PC), 
        .Q(PC_fetch0) );
  regFFD_NBIT32_18 pipeline_fetch1_NPC ( .CK(CLK), .RESET(n9), .ENABLE(
        NPC_LATCH_EN), .D(NPC), .Q(NPC_fetch1) );
  regFFD_NBIT32_17 pipeline_fetch1_PC ( .CK(CLK), .RESET(n9), .ENABLE(
        ir_LATCH_EN), .D(PC_fetch0), .Q(PC_fetch1) );
  MUX21_GENERIC_NBIT32_0 MUX_PC1 ( .A(PC_OUT_i), .B(NPC_fetch1), .SEL(sel_npc), 
        .Y(PC_OUT) );
  regFFD_NBIT32_16 pipeline_fetch_NPC ( .CK(CLK), .RESET(n9), .ENABLE(
        NPC_LATCH_EN), .D(NPC_fetch1), .Q(NPC_fetch) );
  regFFD_NBIT32_15 pipeline_fetch_PC ( .CK(CLK), .RESET(n9), .ENABLE(
        ir_LATCH_EN), .D(PC_fetch1), .Q(PC_fetch) );
  regFFD_NBIT32_14 pipeline_fetch_ir ( .CK(CLK), .RESET(n9), .ENABLE(
        ir_LATCH_EN), .D(IR), .Q(ir_fetch) );
  regFFD_NBIT32_13 pipeline_newpc1 ( .CK(CLK), .RESET(n9), .ENABLE(
        NPC_LATCH_EN), .D(NPC_fetch), .Q(NPC_Dec) );
  regFFD_NBIT32_12 pipeline_pc1 ( .CK(CLK), .RESET(n9), .ENABLE(ir_LATCH_EN), 
        .D(PC_fetch) );
  regFFD_NBIT32_11 pipeline_IR1 ( .CK(CLK), .RESET(n9), .ENABLE(ir_LATCH_EN), 
        .D(ir_fetch), .Q(IR_Dec) );
  IR_DECODE_NBIT32_opBIT6_regBIT5 IR_OP ( .CLK(CLK), .IR_26(IR_Dec[25:0]), 
        .OPCODE(IR_Dec[31:26]), .is_signed(signed_op), .RS1(RS1), .RS2(RS2), 
        .RD(RD), .IMMEDIATE(Imm) );
  windRF_M8_N8_F5_NBIT32 RF ( .CLK(CLK), .RESET(n8), .ENABLE(1'b1), .CALL(
        trap_cs), .RETRN(ret_cs), .BUSin({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .RD1(RF1), .RD2(RF2), .WR(WF1), .ADD_WR(RD_wb), 
        .ADD_RD1(RS1), .ADD_RD2(RS2), .DATAIN(OUT_wb), .OUT1(regA), .OUT2(regB), .wr_signal(wr_signal_wb) );
  FF_0 pipeline_sign2 ( .CLK(CLK), .RESET(n9), .EN(1'b1), .D(signed_op), .Q(
        signed_op_ex) );
  regFFD_NBIT32_10 pipeline_newpc2 ( .CK(CLK), .RESET(n9), .ENABLE(1'b1), .D(
        NPC_Dec), .Q(NPC_ex) );
  regFFD_NBIT32_9 pipeline_A2 ( .CK(CLK), .RESET(n9), .ENABLE(RF1), .D(regA), 
        .Q(regA_ex) );
  regFFD_NBIT32_8 pipeline_B2 ( .CK(CLK), .RESET(n9), .ENABLE(RF2), .D(regB), 
        .Q(regB_ex) );
  regFFD_NBIT32_7 pipeline_IMM2 ( .CK(CLK), .RESET(n9), .ENABLE(
        regImm_LATCH_EN), .D(Imm), .Q(Imm_ex) );
  regFFD_NBIT5_0 pipeline_RD2 ( .CK(CLK), .RESET(n8), .ENABLE(1'b1), .D(RD), 
        .Q(RD_ex) );
  FF_7 pipeline_wr_signal ( .CLK(CLK), .RESET(n9), .EN(1'b1), .D(n12), .Q(
        wr_signal_exe) );
  regFFD_NBIT6_0 pipeline_IR2 ( .CK(CLK), .RESET(n8), .ENABLE(1'b1), .D({
        IR_Dec[31], n1, n2, IR_Dec[28:26]}), .Q(IR_26_ex) );
  regFFD_NBIT32_6 pipeline_LHI2 ( .CK(CLK), .RESET(n9), .ENABLE(1'b1), .D({
        Imm[15:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Q(LHI_ex) );
  MUX21_GENERIC_NBIT32_6 MUX_ALU_A ( .A(NPC_ex), .B(regA_ex), .SEL(S1), .Y(
        input1_ALU) );
  MUX21_GENERIC_NBIT32_5 MUX_ALU_B ( .A(Imm_ex), .B(regB_ex), .SEL(S2), .Y(
        input2_ALU) );
  ALU_N32 ALU_OP ( .CLK(CLK), .FUNC({\instruction_alu[5] , 
        \instruction_alu[4] , \instruction_alu[3] , \instruction_alu[2] , 
        \instruction_alu[1] , \instruction_alu[0] }), .DATA1(input1_ALU), 
        .DATA2(input2_ALU), .OUT_ALU(ALU_out) );
  zero_eval_NBIT32 ZERO_OP ( .\input (regA_ex), .res(is_zero) );
  COND_BT_NBIT32 COND_OP ( .ZERO_BIT(is_zero), .OPCODE_0(IR_26_ex[0]), 
        .branch_op(branch_cond), .con_sign(cond) );
  MUX21_GENERIC_NBIT32_4 MUX_alu_out ( .A(LHI_ex), .B(ALU_out), .SEL(lhi_sel), 
        .Y(ALU_ex) );
  FF_6 pipeline_sign3 ( .CLK(CLK), .RESET(n9), .EN(1'b1), .D(signed_op_ex), 
        .Q(signed_op_mem) );
  regFFD_NBIT32_5 pipeline_newpc3 ( .CK(CLK), .RESET(n9), .ENABLE(1'b1), .D(
        NPC_ex), .Q(NPC_mem) );
  FF_5 pipeline_cond3 ( .CLK(CLK), .RESET(n9), .EN(1'b1), .D(cond), .Q(
        cond_mem) );
  regFFD_NBIT32_4 pipeline_B3 ( .CK(CLK), .RESET(n8), .ENABLE(1'b1), .D(
        regB_ex), .Q(regB_mem) );
  regFFD_NBIT5_2 pipeline_RD3 ( .CK(CLK), .RESET(n8), .ENABLE(1'b1), .D(RD_ex), 
        .Q(RD_mem) );
  FF_4 pipeline_wr_signal2 ( .CLK(CLK), .RESET(n9), .EN(1'b1), .D(
        wr_signal_exe), .Q(wr_signal_mem) );
  regFFD_NBIT6_1 pipeline_IR3 ( .CK(CLK), .RESET(n8), .ENABLE(1'b1), .D(
        IR_26_ex), .Q(IR_26_mem) );
  MUX21_GENERIC_NBIT32_3 MUX_PC ( .A(ALU_ex), .B(NPC_mem), .SEL(sel_npc), .Y(
        PC_OUT_i) );
  load_data LOAD_DATA_OUT ( .data_in(DATA_MEM_OUT), .signed_val(signed_op_mem), 
        .load_op(RM), .load_type(IR_26_mem[1:0]), .data_out(LMD_out) );
  regFFD_NBIT32_3 pipeline_alu4 ( .CK(CLK), .RESET(n8), .ENABLE(1'b1), .D(
        ALU_ex), .Q(ALU_wb) );
  regFFD_NBIT32_2 pipeline_LMD4 ( .CK(CLK), .RESET(n8), .ENABLE(RM), .D(
        LMD_out), .Q(LMD_wb) );
  regFFD_NBIT5_1 pipeline_RD4 ( .CK(CLK), .RESET(n8), .ENABLE(1'b1), .D(RD_mem), .Q(RD_wb) );
  FF_3 pipeline_wr_signal3 ( .CLK(CLK), .RESET(n9), .EN(1'b1), .D(
        wr_signal_mem1), .Q(wr_signal_wb) );
  FF_2 pipeline_WM ( .CLK(CLK), .RESET(n9), .EN(1'b1), .D(WM) );
  FF_1 pipeline_JAL ( .CLK(CLK), .RESET(n9), .EN(1'b1), .D(sel_saved_reg), .Q(
        sel_saved_reg_wb) );
  regFFD_NBIT32_1 pipeline_NPC_wb ( .CK(CLK), .RESET(n8), .ENABLE(1'b1), .D(
        NPC_mem), .Q(NPC_wb) );
  MUX21_GENERIC_NBIT32_2 MUX_WB ( .A(ALU_wb), .B(LMD_wb), .SEL(S3), .Y(
        OUT_data) );
  MUX21_GENERIC_NBIT32_1 MUX_jal ( .A(NPC_wb), .B(OUT_data), .SEL(
        sel_saved_reg_wb), .Y(OUT_wb) );
  DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 add_256 ( .A(PC_fetch0), .SUM(NPC) );
  INV_X1 U3 ( .A(n14), .ZN(n1) );
  CLKBUF_X1 U4 ( .A(IR_Dec[29]), .Z(n2) );
  BUF_X2 U5 ( .A(RST), .Z(n9) );
  BUF_X2 U6 ( .A(RST), .Z(n8) );
  BUF_X1 U7 ( .A(n61), .Z(n3) );
  BUF_X1 U8 ( .A(n61), .Z(n4) );
  BUF_X1 U9 ( .A(N13), .Z(n6) );
  BUF_X1 U10 ( .A(N13), .Z(n5) );
  BUF_X1 U11 ( .A(N13), .Z(n7) );
  NOR4_X1 U12 ( .A1(IR_Dec[21]), .A2(IR_Dec[20]), .A3(IR_Dec[1]), .A4(
        IR_Dec[19]), .ZN(n34) );
  NOR4_X1 U13 ( .A1(IR_Dec[2]), .A2(IR_Dec[28]), .A3(IR_Dec[26]), .A4(
        IR_Dec[25]), .ZN(n36) );
  NAND4_X1 U14 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(n29) );
  NOR3_X1 U15 ( .A1(IR_Dec[22]), .A2(IR_Dec[24]), .A3(IR_Dec[23]), .ZN(n35) );
  NOR3_X1 U16 ( .A1(IR_Dec[3]), .A2(IR_Dec[5]), .A3(IR_Dec[4]), .ZN(n37) );
  NOR4_X1 U17 ( .A1(IR_Dec[9]), .A2(IR_Dec[8]), .A3(IR_Dec[7]), .A4(IR_Dec[6]), 
        .ZN(n38) );
  NAND4_X1 U18 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .ZN(n30) );
  NOR3_X1 U19 ( .A1(IR_Dec[0]), .A2(IR_Dec[11]), .A3(IR_Dec[10]), .ZN(n31) );
  NOR3_X1 U20 ( .A1(IR_Dec[16]), .A2(IR_Dec[18]), .A3(IR_Dec[17]), .ZN(n33) );
  NOR4_X1 U21 ( .A1(IR_Dec[15]), .A2(IR_Dec[14]), .A3(IR_Dec[13]), .A4(
        IR_Dec[12]), .ZN(n32) );
  INV_X1 U22 ( .A(n23), .ZN(n12) );
  INV_X1 U23 ( .A(IR_Dec[31]), .ZN(n13) );
  INV_X1 U24 ( .A(IR_Dec[28]), .ZN(n16) );
  INV_X1 U25 ( .A(n26), .ZN(n15) );
  AOI21_X1 U26 ( .B1(n27), .B2(n28), .A(IR_Dec[27]), .ZN(n26) );
  OAI21_X1 U27 ( .B1(n16), .B2(IR_Dec[26]), .A(n1), .ZN(n28) );
  OR2_X1 U28 ( .A1(n29), .A2(n30), .ZN(n27) );
  AOI21_X1 U29 ( .B1(jump_en), .B2(n21), .A(n11), .ZN(wr_signal_mem1) );
  NAND4_X1 U30 ( .A1(IR_26_mem[1]), .A2(IR_26_mem[0]), .A3(n22), .A4(n10), 
        .ZN(n21) );
  INV_X1 U31 ( .A(wr_signal_mem), .ZN(n11) );
  INV_X1 U32 ( .A(IR_26_mem[2]), .ZN(n10) );
  INV_X1 U33 ( .A(IR_Dec[30]), .ZN(n14) );
  NAND4_X1 U34 ( .A1(IR_26_mem[2]), .A2(IR_26_mem[0]), .A3(IR_26_mem[4]), .A4(
        n39), .ZN(N13) );
  NOR3_X1 U35 ( .A1(IR_26_mem[1]), .A2(IR_26_mem[5]), .A3(IR_26_mem[3]), .ZN(
        n39) );
  AOI22_X1 U36 ( .A1(n51), .A2(instruction_alu[1]), .B1(instruction_alu[2]), 
        .B2(n59), .ZN(n50) );
  INV_X1 U37 ( .A(instruction_alu[1]), .ZN(n59) );
  NOR2_X1 U38 ( .A1(instruction_alu[2]), .A2(n60), .ZN(n51) );
  OR2_X1 U39 ( .A1(cond_mem), .A2(jump_en), .ZN(sel_npc) );
  INV_X1 U40 ( .A(instruction_alu[0]), .ZN(n60) );
  INV_X1 U41 ( .A(sb_op), .ZN(n61) );
  INV_X1 U42 ( .A(instruction_alu[3]), .ZN(n58) );
  NOR2_X1 U43 ( .A1(IR_26_mem[5]), .A2(IR_26_mem[3]), .ZN(n22) );
  OR4_X1 U44 ( .A1(n48), .A2(n49), .A3(WM), .A4(RM), .ZN(DATA_MEM_ENABLE) );
  NOR4_X1 U45 ( .A1(instruction_alu[4]), .A2(n50), .A3(n58), .A4(n57), .ZN(n49) );
  NOR4_X1 U46 ( .A1(n52), .A2(n60), .A3(instruction_alu[5]), .A4(
        instruction_alu[3]), .ZN(n48) );
  INV_X1 U47 ( .A(instruction_alu[5]), .ZN(n57) );
  AND2_X1 U48 ( .A1(IR_26_mem[0]), .A2(jump_en), .ZN(sel_saved_reg) );
  INV_X1 U49 ( .A(n41), .ZN(DATA_MEM_IN[6]) );
  AOI22_X1 U50 ( .A1(n3), .A2(regB_mem[6]), .B1(sb_op), .B2(regB_mem[30]), 
        .ZN(n41) );
  INV_X1 U51 ( .A(n42), .ZN(DATA_MEM_IN[5]) );
  AOI22_X1 U52 ( .A1(n3), .A2(regB_mem[5]), .B1(sb_op), .B2(regB_mem[29]), 
        .ZN(n42) );
  INV_X1 U53 ( .A(n43), .ZN(DATA_MEM_IN[4]) );
  AOI22_X1 U54 ( .A1(n3), .A2(regB_mem[4]), .B1(sb_op), .B2(regB_mem[28]), 
        .ZN(n43) );
  INV_X1 U55 ( .A(n44), .ZN(DATA_MEM_IN[3]) );
  AOI22_X1 U56 ( .A1(n3), .A2(regB_mem[3]), .B1(sb_op), .B2(regB_mem[27]), 
        .ZN(n44) );
  INV_X1 U57 ( .A(n45), .ZN(DATA_MEM_IN[2]) );
  AOI22_X1 U58 ( .A1(n3), .A2(regB_mem[2]), .B1(sb_op), .B2(regB_mem[26]), 
        .ZN(n45) );
  INV_X1 U59 ( .A(n46), .ZN(DATA_MEM_IN[1]) );
  AOI22_X1 U60 ( .A1(sb_op), .A2(regB_mem[25]), .B1(n3), .B2(regB_mem[1]), 
        .ZN(n46) );
  INV_X1 U61 ( .A(n47), .ZN(DATA_MEM_IN[0]) );
  AOI22_X1 U62 ( .A1(sb_op), .A2(regB_mem[24]), .B1(n3), .B2(regB_mem[0]), 
        .ZN(n47) );
  INV_X1 U63 ( .A(n40), .ZN(DATA_MEM_IN[7]) );
  AOI22_X1 U64 ( .A1(n3), .A2(regB_mem[7]), .B1(regB_mem[31]), .B2(sb_op), 
        .ZN(n40) );
  AND2_X1 U65 ( .A1(n4), .A2(regB_mem[31]), .ZN(DATA_MEM_IN[31]) );
  AND2_X1 U66 ( .A1(n4), .A2(regB_mem[30]), .ZN(DATA_MEM_IN[30]) );
  AND2_X1 U67 ( .A1(n4), .A2(regB_mem[29]), .ZN(DATA_MEM_IN[29]) );
  AND2_X1 U68 ( .A1(n4), .A2(regB_mem[28]), .ZN(DATA_MEM_IN[28]) );
  AND2_X1 U69 ( .A1(n4), .A2(regB_mem[27]), .ZN(DATA_MEM_IN[27]) );
  AND2_X1 U70 ( .A1(n4), .A2(regB_mem[26]), .ZN(DATA_MEM_IN[26]) );
  AND2_X1 U71 ( .A1(n4), .A2(regB_mem[25]), .ZN(DATA_MEM_IN[25]) );
  AND2_X1 U72 ( .A1(n4), .A2(regB_mem[24]), .ZN(DATA_MEM_IN[24]) );
  AND2_X1 U73 ( .A1(regB_mem[14]), .A2(n3), .ZN(DATA_MEM_IN[14]) );
  AND2_X1 U74 ( .A1(regB_mem[13]), .A2(n3), .ZN(DATA_MEM_IN[13]) );
  AND2_X1 U75 ( .A1(regB_mem[12]), .A2(n3), .ZN(DATA_MEM_IN[12]) );
  AND2_X1 U76 ( .A1(regB_mem[11]), .A2(n3), .ZN(DATA_MEM_IN[11]) );
  AND2_X1 U77 ( .A1(regB_mem[10]), .A2(n3), .ZN(DATA_MEM_IN[10]) );
  AND2_X1 U78 ( .A1(regB_mem[9]), .A2(n3), .ZN(DATA_MEM_IN[9]) );
  AND2_X1 U79 ( .A1(regB_mem[23]), .A2(n4), .ZN(DATA_MEM_IN[23]) );
  AND2_X1 U84 ( .A1(regB_mem[22]), .A2(n4), .ZN(DATA_MEM_IN[22]) );
  AND2_X1 U85 ( .A1(regB_mem[21]), .A2(n4), .ZN(DATA_MEM_IN[21]) );
  AND2_X1 U86 ( .A1(regB_mem[20]), .A2(n4), .ZN(DATA_MEM_IN[20]) );
  AND2_X1 U87 ( .A1(regB_mem[19]), .A2(n4), .ZN(DATA_MEM_IN[19]) );
  AND2_X1 U88 ( .A1(regB_mem[18]), .A2(n4), .ZN(DATA_MEM_IN[18]) );
  AND2_X1 U89 ( .A1(regB_mem[17]), .A2(n4), .ZN(DATA_MEM_IN[17]) );
  AND2_X1 U90 ( .A1(regB_mem[16]), .A2(n4), .ZN(DATA_MEM_IN[16]) );
  AND2_X1 U91 ( .A1(regB_mem[15]), .A2(n4), .ZN(DATA_MEM_IN[15]) );
  AND2_X1 U92 ( .A1(regB_mem[8]), .A2(n4), .ZN(DATA_MEM_IN[8]) );
endmodule


module DLX_IR_SIZE32_PC_SIZE32 ( CLK, RST, IRAM_ADDRESS, IRAM_ISSUE, 
        IRAM_READY, IRAM_DATA, DRAM_ADDRESS, DRAM_ISSUE, DRAM_READNOTWRITE, 
        DRAM_READY, DRAM_DATA );
  output [31:0] IRAM_ADDRESS;
  input [63:0] IRAM_DATA;
  output [31:0] DRAM_ADDRESS;
  inout [63:0] DRAM_DATA;
  input CLK, RST, IRAM_READY, DRAM_READY;
  output IRAM_ISSUE, DRAM_ISSUE, DRAM_READNOTWRITE;
  wire   signed_unsigned_i, lhi_sel_i, sb_op_i, trap_cs_i, ret_cs_i,
         DATA_MEM_WM_i, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273;
  wire   [31:0] IR;
  wire   [31:0] PC;
  wire   [5:0] ALU_OPCODE_i;
  wire   [31:0] DATA_MEM_IN_i;
  wire   [31:0] dram_data_i;
  tri   [63:0] DRAM_DATA;
  assign IRAM_ADDRESS[31] = 1'b0;
  assign IRAM_ADDRESS[30] = 1'b0;
  assign IRAM_ADDRESS[29] = 1'b0;
  assign IRAM_ADDRESS[28] = 1'b0;
  assign IRAM_ADDRESS[27] = 1'b0;
  assign IRAM_ADDRESS[26] = 1'b0;
  assign IRAM_ADDRESS[25] = 1'b0;
  assign IRAM_ADDRESS[24] = 1'b0;
  assign IRAM_ADDRESS[23] = 1'b0;
  assign IRAM_ADDRESS[22] = 1'b0;
  assign IRAM_ADDRESS[21] = 1'b0;
  assign IRAM_ADDRESS[20] = 1'b0;
  assign IRAM_ADDRESS[19] = 1'b0;
  assign IRAM_ADDRESS[18] = 1'b0;
  assign IRAM_ADDRESS[17] = 1'b0;
  assign IRAM_ADDRESS[16] = 1'b0;
  assign IRAM_ADDRESS[15] = 1'b0;
  assign IRAM_ADDRESS[14] = 1'b0;
  assign IRAM_ADDRESS[13] = 1'b0;
  assign IRAM_ADDRESS[12] = 1'b0;
  assign IRAM_ADDRESS[11] = 1'b0;
  assign IRAM_ADDRESS[10] = 1'b0;
  assign IRAM_ADDRESS[9] = 1'b0;
  assign IRAM_ADDRESS[8] = 1'b0;
  assign IRAM_ADDRESS[7] = 1'b0;
  assign IRAM_ADDRESS[6] = 1'b0;
  assign IRAM_ADDRESS[5] = 1'b0;
  assign IRAM_ADDRESS[4] = 1'b0;
  assign IRAM_ADDRESS[3] = 1'b0;
  assign IRAM_ADDRESS[2] = 1'b0;
  assign IRAM_ADDRESS[1] = 1'b0;
  assign IRAM_ADDRESS[0] = 1'b0;

  DFF_X1 DRAM_READNOTWRITE_reg ( .D(n270), .CK(CLK), .Q(DRAM_READNOTWRITE) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 CU_I ( 
        .Clk(CLK), .Rst(n271), .IR_IN({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .ALU_OPCODE(ALU_OPCODE_i), .signed_unsigned(
        signed_unsigned_i), .lhi_sel(lhi_sel_i), .sb_op(sb_op_i), .s_trap(
        trap_cs_i), .s_ret(ret_cs_i) );
  DATAPTH_NBIT32_REG_BIT5 DTPTH_I ( .CLK(CLK), .RST(n271), .PC({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IR({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .NPC_LATCH_EN(1'b0), .ir_LATCH_EN(1'b0), 
        .signed_op(signed_unsigned_i), .trap_cs(trap_cs_i), .ret_cs(ret_cs_i), 
        .RF1(1'b0), .RF2(1'b0), .WF1(1'b0), .regImm_LATCH_EN(1'b0), .S1(1'b0), 
        .S2(1'b0), .EN2(1'b0), .lhi_sel(lhi_sel_i), .jump_en(1'b0), 
        .branch_cond(1'b0), .sb_op(sb_op_i), .RM(1'b0), .WM(1'b0), .EN3(1'b0), 
        .S3(1'b0), .instruction_alu(ALU_OPCODE_i), .DATA_MEM_ADDR(DRAM_ADDRESS), .DATA_MEM_IN(DATA_MEM_IN_i), .DATA_MEM_OUT(dram_data_i), .DATA_MEM_ENABLE(
        DRAM_ISSUE), .DATA_MEM_WM(DATA_MEM_WM_i) );
  TBUF_X1 \DRAM_DATA_tri[32]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[32]) );
  TBUF_X1 \DRAM_DATA_tri[33]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[33]) );
  TBUF_X1 \DRAM_DATA_tri[34]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[34]) );
  TBUF_X1 \DRAM_DATA_tri[35]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[35]) );
  TBUF_X1 \DRAM_DATA_tri[36]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[36]) );
  TBUF_X1 \DRAM_DATA_tri[37]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[37]) );
  TBUF_X1 \DRAM_DATA_tri[38]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[38]) );
  TBUF_X1 \DRAM_DATA_tri[39]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[39]) );
  TBUF_X1 \DRAM_DATA_tri[40]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[40]) );
  TBUF_X1 \DRAM_DATA_tri[41]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[41]) );
  TBUF_X1 \DRAM_DATA_tri[42]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[42]) );
  TBUF_X1 \DRAM_DATA_tri[43]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[43]) );
  TBUF_X1 \DRAM_DATA_tri[44]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[44]) );
  TBUF_X1 \DRAM_DATA_tri[45]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[45]) );
  TBUF_X1 \DRAM_DATA_tri[46]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[46]) );
  TBUF_X1 \DRAM_DATA_tri[47]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[47]) );
  TBUF_X1 \DRAM_DATA_tri[48]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[48]) );
  TBUF_X1 \DRAM_DATA_tri[49]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[49]) );
  TBUF_X1 \DRAM_DATA_tri[50]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[50]) );
  TBUF_X1 \DRAM_DATA_tri[51]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[51]) );
  TBUF_X1 \DRAM_DATA_tri[52]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[52]) );
  TBUF_X1 \DRAM_DATA_tri[53]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[53]) );
  TBUF_X1 \DRAM_DATA_tri[54]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[54]) );
  TBUF_X1 \DRAM_DATA_tri[55]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[55]) );
  TBUF_X1 \DRAM_DATA_tri[56]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[56]) );
  TBUF_X1 \DRAM_DATA_tri[57]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[57]) );
  TBUF_X1 \DRAM_DATA_tri[58]  ( .A(1'b0), .EN(n267), .Z(DRAM_DATA[58]) );
  TBUF_X1 \DRAM_DATA_tri[59]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[59]) );
  TBUF_X1 \DRAM_DATA_tri[60]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[60]) );
  TBUF_X1 \DRAM_DATA_tri[61]  ( .A(1'b0), .EN(n268), .Z(DRAM_DATA[61]) );
  TBUF_X1 \DRAM_DATA_tri[62]  ( .A(1'b0), .EN(n263), .Z(DRAM_DATA[62]) );
  TBUF_X1 \DRAM_DATA_tri[63]  ( .A(1'b0), .EN(n268), .Z(DRAM_DATA[63]) );
  TBUF_X1 \DRAM_DATA_tri[0]  ( .A(DATA_MEM_IN_i[0]), .EN(n265), .Z(
        DRAM_DATA[0]) );
  TBUF_X1 \DRAM_DATA_tri[1]  ( .A(DATA_MEM_IN_i[1]), .EN(n266), .Z(
        DRAM_DATA[1]) );
  TBUF_X1 \DRAM_DATA_tri[2]  ( .A(DATA_MEM_IN_i[2]), .EN(n264), .Z(
        DRAM_DATA[2]) );
  TBUF_X1 \DRAM_DATA_tri[3]  ( .A(DATA_MEM_IN_i[3]), .EN(n267), .Z(
        DRAM_DATA[3]) );
  TBUF_X1 \DRAM_DATA_tri[4]  ( .A(DATA_MEM_IN_i[4]), .EN(n263), .Z(
        DRAM_DATA[4]) );
  TBUF_X1 \DRAM_DATA_tri[5]  ( .A(DATA_MEM_IN_i[5]), .EN(n267), .Z(
        DRAM_DATA[5]) );
  TBUF_X1 \DRAM_DATA_tri[6]  ( .A(DATA_MEM_IN_i[6]), .EN(n263), .Z(
        DRAM_DATA[6]) );
  TBUF_X1 \DRAM_DATA_tri[7]  ( .A(DATA_MEM_IN_i[7]), .EN(n268), .Z(
        DRAM_DATA[7]) );
  TBUF_X1 \DRAM_DATA_tri[8]  ( .A(DATA_MEM_IN_i[8]), .EN(n263), .Z(
        DRAM_DATA[8]) );
  TBUF_X1 \DRAM_DATA_tri[9]  ( .A(DATA_MEM_IN_i[9]), .EN(n268), .Z(
        DRAM_DATA[9]) );
  TBUF_X1 \DRAM_DATA_tri[10]  ( .A(DATA_MEM_IN_i[10]), .EN(n265), .Z(
        DRAM_DATA[10]) );
  TBUF_X1 \DRAM_DATA_tri[11]  ( .A(DATA_MEM_IN_i[11]), .EN(n265), .Z(
        DRAM_DATA[11]) );
  TBUF_X1 \DRAM_DATA_tri[12]  ( .A(DATA_MEM_IN_i[12]), .EN(n265), .Z(
        DRAM_DATA[12]) );
  TBUF_X1 \DRAM_DATA_tri[13]  ( .A(DATA_MEM_IN_i[13]), .EN(n265), .Z(
        DRAM_DATA[13]) );
  TBUF_X1 \DRAM_DATA_tri[14]  ( .A(DATA_MEM_IN_i[14]), .EN(n265), .Z(
        DRAM_DATA[14]) );
  TBUF_X1 \DRAM_DATA_tri[15]  ( .A(DATA_MEM_IN_i[15]), .EN(n265), .Z(
        DRAM_DATA[15]) );
  TBUF_X1 \DRAM_DATA_tri[16]  ( .A(DATA_MEM_IN_i[16]), .EN(n265), .Z(
        DRAM_DATA[16]) );
  TBUF_X1 \DRAM_DATA_tri[17]  ( .A(DATA_MEM_IN_i[17]), .EN(n265), .Z(
        DRAM_DATA[17]) );
  TBUF_X1 \DRAM_DATA_tri[18]  ( .A(DATA_MEM_IN_i[18]), .EN(n266), .Z(
        DRAM_DATA[18]) );
  TBUF_X1 \DRAM_DATA_tri[19]  ( .A(DATA_MEM_IN_i[19]), .EN(n265), .Z(
        DRAM_DATA[19]) );
  TBUF_X1 \DRAM_DATA_tri[20]  ( .A(DATA_MEM_IN_i[20]), .EN(n265), .Z(
        DRAM_DATA[20]) );
  TBUF_X1 \DRAM_DATA_tri[21]  ( .A(DATA_MEM_IN_i[21]), .EN(n266), .Z(
        DRAM_DATA[21]) );
  TBUF_X1 \DRAM_DATA_tri[22]  ( .A(DATA_MEM_IN_i[22]), .EN(n265), .Z(
        DRAM_DATA[22]) );
  TBUF_X1 \DRAM_DATA_tri[23]  ( .A(DATA_MEM_IN_i[23]), .EN(n266), .Z(
        DRAM_DATA[23]) );
  TBUF_X1 \DRAM_DATA_tri[24]  ( .A(DATA_MEM_IN_i[24]), .EN(n264), .Z(
        DRAM_DATA[24]) );
  TBUF_X1 \DRAM_DATA_tri[25]  ( .A(DATA_MEM_IN_i[25]), .EN(n266), .Z(
        DRAM_DATA[25]) );
  TBUF_X1 \DRAM_DATA_tri[26]  ( .A(DATA_MEM_IN_i[26]), .EN(n264), .Z(
        DRAM_DATA[26]) );
  TBUF_X1 \DRAM_DATA_tri[27]  ( .A(DATA_MEM_IN_i[27]), .EN(n266), .Z(
        DRAM_DATA[27]) );
  TBUF_X1 \DRAM_DATA_tri[28]  ( .A(DATA_MEM_IN_i[28]), .EN(n264), .Z(
        DRAM_DATA[28]) );
  TBUF_X1 \DRAM_DATA_tri[29]  ( .A(DATA_MEM_IN_i[29]), .EN(n266), .Z(
        DRAM_DATA[29]) );
  TBUF_X1 \DRAM_DATA_tri[30]  ( .A(DATA_MEM_IN_i[30]), .EN(n266), .Z(
        DRAM_DATA[30]) );
  TBUF_X1 \DRAM_DATA_tri[31]  ( .A(DATA_MEM_IN_i[31]), .EN(n264), .Z(
        DRAM_DATA[31]) );
  BUF_X1 U198 ( .A(n260), .Z(n263) );
  BUF_X1 U199 ( .A(n261), .Z(n267) );
  BUF_X1 U200 ( .A(n260), .Z(n264) );
  BUF_X1 U201 ( .A(n261), .Z(n266) );
  BUF_X1 U202 ( .A(n260), .Z(n265) );
  BUF_X1 U203 ( .A(n261), .Z(n268) );
  BUF_X1 U204 ( .A(n262), .Z(n269) );
  AND2_X1 U205 ( .A1(DRAM_DATA[63]), .A2(n269), .ZN(dram_data_i[31]) );
  AND2_X1 U206 ( .A1(DRAM_DATA[40]), .A2(n270), .ZN(dram_data_i[8]) );
  AND2_X1 U207 ( .A1(DRAM_DATA[41]), .A2(n270), .ZN(dram_data_i[9]) );
  AND2_X1 U208 ( .A1(DRAM_DATA[42]), .A2(n268), .ZN(dram_data_i[10]) );
  AND2_X1 U209 ( .A1(DRAM_DATA[43]), .A2(n268), .ZN(dram_data_i[11]) );
  AND2_X1 U210 ( .A1(DRAM_DATA[44]), .A2(n268), .ZN(dram_data_i[12]) );
  AND2_X1 U211 ( .A1(DRAM_DATA[45]), .A2(n268), .ZN(dram_data_i[13]) );
  AND2_X1 U212 ( .A1(DRAM_DATA[46]), .A2(n268), .ZN(dram_data_i[14]) );
  AND2_X1 U213 ( .A1(DRAM_DATA[47]), .A2(n268), .ZN(dram_data_i[15]) );
  AND2_X1 U214 ( .A1(DRAM_DATA[52]), .A2(n269), .ZN(dram_data_i[20]) );
  AND2_X1 U215 ( .A1(DRAM_DATA[53]), .A2(n269), .ZN(dram_data_i[21]) );
  AND2_X1 U216 ( .A1(DRAM_DATA[54]), .A2(n269), .ZN(dram_data_i[22]) );
  AND2_X1 U217 ( .A1(DRAM_DATA[55]), .A2(n269), .ZN(dram_data_i[23]) );
  AND2_X1 U218 ( .A1(DRAM_DATA[56]), .A2(n269), .ZN(dram_data_i[24]) );
  AND2_X1 U219 ( .A1(DRAM_DATA[57]), .A2(n269), .ZN(dram_data_i[25]) );
  AND2_X1 U220 ( .A1(DRAM_DATA[58]), .A2(n269), .ZN(dram_data_i[26]) );
  AND2_X1 U221 ( .A1(DRAM_DATA[59]), .A2(n269), .ZN(dram_data_i[27]) );
  AND2_X1 U222 ( .A1(DRAM_DATA[60]), .A2(n269), .ZN(dram_data_i[28]) );
  AND2_X1 U223 ( .A1(DRAM_DATA[61]), .A2(n269), .ZN(dram_data_i[29]) );
  AND2_X1 U224 ( .A1(DRAM_DATA[62]), .A2(n269), .ZN(dram_data_i[30]) );
  AND2_X1 U225 ( .A1(DRAM_DATA[48]), .A2(n268), .ZN(dram_data_i[16]) );
  AND2_X1 U226 ( .A1(DRAM_DATA[49]), .A2(n268), .ZN(dram_data_i[17]) );
  AND2_X1 U227 ( .A1(DRAM_DATA[50]), .A2(n268), .ZN(dram_data_i[18]) );
  AND2_X1 U228 ( .A1(DRAM_DATA[51]), .A2(n269), .ZN(dram_data_i[19]) );
  BUF_X1 U229 ( .A(n272), .Z(n271) );
  BUF_X1 U230 ( .A(RST), .Z(n272) );
  AND2_X1 U231 ( .A1(DRAM_DATA[32]), .A2(n268), .ZN(dram_data_i[0]) );
  AND2_X1 U232 ( .A1(DRAM_DATA[33]), .A2(n268), .ZN(dram_data_i[1]) );
  AND2_X1 U233 ( .A1(DRAM_DATA[34]), .A2(n269), .ZN(dram_data_i[2]) );
  AND2_X1 U234 ( .A1(DRAM_DATA[35]), .A2(n269), .ZN(dram_data_i[3]) );
  AND2_X1 U235 ( .A1(DRAM_DATA[36]), .A2(n270), .ZN(dram_data_i[4]) );
  AND2_X1 U236 ( .A1(DRAM_DATA[37]), .A2(n269), .ZN(dram_data_i[5]) );
  AND2_X1 U237 ( .A1(DRAM_DATA[38]), .A2(n270), .ZN(dram_data_i[6]) );
  AND2_X1 U238 ( .A1(DRAM_DATA[39]), .A2(n270), .ZN(dram_data_i[7]) );
  INV_X1 U239 ( .A(DATA_MEM_WM_i), .ZN(n273) );
  CLKBUF_X1 U336 ( .A(n273), .Z(n260) );
  CLKBUF_X1 U337 ( .A(n273), .Z(n261) );
  CLKBUF_X1 U338 ( .A(n273), .Z(n262) );
  CLKBUF_X1 U339 ( .A(n262), .Z(n270) );
endmodule




    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 ( 
        A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85;

  INV_X1 U2 ( .A(A[2]), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(n2) );
  AND2_X2 U4 ( .A1(n29), .A2(n78), .ZN(n26) );
  AND2_X2 U5 ( .A1(n85), .A2(n84), .ZN(n12) );
  AND2_X2 U6 ( .A1(n12), .A2(n78), .ZN(n15) );
  AND2_X1 U7 ( .A1(n15), .A2(n72), .ZN(n22) );
  AND2_X1 U8 ( .A1(n25), .A2(n24), .ZN(n30) );
  AND3_X1 U9 ( .A1(n8), .A2(A[17]), .A3(n22), .ZN(n3) );
  AND2_X1 U10 ( .A1(A[12]), .A2(A[13]), .ZN(n4) );
  AND2_X1 U11 ( .A1(A[20]), .A2(A[21]), .ZN(n5) );
  NOR2_X1 U12 ( .A1(n69), .A2(n70), .ZN(n6) );
  AND2_X1 U13 ( .A1(A[24]), .A2(A[25]), .ZN(n7) );
  CLKBUF_X1 U14 ( .A(A[16]), .Z(n8) );
  AND4_X1 U15 ( .A1(A[1]), .A2(A[0]), .A3(A[3]), .A4(A[2]), .ZN(n9) );
  AND4_X1 U16 ( .A1(A[1]), .A2(A[0]), .A3(A[3]), .A4(A[2]), .ZN(n85) );
  XOR2_X1 U17 ( .A(A[18]), .B(n3), .Z(SUM[18]) );
  AND2_X1 U18 ( .A1(n5), .A2(n24), .ZN(n10) );
  XOR2_X1 U19 ( .A(A[7]), .B(n11), .Z(SUM[7]) );
  AND2_X1 U20 ( .A1(n40), .A2(A[6]), .ZN(n11) );
  AND2_X2 U21 ( .A1(n23), .A2(n26), .ZN(n28) );
  AND2_X1 U22 ( .A1(n15), .A2(n4), .ZN(n13) );
  CLKBUF_X1 U23 ( .A(n26), .Z(n14) );
  INV_X1 U24 ( .A(n14), .ZN(n27) );
  CLKBUF_X1 U25 ( .A(A[4]), .Z(n16) );
  AND4_X2 U26 ( .A1(A[5]), .A2(A[4]), .A3(A[7]), .A4(A[6]), .ZN(n84) );
  AND3_X1 U27 ( .A1(n64), .A2(n72), .A3(n6), .ZN(n23) );
  AND2_X1 U28 ( .A1(n58), .A2(n26), .ZN(n17) );
  XOR2_X1 U29 ( .A(A[25]), .B(n18), .Z(SUM[25]) );
  AND2_X1 U30 ( .A1(A[24]), .A2(n28), .ZN(n18) );
  AND2_X1 U31 ( .A1(n9), .A2(n84), .ZN(n19) );
  CLKBUF_X1 U32 ( .A(n2), .Z(n20) );
  AND2_X1 U33 ( .A1(n9), .A2(n84), .ZN(n29) );
  AND2_X1 U34 ( .A1(n28), .A2(n7), .ZN(n61) );
  INV_X1 U35 ( .A(n22), .ZN(n71) );
  AND2_X1 U36 ( .A1(n10), .A2(n25), .ZN(n21) );
  NAND2_X1 U37 ( .A1(n26), .A2(n4), .ZN(n76) );
  NAND2_X1 U38 ( .A1(n30), .A2(n5), .ZN(n67) );
  INV_X1 U39 ( .A(n28), .ZN(n63) );
  INV_X1 U40 ( .A(n19), .ZN(n39) );
  AND2_X1 U41 ( .A1(n29), .A2(n78), .ZN(n24) );
  AND2_X1 U42 ( .A1(n72), .A2(n6), .ZN(n25) );
  INV_X1 U43 ( .A(n30), .ZN(n68) );
  INV_X1 U44 ( .A(SUM[0]), .ZN(n31) );
  XOR2_X1 U45 ( .A(A[9]), .B(n32), .Z(SUM[9]) );
  AND2_X1 U46 ( .A1(A[8]), .A2(n19), .ZN(n32) );
  XOR2_X1 U47 ( .A(A[21]), .B(n33), .Z(SUM[21]) );
  AND2_X1 U48 ( .A1(A[20]), .A2(n30), .ZN(n33) );
  XOR2_X1 U49 ( .A(A[17]), .B(n34), .Z(SUM[17]) );
  AND2_X1 U50 ( .A1(A[16]), .A2(n22), .ZN(n34) );
  NOR2_X1 U51 ( .A1(n73), .A2(n74), .ZN(n72) );
  NAND2_X1 U52 ( .A1(A[15]), .A2(A[14]), .ZN(n73) );
  NAND2_X1 U53 ( .A1(A[12]), .A2(A[13]), .ZN(n74) );
  NAND2_X1 U54 ( .A1(n17), .A2(n23), .ZN(n51) );
  NOR2_X1 U55 ( .A1(n59), .A2(n60), .ZN(n58) );
  NAND2_X1 U56 ( .A1(A[27]), .A2(A[26]), .ZN(n59) );
  NAND2_X1 U57 ( .A1(A[24]), .A2(A[25]), .ZN(n60) );
  INV_X1 U58 ( .A(A[30]), .ZN(n53) );
  NOR2_X1 U59 ( .A1(n51), .A2(n54), .ZN(n52) );
  NOR2_X1 U60 ( .A1(n79), .A2(n80), .ZN(n78) );
  NAND2_X1 U61 ( .A1(A[11]), .A2(A[10]), .ZN(n79) );
  NAND2_X1 U62 ( .A1(A[8]), .A2(A[9]), .ZN(n80) );
  NOR2_X1 U63 ( .A1(n65), .A2(n66), .ZN(n64) );
  NAND2_X1 U64 ( .A1(A[23]), .A2(A[22]), .ZN(n65) );
  NAND2_X1 U65 ( .A1(A[20]), .A2(A[21]), .ZN(n66) );
  XOR2_X1 U66 ( .A(A[19]), .B(n35), .Z(SUM[19]) );
  AND2_X1 U67 ( .A1(n3), .A2(A[18]), .ZN(n35) );
  XOR2_X1 U68 ( .A(A[23]), .B(n36), .Z(SUM[23]) );
  AND2_X1 U69 ( .A1(n21), .A2(A[22]), .ZN(n36) );
  XNOR2_X1 U70 ( .A(A[14]), .B(n76), .ZN(SUM[14]) );
  XNOR2_X1 U71 ( .A(A[10]), .B(n83), .ZN(SUM[10]) );
  XNOR2_X1 U72 ( .A(A[22]), .B(n67), .ZN(SUM[22]) );
  XNOR2_X1 U73 ( .A(A[3]), .B(n45), .ZN(SUM[3]) );
  INV_X1 U74 ( .A(n47), .ZN(n46) );
  NAND2_X1 U75 ( .A1(A[19]), .A2(A[18]), .ZN(n69) );
  NAND2_X1 U76 ( .A1(A[16]), .A2(A[17]), .ZN(n70) );
  XNOR2_X1 U77 ( .A(A[5]), .B(n43), .ZN(SUM[5]) );
  INV_X1 U78 ( .A(n42), .ZN(n44) );
  XNOR2_X1 U79 ( .A(A[13]), .B(n77), .ZN(SUM[13]) );
  NAND2_X1 U80 ( .A1(A[12]), .A2(n15), .ZN(n77) );
  OR2_X1 U81 ( .A1(n37), .A2(n42), .ZN(n41) );
  NAND2_X1 U82 ( .A1(A[5]), .A2(A[4]), .ZN(n37) );
  NAND2_X1 U83 ( .A1(A[28]), .A2(A[29]), .ZN(n54) );
  INV_X1 U84 ( .A(A[31]), .ZN(n49) );
  NOR2_X1 U85 ( .A1(n51), .A2(n50), .ZN(n48) );
  INV_X1 U86 ( .A(A[29]), .ZN(n56) );
  NOR2_X1 U87 ( .A1(n51), .A2(n57), .ZN(n55) );
  INV_X1 U88 ( .A(A[28]), .ZN(n57) );
  XNOR2_X1 U89 ( .A(n55), .B(n56), .ZN(SUM[29]) );
  XNOR2_X1 U90 ( .A(n52), .B(n53), .ZN(SUM[30]) );
  XNOR2_X1 U91 ( .A(n48), .B(n49), .ZN(SUM[31]) );
  XNOR2_X1 U92 ( .A(A[26]), .B(n62), .ZN(SUM[26]) );
  XNOR2_X1 U93 ( .A(n51), .B(A[28]), .ZN(SUM[28]) );
  XNOR2_X1 U94 ( .A(A[6]), .B(n41), .ZN(SUM[6]) );
  XOR2_X1 U95 ( .A(A[27]), .B(n38), .Z(SUM[27]) );
  AND2_X1 U96 ( .A1(n61), .A2(A[26]), .ZN(n38) );
  NAND2_X1 U97 ( .A1(n16), .A2(n44), .ZN(n43) );
  XNOR2_X1 U98 ( .A(A[20]), .B(n68), .ZN(SUM[20]) );
  XNOR2_X1 U99 ( .A(n20), .B(n47), .ZN(SUM[2]) );
  XNOR2_X1 U100 ( .A(n8), .B(n71), .ZN(SUM[16]) );
  NAND2_X1 U101 ( .A1(n2), .A2(n46), .ZN(n45) );
  INV_X1 U102 ( .A(A[0]), .ZN(SUM[0]) );
  XNOR2_X1 U103 ( .A(A[12]), .B(n27), .ZN(SUM[12]) );
  NAND2_X1 U104 ( .A1(A[1]), .A2(n31), .ZN(n47) );
  NAND4_X1 U105 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(n42) );
  XNOR2_X1 U106 ( .A(A[24]), .B(n63), .ZN(SUM[24]) );
  XNOR2_X1 U107 ( .A(A[8]), .B(n39), .ZN(SUM[8]) );
  INV_X1 U108 ( .A(n41), .ZN(n40) );
  XNOR2_X1 U109 ( .A(n16), .B(n42), .ZN(SUM[4]) );
  NAND3_X1 U110 ( .A1(A[30]), .A2(A[29]), .A3(A[28]), .ZN(n50) );
  NAND3_X1 U111 ( .A1(A[24]), .A2(A[25]), .A3(n28), .ZN(n62) );
  XOR2_X1 U112 ( .A(A[1]), .B(n31), .Z(SUM[1]) );
  XNOR2_X1 U113 ( .A(A[15]), .B(n75), .ZN(SUM[15]) );
  NAND2_X1 U114 ( .A1(n13), .A2(A[14]), .ZN(n75) );
  XNOR2_X1 U115 ( .A(A[11]), .B(n81), .ZN(SUM[11]) );
  NAND2_X1 U116 ( .A1(n82), .A2(A[10]), .ZN(n81) );
  INV_X1 U117 ( .A(n83), .ZN(n82) );
  NAND3_X1 U118 ( .A1(A[8]), .A2(A[9]), .A3(n12), .ZN(n83) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 ( 
        A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;

  AND2_X1 U2 ( .A1(n46), .A2(n36), .ZN(n17) );
  OR2_X1 U3 ( .A1(n19), .A2(n61), .ZN(n43) );
  INV_X1 U4 ( .A(n68), .ZN(n67) );
  INV_X1 U5 ( .A(n17), .ZN(n89) );
  INV_X1 U6 ( .A(n14), .ZN(n83) );
  AND2_X1 U7 ( .A1(n13), .A2(A[17]), .ZN(n1) );
  AND2_X1 U8 ( .A1(A[19]), .A2(A[18]), .ZN(n2) );
  AND2_X1 U9 ( .A1(A[16]), .A2(A[17]), .ZN(n3) );
  NOR2_X1 U10 ( .A1(n80), .A2(n61), .ZN(n4) );
  AND2_X1 U11 ( .A1(A[24]), .A2(A[25]), .ZN(n5) );
  AND2_X1 U12 ( .A1(n27), .A2(n24), .ZN(n6) );
  AND2_X1 U13 ( .A1(n94), .A2(n95), .ZN(n7) );
  AND2_X1 U14 ( .A1(n94), .A2(n95), .ZN(n8) );
  AND2_X1 U15 ( .A1(n94), .A2(n95), .ZN(n59) );
  BUF_X1 U16 ( .A(n12), .Z(n39) );
  AND4_X1 U17 ( .A1(A[15]), .A2(A[14]), .A3(A[12]), .A4(A[13]), .ZN(n9) );
  AND4_X1 U18 ( .A1(A[15]), .A2(A[14]), .A3(A[12]), .A4(A[13]), .ZN(n30) );
  AND4_X2 U19 ( .A1(A[8]), .A2(A[9]), .A3(A[10]), .A4(A[11]), .ZN(n90) );
  CLKBUF_X1 U20 ( .A(A[2]), .Z(n10) );
  CLKBUF_X1 U21 ( .A(A[1]), .Z(n11) );
  NAND2_X1 U22 ( .A1(n15), .A2(n7), .ZN(n12) );
  CLKBUF_X1 U23 ( .A(A[16]), .Z(n13) );
  AND4_X2 U24 ( .A1(n9), .A2(n90), .A3(n3), .A4(n2), .ZN(n15) );
  AND2_X2 U25 ( .A1(n50), .A2(n8), .ZN(n14) );
  AND4_X1 U26 ( .A1(n90), .A2(n30), .A3(n3), .A4(n2), .ZN(n40) );
  CLKBUF_X1 U27 ( .A(A[4]), .Z(n16) );
  XOR2_X1 U28 ( .A(n29), .B(n18), .Z(SUM[13]) );
  AND2_X1 U29 ( .A1(n35), .A2(n17), .ZN(n18) );
  AND2_X1 U30 ( .A1(n46), .A2(n6), .ZN(n92) );
  NAND2_X1 U31 ( .A1(n15), .A2(n7), .ZN(n19) );
  AND3_X1 U32 ( .A1(A[18]), .A2(n14), .A3(n1), .ZN(n57) );
  NOR2_X1 U33 ( .A1(n71), .A2(n70), .ZN(n69) );
  AND4_X1 U34 ( .A1(A[5]), .A2(A[4]), .A3(A[7]), .A4(A[6]), .ZN(n37) );
  NOR3_X1 U35 ( .A1(n20), .A2(n21), .A3(n43), .ZN(n41) );
  INV_X1 U36 ( .A(A[24]), .ZN(n20) );
  INV_X1 U37 ( .A(A[25]), .ZN(n21) );
  NOR2_X1 U38 ( .A1(n79), .A2(n22), .ZN(n56) );
  INV_X1 U39 ( .A(A[22]), .ZN(n22) );
  AND4_X1 U40 ( .A1(A[11]), .A2(A[9]), .A3(A[8]), .A4(A[10]), .ZN(n36) );
  AND4_X1 U41 ( .A1(A[5]), .A2(A[4]), .A3(A[7]), .A4(A[6]), .ZN(n94) );
  AND4_X1 U42 ( .A1(A[1]), .A2(A[0]), .A3(A[3]), .A4(A[2]), .ZN(n38) );
  AND4_X1 U43 ( .A1(A[1]), .A2(A[0]), .A3(A[3]), .A4(A[2]), .ZN(n95) );
  NAND3_X1 U44 ( .A1(n23), .A2(n66), .A3(A[6]), .ZN(n62) );
  INV_X1 U45 ( .A(n55), .ZN(n23) );
  CLKBUF_X1 U46 ( .A(A[8]), .Z(n24) );
  CLKBUF_X1 U47 ( .A(A[11]), .Z(n25) );
  CLKBUF_X1 U48 ( .A(A[14]), .Z(n26) );
  CLKBUF_X1 U49 ( .A(A[9]), .Z(n27) );
  CLKBUF_X1 U50 ( .A(A[10]), .Z(n28) );
  CLKBUF_X1 U51 ( .A(A[13]), .Z(n29) );
  CLKBUF_X1 U52 ( .A(n24), .Z(n31) );
  AND2_X1 U53 ( .A1(n4), .A2(n32), .ZN(n60) );
  AND2_X1 U54 ( .A1(n5), .A2(A[26]), .ZN(n32) );
  AND2_X2 U55 ( .A1(n37), .A2(n38), .ZN(n46) );
  INV_X1 U56 ( .A(n39), .ZN(n33) );
  AND2_X1 U57 ( .A1(n33), .A2(n34), .ZN(n74) );
  AND2_X1 U58 ( .A1(n42), .A2(A[28]), .ZN(n34) );
  CLKBUF_X1 U59 ( .A(A[12]), .Z(n35) );
  NAND2_X1 U60 ( .A1(n14), .A2(n1), .ZN(n82) );
  OR2_X1 U61 ( .A1(n44), .A2(n12), .ZN(n79) );
  NAND2_X1 U62 ( .A1(n40), .A2(n59), .ZN(n80) );
  XOR2_X1 U63 ( .A(n41), .B(A[26]), .Z(SUM[26]) );
  NAND2_X1 U64 ( .A1(n81), .A2(n42), .ZN(n71) );
  NOR2_X1 U65 ( .A1(n61), .A2(n45), .ZN(n42) );
  NAND2_X1 U66 ( .A1(A[20]), .A2(A[21]), .ZN(n44) );
  OR2_X1 U67 ( .A1(n75), .A2(n76), .ZN(n45) );
  INV_X1 U68 ( .A(A[31]), .ZN(n49) );
  CLKBUF_X1 U69 ( .A(A[0]), .Z(n47) );
  NOR2_X1 U70 ( .A1(n85), .A2(n86), .ZN(n48) );
  XNOR2_X1 U71 ( .A(n69), .B(n49), .ZN(SUM[31]) );
  AND2_X1 U72 ( .A1(n36), .A2(n48), .ZN(n50) );
  XOR2_X1 U73 ( .A(A[25]), .B(n51), .Z(SUM[25]) );
  AND2_X1 U74 ( .A1(A[24]), .A2(n4), .ZN(n51) );
  XOR2_X1 U75 ( .A(A[21]), .B(n52), .Z(SUM[21]) );
  AND2_X1 U76 ( .A1(n81), .A2(A[20]), .ZN(n52) );
  XOR2_X1 U77 ( .A(A[15]), .B(n53), .Z(SUM[15]) );
  AND2_X1 U78 ( .A1(n87), .A2(n26), .ZN(n53) );
  NAND2_X1 U79 ( .A1(A[27]), .A2(A[26]), .ZN(n75) );
  NAND2_X1 U80 ( .A1(A[24]), .A2(A[25]), .ZN(n76) );
  XNOR2_X1 U81 ( .A(n28), .B(n93), .ZN(SUM[10]) );
  XNOR2_X1 U82 ( .A(n26), .B(n88), .ZN(SUM[14]) );
  XOR2_X1 U83 ( .A(n27), .B(n54), .Z(SUM[9]) );
  AND2_X1 U84 ( .A1(n31), .A2(n46), .ZN(n54) );
  OR2_X1 U85 ( .A1(n55), .A2(n64), .ZN(n63) );
  NAND2_X1 U86 ( .A1(A[5]), .A2(A[4]), .ZN(n55) );
  XNOR2_X1 U87 ( .A(A[17]), .B(n84), .ZN(SUM[17]) );
  NAND2_X1 U88 ( .A1(n13), .A2(n14), .ZN(n84) );
  XOR2_X1 U89 ( .A(n74), .B(A[29]), .Z(SUM[29]) );
  NAND2_X1 U90 ( .A1(A[15]), .A2(A[14]), .ZN(n85) );
  NAND2_X1 U91 ( .A1(A[13]), .A2(A[12]), .ZN(n86) );
  XOR2_X1 U92 ( .A(n56), .B(A[23]), .Z(SUM[23]) );
  XOR2_X1 U93 ( .A(A[19]), .B(n57), .Z(SUM[19]) );
  XNOR2_X1 U94 ( .A(n79), .B(A[22]), .ZN(SUM[22]) );
  XNOR2_X1 U95 ( .A(A[18]), .B(n82), .ZN(SUM[18]) );
  XOR2_X1 U96 ( .A(n72), .B(A[30]), .Z(SUM[30]) );
  XNOR2_X1 U97 ( .A(A[5]), .B(n65), .ZN(SUM[5]) );
  INV_X1 U98 ( .A(n64), .ZN(n66) );
  XOR2_X1 U99 ( .A(n31), .B(n46), .Z(SUM[8]) );
  NAND2_X1 U100 ( .A1(A[23]), .A2(A[22]), .ZN(n77) );
  NAND2_X1 U101 ( .A1(A[20]), .A2(A[21]), .ZN(n78) );
  NAND2_X1 U102 ( .A1(A[28]), .A2(A[29]), .ZN(n73) );
  XOR2_X1 U103 ( .A(A[3]), .B(n58), .Z(SUM[3]) );
  AND2_X1 U104 ( .A1(n10), .A2(n67), .ZN(n58) );
  NOR2_X1 U105 ( .A1(n71), .A2(n73), .ZN(n72) );
  XNOR2_X1 U106 ( .A(n71), .B(A[28]), .ZN(SUM[28]) );
  XOR2_X1 U107 ( .A(n60), .B(A[27]), .Z(SUM[27]) );
  XNOR2_X1 U108 ( .A(A[6]), .B(n63), .ZN(SUM[6]) );
  NAND2_X1 U109 ( .A1(n16), .A2(n66), .ZN(n65) );
  OR2_X1 U110 ( .A1(n77), .A2(n78), .ZN(n61) );
  XNOR2_X1 U111 ( .A(n43), .B(A[24]), .ZN(SUM[24]) );
  XNOR2_X1 U112 ( .A(A[20]), .B(n39), .ZN(SUM[20]) );
  INV_X1 U113 ( .A(n80), .ZN(n81) );
  XNOR2_X1 U114 ( .A(n13), .B(n83), .ZN(SUM[16]) );
  XNOR2_X1 U115 ( .A(n35), .B(n89), .ZN(SUM[12]) );
  XNOR2_X1 U116 ( .A(n10), .B(n68), .ZN(SUM[2]) );
  INV_X1 U117 ( .A(n47), .ZN(SUM[0]) );
  NAND2_X1 U118 ( .A1(n11), .A2(n47), .ZN(n68) );
  NAND4_X1 U119 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(n64) );
  XNOR2_X1 U120 ( .A(A[7]), .B(n62), .ZN(SUM[7]) );
  XNOR2_X1 U121 ( .A(n16), .B(n64), .ZN(SUM[4]) );
  NAND3_X1 U122 ( .A1(A[30]), .A2(A[29]), .A3(A[28]), .ZN(n70) );
  XOR2_X1 U123 ( .A(n11), .B(n47), .Z(SUM[1]) );
  INV_X1 U124 ( .A(n88), .ZN(n87) );
  NAND3_X1 U125 ( .A1(n35), .A2(n29), .A3(n17), .ZN(n88) );
  XNOR2_X1 U126 ( .A(n25), .B(n91), .ZN(SUM[11]) );
  NAND2_X1 U127 ( .A1(n92), .A2(n28), .ZN(n91) );
  NAND3_X1 U128 ( .A1(n24), .A2(n27), .A3(n46), .ZN(n93) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_6 ( 
        A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  CLKBUF_X1 U2 ( .A(A[2]), .Z(n1) );
  AND2_X1 U3 ( .A1(n40), .A2(n2), .ZN(n34) );
  AND2_X1 U4 ( .A1(n27), .A2(n3), .ZN(n2) );
  INV_X1 U5 ( .A(n41), .ZN(n3) );
  AND2_X2 U6 ( .A1(n16), .A2(n15), .ZN(n40) );
  AND2_X1 U7 ( .A1(A[8]), .A2(A[9]), .ZN(n4) );
  AND2_X1 U8 ( .A1(A[16]), .A2(A[17]), .ZN(n5) );
  CLKBUF_X1 U9 ( .A(A[8]), .Z(n6) );
  NOR2_X1 U10 ( .A1(n55), .A2(n7), .ZN(n37) );
  OR2_X1 U11 ( .A1(n58), .A2(n76), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n17), .A2(n4), .ZN(n95) );
  BUF_X1 U13 ( .A(n49), .Z(n8) );
  AND3_X1 U14 ( .A1(n11), .A2(n13), .A3(n91), .ZN(n9) );
  AND2_X1 U15 ( .A1(n56), .A2(n85), .ZN(n10) );
  AND2_X1 U16 ( .A1(n56), .A2(n85), .ZN(n23) );
  AND4_X1 U17 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .A4(A[3]), .ZN(n11) );
  AND4_X1 U18 ( .A1(A[1]), .A2(A[0]), .A3(A[2]), .A4(A[3]), .ZN(n97) );
  NAND2_X1 U19 ( .A1(A[8]), .A2(A[9]), .ZN(n12) );
  AND4_X1 U20 ( .A1(A[5]), .A2(A[4]), .A3(A[7]), .A4(A[6]), .ZN(n13) );
  CLKBUF_X1 U21 ( .A(A[4]), .Z(n14) );
  AND4_X1 U22 ( .A1(A[5]), .A2(A[4]), .A3(A[7]), .A4(A[6]), .ZN(n96) );
  NOR2_X1 U23 ( .A1(n92), .A2(n12), .ZN(n15) );
  AND2_X1 U24 ( .A1(n11), .A2(n13), .ZN(n16) );
  AND2_X1 U25 ( .A1(n97), .A2(n96), .ZN(n17) );
  AND2_X1 U26 ( .A1(n97), .A2(n96), .ZN(n57) );
  AND4_X1 U27 ( .A1(n85), .A2(n17), .A3(n4), .A4(n18), .ZN(n49) );
  INV_X1 U28 ( .A(n92), .ZN(n18) );
  AND3_X1 U29 ( .A1(n11), .A2(n13), .A3(n91), .ZN(n25) );
  CLKBUF_X1 U30 ( .A(n16), .Z(n19) );
  XOR2_X1 U31 ( .A(A[26]), .B(n20), .Z(SUM[26]) );
  AND3_X1 U32 ( .A1(A[24]), .A2(A[25]), .A3(n39), .ZN(n20) );
  NAND2_X1 U33 ( .A1(n8), .A2(n21), .ZN(n72) );
  AND2_X1 U34 ( .A1(n50), .A2(n22), .ZN(n21) );
  INV_X1 U35 ( .A(n47), .ZN(n22) );
  CLKBUF_X1 U36 ( .A(A[1]), .Z(n24) );
  INV_X1 U37 ( .A(SUM[0]), .ZN(n26) );
  NAND2_X1 U38 ( .A1(n40), .A2(n27), .ZN(n82) );
  AND2_X1 U39 ( .A1(n85), .A2(n28), .ZN(n27) );
  INV_X1 U40 ( .A(n58), .ZN(n28) );
  XOR2_X1 U41 ( .A(A[11]), .B(n29), .Z(SUM[11]) );
  AND2_X1 U42 ( .A1(n94), .A2(A[10]), .ZN(n29) );
  XOR2_X1 U43 ( .A(A[15]), .B(n30), .Z(SUM[15]) );
  AND2_X1 U44 ( .A1(n88), .A2(A[14]), .ZN(n30) );
  AND2_X1 U45 ( .A1(n49), .A2(n50), .ZN(n31) );
  NOR2_X2 U46 ( .A1(n55), .A2(n58), .ZN(n50) );
  INV_X1 U47 ( .A(n34), .ZN(n81) );
  AND2_X1 U48 ( .A1(n23), .A2(n5), .ZN(n32) );
  CLKBUF_X1 U49 ( .A(n82), .Z(n33) );
  XOR2_X1 U50 ( .A(A[17]), .B(n35), .Z(SUM[17]) );
  AND2_X1 U51 ( .A1(A[16]), .A2(n10), .ZN(n35) );
  AND2_X1 U52 ( .A1(n25), .A2(n85), .ZN(n36) );
  AND2_X1 U53 ( .A1(n36), .A2(n37), .ZN(n77) );
  XOR2_X1 U54 ( .A(A[25]), .B(n38), .Z(SUM[25]) );
  AND2_X1 U55 ( .A1(A[24]), .A2(n31), .ZN(n38) );
  AND2_X1 U56 ( .A1(n36), .A2(n50), .ZN(n39) );
  NAND2_X1 U57 ( .A1(n10), .A2(n5), .ZN(n84) );
  AND2_X1 U58 ( .A1(n57), .A2(n15), .ZN(n56) );
  NAND2_X1 U59 ( .A1(A[20]), .A2(A[21]), .ZN(n41) );
  CLKBUF_X1 U60 ( .A(n1), .Z(n42) );
  XOR2_X1 U61 ( .A(A[19]), .B(n43), .Z(SUM[19]) );
  AND2_X1 U62 ( .A1(n32), .A2(A[18]), .ZN(n43) );
  INV_X1 U63 ( .A(n10), .ZN(n44) );
  NAND2_X1 U64 ( .A1(n31), .A2(n45), .ZN(n71) );
  NOR2_X1 U65 ( .A1(n52), .A2(n47), .ZN(n45) );
  XOR2_X1 U66 ( .A(A[27]), .B(n46), .Z(SUM[27]) );
  AND2_X1 U67 ( .A1(n77), .A2(A[26]), .ZN(n46) );
  OR2_X1 U68 ( .A1(n75), .A2(n76), .ZN(n47) );
  XOR2_X1 U69 ( .A(n73), .B(A[29]), .Z(SUM[29]) );
  XOR2_X1 U70 ( .A(n48), .B(A[21]), .Z(SUM[21]) );
  AND2_X1 U71 ( .A1(A[20]), .A2(n83), .ZN(n48) );
  NAND2_X1 U72 ( .A1(n8), .A2(n50), .ZN(n78) );
  XNOR2_X1 U73 ( .A(n24), .B(SUM[0]), .ZN(SUM[1]) );
  NAND2_X1 U74 ( .A1(A[27]), .A2(A[26]), .ZN(n75) );
  NAND2_X1 U75 ( .A1(A[24]), .A2(A[25]), .ZN(n76) );
  XOR2_X1 U76 ( .A(n51), .B(A[23]), .Z(SUM[23]) );
  AND2_X1 U77 ( .A1(n34), .A2(A[22]), .ZN(n51) );
  XOR2_X1 U78 ( .A(n6), .B(n19), .Z(SUM[8]) );
  XNOR2_X1 U79 ( .A(n81), .B(A[22]), .ZN(SUM[22]) );
  XNOR2_X1 U80 ( .A(n89), .B(A[14]), .ZN(SUM[14]) );
  XNOR2_X1 U81 ( .A(A[28]), .B(n72), .ZN(SUM[28]) );
  XNOR2_X1 U82 ( .A(A[9]), .B(n59), .ZN(SUM[9]) );
  XNOR2_X1 U83 ( .A(A[30]), .B(n71), .ZN(SUM[30]) );
  NOR2_X1 U84 ( .A1(n72), .A2(n74), .ZN(n73) );
  INV_X1 U85 ( .A(A[28]), .ZN(n74) );
  OR2_X1 U86 ( .A1(n98), .A2(n63), .ZN(n62) );
  XNOR2_X1 U87 ( .A(A[13]), .B(n90), .ZN(SUM[13]) );
  NOR2_X1 U88 ( .A1(n86), .A2(n87), .ZN(n85) );
  NAND2_X1 U89 ( .A1(A[15]), .A2(A[14]), .ZN(n86) );
  NAND2_X1 U90 ( .A1(A[12]), .A2(A[13]), .ZN(n87) );
  XNOR2_X1 U91 ( .A(A[18]), .B(n84), .ZN(SUM[18]) );
  NOR2_X1 U92 ( .A1(n92), .A2(n93), .ZN(n91) );
  NAND2_X1 U93 ( .A1(A[11]), .A2(A[10]), .ZN(n92) );
  NAND2_X1 U94 ( .A1(A[8]), .A2(A[9]), .ZN(n93) );
  NAND2_X1 U95 ( .A1(A[28]), .A2(A[29]), .ZN(n52) );
  XOR2_X1 U96 ( .A(A[12]), .B(n40), .Z(SUM[12]) );
  XNOR2_X1 U97 ( .A(A[10]), .B(n95), .ZN(SUM[10]) );
  XNOR2_X1 U98 ( .A(A[3]), .B(n66), .ZN(SUM[3]) );
  INV_X1 U99 ( .A(n68), .ZN(n67) );
  XNOR2_X1 U100 ( .A(A[5]), .B(n64), .ZN(SUM[5]) );
  INV_X1 U101 ( .A(n63), .ZN(n65) );
  NAND2_X1 U102 ( .A1(n53), .A2(n54), .ZN(n58) );
  AND2_X1 U103 ( .A1(A[19]), .A2(A[18]), .ZN(n53) );
  AND2_X1 U104 ( .A1(A[16]), .A2(A[17]), .ZN(n54) );
  NAND2_X1 U105 ( .A1(A[20]), .A2(A[21]), .ZN(n80) );
  NAND2_X1 U106 ( .A1(A[23]), .A2(A[22]), .ZN(n79) );
  OR2_X1 U107 ( .A1(n79), .A2(n80), .ZN(n55) );
  NAND2_X1 U108 ( .A1(A[12]), .A2(n9), .ZN(n90) );
  NAND2_X1 U109 ( .A1(n6), .A2(n19), .ZN(n59) );
  XNOR2_X1 U110 ( .A(A[6]), .B(n62), .ZN(SUM[6]) );
  INV_X1 U111 ( .A(n33), .ZN(n83) );
  XNOR2_X1 U112 ( .A(n82), .B(A[20]), .ZN(SUM[20]) );
  XNOR2_X1 U113 ( .A(A[16]), .B(n44), .ZN(SUM[16]) );
  NAND2_X1 U114 ( .A1(n14), .A2(n65), .ZN(n64) );
  NAND2_X1 U115 ( .A1(A[5]), .A2(A[4]), .ZN(n98) );
  XNOR2_X1 U116 ( .A(n42), .B(n68), .ZN(SUM[2]) );
  NAND2_X1 U117 ( .A1(n1), .A2(n67), .ZN(n66) );
  XNOR2_X1 U118 ( .A(A[24]), .B(n78), .ZN(SUM[24]) );
  INV_X1 U119 ( .A(A[0]), .ZN(SUM[0]) );
  NAND2_X1 U120 ( .A1(n24), .A2(n26), .ZN(n68) );
  NAND4_X1 U121 ( .A1(A[3]), .A2(A[2]), .A3(A[1]), .A4(A[0]), .ZN(n63) );
  XNOR2_X1 U122 ( .A(A[7]), .B(n60), .ZN(SUM[7]) );
  NAND2_X1 U123 ( .A1(n61), .A2(A[6]), .ZN(n60) );
  INV_X1 U124 ( .A(n62), .ZN(n61) );
  XNOR2_X1 U125 ( .A(n14), .B(n63), .ZN(SUM[4]) );
  XNOR2_X1 U126 ( .A(A[31]), .B(n69), .ZN(SUM[31]) );
  NAND2_X1 U127 ( .A1(A[30]), .A2(n70), .ZN(n69) );
  INV_X1 U128 ( .A(n71), .ZN(n70) );
  INV_X1 U129 ( .A(n89), .ZN(n88) );
  NAND3_X1 U130 ( .A1(A[12]), .A2(A[13]), .A3(n9), .ZN(n89) );
  INV_X1 U131 ( .A(n95), .ZN(n94) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_7 ( 
        A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110;

  OR2_X2 U2 ( .A1(n100), .A2(n53), .ZN(n72) );
  OR2_X2 U3 ( .A1(n72), .A2(n73), .ZN(n88) );
  INV_X1 U4 ( .A(n46), .ZN(n1) );
  AND2_X1 U5 ( .A1(n10), .A2(n21), .ZN(n2) );
  CLKBUF_X1 U6 ( .A(n35), .Z(n3) );
  OR2_X1 U7 ( .A1(n76), .A2(n60), .ZN(n4) );
  OR2_X1 U8 ( .A1(n4), .A2(n57), .ZN(n96) );
  CLKBUF_X1 U9 ( .A(A[7]), .Z(n5) );
  BUF_X1 U10 ( .A(A[2]), .Z(n20) );
  CLKBUF_X1 U11 ( .A(A[15]), .Z(n6) );
  CLKBUF_X1 U12 ( .A(A[5]), .Z(n7) );
  CLKBUF_X1 U13 ( .A(A[3]), .Z(n8) );
  CLKBUF_X1 U14 ( .A(A[12]), .Z(n9) );
  CLKBUF_X1 U15 ( .A(A[13]), .Z(n10) );
  CLKBUF_X1 U16 ( .A(A[0]), .Z(n11) );
  CLKBUF_X1 U17 ( .A(A[1]), .Z(n12) );
  CLKBUF_X1 U18 ( .A(A[8]), .Z(n13) );
  CLKBUF_X1 U19 ( .A(n6), .Z(n14) );
  NAND2_X1 U20 ( .A1(n15), .A2(n16), .ZN(n60) );
  AND2_X1 U21 ( .A1(A[19]), .A2(A[18]), .ZN(n15) );
  AND2_X1 U22 ( .A1(A[16]), .A2(A[17]), .ZN(n16) );
  CLKBUF_X1 U23 ( .A(A[10]), .Z(n17) );
  AND4_X1 U24 ( .A1(A[5]), .A2(A[6]), .A3(A[7]), .A4(A[4]), .ZN(n18) );
  AND4_X1 U25 ( .A1(A[5]), .A2(A[4]), .A3(A[7]), .A4(A[6]), .ZN(n109) );
  CLKBUF_X1 U26 ( .A(A[4]), .Z(n19) );
  CLKBUF_X1 U27 ( .A(n9), .Z(n21) );
  CLKBUF_X1 U28 ( .A(A[14]), .Z(n22) );
  CLKBUF_X1 U29 ( .A(A[16]), .Z(n23) );
  INV_X1 U30 ( .A(n27), .ZN(n24) );
  CLKBUF_X1 U31 ( .A(A[6]), .Z(n25) );
  AND4_X1 U32 ( .A1(A[1]), .A2(A[0]), .A3(A[3]), .A4(A[2]), .ZN(n26) );
  AND4_X1 U33 ( .A1(A[1]), .A2(A[0]), .A3(A[3]), .A4(A[2]), .ZN(n110) );
  AND4_X1 U34 ( .A1(A[11]), .A2(A[10]), .A3(A[8]), .A4(A[9]), .ZN(n27) );
  CLKBUF_X1 U35 ( .A(n19), .Z(n28) );
  OR2_X1 U36 ( .A1(n66), .A2(n59), .ZN(n57) );
  NAND2_X1 U37 ( .A1(n26), .A2(n18), .ZN(n29) );
  AND2_X1 U38 ( .A1(n26), .A2(n18), .ZN(n30) );
  INV_X1 U39 ( .A(n43), .ZN(n31) );
  NAND4_X1 U40 ( .A1(A[11]), .A2(A[10]), .A3(A[8]), .A4(A[9]), .ZN(n66) );
  NAND4_X1 U41 ( .A1(A[13]), .A2(A[14]), .A3(A[15]), .A4(A[12]), .ZN(n59) );
  AND4_X1 U42 ( .A1(n49), .A2(n48), .A3(n32), .A4(n27), .ZN(n42) );
  INV_X1 U43 ( .A(n52), .ZN(n32) );
  XOR2_X1 U44 ( .A(A[26]), .B(n3), .Z(SUM[26]) );
  NAND2_X1 U45 ( .A1(n106), .A2(n2), .ZN(n103) );
  OR2_X1 U46 ( .A1(n72), .A2(n33), .ZN(n87) );
  OR2_X1 U47 ( .A1(n73), .A2(n70), .ZN(n33) );
  INV_X1 U48 ( .A(A[31]), .ZN(n39) );
  INV_X1 U49 ( .A(SUM[0]), .ZN(n34) );
  NOR2_X1 U50 ( .A1(n47), .A2(n96), .ZN(n35) );
  NOR2_X1 U51 ( .A1(n36), .A2(n46), .ZN(n67) );
  OR2_X1 U52 ( .A1(n74), .A2(n37), .ZN(n36) );
  INV_X1 U53 ( .A(A[24]), .ZN(n37) );
  OR2_X1 U54 ( .A1(n96), .A2(n55), .ZN(n38) );
  OR2_X1 U55 ( .A1(n96), .A2(n55), .ZN(n95) );
  XNOR2_X1 U56 ( .A(n39), .B(n40), .ZN(SUM[31]) );
  AND2_X1 U57 ( .A1(A[30]), .A2(n86), .ZN(n40) );
  XOR2_X1 U58 ( .A(A[20]), .B(n1), .Z(SUM[20]) );
  XOR2_X1 U59 ( .A(A[11]), .B(n41), .Z(SUM[11]) );
  AND2_X1 U60 ( .A1(n107), .A2(n17), .ZN(n41) );
  NAND2_X1 U61 ( .A1(n30), .A2(n42), .ZN(n99) );
  INV_X1 U62 ( .A(n30), .ZN(n43) );
  INV_X1 U63 ( .A(n101), .ZN(n44) );
  OR2_X1 U64 ( .A1(n57), .A2(n29), .ZN(n100) );
  BUF_X1 U65 ( .A(n99), .Z(n45) );
  OR2_X1 U66 ( .A1(n50), .A2(n57), .ZN(n46) );
  OR2_X1 U67 ( .A1(n91), .A2(n74), .ZN(n47) );
  AND2_X1 U68 ( .A1(n6), .A2(A[14]), .ZN(n48) );
  AND2_X1 U69 ( .A1(n9), .A2(A[13]), .ZN(n49) );
  OR2_X1 U70 ( .A1(n76), .A2(n60), .ZN(n50) );
  CLKBUF_X1 U71 ( .A(A[9]), .Z(n51) );
  NAND2_X1 U72 ( .A1(A[16]), .A2(A[17]), .ZN(n52) );
  OR2_X1 U73 ( .A1(n60), .A2(n74), .ZN(n53) );
  CLKBUF_X1 U74 ( .A(n21), .Z(n54) );
  NAND2_X1 U75 ( .A1(A[20]), .A2(A[21]), .ZN(n55) );
  CLKBUF_X1 U76 ( .A(n13), .Z(n56) );
  OR2_X1 U77 ( .A1(n29), .A2(n24), .ZN(n104) );
  INV_X1 U78 ( .A(A[29]), .ZN(n58) );
  XNOR2_X1 U79 ( .A(n61), .B(n58), .ZN(SUM[29]) );
  NOR2_X1 U80 ( .A1(n88), .A2(n89), .ZN(n61) );
  XOR2_X1 U81 ( .A(A[17]), .B(n62), .Z(SUM[17]) );
  AND2_X1 U82 ( .A1(n23), .A2(n101), .ZN(n62) );
  XOR2_X1 U83 ( .A(n63), .B(A[21]), .Z(SUM[21]) );
  AND2_X1 U84 ( .A1(n97), .A2(A[20]), .ZN(n63) );
  XOR2_X1 U85 ( .A(n64), .B(A[23]), .Z(SUM[23]) );
  AND2_X1 U86 ( .A1(n94), .A2(A[22]), .ZN(n64) );
  XOR2_X1 U87 ( .A(n14), .B(n65), .Z(SUM[15]) );
  AND2_X1 U88 ( .A1(n102), .A2(n22), .ZN(n65) );
  XNOR2_X1 U89 ( .A(n38), .B(A[22]), .ZN(SUM[22]) );
  XNOR2_X1 U90 ( .A(n22), .B(n103), .ZN(SUM[14]) );
  XNOR2_X1 U91 ( .A(n51), .B(n75), .ZN(SUM[9]) );
  NAND2_X1 U92 ( .A1(n56), .A2(n31), .ZN(n75) );
  XOR2_X1 U93 ( .A(n67), .B(A[25]), .Z(SUM[25]) );
  OR2_X1 U94 ( .A1(n68), .A2(n80), .ZN(n79) );
  NAND2_X1 U95 ( .A1(A[5]), .A2(n19), .ZN(n68) );
  XNOR2_X1 U96 ( .A(n8), .B(n83), .ZN(SUM[3]) );
  INV_X1 U97 ( .A(n85), .ZN(n84) );
  NAND2_X1 U98 ( .A1(A[27]), .A2(A[26]), .ZN(n90) );
  XOR2_X1 U99 ( .A(A[19]), .B(n69), .Z(SUM[19]) );
  AND2_X1 U100 ( .A1(n98), .A2(A[18]), .ZN(n69) );
  XNOR2_X1 U101 ( .A(n10), .B(n105), .ZN(SUM[13]) );
  NAND2_X1 U102 ( .A1(n54), .A2(n106), .ZN(n105) );
  XNOR2_X1 U103 ( .A(n25), .B(n79), .ZN(SUM[6]) );
  XNOR2_X1 U104 ( .A(A[18]), .B(n45), .ZN(SUM[18]) );
  XNOR2_X1 U105 ( .A(n7), .B(n81), .ZN(SUM[5]) );
  INV_X1 U106 ( .A(n80), .ZN(n82) );
  XNOR2_X1 U107 ( .A(n108), .B(n17), .ZN(SUM[10]) );
  NAND2_X1 U108 ( .A1(A[28]), .A2(A[29]), .ZN(n70) );
  NAND2_X1 U109 ( .A1(A[23]), .A2(A[22]), .ZN(n92) );
  NAND2_X1 U110 ( .A1(A[20]), .A2(A[21]), .ZN(n93) );
  XOR2_X1 U111 ( .A(A[27]), .B(n71), .Z(SUM[27]) );
  AND2_X1 U112 ( .A1(n35), .A2(A[26]), .ZN(n71) );
  INV_X1 U113 ( .A(A[28]), .ZN(n89) );
  NAND2_X1 U114 ( .A1(A[24]), .A2(A[25]), .ZN(n91) );
  XNOR2_X1 U115 ( .A(n87), .B(A[30]), .ZN(SUM[30]) );
  XNOR2_X1 U116 ( .A(A[28]), .B(n88), .ZN(SUM[28]) );
  OR2_X1 U117 ( .A1(n90), .A2(n91), .ZN(n73) );
  XNOR2_X1 U118 ( .A(n20), .B(n85), .ZN(SUM[2]) );
  OR2_X1 U119 ( .A1(n92), .A2(n93), .ZN(n74) );
  NAND2_X1 U120 ( .A1(n28), .A2(n82), .ZN(n81) );
  NAND2_X1 U121 ( .A1(n110), .A2(n109), .ZN(n76) );
  XNOR2_X1 U122 ( .A(n23), .B(n44), .ZN(SUM[16]) );
  INV_X1 U123 ( .A(n100), .ZN(n101) );
  XNOR2_X1 U124 ( .A(n54), .B(n104), .ZN(SUM[12]) );
  INV_X1 U125 ( .A(n104), .ZN(n106) );
  INV_X1 U126 ( .A(n46), .ZN(n97) );
  XOR2_X1 U127 ( .A(n12), .B(n34), .Z(SUM[1]) );
  XNOR2_X1 U128 ( .A(n56), .B(n43), .ZN(SUM[8]) );
  XNOR2_X1 U129 ( .A(A[24]), .B(n72), .ZN(SUM[24]) );
  NAND2_X1 U130 ( .A1(n20), .A2(n84), .ZN(n83) );
  INV_X1 U131 ( .A(n11), .ZN(SUM[0]) );
  NAND2_X1 U132 ( .A1(n12), .A2(n34), .ZN(n85) );
  NAND4_X1 U133 ( .A1(n20), .A2(n8), .A3(A[1]), .A4(n11), .ZN(n80) );
  XNOR2_X1 U134 ( .A(n5), .B(n77), .ZN(SUM[7]) );
  NAND2_X1 U135 ( .A1(n78), .A2(n25), .ZN(n77) );
  INV_X1 U136 ( .A(n79), .ZN(n78) );
  XNOR2_X1 U137 ( .A(n28), .B(n80), .ZN(SUM[4]) );
  INV_X1 U138 ( .A(n87), .ZN(n86) );
  INV_X1 U139 ( .A(n95), .ZN(n94) );
  INV_X1 U140 ( .A(n99), .ZN(n98) );
  INV_X1 U141 ( .A(n103), .ZN(n102) );
  INV_X1 U142 ( .A(n108), .ZN(n107) );
  NAND3_X1 U143 ( .A1(n13), .A2(n51), .A3(n30), .ZN(n108) );
endmodule



    module dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 ( 
        Clk, Rst, IR_IN, IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, 
        RegB_LATCH_EN, RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
        EQ_COND, .ALU_OPCODE({\ALU_OPCODE[5] , \ALU_OPCODE[4] , 
        \ALU_OPCODE[3] , \ALU_OPCODE[2] , \ALU_OPCODE[1] , \ALU_OPCODE[0] }), 
        signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
        WB_MUX_SEL, RF_WE, lhi_sel, sb_op, s_trap, s_ret );
  input [31:0] IR_IN;
  input Clk, Rst;
  output IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN,
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND,
         \ALU_OPCODE[5] , \ALU_OPCODE[4] , \ALU_OPCODE[3] , \ALU_OPCODE[2] ,
         \ALU_OPCODE[1] , \ALU_OPCODE[0] , signed_unsigned, DRAM_WE,
         LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, WB_MUX_SEL, RF_WE, lhi_sel, sb_op,
         s_trap, s_ret;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26, N40, N41,
         N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407,
         signed_unsigned_i, N717, N718, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n424, n425, n426, n428, n429, n430, n431, n432, n433,
         n434, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n532, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n183,
         n184, n200, n217, n218, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n419, n420, n421, n422, n423, n427, n435, n499, n500, n503, n504,
         n505, n506, n507, n509, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980;
  wire   [5:0] ALU_OPCODE;
  wire   [5:0] aluOpcode1;
  wire   [5:0] aluOpcode2;
  wire   [31:0] iterator_trap;
  wire   [31:0] iterator_ret;
  wire   [31:0] iterator1;
  wire   [31:0] iterator2;
  wire   [5:0] aluOpcode_i;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];
  assign IR_LATCH_EN = 1'b0;
  assign NPC_LATCH_EN = 1'b0;
  assign RegA_LATCH_EN = 1'b0;
  assign RegB_LATCH_EN = 1'b0;
  assign RegIMM_LATCH_EN = 1'b0;
  assign MUXA_SEL = 1'b0;
  assign MUXB_SEL = 1'b0;
  assign ALU_OUTREG_EN = 1'b0;
  assign EQ_COND = 1'b0;
  assign DRAM_WE = 1'b0;
  assign LMD_LATCH_EN = 1'b0;
  assign JUMP_EN = 1'b0;
  assign PC_LATCH_EN = 1'b0;
  assign WB_MUX_SEL = 1'b0;
  assign RF_WE = 1'b0;

  DFFR_X1 \aluOpcode1_reg[5]  ( .D(aluOpcode_i[5]), .CK(Clk), .RN(n774), .Q(
        aluOpcode1[5]) );
  DFFR_X1 \aluOpcode1_reg[4]  ( .D(n565), .CK(Clk), .RN(Rst), .Q(aluOpcode1[4]) );
  DFFR_X1 \aluOpcode1_reg[3]  ( .D(aluOpcode_i[3]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[3]) );
  DFFR_X1 \aluOpcode1_reg[2]  ( .D(aluOpcode_i[2]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[2]) );
  DFFR_X1 \aluOpcode1_reg[1]  ( .D(aluOpcode_i[1]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode1[1]) );
  DFFR_X1 \aluOpcode1_reg[0]  ( .D(aluOpcode_i[0]), .CK(Clk), .RN(n774), .Q(
        aluOpcode1[0]) );
  DFFR_X1 \aluOpcode2_reg[5]  ( .D(aluOpcode1[5]), .CK(Clk), .RN(n774), .Q(
        aluOpcode2[5]) );
  DFFR_X1 \aluOpcode2_reg[4]  ( .D(aluOpcode1[4]), .CK(Clk), .RN(n774), .Q(
        aluOpcode2[4]) );
  DFFR_X1 \aluOpcode2_reg[3]  ( .D(aluOpcode1[3]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[3]) );
  DFFR_X1 \aluOpcode2_reg[2]  ( .D(aluOpcode1[2]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[2]) );
  DFFR_X1 \aluOpcode2_reg[1]  ( .D(aluOpcode1[1]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[1]) );
  DFFR_X1 \aluOpcode2_reg[0]  ( .D(aluOpcode1[0]), .CK(Clk), .RN(Rst), .Q(
        aluOpcode2[0]) );
  DFFR_X1 \aluOpcode3_reg[4]  ( .D(aluOpcode2[4]), .CK(Clk), .RN(n774), .Q(
        ALU_OPCODE[4]) );
  DFFR_X1 \aluOpcode3_reg[3]  ( .D(aluOpcode2[3]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[3]) );
  DFFR_X1 \aluOpcode3_reg[2]  ( .D(aluOpcode2[2]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[2]) );
  DFFR_X1 \aluOpcode3_reg[1]  ( .D(aluOpcode2[1]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[1]) );
  DFFR_X1 \aluOpcode3_reg[0]  ( .D(aluOpcode2[0]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[0]) );
  DFF_X1 \iterator_trap_reg[0]  ( .D(n507), .CK(Clk), .Q(iterator_trap[0]), 
        .QN(n323) );
  DFF_X1 s_trap_reg ( .D(n434), .CK(Clk), .Q(s_trap), .QN(n424) );
  DFF_X1 \iterator_trap_reg[30]  ( .D(n465), .CK(Clk), .Q(iterator_trap[30]), 
        .QN(n353) );
  DFF_X1 \iterator_trap_reg[29]  ( .D(n464), .CK(Clk), .Q(iterator_trap[29]), 
        .QN(n352) );
  DFF_X1 \iterator_trap_reg[28]  ( .D(n463), .CK(Clk), .Q(iterator_trap[28]), 
        .QN(n351) );
  DFF_X1 \iterator_trap_reg[27]  ( .D(n462), .CK(Clk), .Q(iterator_trap[27]), 
        .QN(n350) );
  DFF_X1 \iterator_trap_reg[26]  ( .D(n461), .CK(Clk), .Q(iterator_trap[26]), 
        .QN(n349) );
  DFF_X1 \iterator_trap_reg[25]  ( .D(n460), .CK(Clk), .Q(iterator_trap[25]), 
        .QN(n348) );
  DFF_X1 \iterator_trap_reg[24]  ( .D(n459), .CK(Clk), .Q(iterator_trap[24]), 
        .QN(n347) );
  DFF_X1 \iterator_trap_reg[23]  ( .D(n458), .CK(Clk), .Q(iterator_trap[23]), 
        .QN(n346) );
  DFF_X1 \iterator_trap_reg[22]  ( .D(n457), .CK(Clk), .Q(iterator_trap[22]), 
        .QN(n345) );
  DFF_X1 \iterator_trap_reg[21]  ( .D(n456), .CK(Clk), .Q(iterator_trap[21]), 
        .QN(n344) );
  DFF_X1 \iterator_trap_reg[20]  ( .D(n455), .CK(Clk), .Q(iterator_trap[20]), 
        .QN(n343) );
  DFF_X1 \iterator_trap_reg[19]  ( .D(n454), .CK(Clk), .Q(iterator_trap[19]), 
        .QN(n342) );
  DFF_X1 \iterator_trap_reg[18]  ( .D(n453), .CK(Clk), .Q(iterator_trap[18]), 
        .QN(n341) );
  DFF_X1 \iterator_trap_reg[17]  ( .D(n452), .CK(Clk), .Q(iterator_trap[17]), 
        .QN(n340) );
  DFF_X1 \iterator_trap_reg[16]  ( .D(n451), .CK(Clk), .Q(iterator_trap[16]), 
        .QN(n339) );
  DFF_X1 \iterator_trap_reg[15]  ( .D(n450), .CK(Clk), .Q(iterator_trap[15]), 
        .QN(n338) );
  DFF_X1 \iterator_trap_reg[14]  ( .D(n449), .CK(Clk), .Q(iterator_trap[14]), 
        .QN(n337) );
  DFF_X1 \iterator_trap_reg[13]  ( .D(n448), .CK(Clk), .Q(iterator_trap[13]), 
        .QN(n336) );
  DFF_X1 \iterator_trap_reg[12]  ( .D(n447), .CK(Clk), .Q(iterator_trap[12]), 
        .QN(n335) );
  DFF_X1 \iterator_trap_reg[11]  ( .D(n446), .CK(Clk), .Q(iterator_trap[11]), 
        .QN(n334) );
  DFF_X1 \iterator_trap_reg[10]  ( .D(n445), .CK(Clk), .Q(iterator_trap[10]), 
        .QN(n333) );
  DFF_X1 \iterator_trap_reg[9]  ( .D(n444), .CK(Clk), .Q(iterator_trap[9]), 
        .QN(n332) );
  DFF_X1 \iterator_trap_reg[8]  ( .D(n443), .CK(Clk), .Q(iterator_trap[8]), 
        .QN(n331) );
  DFF_X1 \iterator_trap_reg[7]  ( .D(n442), .CK(Clk), .Q(iterator_trap[7]), 
        .QN(n330) );
  DFF_X1 \iterator_trap_reg[6]  ( .D(n441), .CK(Clk), .Q(iterator_trap[6]), 
        .QN(n329) );
  DFF_X1 \iterator_trap_reg[5]  ( .D(n440), .CK(Clk), .Q(iterator_trap[5]), 
        .QN(n328) );
  DFF_X1 \iterator_trap_reg[4]  ( .D(n439), .CK(Clk), .Q(iterator_trap[4]), 
        .QN(n327) );
  DFF_X1 \iterator_trap_reg[3]  ( .D(n438), .CK(Clk), .Q(iterator_trap[3]), 
        .QN(n326) );
  DFF_X1 \iterator_trap_reg[2]  ( .D(n437), .CK(Clk), .Q(iterator_trap[2]), 
        .QN(n325) );
  DFF_X1 \iterator_trap_reg[1]  ( .D(n436), .CK(Clk), .Q(iterator_trap[1]), 
        .QN(n324) );
  DFF_X1 \iterator_trap_reg[31]  ( .D(n466), .CK(Clk), .Q(iterator_trap[31]), 
        .QN(n354) );
  DFF_X1 \iterator_ret_reg[0]  ( .D(n467), .CK(Clk), .Q(iterator_ret[0]), .QN(
        n355) );
  DFF_X1 s_ret_reg ( .D(n433), .CK(Clk), .Q(s_ret), .QN(n425) );
  DFF_X1 \iterator_ret_reg[30]  ( .D(n497), .CK(Clk), .Q(iterator_ret[30]), 
        .QN(n385) );
  DFF_X1 \iterator_ret_reg[29]  ( .D(n496), .CK(Clk), .Q(iterator_ret[29]), 
        .QN(n384) );
  DFF_X1 \iterator_ret_reg[28]  ( .D(n495), .CK(Clk), .Q(iterator_ret[28]), 
        .QN(n383) );
  DFF_X1 \iterator_ret_reg[27]  ( .D(n494), .CK(Clk), .Q(iterator_ret[27]), 
        .QN(n382) );
  DFF_X1 \iterator_ret_reg[26]  ( .D(n493), .CK(Clk), .Q(iterator_ret[26]), 
        .QN(n381) );
  DFF_X1 \iterator_ret_reg[25]  ( .D(n492), .CK(Clk), .Q(iterator_ret[25]), 
        .QN(n380) );
  DFF_X1 \iterator_ret_reg[24]  ( .D(n491), .CK(Clk), .Q(iterator_ret[24]), 
        .QN(n379) );
  DFF_X1 \iterator_ret_reg[23]  ( .D(n490), .CK(Clk), .Q(iterator_ret[23]), 
        .QN(n378) );
  DFF_X1 \iterator_ret_reg[22]  ( .D(n489), .CK(Clk), .Q(iterator_ret[22]), 
        .QN(n377) );
  DFF_X1 \iterator_ret_reg[21]  ( .D(n488), .CK(Clk), .Q(iterator_ret[21]), 
        .QN(n376) );
  DFF_X1 \iterator_ret_reg[20]  ( .D(n487), .CK(Clk), .Q(iterator_ret[20]), 
        .QN(n375) );
  DFF_X1 \iterator_ret_reg[19]  ( .D(n486), .CK(Clk), .Q(iterator_ret[19]), 
        .QN(n374) );
  DFF_X1 \iterator_ret_reg[18]  ( .D(n485), .CK(Clk), .Q(iterator_ret[18]), 
        .QN(n373) );
  DFF_X1 \iterator_ret_reg[17]  ( .D(n484), .CK(Clk), .Q(iterator_ret[17]), 
        .QN(n372) );
  DFF_X1 \iterator_ret_reg[16]  ( .D(n483), .CK(Clk), .Q(iterator_ret[16]), 
        .QN(n371) );
  DFF_X1 \iterator_ret_reg[15]  ( .D(n482), .CK(Clk), .Q(iterator_ret[15]), 
        .QN(n370) );
  DFF_X1 \iterator_ret_reg[14]  ( .D(n481), .CK(Clk), .Q(iterator_ret[14]), 
        .QN(n369) );
  DFF_X1 \iterator_ret_reg[13]  ( .D(n480), .CK(Clk), .Q(iterator_ret[13]), 
        .QN(n368) );
  DFF_X1 \iterator_ret_reg[12]  ( .D(n479), .CK(Clk), .Q(iterator_ret[12]), 
        .QN(n367) );
  DFF_X1 \iterator_ret_reg[11]  ( .D(n478), .CK(Clk), .Q(iterator_ret[11]), 
        .QN(n366) );
  DFF_X1 \iterator_ret_reg[10]  ( .D(n477), .CK(Clk), .Q(iterator_ret[10]), 
        .QN(n365) );
  DFF_X1 \iterator_ret_reg[9]  ( .D(n476), .CK(Clk), .Q(iterator_ret[9]), .QN(
        n364) );
  DFF_X1 \iterator_ret_reg[8]  ( .D(n475), .CK(Clk), .Q(iterator_ret[8]), .QN(
        n363) );
  DFF_X1 \iterator_ret_reg[7]  ( .D(n474), .CK(Clk), .Q(iterator_ret[7]), .QN(
        n362) );
  DFF_X1 \iterator_ret_reg[6]  ( .D(n473), .CK(Clk), .Q(iterator_ret[6]), .QN(
        n361) );
  DFF_X1 \iterator_ret_reg[5]  ( .D(n472), .CK(Clk), .Q(iterator_ret[5]), .QN(
        n360) );
  DFF_X1 \iterator_ret_reg[4]  ( .D(n471), .CK(Clk), .Q(iterator_ret[4]), .QN(
        n359) );
  DFF_X1 \iterator_ret_reg[3]  ( .D(n470), .CK(Clk), .Q(iterator_ret[3]), .QN(
        n358) );
  DFF_X1 \iterator_ret_reg[2]  ( .D(n469), .CK(Clk), .Q(iterator_ret[2]), .QN(
        n357) );
  DFF_X1 \iterator_ret_reg[1]  ( .D(n468), .CK(Clk), .Q(iterator_ret[1]), .QN(
        n356) );
  DFF_X1 \iterator_ret_reg[31]  ( .D(n498), .CK(Clk), .Q(iterator_ret[31]), 
        .QN(n386) );
  DFF_X1 \iterator1_reg[0]  ( .D(n612), .CK(Clk), .Q(iterator1[0]), .QN(n513)
         );
  DFF_X1 \iterator1_reg[30]  ( .D(n582), .CK(Clk), .Q(iterator1[30]), .QN(n579) );
  DFF_X1 \iterator1_reg[29]  ( .D(n583), .CK(Clk), .Q(iterator1[29]), .QN(n578) );
  DFF_X1 \iterator1_reg[28]  ( .D(n584), .CK(Clk), .Q(iterator1[28]), .QN(n577) );
  DFF_X1 \iterator1_reg[27]  ( .D(n585), .CK(Clk), .Q(iterator1[27]), .QN(n576) );
  DFF_X1 \iterator1_reg[26]  ( .D(n586), .CK(Clk), .Q(iterator1[26]), .QN(n575) );
  DFF_X1 \iterator1_reg[25]  ( .D(n587), .CK(Clk), .Q(iterator1[25]), .QN(n574) );
  DFF_X1 \iterator1_reg[24]  ( .D(n588), .CK(Clk), .Q(iterator1[24]), .QN(n573) );
  DFF_X1 \iterator1_reg[23]  ( .D(n589), .CK(Clk), .Q(iterator1[23]), .QN(n572) );
  DFF_X1 \iterator1_reg[22]  ( .D(n590), .CK(Clk), .Q(iterator1[22]), .QN(n571) );
  DFF_X1 \iterator1_reg[21]  ( .D(n591), .CK(Clk), .Q(iterator1[21]), .QN(n570) );
  DFF_X1 \iterator1_reg[20]  ( .D(n592), .CK(Clk), .Q(iterator1[20]), .QN(n569) );
  DFF_X1 \iterator1_reg[19]  ( .D(n593), .CK(Clk), .Q(iterator1[19]), .QN(n568) );
  DFF_X1 \iterator1_reg[18]  ( .D(n594), .CK(Clk), .Q(iterator1[18]), .QN(n531) );
  DFF_X1 \iterator1_reg[17]  ( .D(n595), .CK(Clk), .Q(iterator1[17]), .QN(n530) );
  DFF_X1 \iterator1_reg[16]  ( .D(n596), .CK(Clk), .Q(iterator1[16]), .QN(n529) );
  DFF_X1 \iterator1_reg[15]  ( .D(n597), .CK(Clk), .Q(iterator1[15]), .QN(n528) );
  DFF_X1 \iterator1_reg[14]  ( .D(n598), .CK(Clk), .Q(iterator1[14]), .QN(n527) );
  DFF_X1 \iterator1_reg[13]  ( .D(n599), .CK(Clk), .Q(iterator1[13]), .QN(n526) );
  DFF_X1 \iterator1_reg[12]  ( .D(n600), .CK(Clk), .Q(iterator1[12]), .QN(n525) );
  DFF_X1 \iterator1_reg[11]  ( .D(n601), .CK(Clk), .Q(iterator1[11]), .QN(n524) );
  DFF_X1 \iterator1_reg[10]  ( .D(n602), .CK(Clk), .Q(iterator1[10]), .QN(n523) );
  DFF_X1 \iterator1_reg[9]  ( .D(n603), .CK(Clk), .Q(iterator1[9]), .QN(n522)
         );
  DFF_X1 \iterator1_reg[8]  ( .D(n604), .CK(Clk), .Q(iterator1[8]), .QN(n521)
         );
  DFF_X1 \iterator1_reg[7]  ( .D(n605), .CK(Clk), .Q(iterator1[7]), .QN(n520)
         );
  DFF_X1 \iterator1_reg[6]  ( .D(n606), .CK(Clk), .Q(iterator1[6]), .QN(n519)
         );
  DFF_X1 \iterator1_reg[5]  ( .D(n607), .CK(Clk), .Q(iterator1[5]), .QN(n518)
         );
  DFF_X1 \iterator1_reg[4]  ( .D(n608), .CK(Clk), .Q(iterator1[4]), .QN(n517)
         );
  DFF_X1 \iterator1_reg[3]  ( .D(n609), .CK(Clk), .Q(iterator1[3]), .QN(n516)
         );
  DFF_X1 \iterator1_reg[2]  ( .D(n610), .CK(Clk), .Q(iterator1[2]), .QN(n515)
         );
  DFF_X1 \iterator1_reg[1]  ( .D(n611), .CK(Clk), .Q(iterator1[1]), .QN(n514)
         );
  DFF_X1 \iterator1_reg[31]  ( .D(n581), .CK(Clk), .Q(iterator1[31]), .QN(n580) );
  DFF_X1 \iterator2_reg[0]  ( .D(n509), .CK(Clk), .Q(iterator2[0]), .QN(n387)
         );
  DFF_X1 sig3_reg ( .D(n532), .CK(Clk), .Q(n503) );
  DFF_X1 \iterator2_reg[30]  ( .D(n563), .CK(Clk), .Q(iterator2[30]), .QN(n417) );
  DFF_X1 \iterator2_reg[29]  ( .D(n562), .CK(Clk), .Q(iterator2[29]), .QN(n416) );
  DFF_X1 \iterator2_reg[28]  ( .D(n561), .CK(Clk), .Q(iterator2[28]), .QN(n415) );
  DFF_X1 \iterator2_reg[27]  ( .D(n560), .CK(Clk), .Q(iterator2[27]), .QN(n414) );
  DFF_X1 \iterator2_reg[26]  ( .D(n559), .CK(Clk), .Q(iterator2[26]), .QN(n413) );
  DFF_X1 \iterator2_reg[25]  ( .D(n558), .CK(Clk), .Q(iterator2[25]), .QN(n412) );
  DFF_X1 \iterator2_reg[24]  ( .D(n557), .CK(Clk), .Q(iterator2[24]), .QN(n411) );
  DFF_X1 \iterator2_reg[23]  ( .D(n556), .CK(Clk), .Q(iterator2[23]), .QN(n410) );
  DFF_X1 \iterator2_reg[22]  ( .D(n555), .CK(Clk), .Q(iterator2[22]), .QN(n409) );
  DFF_X1 \iterator2_reg[21]  ( .D(n554), .CK(Clk), .Q(iterator2[21]), .QN(n408) );
  DFF_X1 \iterator2_reg[20]  ( .D(n553), .CK(Clk), .Q(iterator2[20]), .QN(n407) );
  DFF_X1 \iterator2_reg[19]  ( .D(n552), .CK(Clk), .Q(iterator2[19]), .QN(n406) );
  DFF_X1 \iterator2_reg[18]  ( .D(n551), .CK(Clk), .Q(iterator2[18]), .QN(n405) );
  DFF_X1 \iterator2_reg[17]  ( .D(n550), .CK(Clk), .Q(iterator2[17]), .QN(n404) );
  DFF_X1 \iterator2_reg[16]  ( .D(n549), .CK(Clk), .Q(iterator2[16]), .QN(n403) );
  DFF_X1 \iterator2_reg[15]  ( .D(n548), .CK(Clk), .Q(iterator2[15]), .QN(n402) );
  DFF_X1 \iterator2_reg[14]  ( .D(n547), .CK(Clk), .Q(iterator2[14]), .QN(n401) );
  DFF_X1 \iterator2_reg[13]  ( .D(n546), .CK(Clk), .Q(iterator2[13]), .QN(n400) );
  DFF_X1 \iterator2_reg[12]  ( .D(n545), .CK(Clk), .Q(iterator2[12]), .QN(n399) );
  DFF_X1 \iterator2_reg[11]  ( .D(n544), .CK(Clk), .Q(iterator2[11]), .QN(n398) );
  DFF_X1 \iterator2_reg[10]  ( .D(n543), .CK(Clk), .Q(iterator2[10]), .QN(n397) );
  DFF_X1 \iterator2_reg[9]  ( .D(n542), .CK(Clk), .Q(iterator2[9]), .QN(n396)
         );
  DFF_X1 \iterator2_reg[8]  ( .D(n541), .CK(Clk), .Q(iterator2[8]), .QN(n395)
         );
  DFF_X1 \iterator2_reg[7]  ( .D(n540), .CK(Clk), .Q(iterator2[7]), .QN(n394)
         );
  DFF_X1 \iterator2_reg[6]  ( .D(n539), .CK(Clk), .Q(iterator2[6]), .QN(n393)
         );
  DFF_X1 \iterator2_reg[5]  ( .D(n538), .CK(Clk), .Q(iterator2[5]), .QN(n392)
         );
  DFF_X1 \iterator2_reg[4]  ( .D(n537), .CK(Clk), .Q(iterator2[4]), .QN(n391)
         );
  DFF_X1 \iterator2_reg[3]  ( .D(n536), .CK(Clk), .Q(iterator2[3]), .QN(n390)
         );
  DFF_X1 \iterator2_reg[2]  ( .D(n535), .CK(Clk), .Q(iterator2[2]), .QN(n389)
         );
  DFF_X1 \iterator2_reg[1]  ( .D(n534), .CK(Clk), .Q(iterator2[1]), .QN(n388)
         );
  DFF_X1 sb_op_reg ( .D(n431), .CK(Clk), .Q(sb_op), .QN(n426) );
  DFF_X1 \iterator2_reg[31]  ( .D(n564), .CK(Clk), .Q(iterator2[31]), .QN(n418) );
  DLH_X1 signed_unsigned_i_reg ( .G(N717), .D(N718), .Q(signed_unsigned_i) );
  DFF_X1 signed_unsigned_1_reg ( .D(n430), .CK(Clk), .QN(n504) );
  DFF_X1 signed_unsigned_2_reg ( .D(n429), .CK(Clk), .QN(n505) );
  DFF_X1 signed_unsigned_3_reg ( .D(n428), .CK(Clk), .Q(signed_unsigned), .QN(
        n506) );
  NOR4_X2 U235 ( .A1(n976), .A2(n980), .A3(IR_IN_29), .A4(IR_IN_31), .ZN(n244)
         );
  NOR4_X2 U277 ( .A1(IR_IN[6]), .A2(IR_IN[10]), .A3(n307), .A4(n499), .ZN(n245) );
  NAND3_X1 U463 ( .A1(n241), .A2(n242), .A3(n243), .ZN(aluOpcode_i[5]) );
  NAND3_X1 U479 ( .A1(n263), .A2(n950), .A3(n264), .ZN(aluOpcode_i[2]) );
  NAND3_X1 U480 ( .A1(n239), .A2(n971), .A3(n277), .ZN(n270) );
  NAND3_X1 U481 ( .A1(n291), .A2(n200), .A3(n217), .ZN(n290) );
  NAND3_X1 U482 ( .A1(n248), .A2(n954), .A3(n268), .ZN(n299) );
  NAND3_X1 U483 ( .A1(n217), .A2(n303), .A3(n281), .ZN(n294) );
  NAND3_X1 U484 ( .A1(n304), .A2(n963), .A3(n305), .ZN(N718) );
  NAND3_X1 U485 ( .A1(n256), .A2(n242), .A3(n314), .ZN(n309) );
  NAND3_X1 U486 ( .A1(n976), .A2(n980), .A3(n320), .ZN(n255) );
  NAND3_X1 U487 ( .A1(n955), .A2(n957), .A3(n322), .ZN(n268) );
  NAND3_X1 U488 ( .A1(n322), .A2(n957), .A3(IR_IN[2]), .ZN(n259) );
  NAND3_X1 U490 ( .A1(n976), .A2(n980), .A3(IR_IN_31), .ZN(n319) );
  NAND3_X1 U491 ( .A1(n979), .A2(n980), .A3(IR_IN_28), .ZN(n292) );
  NAND3_X1 U492 ( .A1(n320), .A2(n980), .A3(IR_IN_28), .ZN(n217) );
  NAND3_X1 U493 ( .A1(n322), .A2(n955), .A3(IR_IN[3]), .ZN(n248) );
  NAND3_X1 U494 ( .A1(n308), .A2(n980), .A3(n289), .ZN(n307) );
  NAND3_X1 U495 ( .A1(IR_IN_30), .A2(n976), .A3(n320), .ZN(n281) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 add_217 ( 
        .A(iterator_trap), .SUM({N71, N70, N69, N68, N67, N66, N65, N64, N63, 
        N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, 
        N48, N47, N46, N45, N44, N43, N42, N41, N40}) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 add_236 ( 
        .A(iterator_ret), .SUM({N182, N181, N180, N179, N178, N177, N176, N175, 
        N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151}) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_6 add_277 ( 
        .A(iterator2), .SUM({N407, N406, N405, N404, N403, N402, N401, N400, 
        N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, 
        N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376}) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_7 add_256 ( 
        .A(iterator1), .SUM({N294, N293, N292, N291, N290, N289, N288, N287, 
        N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, 
        N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263}) );
  DFFR_X1 \aluOpcode3_reg[5]  ( .D(aluOpcode2[5]), .CK(Clk), .RN(Rst), .Q(
        ALU_OPCODE[5]) );
  DFF_X1 sig1_reg ( .D(n567), .CK(Clk), .QN(n941) );
  DFF_X1 sig2_reg ( .D(n566), .CK(Clk), .QN(n897) );
  DFF_X1 sig4_reg ( .D(n613), .CK(Clk), .QN(n860) );
  DFF_X1 lhi_sel_reg ( .D(n432), .CK(Clk), .Q(lhi_sel), .QN(n773) );
  AND2_X1 U3 ( .A1(n826), .A2(n759), .ZN(n614) );
  INV_X1 U4 ( .A(n614), .ZN(n615) );
  INV_X1 U5 ( .A(n708), .ZN(n616) );
  INV_X1 U6 ( .A(n705), .ZN(n617) );
  AND3_X1 U7 ( .A1(n618), .A2(n619), .A3(n620), .ZN(n904) );
  AND4_X1 U8 ( .A1(n903), .A2(n912), .A3(n911), .A4(n913), .ZN(n618) );
  AND4_X1 U9 ( .A1(n921), .A2(n920), .A3(n919), .A4(n918), .ZN(n619) );
  AND4_X1 U10 ( .A1(n925), .A2(n924), .A3(n923), .A4(n922), .ZN(n620) );
  AND2_X1 U11 ( .A1(n635), .A2(n771), .ZN(n621) );
  BUF_X1 U12 ( .A(n816), .Z(n755) );
  INV_X1 U13 ( .A(N389), .ZN(n797) );
  BUF_X1 U14 ( .A(n816), .Z(n754) );
  BUF_X1 U15 ( .A(n816), .Z(n753) );
  BUF_X1 U16 ( .A(n625), .Z(n758) );
  BUF_X1 U17 ( .A(n625), .Z(n756) );
  BUF_X2 U18 ( .A(n899), .Z(n731) );
  BUF_X1 U19 ( .A(n942), .Z(n771) );
  INV_X1 U20 ( .A(N50), .ZN(n918) );
  BUF_X1 U21 ( .A(n942), .Z(n770) );
  INV_X1 U22 ( .A(N60), .ZN(n928) );
  INV_X1 U23 ( .A(n713), .ZN(n622) );
  INV_X1 U24 ( .A(n715), .ZN(n623) );
  INV_X1 U25 ( .A(n747), .ZN(n624) );
  AND2_X1 U26 ( .A1(n818), .A2(n774), .ZN(n625) );
  AND2_X1 U27 ( .A1(N41), .A2(n717), .ZN(n626) );
  AND3_X1 U28 ( .A1(N378), .A2(N377), .A3(N376), .ZN(n627) );
  BUF_X1 U29 ( .A(n942), .Z(n769) );
  OR2_X1 U30 ( .A1(N164), .A2(N167), .ZN(n628) );
  AND2_X1 U31 ( .A1(n839), .A2(n841), .ZN(n629) );
  MUX2_X1 U32 ( .A(n768), .B(n900), .S(n639), .Z(n467) );
  BUF_X1 U33 ( .A(n631), .Z(n636) );
  AND2_X1 U34 ( .A1(n908), .A2(n771), .ZN(n630) );
  BUF_X1 U35 ( .A(n647), .Z(n631) );
  CLKBUF_X1 U36 ( .A(N172), .Z(n632) );
  INV_X1 U37 ( .A(N182), .ZN(n633) );
  CLKBUF_X1 U38 ( .A(N173), .Z(n634) );
  NAND2_X1 U39 ( .A1(n744), .A2(n626), .ZN(n635) );
  AND4_X2 U40 ( .A1(n905), .A2(n904), .A3(n907), .A4(n906), .ZN(n744) );
  NAND3_X1 U41 ( .A1(n842), .A2(n840), .A3(n629), .ZN(n820) );
  OR2_X1 U42 ( .A1(N277), .A2(N279), .ZN(n637) );
  OR2_X1 U43 ( .A1(N58), .A2(N60), .ZN(n638) );
  INV_X1 U44 ( .A(n355), .ZN(n639) );
  CLKBUF_X1 U45 ( .A(N175), .Z(n640) );
  AND4_X1 U46 ( .A1(n641), .A2(n876), .A3(n642), .A4(n643), .ZN(n864) );
  INV_X1 U47 ( .A(N160), .ZN(n641) );
  INV_X1 U48 ( .A(N162), .ZN(n642) );
  INV_X1 U49 ( .A(N163), .ZN(n643) );
  OAI22_X1 U50 ( .A1(n660), .A2(n797), .B1(n754), .B2(n400), .ZN(n546) );
  OAI22_X1 U51 ( .A1(n660), .A2(n809), .B1(n753), .B2(n412), .ZN(n558) );
  OAI22_X1 U52 ( .A1(n700), .A2(n928), .B1(n769), .B2(n343), .ZN(n455) );
  OAI22_X1 U53 ( .A1(n700), .A2(n918), .B1(n770), .B2(n333), .ZN(n445) );
  OAI22_X1 U54 ( .A1(n696), .A2(n857), .B1(n756), .B2(n577), .ZN(n584) );
  INV_X2 U55 ( .A(N291), .ZN(n857) );
  OAI22_X1 U56 ( .A1(n671), .A2(n837), .B1(n758), .B2(n521), .ZN(n604) );
  OAI22_X1 U57 ( .A1(n719), .A2(n786), .B1(n755), .B2(n389), .ZN(n535) );
  INV_X2 U58 ( .A(N378), .ZN(n786) );
  OAI22_X1 U59 ( .A1(n695), .A2(n909), .B1(n771), .B2(n354), .ZN(n466) );
  CLKBUF_X1 U60 ( .A(N285), .Z(n644) );
  AND2_X1 U61 ( .A1(n908), .A2(n771), .ZN(n645) );
  BUF_X1 U62 ( .A(n631), .Z(n727) );
  CLKBUF_X1 U63 ( .A(N277), .Z(n646) );
  OAI21_X1 U64 ( .B1(n895), .B2(n639), .A(n763), .ZN(n647) );
  CLKBUF_X1 U65 ( .A(n883), .Z(n648) );
  CLKBUF_X1 U66 ( .A(N58), .Z(n649) );
  OR2_X1 U67 ( .A1(n783), .A2(n707), .ZN(n650) );
  NAND4_X1 U68 ( .A1(n884), .A2(n648), .A3(n882), .A4(n881), .ZN(n651) );
  OR2_X1 U69 ( .A1(n783), .A2(n707), .ZN(n781) );
  NOR2_X1 U70 ( .A1(n653), .A2(n654), .ZN(n652) );
  NAND4_X1 U71 ( .A1(n673), .A2(n800), .A3(n799), .A4(n798), .ZN(n653) );
  OR4_X2 U72 ( .A1(n777), .A2(N385), .A3(N384), .A4(N383), .ZN(n654) );
  AND4_X1 U73 ( .A1(n794), .A2(n795), .A3(n796), .A4(n797), .ZN(n673) );
  NOR3_X1 U74 ( .A1(N166), .A2(N165), .A3(n628), .ZN(n865) );
  NOR3_X1 U75 ( .A1(n820), .A2(N278), .A3(n637), .ZN(n824) );
  INV_X1 U76 ( .A(n658), .ZN(n655) );
  CLKBUF_X1 U77 ( .A(N284), .Z(n656) );
  CLKBUF_X1 U78 ( .A(N177), .Z(n657) );
  AND2_X1 U79 ( .A1(n781), .A2(n755), .ZN(n658) );
  AND2_X1 U80 ( .A1(n650), .A2(n755), .ZN(n749) );
  BUF_X1 U81 ( .A(n631), .Z(n728) );
  CLKBUF_X1 U82 ( .A(n744), .Z(n659) );
  NOR2_X1 U83 ( .A1(N292), .A2(N291), .ZN(n720) );
  INV_X1 U84 ( .A(n704), .ZN(n660) );
  INV_X1 U85 ( .A(n704), .ZN(n718) );
  CLKBUF_X1 U86 ( .A(n690), .Z(n661) );
  INV_X1 U87 ( .A(n706), .ZN(n662) );
  OR2_X1 U88 ( .A1(n763), .A2(n897), .ZN(n663) );
  NAND2_X1 U89 ( .A1(n663), .A2(n636), .ZN(n566) );
  INV_X1 U90 ( .A(n768), .ZN(n767) );
  BUF_X1 U91 ( .A(n899), .Z(n664) );
  AND3_X1 U92 ( .A1(n742), .A2(n859), .A3(n720), .ZN(n665) );
  CLKBUF_X1 U93 ( .A(N397), .Z(n666) );
  OR2_X1 U94 ( .A1(N285), .A2(N284), .ZN(n667) );
  NAND2_X1 U95 ( .A1(n744), .A2(n626), .ZN(n908) );
  AND2_X1 U96 ( .A1(n864), .A2(n863), .ZN(n668) );
  AND2_X1 U97 ( .A1(n865), .A2(n668), .ZN(n680) );
  CLKBUF_X1 U98 ( .A(n665), .Z(n669) );
  AND4_X1 U99 ( .A1(n867), .A2(N153), .A3(n894), .A4(n893), .ZN(n670) );
  AND4_X1 U100 ( .A1(n894), .A2(n633), .A3(N153), .A4(n893), .ZN(n739) );
  NOR3_X1 U101 ( .A1(n902), .A2(N59), .A3(n638), .ZN(n905) );
  INV_X1 U102 ( .A(n614), .ZN(n671) );
  NOR2_X1 U103 ( .A1(N393), .A2(N396), .ZN(n672) );
  INV_X1 U104 ( .A(n749), .ZN(n674) );
  INV_X1 U105 ( .A(n658), .ZN(n675) );
  INV_X1 U106 ( .A(n748), .ZN(n676) );
  CLKBUF_X1 U107 ( .A(N398), .Z(n677) );
  NOR3_X1 U108 ( .A1(N173), .A2(N175), .A3(N172), .ZN(n698) );
  CLKBUF_X1 U109 ( .A(n686), .Z(n678) );
  CLKBUF_X1 U110 ( .A(N399), .Z(n679) );
  NAND3_X1 U111 ( .A1(n803), .A2(n802), .A3(n672), .ZN(n778) );
  NOR2_X1 U112 ( .A1(n661), .A2(n651), .ZN(n681) );
  OR2_X1 U113 ( .A1(n774), .A2(n773), .ZN(n682) );
  NAND2_X1 U114 ( .A1(n829), .A2(n682), .ZN(n432) );
  CLKBUF_X1 U115 ( .A(n783), .Z(n683) );
  AND2_X1 U116 ( .A1(n684), .A2(n685), .ZN(n779) );
  AND4_X1 U117 ( .A1(n808), .A2(n809), .A3(n810), .A4(n811), .ZN(n684) );
  NOR3_X1 U118 ( .A1(N405), .A2(N406), .A3(N404), .ZN(n685) );
  AND3_X1 U119 ( .A1(n823), .A2(n825), .A3(n824), .ZN(n686) );
  INV_X1 U120 ( .A(n748), .ZN(n687) );
  INV_X1 U121 ( .A(n658), .ZN(n688) );
  NOR3_X1 U122 ( .A1(n667), .A2(N286), .A3(n821), .ZN(n823) );
  NOR4_X1 U123 ( .A1(N176), .A2(N177), .A3(N178), .A4(N179), .ZN(n693) );
  AND2_X1 U124 ( .A1(n686), .A2(n665), .ZN(n689) );
  NOR2_X1 U125 ( .A1(n690), .A2(n691), .ZN(n722) );
  NAND2_X1 U126 ( .A1(n698), .A2(n887), .ZN(n690) );
  NAND4_X1 U127 ( .A1(n884), .A2(n883), .A3(n882), .A4(n881), .ZN(n691) );
  CLKBUF_X1 U128 ( .A(n887), .Z(n692) );
  AND4_X1 U129 ( .A1(n891), .A2(n892), .A3(n890), .A4(n889), .ZN(n738) );
  INV_X1 U130 ( .A(n747), .ZN(n694) );
  INV_X1 U131 ( .A(n706), .ZN(n695) );
  INV_X1 U132 ( .A(n715), .ZN(n696) );
  CLKBUF_X1 U133 ( .A(N286), .Z(n697) );
  NAND2_X1 U134 ( .A1(n689), .A2(n711), .ZN(n699) );
  INV_X1 U135 ( .A(n645), .ZN(n700) );
  NOR4_X1 U136 ( .A1(n778), .A2(N397), .A3(N398), .A4(N399), .ZN(n780) );
  AND3_X1 U137 ( .A1(n722), .A2(n739), .A3(n693), .ZN(n701) );
  INV_X1 U138 ( .A(n714), .ZN(n702) );
  OR2_X1 U139 ( .A1(n769), .A2(n941), .ZN(n703) );
  NAND2_X1 U140 ( .A1(n734), .A2(n703), .ZN(n567) );
  AND2_X1 U141 ( .A1(n755), .A2(n650), .ZN(n704) );
  NAND3_X1 U142 ( .A1(n779), .A2(n652), .A3(n780), .ZN(n783) );
  AND2_X1 U143 ( .A1(n635), .A2(n771), .ZN(n705) );
  AND2_X1 U144 ( .A1(n908), .A2(n771), .ZN(n706) );
  AND2_X1 U145 ( .A1(n635), .A2(n771), .ZN(n708) );
  NAND2_X1 U146 ( .A1(n782), .A2(n627), .ZN(n707) );
  AND2_X1 U147 ( .A1(n862), .A2(n680), .ZN(n709) );
  NAND2_X1 U148 ( .A1(n710), .A2(n711), .ZN(n826) );
  AND2_X1 U149 ( .A1(n686), .A2(n822), .ZN(n710) );
  NOR2_X1 U150 ( .A1(n723), .A2(N294), .ZN(n711) );
  CLKBUF_X1 U151 ( .A(N406), .Z(n712) );
  AND2_X1 U152 ( .A1(n699), .A2(n759), .ZN(n713) );
  AND2_X1 U153 ( .A1(n699), .A2(n759), .ZN(n714) );
  AND2_X1 U154 ( .A1(n826), .A2(n759), .ZN(n715) );
  INV_X1 U155 ( .A(n713), .ZN(n716) );
  INV_X1 U156 ( .A(n323), .ZN(n717) );
  INV_X1 U157 ( .A(n704), .ZN(n719) );
  INV_X1 U158 ( .A(n749), .ZN(n750) );
  INV_X1 U159 ( .A(n749), .ZN(n751) );
  AND3_X1 U160 ( .A1(n742), .A2(n859), .A3(n720), .ZN(n822) );
  OR2_X1 U161 ( .A1(n756), .A2(n860), .ZN(n721) );
  NAND2_X1 U162 ( .A1(n721), .A2(n741), .ZN(n613) );
  AND3_X1 U163 ( .A1(n670), .A2(n738), .A3(n681), .ZN(n862) );
  NAND3_X1 U164 ( .A1(N265), .A2(N264), .A3(N263), .ZN(n723) );
  NAND2_X1 U165 ( .A1(n669), .A2(n678), .ZN(n828) );
  NAND2_X1 U166 ( .A1(n701), .A2(n680), .ZN(n895) );
  INV_X1 U167 ( .A(n708), .ZN(n724) );
  INV_X1 U168 ( .A(n630), .ZN(n725) );
  BUF_X1 U169 ( .A(n898), .Z(n763) );
  BUF_X1 U170 ( .A(n898), .Z(n765) );
  BUF_X1 U171 ( .A(n898), .Z(n764) );
  OAI22_X1 U172 ( .A1(n962), .A2(n974), .B1(n968), .B2(n255), .ZN(n296) );
  INV_X1 U173 ( .A(n255), .ZN(n973) );
  NAND2_X1 U174 ( .A1(n968), .A2(n966), .ZN(n184) );
  INV_X1 U175 ( .A(n303), .ZN(n975) );
  NAND2_X1 U176 ( .A1(n962), .A2(n968), .ZN(n283) );
  INV_X1 U177 ( .A(n275), .ZN(n962) );
  NAND4_X1 U178 ( .A1(n963), .A2(n965), .A3(n945), .A4(n183), .ZN(n565) );
  NAND2_X1 U179 ( .A1(n977), .A2(n184), .ZN(n183) );
  AND3_X1 U180 ( .A1(n965), .A2(n262), .A3(n251), .ZN(n263) );
  INV_X1 U181 ( .A(n309), .ZN(n963) );
  INV_X1 U182 ( .A(n258), .ZN(n948) );
  INV_X1 U183 ( .A(n271), .ZN(n969) );
  BUF_X1 U184 ( .A(n625), .Z(n757) );
  AND2_X1 U185 ( .A1(n854), .A2(n853), .ZN(n726) );
  AOI211_X1 U186 ( .C1(n283), .C2(n972), .A(n960), .B(n423), .ZN(n241) );
  INV_X1 U187 ( .A(n304), .ZN(n960) );
  INV_X1 U188 ( .A(n281), .ZN(n972) );
  OAI21_X1 U189 ( .B1(n291), .B2(n968), .A(n239), .ZN(n423) );
  NOR2_X1 U190 ( .A1(n279), .A2(n257), .ZN(n267) );
  INV_X1 U191 ( .A(n775), .ZN(n774) );
  NOR2_X1 U192 ( .A1(n291), .A2(n218), .ZN(n280) );
  OAI21_X1 U193 ( .B1(n248), .B2(n302), .A(n284), .ZN(n258) );
  NAND2_X1 U194 ( .A1(n245), .A2(n435), .ZN(n262) );
  OAI22_X1 U195 ( .A1(n267), .A2(n248), .B1(n954), .B2(n247), .ZN(n435) );
  INV_X1 U196 ( .A(n245), .ZN(n959) );
  AOI21_X1 U197 ( .B1(n289), .B2(n978), .A(n427), .ZN(n251) );
  INV_X1 U198 ( .A(n280), .ZN(n971) );
  AOI22_X1 U199 ( .A1(n278), .A2(n279), .B1(n961), .B2(n975), .ZN(n277) );
  NOR2_X1 U200 ( .A1(n959), .A2(n259), .ZN(n278) );
  AOI221_X1 U201 ( .B1(n951), .B2(n298), .C1(n257), .C2(n299), .A(n300), .ZN(
        n297) );
  INV_X1 U202 ( .A(n247), .ZN(n951) );
  NOR4_X1 U203 ( .A1(n301), .A2(n958), .A3(n957), .A4(n302), .ZN(n300) );
  AOI211_X1 U204 ( .C1(n978), .C2(n266), .A(n280), .B(n315), .ZN(n314) );
  AOI21_X1 U205 ( .B1(n254), .B2(n968), .A(n974), .ZN(n315) );
  NOR2_X1 U206 ( .A1(n292), .A2(n964), .ZN(n427) );
  INV_X1 U207 ( .A(n184), .ZN(n964) );
  AOI21_X1 U208 ( .B1(n970), .B2(n975), .A(n288), .ZN(n242) );
  INV_X1 U209 ( .A(n217), .ZN(n978) );
  NAND4_X1 U210 ( .A1(n241), .A2(n945), .A3(n251), .A4(n949), .ZN(
        aluOpcode_i[3]) );
  INV_X1 U211 ( .A(n252), .ZN(n949) );
  OAI221_X1 U212 ( .B1(n959), .B2(n253), .C1(n254), .C2(n255), .A(n256), .ZN(
        n252) );
  AOI21_X1 U213 ( .B1(n257), .B2(n956), .A(n258), .ZN(n253) );
  OAI21_X1 U214 ( .B1(n966), .B2(n292), .A(n293), .ZN(n287) );
  INV_X1 U215 ( .A(n218), .ZN(n970) );
  INV_X1 U216 ( .A(n254), .ZN(n961) );
  AOI222_X1 U217 ( .A1(n244), .A2(n970), .B1(n245), .B2(n246), .C1(n977), .C2(
        n184), .ZN(n243) );
  OAI211_X1 U218 ( .C1(n247), .C2(n248), .A(n249), .B(n250), .ZN(n246) );
  NAND4_X1 U219 ( .A1(n263), .A2(n241), .A3(n310), .A4(n311), .ZN(N717) );
  AOI21_X1 U220 ( .B1(n245), .B2(n313), .A(n309), .ZN(n310) );
  NOR4_X1 U221 ( .A1(n978), .A2(n244), .A3(n973), .A4(n312), .ZN(n311) );
  NAND4_X1 U222 ( .A1(n946), .A2(n948), .A3(n268), .A4(n248), .ZN(n313) );
  NAND2_X1 U223 ( .A1(n254), .A2(n966), .ZN(n266) );
  INV_X1 U224 ( .A(n200), .ZN(n977) );
  NAND2_X1 U225 ( .A1(n944), .A2(n979), .ZN(n291) );
  NAND4_X1 U226 ( .A1(n271), .A2(n272), .A3(n273), .A4(n274), .ZN(
        aluOpcode_i[1]) );
  AOI22_X1 U227 ( .A1(n245), .A2(n282), .B1(n244), .B2(n283), .ZN(n273) );
  AOI211_X1 U228 ( .C1(n973), .C2(n275), .A(n276), .B(n270), .ZN(n274) );
  OAI211_X1 U229 ( .C1(n267), .C2(n248), .A(n284), .B(n947), .ZN(n282) );
  OR2_X1 U230 ( .A1(n259), .A2(n302), .ZN(n269) );
  INV_X1 U231 ( .A(n259), .ZN(n956) );
  NAND2_X1 U232 ( .A1(n254), .A2(n218), .ZN(n275) );
  NAND2_X1 U233 ( .A1(n289), .A2(n290), .ZN(n271) );
  INV_X1 U234 ( .A(n298), .ZN(n954) );
  INV_X1 U236 ( .A(n419), .ZN(n946) );
  OAI211_X1 U237 ( .C1(n267), .C2(n259), .A(n250), .B(n947), .ZN(n419) );
  INV_X1 U238 ( .A(n260), .ZN(n945) );
  OAI21_X1 U239 ( .B1(n261), .B2(n959), .A(n262), .ZN(n260) );
  INV_X1 U240 ( .A(n420), .ZN(n947) );
  OAI221_X1 U241 ( .B1(n268), .B2(n302), .C1(n267), .C2(n954), .A(n421), .ZN(
        n420) );
  AND2_X1 U242 ( .A1(n269), .A2(n249), .ZN(n421) );
  INV_X1 U243 ( .A(n270), .ZN(n950) );
  AOI222_X1 U244 ( .A1(n244), .A2(n970), .B1(n245), .B2(n265), .C1(n973), .C2(
        n266), .ZN(n264) );
  OAI21_X1 U245 ( .B1(n267), .B2(n268), .A(n269), .ZN(n265) );
  INV_X1 U246 ( .A(n500), .ZN(n965) );
  OAI211_X1 U247 ( .C1(n966), .C2(n281), .A(n293), .B(n272), .ZN(n500) );
  AOI221_X1 U248 ( .B1(n978), .B2(n289), .C1(n961), .C2(n977), .A(n306), .ZN(
        n305) );
  AOI21_X1 U249 ( .B1(n946), .B2(n261), .A(n307), .ZN(n306) );
  INV_X1 U250 ( .A(n244), .ZN(n974) );
  NAND2_X1 U251 ( .A1(n317), .A2(n976), .ZN(n303) );
  NAND2_X1 U252 ( .A1(n285), .A2(n286), .ZN(aluOpcode_i[0]) );
  AOI221_X1 U253 ( .B1(n961), .B2(n294), .C1(n245), .C2(n295), .A(n296), .ZN(
        n285) );
  NOR4_X1 U254 ( .A1(n287), .A2(n969), .A3(n288), .A4(n280), .ZN(n286) );
  NAND4_X1 U255 ( .A1(n261), .A2(n250), .A3(n269), .A4(n297), .ZN(n295) );
  AOI22_X1 U256 ( .A1(n316), .A2(n973), .B1(n318), .B2(n970), .ZN(n256) );
  OAI21_X1 U257 ( .B1(n979), .B2(n319), .A(n255), .ZN(n318) );
  OAI22_X1 U258 ( .A1(n218), .A2(n281), .B1(n966), .B2(n200), .ZN(n276) );
  OAI22_X1 U259 ( .A1(n505), .A2(n775), .B1(Rst), .B2(n506), .ZN(n428) );
  OAI22_X1 U260 ( .A1(n504), .A2(n775), .B1(n505), .B2(Rst), .ZN(n429) );
  OAI21_X1 U261 ( .B1(n504), .B2(Rst), .A(n240), .ZN(n430) );
  NAND2_X1 U262 ( .A1(signed_unsigned_i), .A2(Rst), .ZN(n240) );
  OR3_X1 U263 ( .A1(IR_IN[9]), .A2(IR_IN[8]), .A3(IR_IN[7]), .ZN(n499) );
  OAI211_X1 U264 ( .C1(n279), .C2(n321), .A(n322), .B(IR_IN[3]), .ZN(n284) );
  NOR2_X1 U265 ( .A1(n955), .A2(n302), .ZN(n321) );
  NOR3_X1 U266 ( .A1(n962), .A2(IR_IN_31), .A3(IR_IN_28), .ZN(n312) );
  NAND4_X1 U267 ( .A1(n257), .A2(n301), .A3(IR_IN[3]), .A4(IR_IN[5]), .ZN(n250) );
  NAND4_X1 U268 ( .A1(IR_IN_28), .A2(n320), .A3(n289), .A4(IR_IN_30), .ZN(n293) );
  NAND4_X1 U269 ( .A1(IR_IN_28), .A2(n320), .A3(n316), .A4(IR_IN_30), .ZN(n272) );
  NAND2_X1 U270 ( .A1(IR_IN_30), .A2(n308), .ZN(n200) );
  NAND4_X1 U271 ( .A1(IR_IN[4]), .A2(IR_IN[3]), .A3(n422), .A4(IR_IN[5]), .ZN(
        n249) );
  AOI22_X1 U272 ( .A1(IR_IN[2]), .A2(n302), .B1(n247), .B2(n955), .ZN(n422) );
  INV_X1 U273 ( .A(Rst), .ZN(n775) );
  NAND2_X1 U274 ( .A1(IR_IN[0]), .A2(n953), .ZN(n261) );
  INV_X1 U275 ( .A(n268), .ZN(n953) );
  AND3_X1 U276 ( .A1(IR_IN_28), .A2(n316), .A3(n317), .ZN(n288) );
  NOR2_X1 U278 ( .A1(IR_IN_26), .A2(IR_IN_27), .ZN(n289) );
  NAND2_X1 U279 ( .A1(IR_IN[0]), .A2(n952), .ZN(n302) );
  INV_X1 U280 ( .A(IR_IN[2]), .ZN(n955) );
  NAND2_X1 U281 ( .A1(IR_IN_27), .A2(n967), .ZN(n254) );
  NAND2_X1 U282 ( .A1(IR_IN_27), .A2(IR_IN_26), .ZN(n218) );
  INV_X1 U283 ( .A(IR_IN_30), .ZN(n980) );
  NAND2_X1 U284 ( .A1(IR_IN[1]), .A2(IR_IN[0]), .ZN(n247) );
  NOR2_X1 U285 ( .A1(n952), .A2(IR_IN[0]), .ZN(n257) );
  INV_X1 U286 ( .A(IR_IN_28), .ZN(n976) );
  NOR2_X1 U287 ( .A1(n979), .A2(IR_IN_31), .ZN(n320) );
  INV_X1 U288 ( .A(IR_IN_29), .ZN(n979) );
  NOR2_X1 U289 ( .A1(n967), .A2(IR_IN_27), .ZN(n316) );
  NOR2_X1 U290 ( .A1(IR_IN[1]), .A2(IR_IN[0]), .ZN(n279) );
  NOR2_X1 U291 ( .A1(n958), .A2(IR_IN[4]), .ZN(n322) );
  INV_X1 U292 ( .A(IR_IN[3]), .ZN(n957) );
  INV_X1 U293 ( .A(IR_IN_26), .ZN(n967) );
  INV_X1 U294 ( .A(IR_IN[1]), .ZN(n952) );
  INV_X1 U295 ( .A(IR_IN[5]), .ZN(n958) );
  AND2_X1 U296 ( .A1(IR_IN[4]), .A2(n955), .ZN(n301) );
  NOR4_X1 U297 ( .A1(n955), .A2(IR_IN[3]), .A3(IR_IN[4]), .A4(IR_IN[5]), .ZN(
        n298) );
  NOR3_X1 U298 ( .A1(IR_IN_29), .A2(IR_IN_31), .A3(IR_IN_28), .ZN(n308) );
  AOI22_X1 U299 ( .A1(n975), .A2(n961), .B1(IR_IN_31), .B2(n427), .ZN(n304) );
  AND3_X1 U300 ( .A1(IR_IN_31), .A2(IR_IN_30), .A3(IR_IN_29), .ZN(n317) );
  BUF_X1 U301 ( .A(n899), .Z(n729) );
  BUF_X1 U302 ( .A(n899), .Z(n730) );
  INV_X1 U303 ( .A(n630), .ZN(n732) );
  INV_X1 U304 ( .A(n708), .ZN(n733) );
  INV_X1 U305 ( .A(n645), .ZN(n734) );
  INV_X1 U306 ( .A(n705), .ZN(n735) );
  INV_X1 U307 ( .A(n705), .ZN(n736) );
  INV_X1 U308 ( .A(n621), .ZN(n737) );
  AND4_X1 U309 ( .A1(n937), .A2(n938), .A3(n909), .A4(N42), .ZN(n907) );
  INV_X1 U310 ( .A(n714), .ZN(n740) );
  INV_X1 U311 ( .A(n715), .ZN(n741) );
  INV_X1 U312 ( .A(n614), .ZN(n743) );
  INV_X1 U313 ( .A(n745), .ZN(n760) );
  INV_X1 U314 ( .A(n713), .ZN(n761) );
  INV_X1 U315 ( .A(n745), .ZN(n762) );
  AND2_X1 U316 ( .A1(n826), .A2(n759), .ZN(n747) );
  AND4_X1 U317 ( .A1(n933), .A2(n934), .A3(n935), .A4(n936), .ZN(n906) );
  AND3_X1 U318 ( .A1(n856), .A2(n855), .A3(n726), .ZN(n742) );
  AND2_X1 U319 ( .A1(n826), .A2(n759), .ZN(n745) );
  INV_X1 U320 ( .A(n513), .ZN(n746) );
  INV_X1 U321 ( .A(n658), .ZN(n752) );
  AND2_X1 U322 ( .A1(n781), .A2(n755), .ZN(n748) );
  INV_X1 U323 ( .A(n647), .ZN(n768) );
  CLKBUF_X1 U324 ( .A(n625), .Z(n759) );
  CLKBUF_X1 U325 ( .A(n898), .Z(n766) );
  INV_X1 U326 ( .A(n319), .ZN(n944) );
  NAND3_X1 U327 ( .A1(IR_IN_29), .A2(n289), .A3(n944), .ZN(n239) );
  INV_X1 U328 ( .A(n316), .ZN(n966) );
  INV_X1 U329 ( .A(n289), .ZN(n968) );
  INV_X1 U330 ( .A(n239), .ZN(n776) );
  OAI21_X1 U331 ( .B1(n503), .B2(n776), .A(n774), .ZN(n817) );
  INV_X1 U332 ( .A(n817), .ZN(n816) );
  INV_X1 U333 ( .A(N379), .ZN(n787) );
  INV_X1 U334 ( .A(N380), .ZN(n788) );
  INV_X1 U335 ( .A(N381), .ZN(n789) );
  INV_X1 U336 ( .A(N382), .ZN(n790) );
  NAND4_X1 U337 ( .A1(n787), .A2(n788), .A3(n789), .A4(n790), .ZN(n777) );
  INV_X1 U338 ( .A(N386), .ZN(n794) );
  INV_X1 U339 ( .A(N387), .ZN(n795) );
  INV_X1 U340 ( .A(N388), .ZN(n796) );
  INV_X1 U341 ( .A(N393), .ZN(n801) );
  INV_X1 U342 ( .A(N394), .ZN(n802) );
  INV_X1 U343 ( .A(N395), .ZN(n803) );
  INV_X1 U344 ( .A(N396), .ZN(n804) );
  INV_X1 U345 ( .A(N400), .ZN(n808) );
  INV_X1 U346 ( .A(N401), .ZN(n809) );
  INV_X1 U347 ( .A(N402), .ZN(n810) );
  INV_X1 U348 ( .A(N403), .ZN(n811) );
  INV_X1 U349 ( .A(N407), .ZN(n782) );
  OAI22_X1 U350 ( .A1(n676), .A2(n782), .B1(n418), .B2(n755), .ZN(n564) );
  OAI211_X1 U351 ( .C1(N378), .C2(n683), .A(n748), .B(n782), .ZN(n784) );
  OAI21_X1 U352 ( .B1(n426), .B2(n774), .A(n784), .ZN(n431) );
  INV_X1 U353 ( .A(N377), .ZN(n785) );
  OAI22_X1 U354 ( .A1(n785), .A2(n750), .B1(n388), .B2(n755), .ZN(n534) );
  OAI22_X1 U355 ( .A1(n750), .A2(n787), .B1(n390), .B2(n755), .ZN(n536) );
  OAI22_X1 U356 ( .A1(n660), .A2(n788), .B1(n391), .B2(n755), .ZN(n537) );
  OAI22_X1 U357 ( .A1(n687), .A2(n789), .B1(n392), .B2(n755), .ZN(n538) );
  OAI22_X1 U358 ( .A1(n687), .A2(n790), .B1(n393), .B2(n755), .ZN(n539) );
  INV_X1 U359 ( .A(N383), .ZN(n791) );
  OAI22_X1 U360 ( .A1(n718), .A2(n791), .B1(n394), .B2(n755), .ZN(n540) );
  INV_X1 U361 ( .A(N384), .ZN(n792) );
  OAI22_X1 U362 ( .A1(n688), .A2(n792), .B1(n395), .B2(n755), .ZN(n541) );
  INV_X1 U363 ( .A(N385), .ZN(n793) );
  OAI22_X1 U364 ( .A1(n751), .A2(n793), .B1(n396), .B2(n755), .ZN(n542) );
  OAI22_X1 U365 ( .A1(n687), .A2(n794), .B1(n397), .B2(n754), .ZN(n543) );
  OAI22_X1 U366 ( .A1(n676), .A2(n795), .B1(n398), .B2(n754), .ZN(n544) );
  OAI22_X1 U367 ( .A1(n688), .A2(n796), .B1(n399), .B2(n754), .ZN(n545) );
  INV_X1 U368 ( .A(N390), .ZN(n798) );
  OAI22_X1 U369 ( .A1(n655), .A2(n798), .B1(n401), .B2(n754), .ZN(n547) );
  INV_X1 U370 ( .A(N391), .ZN(n799) );
  OAI22_X1 U371 ( .A1(n751), .A2(n799), .B1(n402), .B2(n754), .ZN(n548) );
  INV_X1 U372 ( .A(N392), .ZN(n800) );
  OAI22_X1 U373 ( .A1(n719), .A2(n800), .B1(n403), .B2(n754), .ZN(n549) );
  OAI22_X1 U374 ( .A1(n752), .A2(n801), .B1(n404), .B2(n754), .ZN(n550) );
  OAI22_X1 U375 ( .A1(n718), .A2(n802), .B1(n405), .B2(n754), .ZN(n551) );
  OAI22_X1 U376 ( .A1(n750), .A2(n803), .B1(n406), .B2(n754), .ZN(n552) );
  OAI22_X1 U377 ( .A1(n655), .A2(n804), .B1(n407), .B2(n754), .ZN(n553) );
  INV_X1 U378 ( .A(n666), .ZN(n805) );
  OAI22_X1 U379 ( .A1(n675), .A2(n805), .B1(n408), .B2(n753), .ZN(n554) );
  INV_X1 U380 ( .A(n677), .ZN(n806) );
  OAI22_X1 U381 ( .A1(n806), .A2(n674), .B1(n409), .B2(n753), .ZN(n555) );
  INV_X1 U382 ( .A(n679), .ZN(n807) );
  OAI22_X1 U383 ( .A1(n752), .A2(n807), .B1(n410), .B2(n753), .ZN(n556) );
  OAI22_X1 U384 ( .A1(n751), .A2(n808), .B1(n411), .B2(n753), .ZN(n557) );
  OAI22_X1 U385 ( .A1(n675), .A2(n810), .B1(n413), .B2(n753), .ZN(n559) );
  OAI22_X1 U386 ( .A1(n718), .A2(n811), .B1(n414), .B2(n753), .ZN(n560) );
  INV_X1 U387 ( .A(N404), .ZN(n812) );
  OAI22_X1 U388 ( .A1(n812), .A2(n674), .B1(n415), .B2(n753), .ZN(n561) );
  INV_X1 U389 ( .A(N405), .ZN(n813) );
  OAI22_X1 U390 ( .A1(n676), .A2(n813), .B1(n416), .B2(n753), .ZN(n562) );
  INV_X1 U391 ( .A(n712), .ZN(n814) );
  OAI22_X1 U392 ( .A1(n719), .A2(n814), .B1(n417), .B2(n753), .ZN(n563) );
  INV_X1 U393 ( .A(n503), .ZN(n815) );
  OAI21_X1 U394 ( .B1(n753), .B2(n815), .A(n674), .ZN(n532) );
  MUX2_X1 U395 ( .A(n817), .B(n658), .S(n387), .Z(n509) );
  OAI21_X1 U396 ( .B1(n218), .B2(n217), .A(n860), .ZN(n818) );
  INV_X1 U397 ( .A(N266), .ZN(n832) );
  INV_X1 U398 ( .A(N267), .ZN(n833) );
  INV_X1 U399 ( .A(N268), .ZN(n834) );
  INV_X1 U400 ( .A(N269), .ZN(n835) );
  NAND4_X1 U401 ( .A1(n832), .A2(n833), .A3(n834), .A4(n835), .ZN(n819) );
  NOR4_X1 U402 ( .A1(n819), .A2(N272), .A3(N271), .A4(N270), .ZN(n825) );
  INV_X1 U403 ( .A(N273), .ZN(n839) );
  INV_X1 U404 ( .A(N274), .ZN(n840) );
  INV_X1 U405 ( .A(N275), .ZN(n841) );
  INV_X1 U406 ( .A(N276), .ZN(n842) );
  INV_X1 U407 ( .A(N280), .ZN(n846) );
  INV_X1 U408 ( .A(N281), .ZN(n847) );
  INV_X1 U409 ( .A(N282), .ZN(n848) );
  INV_X1 U410 ( .A(N283), .ZN(n849) );
  NAND4_X1 U411 ( .A1(n849), .A2(n847), .A3(n848), .A4(n846), .ZN(n821) );
  INV_X1 U412 ( .A(N287), .ZN(n853) );
  INV_X1 U413 ( .A(N288), .ZN(n854) );
  INV_X1 U414 ( .A(N289), .ZN(n855) );
  INV_X1 U415 ( .A(N290), .ZN(n856) );
  INV_X1 U416 ( .A(N294), .ZN(n827) );
  OAI22_X1 U417 ( .A1(n622), .A2(n827), .B1(n580), .B2(n758), .ZN(n581) );
  OAI211_X1 U418 ( .C1(N265), .C2(n828), .A(n747), .B(n827), .ZN(n829) );
  INV_X1 U419 ( .A(N264), .ZN(n830) );
  OAI22_X1 U420 ( .A1(n830), .A2(n760), .B1(n514), .B2(n758), .ZN(n611) );
  INV_X1 U421 ( .A(N265), .ZN(n831) );
  OAI22_X1 U422 ( .A1(n831), .A2(n761), .B1(n515), .B2(n758), .ZN(n610) );
  OAI22_X1 U423 ( .A1(n623), .A2(n832), .B1(n516), .B2(n758), .ZN(n609) );
  OAI22_X1 U424 ( .A1(n694), .A2(n833), .B1(n517), .B2(n758), .ZN(n608) );
  OAI22_X1 U425 ( .A1(n743), .A2(n834), .B1(n518), .B2(n758), .ZN(n607) );
  OAI22_X1 U426 ( .A1(n716), .A2(n835), .B1(n519), .B2(n758), .ZN(n606) );
  INV_X1 U427 ( .A(N270), .ZN(n836) );
  OAI22_X1 U428 ( .A1(n624), .A2(n836), .B1(n520), .B2(n758), .ZN(n605) );
  INV_X1 U429 ( .A(N271), .ZN(n837) );
  INV_X1 U430 ( .A(N272), .ZN(n838) );
  OAI22_X1 U431 ( .A1(n762), .A2(n838), .B1(n522), .B2(n758), .ZN(n603) );
  OAI22_X1 U432 ( .A1(n694), .A2(n839), .B1(n523), .B2(n758), .ZN(n602) );
  OAI22_X1 U433 ( .A1(n702), .A2(n840), .B1(n524), .B2(n757), .ZN(n601) );
  OAI22_X1 U434 ( .A1(n702), .A2(n841), .B1(n525), .B2(n757), .ZN(n600) );
  OAI22_X1 U435 ( .A1(n696), .A2(n842), .B1(n526), .B2(n757), .ZN(n599) );
  INV_X1 U436 ( .A(n646), .ZN(n843) );
  OAI22_X1 U437 ( .A1(n716), .A2(n843), .B1(n527), .B2(n757), .ZN(n598) );
  INV_X1 U438 ( .A(N278), .ZN(n844) );
  OAI22_X1 U439 ( .A1(n761), .A2(n844), .B1(n528), .B2(n757), .ZN(n597) );
  INV_X1 U440 ( .A(N279), .ZN(n845) );
  OAI22_X1 U441 ( .A1(n740), .A2(n845), .B1(n529), .B2(n757), .ZN(n596) );
  OAI22_X1 U442 ( .A1(n741), .A2(n846), .B1(n530), .B2(n757), .ZN(n595) );
  OAI22_X1 U443 ( .A1(n716), .A2(n847), .B1(n531), .B2(n757), .ZN(n594) );
  OAI22_X1 U444 ( .A1(n671), .A2(n848), .B1(n568), .B2(n757), .ZN(n593) );
  OAI22_X1 U445 ( .A1(n740), .A2(n849), .B1(n569), .B2(n757), .ZN(n592) );
  INV_X1 U446 ( .A(n656), .ZN(n850) );
  OAI22_X1 U447 ( .A1(n762), .A2(n850), .B1(n570), .B2(n756), .ZN(n591) );
  INV_X1 U448 ( .A(n644), .ZN(n851) );
  OAI22_X1 U449 ( .A1(n624), .A2(n851), .B1(n571), .B2(n756), .ZN(n590) );
  INV_X1 U450 ( .A(n697), .ZN(n852) );
  OAI22_X1 U451 ( .A1(n760), .A2(n852), .B1(n572), .B2(n756), .ZN(n589) );
  OAI22_X1 U452 ( .A1(n702), .A2(n853), .B1(n573), .B2(n756), .ZN(n588) );
  OAI22_X1 U453 ( .A1(n622), .A2(n854), .B1(n574), .B2(n756), .ZN(n587) );
  OAI22_X1 U454 ( .A1(n743), .A2(n855), .B1(n575), .B2(n756), .ZN(n586) );
  OAI22_X1 U455 ( .A1(n702), .A2(n856), .B1(n576), .B2(n756), .ZN(n585) );
  INV_X1 U456 ( .A(N292), .ZN(n858) );
  OAI22_X1 U457 ( .A1(n615), .A2(n858), .B1(n578), .B2(n756), .ZN(n583) );
  INV_X1 U458 ( .A(N293), .ZN(n859) );
  OAI22_X1 U459 ( .A1(n615), .A2(n859), .B1(n579), .B2(n756), .ZN(n582) );
  OAI22_X1 U460 ( .A1(n746), .A2(n740), .B1(n513), .B2(n757), .ZN(n612) );
  INV_X1 U461 ( .A(N159), .ZN(n875) );
  INV_X1 U462 ( .A(N158), .ZN(n874) );
  INV_X1 U489 ( .A(N157), .ZN(n873) );
  INV_X1 U496 ( .A(N156), .ZN(n872) );
  NAND4_X1 U497 ( .A1(n875), .A2(n874), .A3(n873), .A4(n872), .ZN(n861) );
  NOR4_X1 U498 ( .A1(n861), .A2(N152), .A3(N154), .A4(N155), .ZN(n863) );
  INV_X1 U499 ( .A(N171), .ZN(n884) );
  INV_X1 U500 ( .A(N170), .ZN(n883) );
  INV_X1 U501 ( .A(N169), .ZN(n882) );
  INV_X1 U502 ( .A(N168), .ZN(n881) );
  INV_X1 U503 ( .A(n640), .ZN(n888) );
  INV_X1 U504 ( .A(N174), .ZN(n887) );
  INV_X1 U505 ( .A(n634), .ZN(n886) );
  INV_X1 U506 ( .A(n632), .ZN(n885) );
  INV_X1 U507 ( .A(N179), .ZN(n892) );
  INV_X1 U508 ( .A(N178), .ZN(n891) );
  INV_X1 U509 ( .A(n657), .ZN(n890) );
  INV_X1 U510 ( .A(N176), .ZN(n889) );
  INV_X1 U511 ( .A(N182), .ZN(n867) );
  INV_X1 U512 ( .A(N181), .ZN(n894) );
  INV_X1 U513 ( .A(N180), .ZN(n893) );
  OAI21_X1 U514 ( .B1(n200), .B2(n968), .A(n897), .ZN(n866) );
  NAND2_X1 U515 ( .A1(n866), .A2(n774), .ZN(n900) );
  INV_X1 U516 ( .A(n900), .ZN(n898) );
  OAI21_X1 U517 ( .B1(n639), .B2(n895), .A(n763), .ZN(n899) );
  OAI22_X1 U518 ( .A1(n730), .A2(n867), .B1(n386), .B2(n763), .ZN(n498) );
  INV_X1 U519 ( .A(N152), .ZN(n868) );
  OAI22_X1 U520 ( .A1(n636), .A2(n868), .B1(n356), .B2(n766), .ZN(n468) );
  INV_X1 U521 ( .A(N153), .ZN(n869) );
  OAI22_X1 U522 ( .A1(n869), .A2(n728), .B1(n357), .B2(n765), .ZN(n469) );
  INV_X1 U523 ( .A(N154), .ZN(n870) );
  OAI22_X1 U524 ( .A1(n767), .A2(n870), .B1(n358), .B2(n765), .ZN(n470) );
  INV_X1 U525 ( .A(N155), .ZN(n871) );
  OAI22_X1 U526 ( .A1(n728), .A2(n871), .B1(n359), .B2(n765), .ZN(n471) );
  OAI22_X1 U527 ( .A1(n731), .A2(n872), .B1(n360), .B2(n765), .ZN(n472) );
  OAI22_X1 U528 ( .A1(n731), .A2(n873), .B1(n361), .B2(n765), .ZN(n473) );
  OAI22_X1 U529 ( .A1(n767), .A2(n874), .B1(n362), .B2(n765), .ZN(n474) );
  OAI22_X1 U530 ( .A1(n767), .A2(n875), .B1(n363), .B2(n765), .ZN(n475) );
  OAI22_X1 U531 ( .A1(n767), .A2(n641), .B1(n364), .B2(n765), .ZN(n476) );
  INV_X1 U532 ( .A(N161), .ZN(n876) );
  OAI22_X1 U533 ( .A1(n727), .A2(n876), .B1(n365), .B2(n765), .ZN(n477) );
  OAI22_X1 U534 ( .A1(n767), .A2(n642), .B1(n366), .B2(n765), .ZN(n478) );
  OAI22_X1 U535 ( .A1(n727), .A2(n643), .B1(n367), .B2(n765), .ZN(n479) );
  INV_X1 U536 ( .A(N164), .ZN(n877) );
  OAI22_X1 U537 ( .A1(n731), .A2(n877), .B1(n368), .B2(n764), .ZN(n480) );
  INV_X1 U538 ( .A(N165), .ZN(n878) );
  OAI22_X1 U539 ( .A1(n729), .A2(n878), .B1(n369), .B2(n764), .ZN(n481) );
  INV_X1 U540 ( .A(N166), .ZN(n879) );
  OAI22_X1 U541 ( .A1(n731), .A2(n879), .B1(n370), .B2(n764), .ZN(n482) );
  INV_X1 U542 ( .A(N167), .ZN(n880) );
  OAI22_X1 U543 ( .A1(n730), .A2(n880), .B1(n371), .B2(n764), .ZN(n483) );
  OAI22_X1 U544 ( .A1(n728), .A2(n881), .B1(n372), .B2(n764), .ZN(n484) );
  OAI22_X1 U545 ( .A1(n664), .A2(n882), .B1(n373), .B2(n764), .ZN(n485) );
  OAI22_X1 U546 ( .A1(n636), .A2(n648), .B1(n374), .B2(n764), .ZN(n486) );
  OAI22_X1 U547 ( .A1(n664), .A2(n884), .B1(n375), .B2(n764), .ZN(n487) );
  OAI22_X1 U548 ( .A1(n731), .A2(n885), .B1(n376), .B2(n764), .ZN(n488) );
  OAI22_X1 U549 ( .A1(n730), .A2(n886), .B1(n377), .B2(n764), .ZN(n489) );
  OAI22_X1 U550 ( .A1(n727), .A2(n692), .B1(n378), .B2(n763), .ZN(n490) );
  OAI22_X1 U551 ( .A1(n729), .A2(n888), .B1(n379), .B2(n764), .ZN(n491) );
  OAI22_X1 U552 ( .A1(n729), .A2(n889), .B1(n380), .B2(n763), .ZN(n492) );
  OAI22_X1 U553 ( .A1(n730), .A2(n890), .B1(n381), .B2(n763), .ZN(n493) );
  OAI22_X1 U554 ( .A1(n729), .A2(n891), .B1(n382), .B2(n763), .ZN(n494) );
  OAI22_X1 U555 ( .A1(n731), .A2(n892), .B1(n383), .B2(n763), .ZN(n495) );
  OAI22_X1 U556 ( .A1(n664), .A2(n893), .B1(n384), .B2(n763), .ZN(n496) );
  OAI22_X1 U557 ( .A1(n664), .A2(n894), .B1(n385), .B2(n763), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n709), .A2(n763), .ZN(n896) );
  OAI22_X1 U559 ( .A1(N151), .A2(n896), .B1(n425), .B2(n774), .ZN(n433) );
  OAI21_X1 U560 ( .B1(n200), .B2(n966), .A(n941), .ZN(n901) );
  NAND2_X1 U561 ( .A1(n901), .A2(n774), .ZN(n943) );
  INV_X1 U562 ( .A(n943), .ZN(n942) );
  INV_X1 U563 ( .A(N42), .ZN(n910) );
  INV_X1 U564 ( .A(N64), .ZN(n932) );
  INV_X1 U565 ( .A(N63), .ZN(n931) );
  INV_X1 U566 ( .A(N62), .ZN(n930) );
  INV_X1 U567 ( .A(N61), .ZN(n929) );
  NAND4_X1 U568 ( .A1(n932), .A2(n931), .A3(n930), .A4(n929), .ZN(n902) );
  INV_X1 U569 ( .A(N45), .ZN(n913) );
  INV_X1 U570 ( .A(N44), .ZN(n912) );
  INV_X1 U571 ( .A(N43), .ZN(n911) );
  NOR4_X1 U572 ( .A1(N46), .A2(N47), .A3(N48), .A4(N49), .ZN(n903) );
  INV_X1 U573 ( .A(N53), .ZN(n921) );
  INV_X1 U574 ( .A(N52), .ZN(n920) );
  INV_X1 U575 ( .A(N51), .ZN(n919) );
  INV_X1 U576 ( .A(N57), .ZN(n925) );
  INV_X1 U577 ( .A(N56), .ZN(n924) );
  INV_X1 U578 ( .A(N55), .ZN(n923) );
  INV_X1 U579 ( .A(N54), .ZN(n922) );
  INV_X1 U580 ( .A(N71), .ZN(n909) );
  INV_X1 U581 ( .A(N41), .ZN(n939) );
  OAI22_X1 U582 ( .A1(n939), .A2(n725), .B1(n324), .B2(n771), .ZN(n436) );
  OAI22_X1 U583 ( .A1(n910), .A2(n725), .B1(n325), .B2(n771), .ZN(n437) );
  OAI22_X1 U584 ( .A1(n735), .A2(n911), .B1(n326), .B2(n771), .ZN(n438) );
  OAI22_X1 U585 ( .A1(n736), .A2(n912), .B1(n327), .B2(n771), .ZN(n439) );
  OAI22_X1 U586 ( .A1(n734), .A2(n913), .B1(n328), .B2(n771), .ZN(n440) );
  INV_X1 U587 ( .A(N46), .ZN(n914) );
  OAI22_X1 U588 ( .A1(n733), .A2(n914), .B1(n329), .B2(n771), .ZN(n441) );
  INV_X1 U589 ( .A(N47), .ZN(n915) );
  OAI22_X1 U590 ( .A1(n732), .A2(n915), .B1(n330), .B2(n771), .ZN(n442) );
  INV_X1 U591 ( .A(N48), .ZN(n916) );
  OAI22_X1 U592 ( .A1(n662), .A2(n916), .B1(n331), .B2(n771), .ZN(n443) );
  INV_X1 U593 ( .A(N49), .ZN(n917) );
  OAI22_X1 U594 ( .A1(n724), .A2(n917), .B1(n332), .B2(n771), .ZN(n444) );
  OAI22_X1 U595 ( .A1(n735), .A2(n919), .B1(n334), .B2(n770), .ZN(n446) );
  OAI22_X1 U596 ( .A1(n662), .A2(n920), .B1(n335), .B2(n770), .ZN(n447) );
  OAI22_X1 U597 ( .A1(n736), .A2(n921), .B1(n336), .B2(n770), .ZN(n448) );
  OAI22_X1 U598 ( .A1(n737), .A2(n922), .B1(n337), .B2(n770), .ZN(n449) );
  OAI22_X1 U599 ( .A1(n734), .A2(n923), .B1(n338), .B2(n770), .ZN(n450) );
  OAI22_X1 U600 ( .A1(n617), .A2(n924), .B1(n339), .B2(n770), .ZN(n451) );
  OAI22_X1 U601 ( .A1(n700), .A2(n925), .B1(n340), .B2(n770), .ZN(n452) );
  INV_X1 U602 ( .A(n649), .ZN(n926) );
  OAI22_X1 U603 ( .A1(n737), .A2(n926), .B1(n341), .B2(n770), .ZN(n453) );
  INV_X1 U604 ( .A(N59), .ZN(n927) );
  OAI22_X1 U605 ( .A1(n733), .A2(n927), .B1(n342), .B2(n770), .ZN(n454) );
  OAI22_X1 U606 ( .A1(n662), .A2(n929), .B1(n344), .B2(n769), .ZN(n456) );
  OAI22_X1 U607 ( .A1(n616), .A2(n930), .B1(n345), .B2(n769), .ZN(n457) );
  OAI22_X1 U608 ( .A1(n695), .A2(n931), .B1(n346), .B2(n769), .ZN(n458) );
  OAI22_X1 U609 ( .A1(n616), .A2(n932), .B1(n347), .B2(n770), .ZN(n459) );
  INV_X1 U610 ( .A(N65), .ZN(n933) );
  OAI22_X1 U611 ( .A1(n732), .A2(n933), .B1(n348), .B2(n769), .ZN(n460) );
  INV_X1 U612 ( .A(N66), .ZN(n934) );
  OAI22_X1 U613 ( .A1(n695), .A2(n934), .B1(n349), .B2(n769), .ZN(n461) );
  INV_X1 U614 ( .A(N67), .ZN(n935) );
  OAI22_X1 U615 ( .A1(n737), .A2(n935), .B1(n350), .B2(n769), .ZN(n462) );
  INV_X1 U616 ( .A(N68), .ZN(n936) );
  OAI22_X1 U617 ( .A1(n732), .A2(n936), .B1(n351), .B2(n769), .ZN(n463) );
  INV_X1 U618 ( .A(N69), .ZN(n937) );
  OAI22_X1 U619 ( .A1(n724), .A2(n937), .B1(n352), .B2(n769), .ZN(n464) );
  INV_X1 U620 ( .A(N70), .ZN(n938) );
  OAI22_X1 U621 ( .A1(n617), .A2(n938), .B1(n353), .B2(n769), .ZN(n465) );
  NAND4_X1 U622 ( .A1(N40), .A2(n769), .A3(n659), .A4(n939), .ZN(n940) );
  OAI21_X1 U623 ( .B1(n424), .B2(n774), .A(n940), .ZN(n434) );
  MUX2_X1 U624 ( .A(n943), .B(n621), .S(n323), .Z(n507) );
endmodule


module regFFD_NBIT32_0 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n65) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n66) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n67) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n68) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n69) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n70) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n71) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n72) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n73) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n74) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n75) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n76) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n77) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n78) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n79) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n80) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n81) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n82) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n83) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n84) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n85) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n86) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n87) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n88) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n89) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n90) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n91) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n92) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n93) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n94) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n95) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n96) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n96), .B2(ENABLE), .A(n39), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n39) );
  OAI21_X1 U7 ( .B1(n95), .B2(ENABLE), .A(n40), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n40) );
  OAI21_X1 U9 ( .B1(n94), .B2(ENABLE), .A(n41), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n41) );
  OAI21_X1 U11 ( .B1(n93), .B2(ENABLE), .A(n43), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n43) );
  OAI21_X1 U13 ( .B1(n92), .B2(ENABLE), .A(n44), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n91), .B2(ENABLE), .A(n45), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n45) );
  OAI21_X1 U17 ( .B1(n90), .B2(ENABLE), .A(n46), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n46) );
  OAI21_X1 U19 ( .B1(n89), .B2(ENABLE), .A(n47), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n47) );
  OAI21_X1 U21 ( .B1(n88), .B2(ENABLE), .A(n48), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n48) );
  OAI21_X1 U23 ( .B1(n87), .B2(ENABLE), .A(n49), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n49) );
  OAI21_X1 U25 ( .B1(n86), .B2(ENABLE), .A(n50), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n50) );
  OAI21_X1 U27 ( .B1(n85), .B2(ENABLE), .A(n51), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n51) );
  OAI21_X1 U29 ( .B1(n84), .B2(ENABLE), .A(n52), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n52) );
  OAI21_X1 U31 ( .B1(n83), .B2(ENABLE), .A(n54), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n82), .B2(ENABLE), .A(n55), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n55) );
  OAI21_X1 U35 ( .B1(n81), .B2(ENABLE), .A(n56), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n56) );
  OAI21_X1 U37 ( .B1(n80), .B2(ENABLE), .A(n57), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n57) );
  OAI21_X1 U39 ( .B1(n79), .B2(ENABLE), .A(n58), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n58) );
  OAI21_X1 U41 ( .B1(n78), .B2(ENABLE), .A(n59), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n59) );
  OAI21_X1 U43 ( .B1(n77), .B2(ENABLE), .A(n60), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n60) );
  OAI21_X1 U45 ( .B1(n76), .B2(ENABLE), .A(n61), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n61) );
  OAI21_X1 U47 ( .B1(n75), .B2(ENABLE), .A(n62), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n62) );
  OAI21_X1 U49 ( .B1(n74), .B2(ENABLE), .A(n63), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n63) );
  OAI21_X1 U51 ( .B1(n73), .B2(ENABLE), .A(n33), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U53 ( .B1(n72), .B2(ENABLE), .A(n34), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n34) );
  OAI21_X1 U55 ( .B1(n71), .B2(ENABLE), .A(n35), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n35) );
  OAI21_X1 U57 ( .B1(n70), .B2(ENABLE), .A(n36), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n36) );
  OAI21_X1 U59 ( .B1(n69), .B2(ENABLE), .A(n37), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n37) );
  OAI21_X1 U61 ( .B1(n68), .B2(ENABLE), .A(n38), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n38) );
  OAI21_X1 U63 ( .B1(n67), .B2(ENABLE), .A(n42), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n42) );
  OAI21_X1 U65 ( .B1(n66), .B2(ENABLE), .A(n53), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n65), .B2(ENABLE), .A(n64), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n64) );
endmodule


module regFFD_NBIT32_19 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module regFFD_NBIT32_18 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_767 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_766 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0 UIV ( .A(S), .Y(SB) );
  ND2_0 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_767 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_766 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_255 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_765 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_764 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_763 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_255 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_255 UIV ( .A(S), .Y(SB) );
  ND2_765 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_764 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_763 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_254 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_762 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_761 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_760 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_254 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_254 UIV ( .A(S), .Y(SB) );
  ND2_762 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_761 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_760 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_253 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_759 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_758 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_757 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_253 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_253 UIV ( .A(S), .Y(SB) );
  ND2_759 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_758 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_757 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_252 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_756 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_755 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_754 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_252 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_252 UIV ( .A(S), .Y(SB) );
  ND2_756 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_755 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_754 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_251 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_753 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_752 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_751 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_251 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_251 UIV ( .A(S), .Y(SB) );
  ND2_753 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_752 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_751 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_250 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_750 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_749 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_748 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_250 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_250 UIV ( .A(S), .Y(SB) );
  ND2_750 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_749 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_748 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_249 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_747 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_746 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_745 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_249 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_249 UIV ( .A(S), .Y(SB) );
  ND2_747 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_746 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_745 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_248 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_744 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_743 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_742 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_248 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_248 UIV ( .A(S), .Y(SB) );
  ND2_744 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_743 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_742 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_247 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_741 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_740 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_739 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_247 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_247 UIV ( .A(S), .Y(SB) );
  ND2_741 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_740 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_739 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_246 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_738 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_737 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_736 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_246 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_246 UIV ( .A(S), .Y(SB) );
  ND2_738 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_737 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_736 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_245 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_735 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_734 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_733 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_245 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_245 UIV ( .A(S), .Y(SB) );
  ND2_735 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_734 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_733 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_244 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_732 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_731 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_730 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_244 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_244 UIV ( .A(S), .Y(SB) );
  ND2_732 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_731 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_730 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_243 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_729 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_728 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_727 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_243 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_243 UIV ( .A(S), .Y(SB) );
  ND2_729 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_728 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_727 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_242 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_726 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_725 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_724 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_242 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_242 UIV ( .A(S), .Y(SB) );
  ND2_726 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_725 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_724 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_241 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_723 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_722 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_721 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_241 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_241 UIV ( .A(S), .Y(SB) );
  ND2_723 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_722 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_721 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_240 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_720 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_719 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_718 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_240 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_240 UIV ( .A(S), .Y(SB) );
  ND2_720 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_719 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_718 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_239 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_717 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_716 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_715 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_239 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_239 UIV ( .A(S), .Y(SB) );
  ND2_717 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_716 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_715 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_238 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_714 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_713 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_712 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_238 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_238 UIV ( .A(S), .Y(SB) );
  ND2_714 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_713 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_712 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_237 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_711 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_710 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_709 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_237 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_237 UIV ( .A(S), .Y(SB) );
  ND2_711 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_710 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_709 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_236 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_708 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_707 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_706 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_236 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_236 UIV ( .A(S), .Y(SB) );
  ND2_708 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_707 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_706 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_235 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_705 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_704 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_703 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_235 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_235 UIV ( .A(S), .Y(SB) );
  ND2_705 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_704 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_703 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_234 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_702 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_701 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_700 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_234 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_234 UIV ( .A(S), .Y(SB) );
  ND2_702 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_701 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_700 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_233 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_699 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_698 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_697 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_233 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_233 UIV ( .A(S), .Y(SB) );
  ND2_699 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_698 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_697 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_232 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_696 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_695 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_694 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_232 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_232 UIV ( .A(S), .Y(SB) );
  ND2_696 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_695 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_694 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_231 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_693 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_692 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_691 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_231 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_231 UIV ( .A(S), .Y(SB) );
  ND2_693 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_692 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_691 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_230 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_690 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_689 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_688 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_230 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_230 UIV ( .A(S), .Y(SB) );
  ND2_690 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_689 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_688 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_229 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_687 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_686 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_685 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_229 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_229 UIV ( .A(S), .Y(SB) );
  ND2_687 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_686 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_685 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_228 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_684 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_683 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_682 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_228 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_228 UIV ( .A(S), .Y(SB) );
  ND2_684 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_683 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_682 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_227 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_681 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_680 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_679 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_227 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_227 UIV ( .A(S), .Y(SB) );
  ND2_681 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_680 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_679 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_226 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_678 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_677 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_676 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_226 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_226 UIV ( .A(S), .Y(SB) );
  ND2_678 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_677 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_676 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_225 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_675 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_674 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_673 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_225 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_225 UIV ( .A(S), .Y(SB) );
  ND2_675 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_674 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_673 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n4, n5, n6;

  MUX21_0 gen1_0 ( .A(A[0]), .B(B[0]), .S(n6), .Y(Y[0]) );
  MUX21_255 gen1_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_254 gen1_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_253 gen1_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_252 gen1_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_251 gen1_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_250 gen1_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_249 gen1_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_248 gen1_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_247 gen1_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_246 gen1_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_245 gen1_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_244 gen1_12 ( .A(A[12]), .B(B[12]), .S(n4), .Y(Y[12]) );
  MUX21_243 gen1_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_242 gen1_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_241 gen1_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_240 gen1_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_239 gen1_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_238 gen1_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_237 gen1_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_236 gen1_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_235 gen1_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_234 gen1_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_233 gen1_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_232 gen1_24 ( .A(A[24]), .B(B[24]), .S(n5), .Y(Y[24]) );
  MUX21_231 gen1_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_230 gen1_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_229 gen1_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_228 gen1_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_227 gen1_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_226 gen1_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_225 gen1_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n4) );
  BUF_X1 U2 ( .A(SEL), .Z(n5) );
  BUF_X1 U3 ( .A(SEL), .Z(n6) );
endmodule


module regFFD_NBIT32_17 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module regFFD_NBIT32_16 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module regFFD_NBIT32_15 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module regFFD_NBIT32_14 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module regFFD_NBIT32_13 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module regFFD_NBIT32_12 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module sign_eval_N_in5_N_out32 ( IR_out, signed_val, Immediate );
  input [4:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   N0, n2;
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];
  assign Immediate[5] = N0;
  assign Immediate[6] = N0;
  assign Immediate[7] = N0;
  assign Immediate[8] = N0;
  assign Immediate[9] = N0;
  assign Immediate[10] = N0;
  assign Immediate[11] = N0;
  assign Immediate[12] = N0;
  assign Immediate[13] = N0;
  assign Immediate[14] = N0;
  assign Immediate[15] = N0;
  assign Immediate[16] = N0;
  assign Immediate[17] = N0;
  assign Immediate[18] = N0;
  assign Immediate[19] = N0;
  assign Immediate[20] = N0;
  assign Immediate[21] = N0;
  assign Immediate[22] = N0;
  assign Immediate[23] = N0;
  assign Immediate[24] = N0;
  assign Immediate[25] = N0;
  assign Immediate[26] = N0;
  assign Immediate[27] = N0;
  assign Immediate[28] = N0;
  assign Immediate[29] = N0;
  assign Immediate[30] = N0;
  assign Immediate[31] = N0;

  NOR2_X1 U1 ( .A1(signed_val), .A2(n2), .ZN(N0) );
  INV_X1 U2 ( .A(IR_out[4]), .ZN(n2) );
endmodule


module sign_eval_N_in16_N_out32 ( IR_out, signed_val, Immediate );
  input [15:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   N0, n2;
  assign Immediate[15] = IR_out[15];
  assign Immediate[14] = IR_out[14];
  assign Immediate[13] = IR_out[13];
  assign Immediate[12] = IR_out[12];
  assign Immediate[11] = IR_out[11];
  assign Immediate[10] = IR_out[10];
  assign Immediate[9] = IR_out[9];
  assign Immediate[8] = IR_out[8];
  assign Immediate[7] = IR_out[7];
  assign Immediate[6] = IR_out[6];
  assign Immediate[5] = IR_out[5];
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];
  assign Immediate[16] = N0;
  assign Immediate[17] = N0;
  assign Immediate[18] = N0;
  assign Immediate[19] = N0;
  assign Immediate[20] = N0;
  assign Immediate[21] = N0;
  assign Immediate[22] = N0;
  assign Immediate[23] = N0;
  assign Immediate[24] = N0;
  assign Immediate[25] = N0;
  assign Immediate[26] = N0;
  assign Immediate[27] = N0;
  assign Immediate[28] = N0;
  assign Immediate[29] = N0;
  assign Immediate[30] = N0;
  assign Immediate[31] = N0;

  NOR2_X1 U1 ( .A1(signed_val), .A2(n2), .ZN(N0) );
  INV_X1 U2 ( .A(IR_out[15]), .ZN(n2) );
endmodule


module sign_eval_N_in26_N_out32 ( IR_out, signed_val, Immediate );
  input [25:0] IR_out;
  output [31:0] Immediate;
  input signed_val;
  wire   N0, n2;
  assign Immediate[25] = IR_out[25];
  assign Immediate[24] = IR_out[24];
  assign Immediate[23] = IR_out[23];
  assign Immediate[22] = IR_out[22];
  assign Immediate[21] = IR_out[21];
  assign Immediate[20] = IR_out[20];
  assign Immediate[19] = IR_out[19];
  assign Immediate[18] = IR_out[18];
  assign Immediate[17] = IR_out[17];
  assign Immediate[16] = IR_out[16];
  assign Immediate[15] = IR_out[15];
  assign Immediate[14] = IR_out[14];
  assign Immediate[13] = IR_out[13];
  assign Immediate[12] = IR_out[12];
  assign Immediate[11] = IR_out[11];
  assign Immediate[10] = IR_out[10];
  assign Immediate[9] = IR_out[9];
  assign Immediate[8] = IR_out[8];
  assign Immediate[7] = IR_out[7];
  assign Immediate[6] = IR_out[6];
  assign Immediate[5] = IR_out[5];
  assign Immediate[4] = IR_out[4];
  assign Immediate[3] = IR_out[3];
  assign Immediate[2] = IR_out[2];
  assign Immediate[1] = IR_out[1];
  assign Immediate[0] = IR_out[0];
  assign Immediate[26] = N0;
  assign Immediate[27] = N0;
  assign Immediate[28] = N0;
  assign Immediate[29] = N0;
  assign Immediate[30] = N0;
  assign Immediate[31] = N0;

  NOR2_X1 U1 ( .A1(signed_val), .A2(n2), .ZN(N0) );
  INV_X1 U2 ( .A(IR_out[25]), .ZN(n2) );
endmodule


module IR_DECODE_NBIT32_opBIT6_regBIT5 ( CLK, IR_26, OPCODE, is_signed, RS1, 
        RS2, RD, IMMEDIATE );
  input [25:0] IR_26;
  input [5:0] OPCODE;
  output [4:0] RS1;
  output [4:0] RS2;
  output [4:0] RD;
  output [31:0] IMMEDIATE;
  input CLK, is_signed;
  wire   N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38;
  wire   [31:0] IMMEDIATE_16;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;
  assign N133 = IR_26[21];
  assign N134 = IR_26[22];
  assign N135 = IR_26[23];
  assign N136 = IR_26[24];
  assign N137 = IR_26[25];
  assign N138 = IR_26[16];
  assign N139 = IR_26[17];
  assign N140 = IR_26[18];
  assign N141 = IR_26[19];
  assign N142 = IR_26[20];

  DLH_X1 \RD_reg[4]  ( .G(CLK), .D(n34), .Q(RD[4]) );
  DLH_X1 \RD_reg[3]  ( .G(CLK), .D(n35), .Q(RD[3]) );
  DLH_X1 \RD_reg[2]  ( .G(CLK), .D(n36), .Q(RD[2]) );
  DLH_X1 \RD_reg[1]  ( .G(CLK), .D(n37), .Q(RD[1]) );
  DLH_X1 \RD_reg[0]  ( .G(CLK), .D(n38), .Q(RD[0]) );
  DLH_X1 \IMMEDIATE_reg[31]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[31]) );
  DLH_X1 \IMMEDIATE_reg[30]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[30]) );
  DLH_X1 \IMMEDIATE_reg[29]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[29]) );
  DLH_X1 \IMMEDIATE_reg[28]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[28]) );
  DLH_X1 \IMMEDIATE_reg[27]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[27]) );
  DLH_X1 \IMMEDIATE_reg[26]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[26]) );
  DLH_X1 \IMMEDIATE_reg[25]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[25]) );
  DLH_X1 \IMMEDIATE_reg[24]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[24]) );
  DLH_X1 \IMMEDIATE_reg[23]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[23]) );
  DLH_X1 \IMMEDIATE_reg[22]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[22]) );
  DLH_X1 \IMMEDIATE_reg[21]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[21]) );
  DLH_X1 \IMMEDIATE_reg[20]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[20]) );
  DLH_X1 \IMMEDIATE_reg[19]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[19]) );
  DLH_X1 \IMMEDIATE_reg[18]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[18]) );
  DLH_X1 \IMMEDIATE_reg[17]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[17]) );
  DLH_X1 \IMMEDIATE_reg[16]  ( .G(CLK), .D(n33), .Q(IMMEDIATE[16]) );
  DLH_X1 \IMMEDIATE_reg[15]  ( .G(CLK), .D(n18), .Q(IMMEDIATE[15]) );
  DLH_X1 \IMMEDIATE_reg[14]  ( .G(CLK), .D(n17), .Q(IMMEDIATE[14]) );
  DLH_X1 \IMMEDIATE_reg[13]  ( .G(CLK), .D(n16), .Q(IMMEDIATE[13]) );
  DLH_X1 \IMMEDIATE_reg[12]  ( .G(CLK), .D(n15), .Q(IMMEDIATE[12]) );
  DLH_X1 \IMMEDIATE_reg[11]  ( .G(CLK), .D(n14), .Q(IMMEDIATE[11]) );
  DLH_X1 \IMMEDIATE_reg[10]  ( .G(CLK), .D(n13), .Q(IMMEDIATE[10]) );
  DLH_X1 \IMMEDIATE_reg[9]  ( .G(CLK), .D(n12), .Q(IMMEDIATE[9]) );
  DLH_X1 \IMMEDIATE_reg[8]  ( .G(CLK), .D(n11), .Q(IMMEDIATE[8]) );
  DLH_X1 \IMMEDIATE_reg[7]  ( .G(CLK), .D(n10), .Q(IMMEDIATE[7]) );
  DLH_X1 \IMMEDIATE_reg[6]  ( .G(CLK), .D(n9), .Q(IMMEDIATE[6]) );
  DLH_X1 \IMMEDIATE_reg[5]  ( .G(CLK), .D(n8), .Q(IMMEDIATE[5]) );
  DLH_X1 \IMMEDIATE_reg[4]  ( .G(CLK), .D(n7), .Q(IMMEDIATE[4]) );
  DLH_X1 \IMMEDIATE_reg[3]  ( .G(CLK), .D(n6), .Q(IMMEDIATE[3]) );
  DLH_X1 \IMMEDIATE_reg[2]  ( .G(CLK), .D(n5), .Q(IMMEDIATE[2]) );
  DLH_X1 \IMMEDIATE_reg[1]  ( .G(CLK), .D(n4), .Q(IMMEDIATE[1]) );
  DLH_X1 \IMMEDIATE_reg[0]  ( .G(CLK), .D(n3), .Q(IMMEDIATE[0]) );
  DLH_X1 \RS1_reg[4]  ( .G(CLK), .D(N137), .Q(RS1[4]) );
  DLH_X1 \RS1_reg[3]  ( .G(CLK), .D(N136), .Q(RS1[3]) );
  DLH_X1 \RS1_reg[2]  ( .G(CLK), .D(N135), .Q(RS1[2]) );
  DLH_X1 \RS1_reg[1]  ( .G(CLK), .D(N134), .Q(RS1[1]) );
  DLH_X1 \RS1_reg[0]  ( .G(CLK), .D(N133), .Q(RS1[0]) );
  DLH_X1 \RS2_reg[4]  ( .G(CLK), .D(N142), .Q(RS2[4]) );
  DLH_X1 \RS2_reg[3]  ( .G(CLK), .D(N141), .Q(RS2[3]) );
  DLH_X1 \RS2_reg[2]  ( .G(CLK), .D(N140), .Q(RS2[2]) );
  DLH_X1 \RS2_reg[1]  ( .G(CLK), .D(N139), .Q(RS2[1]) );
  DLH_X1 \RS2_reg[0]  ( .G(CLK), .D(N138), .Q(RS2[0]) );
  sign_eval_N_in5_N_out32 SIGN_EXTENSION_imm5 ( .IR_out(IR_26[15:11]), 
        .signed_val(is_signed) );
  sign_eval_N_in16_N_out32 SIGN_EXTENSION_imm16 ( .IR_out(IR_26[15:0]), 
        .signed_val(is_signed), .Immediate({IMMEDIATE_16[31], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, IMMEDIATE_16[15:0]}) );
  sign_eval_N_in26_N_out32 SIGN_EXTENSION_imm26 ( .IR_out({N137, N136, N135, 
        N134, N133, N142, N141, N140, N139, N138, IR_26[15:0]}), .signed_val(
        1'b0) );
  INV_X1 U3 ( .A(n31), .ZN(n20) );
  INV_X1 U4 ( .A(n31), .ZN(n21) );
  OR2_X2 U5 ( .A1(n29), .A2(n28), .ZN(n31) );
  OR2_X2 U6 ( .A1(n29), .A2(n28), .ZN(n22) );
  INV_X1 U7 ( .A(n30), .ZN(n33) );
  NOR2_X1 U8 ( .A1(OPCODE[5]), .A2(OPCODE[3]), .ZN(n25) );
  NAND2_X1 U9 ( .A1(n27), .A2(n26), .ZN(n28) );
  INV_X1 U10 ( .A(OPCODE[1]), .ZN(n26) );
  INV_X1 U11 ( .A(OPCODE[0]), .ZN(n27) );
  INV_X1 U12 ( .A(OPCODE[2]), .ZN(n23) );
  INV_X1 U13 ( .A(OPCODE[4]), .ZN(n24) );
  NAND3_X1 U14 ( .A1(n25), .A2(n24), .A3(n23), .ZN(n29) );
  AND2_X1 U15 ( .A1(IMMEDIATE_16[0]), .A2(n22), .ZN(n3) );
  AND2_X1 U16 ( .A1(IMMEDIATE_16[1]), .A2(n22), .ZN(n4) );
  AND2_X1 U17 ( .A1(IMMEDIATE_16[2]), .A2(n22), .ZN(n5) );
  AND2_X1 U18 ( .A1(IMMEDIATE_16[3]), .A2(n22), .ZN(n6) );
  AND2_X1 U19 ( .A1(IMMEDIATE_16[4]), .A2(n22), .ZN(n7) );
  AND2_X1 U20 ( .A1(IMMEDIATE_16[5]), .A2(n22), .ZN(n8) );
  AND2_X1 U21 ( .A1(IMMEDIATE_16[6]), .A2(n22), .ZN(n9) );
  AND2_X1 U22 ( .A1(IMMEDIATE_16[7]), .A2(n22), .ZN(n10) );
  AND2_X1 U23 ( .A1(IMMEDIATE_16[8]), .A2(n22), .ZN(n11) );
  AND2_X1 U24 ( .A1(IMMEDIATE_16[9]), .A2(n22), .ZN(n12) );
  AND2_X1 U25 ( .A1(IMMEDIATE_16[10]), .A2(n22), .ZN(n13) );
  AND2_X1 U26 ( .A1(IMMEDIATE_16[11]), .A2(n22), .ZN(n14) );
  AND2_X1 U27 ( .A1(IMMEDIATE_16[12]), .A2(n22), .ZN(n15) );
  AND2_X1 U28 ( .A1(IMMEDIATE_16[13]), .A2(n22), .ZN(n16) );
  AND2_X1 U29 ( .A1(IMMEDIATE_16[14]), .A2(n22), .ZN(n17) );
  AND2_X1 U30 ( .A1(IMMEDIATE_16[15]), .A2(n22), .ZN(n18) );
  NAND2_X1 U31 ( .A1(n31), .A2(IMMEDIATE_16[31]), .ZN(n30) );
  INV_X1 U32 ( .A(n31), .ZN(n32) );
  MUX2_X1 U33 ( .A(N138), .B(IR_26[11]), .S(n32), .Z(n38) );
  MUX2_X1 U34 ( .A(N139), .B(IR_26[12]), .S(n32), .Z(n37) );
  MUX2_X1 U35 ( .A(N140), .B(IR_26[13]), .S(n20), .Z(n36) );
  MUX2_X1 U36 ( .A(N141), .B(IR_26[14]), .S(n21), .Z(n35) );
  MUX2_X1 U37 ( .A(N142), .B(IR_26[15]), .S(n20), .Z(n34) );
endmodule


module windRF_M8_N8_F5_NBIT32 ( CLK, RESET, ENABLE, CALL, RETRN, FILL, SPILL, 
        BUSin, BUSout, RD1, RD2, WR, ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, 
        OUT2, wr_signal );
  input [31:0] BUSin;
  output [31:0] BUSout;
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, CALL, RETRN, RD1, RD2, WR, wr_signal;
  output FILL, SPILL;
  wire   N2167, N2168, N2169, N2170, N2171, N2172, N2173, N8431, N8432, N8433,
         N8434, N8435, N8436, N8437, N8575, N8576, N8577, N8578, N8579, N8580,
         N8581, N8702, N8703, N8704, N8705, N8706, N8707, N8708, N8709, N8710,
         N8711, N8712, N8713, N8714, N8715, N8716, N8717, N8718, N8719, N8720,
         N8721, N8722, N8723, N8724, N8725, N8726, N8727, N8728, N8729, N8730,
         N8731, N8732, N8733, N8734, N8735, N8736, N8737, N8738, N8739, N8740,
         N8741, N8742, N8743, N8744, N8745, N8746, N8747, N8748, N8749, N8750,
         N8751, N8752, N8753, N8754, N8755, N8756, N8757, N8758, N8759, N8760,
         N8761, N8762, N8763, N8764, N8765, N8766, N8767, \U3/U97/Z_4 ,
         \U3/U97/Z_5 , \U3/U97/Z_6 , \U3/U98/Z_4 , \U3/U98/Z_5 , \U3/U98/Z_6 ,
         \U3/U99/Z_4 , \U3/U99/Z_5 , \U3/U99/Z_6 , n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2935, n2936, n2937, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n141, n142, n143, n153, n154, n155, n165, n166, n167, n177,
         n178, n179, n189, n190, n191, n201, n202, n203, n213, n214, n215,
         n225, n226, n227, n237, n238, n239, n249, n250, n251, n261, n262,
         n263, n273, n274, n275, n285, n286, n287, n297, n298, n299, n309,
         n310, n311, n321, n322, n323, n333, n334, n335, n345, n346, n347,
         n357, n358, n359, n369, n370, n371, n381, n382, n383, n393, n394,
         n395, n405, n406, n407, n417, n418, n419, n429, n430, n431, n441,
         n442, n443, n453, n454, n455, n465, n466, n467, n477, n478, n479,
         n489, n490, n491, n501, n502, n503, n513, n514, n515, n868, n871,
         n872, n875, n876, n879, n880, n883, n884, n887, n888, n891, n892,
         n895, n896, n899, n900, n903, n904, n907, n908, n911, n912, n915,
         n916, n919, n920, n923, n924, n927, n928, n929, n931, n932, n933,
         n935, n936, n937, n939, n940, n941, n943, n944, n945, n947, n948,
         n949, n951, n952, n953, n955, n956, n957, n959, n960, n961, n963,
         n964, n965, n967, n968, n969, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1029, n1041, n1042, n1043, n1053, n1054, n1055, n1065, n1066,
         n1067, n1077, n1078, n1079, n1089, n1090, n1091, n1101, n1102, n1103,
         n1113, n1114, n1115, n1125, n1126, n1127, n1137, n1138, n1139, n1149,
         n1150, n1151, n1161, n1162, n1163, n1173, n1174, n1175, n1185, n1186,
         n1187, n1197, n1198, n1199, n1209, n1210, n1211, n1221, n1222, n1223,
         n1233, n1234, n1235, n1245, n1246, n1247, n1257, n1258, n1259, n1269,
         n1270, n1271, n1281, n1282, n1283, n1293, n1294, n1295, n1305, n1306,
         n1307, n1317, n1318, n1319, n1329, n1330, n1331, n1341, n1342, n1343,
         n1385, n1386, n1387, n1397, n1398, n1399, n1409, n1442, n1443, n1735,
         n1739, n1743, n1747, n1751, n1755, n1759, n1763, n1767, n1771, n1775,
         n1779, n1783, n1787, n1791, n1795, n1799, n1803, n1807, n1811, n1815,
         n1819, n1823, n1827, n1831, n1835, n1839, n1843, n1847, n1851, n1855,
         n1859, n1868, n1869, n1870, n1871, n1880, n1881, n1882, n1883, n1892,
         n1893, n1894, n1895, n1904, n1905, n1906, n1907, n1916, n1917, n1918,
         n1919, n1928, n1929, n1930, n1931, n1940, n1941, n1942, n1943, n1952,
         n1953, n1954, n1955, n1964, n1965, n1966, n1967, n1976, n1977, n1978,
         n1979, n1988, n1989, n1990, n1991, n2000, n2001, n2002, n2003, n2012,
         n2013, n2014, n2015, n2024, n2025, n2026, n2027, n2036, n2037, n2038,
         n2039, n2048, n2049, n2082, n2083, n2093, n2094, n2095, n2105, n2106,
         n2107, n2149, n2150, n2151, n2161, n2162, n2163, n2173, n2174, n2175,
         n2217, n2218, n2219, n2229, n2230, n2231, n2241, n2242, n2243, n2253,
         n2254, n2255, n2265, n2266, n2267, n2277, n2278, n2279, n2289, n2290,
         n2291, n2301, n2302, n2303, n2313, n2314, n2315, n2325, n2326, n2327,
         n2337, n2338, n2339, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2494, n2496, n2498, n2500, n2566, n2568, n2570, n2571, n2573,
         n2574, n2576, n2578, n2580, n2582, n2584, n2586, n2588, n2597, n2599,
         n2615, n2617, n2698, n2715, n2716, n2717, n2719, n2721, n2723, n2725,
         n2730, n2735, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6044, n6140, n6236, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9311, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9696,
         n9697, n9698, n9699, n9700, n9701, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, \r486/n4 ,
         \r486/carry[4] , \r486/carry[5] , \r486/A[3] , \r480/n4 ,
         \r480/carry[4] , \r480/carry[5] , \r480/A[3] , \r472/n4 ,
         \r472/carry[4] , \r472/carry[5] , \r472/B[3] , n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518;
  assign SPILL = 1'b0;
  assign BUSout[31] = 1'b0;
  assign BUSout[30] = 1'b0;
  assign BUSout[29] = 1'b0;
  assign BUSout[28] = 1'b0;
  assign BUSout[27] = 1'b0;
  assign BUSout[26] = 1'b0;
  assign BUSout[25] = 1'b0;
  assign BUSout[24] = 1'b0;
  assign BUSout[23] = 1'b0;
  assign BUSout[22] = 1'b0;
  assign BUSout[21] = 1'b0;
  assign BUSout[20] = 1'b0;
  assign BUSout[19] = 1'b0;
  assign BUSout[18] = 1'b0;
  assign BUSout[17] = 1'b0;
  assign BUSout[16] = 1'b0;
  assign BUSout[15] = 1'b0;
  assign BUSout[14] = 1'b0;
  assign BUSout[13] = 1'b0;
  assign BUSout[12] = 1'b0;
  assign BUSout[11] = 1'b0;
  assign BUSout[10] = 1'b0;
  assign BUSout[9] = 1'b0;
  assign BUSout[8] = 1'b0;
  assign BUSout[7] = 1'b0;
  assign BUSout[6] = 1'b0;
  assign BUSout[5] = 1'b0;
  assign BUSout[4] = 1'b0;
  assign BUSout[3] = 1'b0;
  assign BUSout[2] = 1'b0;
  assign BUSout[1] = 1'b0;
  assign BUSout[0] = 1'b0;
  assign N2167 = ADD_WR[0];
  assign N2168 = ADD_WR[1];
  assign N2169 = ADD_WR[2];
  assign N8431 = ADD_RD1[0];
  assign N8432 = ADD_RD1[1];
  assign N8433 = ADD_RD1[2];
  assign N8575 = ADD_RD2[0];
  assign N8576 = ADD_RD2[1];
  assign N8577 = ADD_RD2[2];
  assign FILL = 1'b0;

  DFFR_X1 \CWP_reg[6]  ( .D(n9132), .CK(CLK), .RN(n12662), .QN(n2935) );
  DFFR_X1 \CWP_reg[4]  ( .D(n12778), .CK(CLK), .RN(n12662), .Q(n10625), .QN(
        n2937) );
  DFFR_X1 \CWP_reg[5]  ( .D(n9133), .CK(CLK), .RN(n12662), .Q(n10626), .QN(
        n2936) );
  DFFR_X1 \REGISTERS_reg[0][31]  ( .D(n6316), .CK(CLK), .RN(n12655), .QN(n1871) );
  DFFR_X1 \REGISTERS_reg[0][30]  ( .D(n6317), .CK(CLK), .RN(n12618), .QN(n1883) );
  DFFR_X1 \REGISTERS_reg[0][29]  ( .D(n6318), .CK(CLK), .RN(n12604), .QN(n1895) );
  DFFR_X1 \REGISTERS_reg[0][28]  ( .D(n6319), .CK(CLK), .RN(n12611), .QN(n1907) );
  DFFR_X1 \REGISTERS_reg[0][27]  ( .D(n6320), .CK(CLK), .RN(n12582), .QN(n1919) );
  DFFR_X1 \REGISTERS_reg[0][26]  ( .D(n6321), .CK(CLK), .RN(n12560), .QN(n1931) );
  DFFR_X1 \REGISTERS_reg[0][25]  ( .D(n6322), .CK(CLK), .RN(n12538), .QN(n1943) );
  DFFR_X1 \REGISTERS_reg[0][24]  ( .D(n6323), .CK(CLK), .RN(n12512), .QN(n1955) );
  DFFR_X1 \REGISTERS_reg[0][23]  ( .D(n6324), .CK(CLK), .RN(n12626), .QN(n1967) );
  DFFR_X1 \REGISTERS_reg[0][22]  ( .D(n6325), .CK(CLK), .RN(n12485), .QN(n1979) );
  DFFR_X1 \REGISTERS_reg[0][21]  ( .D(n6326), .CK(CLK), .RN(n12523), .QN(n1991) );
  DFFR_X1 \REGISTERS_reg[0][20]  ( .D(n6327), .CK(CLK), .RN(n12498), .QN(n2003) );
  DFFR_X1 \REGISTERS_reg[0][19]  ( .D(n6328), .CK(CLK), .RN(n12589), .QN(n2015) );
  DFFR_X1 \REGISTERS_reg[0][18]  ( .D(n6329), .CK(CLK), .RN(n12440), .QN(n2027) );
  DFFR_X1 \REGISTERS_reg[0][17]  ( .D(n6330), .CK(CLK), .RN(n12447), .QN(n2039) );
  DFFR_X1 \REGISTERS_reg[0][16]  ( .D(n6331), .CK(CLK), .RN(n12499), .QN(n2083) );
  DFFR_X1 \REGISTERS_reg[0][15]  ( .D(n6332), .CK(CLK), .RN(n12633), .QN(n2095) );
  DFFR_X1 \REGISTERS_reg[0][14]  ( .D(n6333), .CK(CLK), .RN(n12461), .QN(n2107) );
  DFFR_X1 \REGISTERS_reg[0][13]  ( .D(n6334), .CK(CLK), .RN(n12468), .QN(n2151) );
  DFFR_X1 \REGISTERS_reg[0][12]  ( .D(n6335), .CK(CLK), .RN(n12476), .QN(n2163) );
  DFFR_X1 \REGISTERS_reg[0][11]  ( .D(n6336), .CK(CLK), .RN(n12567), .QN(n2175) );
  DFFR_X1 \REGISTERS_reg[0][10]  ( .D(n6337), .CK(CLK), .RN(n12545), .QN(n2219) );
  DFFR_X1 \REGISTERS_reg[0][9]  ( .D(n6338), .CK(CLK), .RN(n12552), .QN(n2231)
         );
  DFFR_X1 \REGISTERS_reg[0][8]  ( .D(n6339), .CK(CLK), .RN(n12530), .QN(n2243)
         );
  DFFR_X1 \REGISTERS_reg[0][7]  ( .D(n6340), .CK(CLK), .RN(n12640), .QN(n2255)
         );
  DFFR_X1 \REGISTERS_reg[0][6]  ( .D(n6341), .CK(CLK), .RN(n12596), .QN(n2267)
         );
  DFFR_X1 \REGISTERS_reg[0][5]  ( .D(n6342), .CK(CLK), .RN(n12483), .QN(n2279)
         );
  DFFR_X1 \REGISTERS_reg[0][4]  ( .D(n6343), .CK(CLK), .RN(n12490), .QN(n2291)
         );
  DFFR_X1 \REGISTERS_reg[0][3]  ( .D(n6344), .CK(CLK), .RN(n12574), .QN(n2303)
         );
  DFFR_X1 \REGISTERS_reg[0][2]  ( .D(n6345), .CK(CLK), .RN(n12505), .QN(n2315)
         );
  DFFR_X1 \REGISTERS_reg[0][1]  ( .D(n6346), .CK(CLK), .RN(n12433), .QN(n2327)
         );
  DFFR_X1 \REGISTERS_reg[0][0]  ( .D(n6347), .CK(CLK), .RN(n12648), .QN(n2339)
         );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n6348), .CK(CLK), .RN(n12655), .QN(n143)
         );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n6349), .CK(CLK), .RN(n12618), .QN(n155)
         );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n6350), .CK(CLK), .RN(n12604), .QN(n167)
         );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n6351), .CK(CLK), .RN(n12611), .QN(n179)
         );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n6352), .CK(CLK), .RN(n12582), .QN(n191)
         );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n6353), .CK(CLK), .RN(n12560), .QN(n203)
         );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n6354), .CK(CLK), .RN(n12538), .QN(n215)
         );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n6355), .CK(CLK), .RN(n12512), .QN(n227)
         );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n6356), .CK(CLK), .RN(n12626), .QN(n239)
         );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n6357), .CK(CLK), .RN(n12484), .QN(n251)
         );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n6358), .CK(CLK), .RN(n12523), .QN(n263)
         );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n6359), .CK(CLK), .RN(n12498), .QN(n275)
         );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n6360), .CK(CLK), .RN(n12589), .QN(n287)
         );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n6361), .CK(CLK), .RN(n12440), .QN(n299)
         );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n6362), .CK(CLK), .RN(n12447), .QN(n311)
         );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n6363), .CK(CLK), .RN(n12498), .QN(n323)
         );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n6364), .CK(CLK), .RN(n12633), .QN(n335)
         );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n6365), .CK(CLK), .RN(n12461), .QN(n347)
         );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n6366), .CK(CLK), .RN(n12468), .QN(n359)
         );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n6367), .CK(CLK), .RN(n12476), .QN(n371)
         );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n6368), .CK(CLK), .RN(n12567), .QN(n383)
         );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n6369), .CK(CLK), .RN(n12545), .QN(n395)
         );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n6370), .CK(CLK), .RN(n12552), .QN(n407)
         );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n6371), .CK(CLK), .RN(n12530), .QN(n419)
         );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n6372), .CK(CLK), .RN(n12640), .QN(n431)
         );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n6373), .CK(CLK), .RN(n12596), .QN(n443)
         );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n6374), .CK(CLK), .RN(n12483), .QN(n455)
         );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n6375), .CK(CLK), .RN(n12490), .QN(n467)
         );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n6376), .CK(CLK), .RN(n12574), .QN(n479)
         );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n6377), .CK(CLK), .RN(n12505), .QN(n491)
         );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n6378), .CK(CLK), .RN(n12433), .QN(n503)
         );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n6379), .CK(CLK), .RN(n12648), .QN(n515)
         );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n6380), .CK(CLK), .RN(n12655), .QN(
        n12780) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n6381), .CK(CLK), .RN(n12618), .QN(
        n12781) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n6382), .CK(CLK), .RN(n12604), .QN(
        n12782) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n6383), .CK(CLK), .RN(n12611), .QN(n1043) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n6384), .CK(CLK), .RN(n12582), .QN(n1055) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n6385), .CK(CLK), .RN(n12560), .QN(n1067) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n6386), .CK(CLK), .RN(n12538), .QN(n1079) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n6387), .CK(CLK), .RN(n12512), .QN(n1091) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n6388), .CK(CLK), .RN(n12626), .QN(n1103) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n6389), .CK(CLK), .RN(n12483), .QN(n1115) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n6390), .CK(CLK), .RN(n12523), .QN(n1127) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n6391), .CK(CLK), .RN(n12498), .QN(n1139) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n6392), .CK(CLK), .RN(n12589), .QN(n1151) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n6393), .CK(CLK), .RN(n12440), .QN(n1163) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n6394), .CK(CLK), .RN(n12447), .QN(n1175) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n6395), .CK(CLK), .RN(n12497), .QN(n1187) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n6396), .CK(CLK), .RN(n12633), .QN(n1199) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n6397), .CK(CLK), .RN(n12461), .QN(n1211) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n6398), .CK(CLK), .RN(n12468), .QN(n1223) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n6399), .CK(CLK), .RN(n12476), .QN(n1235) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n6400), .CK(CLK), .RN(n12567), .QN(n1247) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n6401), .CK(CLK), .RN(n12545), .QN(n1259) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n6402), .CK(CLK), .RN(n12552), .QN(n1271)
         );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n6403), .CK(CLK), .RN(n12530), .QN(n1283)
         );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n6404), .CK(CLK), .RN(n12640), .QN(n1295)
         );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n6405), .CK(CLK), .RN(n12596), .QN(n1307)
         );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n6406), .CK(CLK), .RN(n12483), .QN(n1319)
         );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n6407), .CK(CLK), .RN(n12490), .QN(n1331)
         );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n6408), .CK(CLK), .RN(n12574), .QN(n1343)
         );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n6409), .CK(CLK), .RN(n12505), .QN(n1387)
         );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n6410), .CK(CLK), .RN(n12433), .QN(n1399)
         );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n6411), .CK(CLK), .RN(n12648), .QN(n1443)
         );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n6412), .CK(CLK), .RN(n12655), .QN(n1870) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n6413), .CK(CLK), .RN(n12618), .QN(n1882) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n6414), .CK(CLK), .RN(n12604), .QN(n1894) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n6415), .CK(CLK), .RN(n12611), .QN(n1906) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n6416), .CK(CLK), .RN(n12582), .QN(n1918) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n6417), .CK(CLK), .RN(n12560), .QN(n1930) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n6418), .CK(CLK), .RN(n12538), .QN(n1942) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n6419), .CK(CLK), .RN(n12512), .QN(n1954) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n6420), .CK(CLK), .RN(n12626), .QN(n1966) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n6421), .CK(CLK), .RN(n12482), .QN(n1978) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n6422), .CK(CLK), .RN(n12523), .QN(n1990) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n6423), .CK(CLK), .RN(n12498), .QN(n2002) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n6424), .CK(CLK), .RN(n12589), .QN(n2014) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n6425), .CK(CLK), .RN(n12440), .QN(n2026) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n6426), .CK(CLK), .RN(n12447), .QN(n2038) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n6427), .CK(CLK), .RN(n12496), .QN(n2082) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n6428), .CK(CLK), .RN(n12633), .QN(n2094) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n6429), .CK(CLK), .RN(n12461), .QN(n2106) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n6430), .CK(CLK), .RN(n12468), .QN(n2150) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n6431), .CK(CLK), .RN(n12476), .QN(n2162) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n6432), .CK(CLK), .RN(n12567), .QN(n2174) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n6433), .CK(CLK), .RN(n12545), .QN(n2218) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n6434), .CK(CLK), .RN(n12552), .QN(n2230)
         );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n6435), .CK(CLK), .RN(n12530), .QN(n2242)
         );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n6436), .CK(CLK), .RN(n12640), .QN(n2254)
         );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n6437), .CK(CLK), .RN(n12596), .QN(n2266)
         );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n6438), .CK(CLK), .RN(n12483), .QN(n2278)
         );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n6439), .CK(CLK), .RN(n12490), .QN(n2290)
         );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n6440), .CK(CLK), .RN(n12574), .QN(n2302)
         );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n6441), .CK(CLK), .RN(n12505), .QN(n2314)
         );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n6442), .CK(CLK), .RN(n12433), .QN(n2326)
         );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n6443), .CK(CLK), .RN(n12648), .QN(n2338)
         );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n6444), .CK(CLK), .RN(n12655), .QN(n142)
         );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n6445), .CK(CLK), .RN(n12619), .QN(n154)
         );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n6446), .CK(CLK), .RN(n12604), .QN(n166)
         );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n6447), .CK(CLK), .RN(n12611), .QN(n178)
         );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n6448), .CK(CLK), .RN(n12582), .QN(n190)
         );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n6449), .CK(CLK), .RN(n12560), .QN(n202)
         );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n6450), .CK(CLK), .RN(n12538), .QN(n214)
         );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n6451), .CK(CLK), .RN(n12513), .QN(n226)
         );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n6452), .CK(CLK), .RN(n12626), .QN(n238)
         );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n6453), .CK(CLK), .RN(n12474), .QN(n250)
         );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n6454), .CK(CLK), .RN(n12523), .QN(n262)
         );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n6455), .CK(CLK), .RN(n12498), .QN(n274)
         );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n6456), .CK(CLK), .RN(n12589), .QN(n286)
         );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n6457), .CK(CLK), .RN(n12440), .QN(n298)
         );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n6458), .CK(CLK), .RN(n12448), .QN(n310)
         );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n6459), .CK(CLK), .RN(n12495), .QN(n322)
         );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n6460), .CK(CLK), .RN(n12633), .QN(n334)
         );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n6461), .CK(CLK), .RN(n12461), .QN(n346)
         );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n6462), .CK(CLK), .RN(n12469), .QN(n358)
         );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n6463), .CK(CLK), .RN(n12476), .QN(n370)
         );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n6464), .CK(CLK), .RN(n12567), .QN(n382)
         );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n6465), .CK(CLK), .RN(n12545), .QN(n394)
         );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n6466), .CK(CLK), .RN(n12553), .QN(n406)
         );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n6467), .CK(CLK), .RN(n12531), .QN(n418)
         );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n6468), .CK(CLK), .RN(n12641), .QN(n430)
         );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n6469), .CK(CLK), .RN(n12597), .QN(n442)
         );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n6470), .CK(CLK), .RN(n12483), .QN(n454)
         );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n6471), .CK(CLK), .RN(n12491), .QN(n466)
         );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n6472), .CK(CLK), .RN(n12575), .QN(n478)
         );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n6473), .CK(CLK), .RN(n12505), .QN(n490)
         );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n6474), .CK(CLK), .RN(n12433), .QN(n502)
         );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n6475), .CK(CLK), .RN(n12648), .QN(n514)
         );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n6476), .CK(CLK), .RN(n12655), .QN(
        n12783) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n6477), .CK(CLK), .RN(n12619), .QN(
        n12784) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n6478), .CK(CLK), .RN(n12604), .QN(
        n12785) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n6479), .CK(CLK), .RN(n12611), .QN(n1042) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n6480), .CK(CLK), .RN(n12582), .QN(n1054) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n6481), .CK(CLK), .RN(n12560), .QN(n1066) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n6482), .CK(CLK), .RN(n12538), .QN(n1078) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n6483), .CK(CLK), .RN(n12513), .QN(n1090) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n6484), .CK(CLK), .RN(n12626), .QN(n1102) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n6485), .CK(CLK), .RN(n12516), .QN(n1114) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n6486), .CK(CLK), .RN(n12523), .QN(n1126) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n6487), .CK(CLK), .RN(n12498), .QN(n1138) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n6488), .CK(CLK), .RN(n12589), .QN(n1150) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n6489), .CK(CLK), .RN(n12440), .QN(n1162) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n6490), .CK(CLK), .RN(n12448), .QN(n1174) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n6491), .CK(CLK), .RN(n12494), .QN(n1186) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n6492), .CK(CLK), .RN(n12633), .QN(n1198) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n6493), .CK(CLK), .RN(n12461), .QN(n1210) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n6494), .CK(CLK), .RN(n12469), .QN(n1222) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n6495), .CK(CLK), .RN(n12476), .QN(n1234) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n6496), .CK(CLK), .RN(n12567), .QN(n1246) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n6497), .CK(CLK), .RN(n12545), .QN(n1258) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n6498), .CK(CLK), .RN(n12553), .QN(n1270)
         );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n6499), .CK(CLK), .RN(n12531), .QN(n1282)
         );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n6500), .CK(CLK), .RN(n12641), .QN(n1294)
         );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n6501), .CK(CLK), .RN(n12597), .QN(n1306)
         );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n6502), .CK(CLK), .RN(n12483), .QN(n1318)
         );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n6503), .CK(CLK), .RN(n12491), .QN(n1330)
         );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n6504), .CK(CLK), .RN(n12575), .QN(n1342)
         );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n6505), .CK(CLK), .RN(n12505), .QN(n1386)
         );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n6506), .CK(CLK), .RN(n12433), .QN(n1398)
         );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n6507), .CK(CLK), .RN(n12648), .QN(n1442)
         );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n6508), .CK(CLK), .RN(n12655), .QN(n1869) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n6509), .CK(CLK), .RN(n12619), .QN(n1881) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n6510), .CK(CLK), .RN(n12604), .QN(n1893) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n6511), .CK(CLK), .RN(n12611), .QN(n1905) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n6512), .CK(CLK), .RN(n12582), .QN(n1917) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n6513), .CK(CLK), .RN(n12560), .QN(n1929) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n6514), .CK(CLK), .RN(n12538), .QN(n1941) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n6515), .CK(CLK), .RN(n12513), .QN(n1953) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n6516), .CK(CLK), .RN(n12626), .QN(n1965) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n6517), .CK(CLK), .RN(n12473), .QN(n1977) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n6518), .CK(CLK), .RN(n12523), .QN(n1989) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n6519), .CK(CLK), .RN(n12498), .QN(n2001) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n6520), .CK(CLK), .RN(n12589), .QN(n2013) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n6521), .CK(CLK), .RN(n12440), .QN(n2025) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n6522), .CK(CLK), .RN(n12448), .QN(n2037) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n6523), .CK(CLK), .RN(n12493), .QN(n2049) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n6524), .CK(CLK), .RN(n12633), .QN(n2093) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n6525), .CK(CLK), .RN(n12461), .QN(n2105) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n6526), .CK(CLK), .RN(n12469), .QN(n2149) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n6527), .CK(CLK), .RN(n12476), .QN(n2161) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n6528), .CK(CLK), .RN(n12567), .QN(n2173) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n6529), .CK(CLK), .RN(n12545), .QN(n2217) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n6530), .CK(CLK), .RN(n12553), .QN(n2229)
         );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n6531), .CK(CLK), .RN(n12531), .QN(n2241)
         );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n6532), .CK(CLK), .RN(n12641), .QN(n2253)
         );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n6533), .CK(CLK), .RN(n12597), .QN(n2265)
         );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n6534), .CK(CLK), .RN(n12483), .QN(n2277)
         );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n6535), .CK(CLK), .RN(n12491), .QN(n2289)
         );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n6536), .CK(CLK), .RN(n12575), .QN(n2301)
         );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n6537), .CK(CLK), .RN(n12505), .QN(n2313)
         );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n6538), .CK(CLK), .RN(n12433), .QN(n2325)
         );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n6539), .CK(CLK), .RN(n12648), .QN(n2337)
         );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n6540), .CK(CLK), .RN(n12655), .QN(n141)
         );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n6541), .CK(CLK), .RN(n12619), .QN(n153)
         );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n6542), .CK(CLK), .RN(n12604), .QN(n165)
         );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n6543), .CK(CLK), .RN(n12611), .QN(n177)
         );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n6544), .CK(CLK), .RN(n12582), .QN(n189)
         );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n6545), .CK(CLK), .RN(n12560), .QN(n201)
         );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n6546), .CK(CLK), .RN(n12538), .QN(n213)
         );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n6547), .CK(CLK), .RN(n12513), .QN(n225)
         );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n6548), .CK(CLK), .RN(n12626), .QN(n237)
         );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n6549), .CK(CLK), .RN(n12472), .QN(n249)
         );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n6550), .CK(CLK), .RN(n12523), .QN(n261)
         );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n6551), .CK(CLK), .RN(n12498), .QN(n273)
         );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n6552), .CK(CLK), .RN(n12589), .QN(n285)
         );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n6553), .CK(CLK), .RN(n12440), .QN(n297)
         );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n6554), .CK(CLK), .RN(n12448), .QN(n309)
         );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n6555), .CK(CLK), .RN(n12492), .QN(n321)
         );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n6556), .CK(CLK), .RN(n12633), .QN(n333)
         );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n6557), .CK(CLK), .RN(n12461), .QN(n345)
         );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n6558), .CK(CLK), .RN(n12469), .QN(n357)
         );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n6559), .CK(CLK), .RN(n12476), .QN(n369)
         );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n6560), .CK(CLK), .RN(n12567), .QN(n381)
         );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n6561), .CK(CLK), .RN(n12545), .QN(n393)
         );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n6562), .CK(CLK), .RN(n12553), .QN(n405)
         );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n6563), .CK(CLK), .RN(n12531), .QN(n417)
         );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n6564), .CK(CLK), .RN(n12641), .QN(n429)
         );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n6565), .CK(CLK), .RN(n12597), .QN(n441)
         );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n6566), .CK(CLK), .RN(n12483), .QN(n453)
         );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n6567), .CK(CLK), .RN(n12491), .QN(n465)
         );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n6568), .CK(CLK), .RN(n12575), .QN(n477)
         );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n6569), .CK(CLK), .RN(n12505), .QN(n489)
         );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n6570), .CK(CLK), .RN(n12433), .QN(n501)
         );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n6571), .CK(CLK), .RN(n12648), .QN(n513)
         );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n6572), .CK(CLK), .RN(n12656), .QN(
        n12786) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n6573), .CK(CLK), .RN(n12619), .QN(
        n12787) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n6574), .CK(CLK), .RN(n12604), .QN(n1029) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n6575), .CK(CLK), .RN(n12612), .QN(n1041) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n6576), .CK(CLK), .RN(n12582), .QN(n1053) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n6577), .CK(CLK), .RN(n12560), .QN(n1065) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n6578), .CK(CLK), .RN(n12538), .QN(n1077) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n6579), .CK(CLK), .RN(n12513), .QN(n1089) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n6580), .CK(CLK), .RN(n12626), .QN(n1101) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n6581), .CK(CLK), .RN(n12471), .QN(n1113) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n6582), .CK(CLK), .RN(n12524), .QN(n1125) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n6583), .CK(CLK), .RN(n12498), .QN(n1137) );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n6584), .CK(CLK), .RN(n12590), .QN(n1149) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n6585), .CK(CLK), .RN(n12441), .QN(n1161) );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n6586), .CK(CLK), .RN(n12448), .QN(n1173) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n6587), .CK(CLK), .RN(n12491), .QN(n1185) );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n6588), .CK(CLK), .RN(n12634), .QN(n1197) );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n6589), .CK(CLK), .RN(n12462), .QN(n1209) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n6590), .CK(CLK), .RN(n12469), .QN(n1221) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n6591), .CK(CLK), .RN(n12476), .QN(n1233) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n6592), .CK(CLK), .RN(n12568), .QN(n1245) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n6593), .CK(CLK), .RN(n12546), .QN(n1257) );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n6594), .CK(CLK), .RN(n12553), .QN(n1269)
         );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n6595), .CK(CLK), .RN(n12531), .QN(n1281)
         );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n6596), .CK(CLK), .RN(n12641), .QN(n1293)
         );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n6597), .CK(CLK), .RN(n12597), .QN(n1305)
         );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n6598), .CK(CLK), .RN(n12484), .QN(n1317)
         );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n6599), .CK(CLK), .RN(n12491), .QN(n1329)
         );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n6600), .CK(CLK), .RN(n12575), .QN(n1341)
         );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n6601), .CK(CLK), .RN(n12506), .QN(n1385)
         );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n6602), .CK(CLK), .RN(n12433), .QN(n1397)
         );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n6603), .CK(CLK), .RN(n12648), .QN(n1409)
         );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n6604), .CK(CLK), .RN(n12656), .QN(n871)
         );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n6605), .CK(CLK), .RN(n12619), .QN(n875)
         );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n6606), .CK(CLK), .RN(n12604), .QN(n879)
         );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n6607), .CK(CLK), .RN(n12612), .QN(n883)
         );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n6608), .CK(CLK), .RN(n12582), .QN(n887)
         );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n6609), .CK(CLK), .RN(n12560), .QN(n891)
         );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n6610), .CK(CLK), .RN(n12538), .QN(n895)
         );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n6611), .CK(CLK), .RN(n12513), .QN(n899)
         );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n6612), .CK(CLK), .RN(n12626), .QN(n903)
         );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n6613), .CK(CLK), .RN(n12470), .QN(n907)
         );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n6614), .CK(CLK), .RN(n12524), .QN(n911)
         );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n6615), .CK(CLK), .RN(n12498), .QN(n915)
         );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n6616), .CK(CLK), .RN(n12590), .QN(n919)
         );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n6617), .CK(CLK), .RN(n12441), .QN(n923)
         );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n6618), .CK(CLK), .RN(n12448), .QN(n927)
         );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n6619), .CK(CLK), .RN(n12490), .QN(n931)
         );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n6620), .CK(CLK), .RN(n12634), .QN(n935)
         );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n6621), .CK(CLK), .RN(n12462), .QN(n939)
         );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n6622), .CK(CLK), .RN(n12469), .QN(n943)
         );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n6623), .CK(CLK), .RN(n12476), .QN(n947)
         );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n6624), .CK(CLK), .RN(n12568), .QN(n951)
         );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n6625), .CK(CLK), .RN(n12546), .QN(n955)
         );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n6626), .CK(CLK), .RN(n12553), .QN(n959)
         );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n6627), .CK(CLK), .RN(n12531), .QN(n963)
         );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n6628), .CK(CLK), .RN(n12641), .QN(n967)
         );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n6629), .CK(CLK), .RN(n12597), .QN(n971)
         );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n6630), .CK(CLK), .RN(n12484), .QN(n975)
         );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n6631), .CK(CLK), .RN(n12491), .QN(n979)
         );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n6632), .CK(CLK), .RN(n12575), .QN(n983)
         );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n6633), .CK(CLK), .RN(n12506), .QN(n987)
         );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n6634), .CK(CLK), .RN(n12433), .QN(n991)
         );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n6635), .CK(CLK), .RN(n12648), .QN(n995)
         );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n6636), .CK(CLK), .RN(n12656), .QN(
        n1735) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n6637), .CK(CLK), .RN(n12619), .QN(
        n1739) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n6638), .CK(CLK), .RN(n12604), .QN(
        n1743) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n6639), .CK(CLK), .RN(n12612), .QN(
        n1747) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n6640), .CK(CLK), .RN(n12582), .QN(
        n1751) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n6641), .CK(CLK), .RN(n12560), .QN(
        n1755) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n6642), .CK(CLK), .RN(n12538), .QN(
        n1759) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n6643), .CK(CLK), .RN(n12513), .QN(
        n1763) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n6644), .CK(CLK), .RN(n12626), .QN(
        n1767) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n6645), .CK(CLK), .RN(n12486), .QN(
        n1771) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n6646), .CK(CLK), .RN(n12524), .QN(
        n1775) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n6647), .CK(CLK), .RN(n12498), .QN(
        n1779) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n6648), .CK(CLK), .RN(n12590), .QN(
        n1783) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n6649), .CK(CLK), .RN(n12441), .QN(
        n1787) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n6650), .CK(CLK), .RN(n12448), .QN(
        n1791) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n6651), .CK(CLK), .RN(n12500), .QN(
        n1795) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n6652), .CK(CLK), .RN(n12634), .QN(
        n1799) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n6653), .CK(CLK), .RN(n12462), .QN(
        n1803) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n6654), .CK(CLK), .RN(n12469), .QN(
        n1807) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n6655), .CK(CLK), .RN(n12476), .QN(
        n1811) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n6656), .CK(CLK), .RN(n12568), .QN(
        n1815) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n6657), .CK(CLK), .RN(n12546), .QN(
        n1819) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n6658), .CK(CLK), .RN(n12553), .QN(n1823) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n6659), .CK(CLK), .RN(n12531), .QN(n1827) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n6660), .CK(CLK), .RN(n12641), .QN(n1831) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n6661), .CK(CLK), .RN(n12597), .QN(n1835) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n6662), .CK(CLK), .RN(n12484), .QN(n1839) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n6663), .CK(CLK), .RN(n12491), .QN(n1843) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n6664), .CK(CLK), .RN(n12575), .QN(n1847) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n6665), .CK(CLK), .RN(n12506), .QN(n1851) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n6666), .CK(CLK), .RN(n12433), .QN(n1855) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n6667), .CK(CLK), .RN(n12648), .QN(n1859) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n6700), .CK(CLK), .RN(n12656), .QN(
        n5736) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n6701), .CK(CLK), .RN(n12619), .QN(
        n5768) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n6702), .CK(CLK), .RN(n12605), .QN(
        n5800) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n6703), .CK(CLK), .RN(n12612), .QN(
        n5832) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n6704), .CK(CLK), .RN(n12583), .QN(
        n5864) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n6705), .CK(CLK), .RN(n12561), .QN(
        n5896) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n6706), .CK(CLK), .RN(n12539), .QN(
        n5928) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n6707), .CK(CLK), .RN(n12513), .QN(
        n5992) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n6708), .CK(CLK), .RN(n12627), .QN(
        n6309) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n6709), .CK(CLK), .RN(n12517), .QN(
        n9159) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n6710), .CK(CLK), .RN(n12524), .QN(
        n9191) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n6711), .CK(CLK), .RN(n12499), .QN(
        n9255) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n6712), .CK(CLK), .RN(n12590), .QN(
        n9589) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n6713), .CK(CLK), .RN(n12441), .QN(
        n9621) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n6714), .CK(CLK), .RN(n12448), .QN(
        n9653) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n6715), .CK(CLK), .RN(n12455), .QN(
        n10015) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n6716), .CK(CLK), .RN(n12634), .QN(
        n10047) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n6717), .CK(CLK), .RN(n12462), .QN(
        n10079) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n6718), .CK(CLK), .RN(n12469), .QN(
        n10111) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n6719), .CK(CLK), .RN(n12477), .QN(
        n10143) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n6720), .CK(CLK), .RN(n12568), .QN(
        n10175) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n6721), .CK(CLK), .RN(n12546), .QN(
        n10209) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n6722), .CK(CLK), .RN(n12553), .QN(
        n10241) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n6723), .CK(CLK), .RN(n12531), .QN(
        n10273) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n6724), .CK(CLK), .RN(n12641), .QN(
        n10308) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n6725), .CK(CLK), .RN(n12597), .QN(
        n10340) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n6726), .CK(CLK), .RN(n12484), .QN(
        n10372) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n6727), .CK(CLK), .RN(n12491), .QN(
        n10407) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n6728), .CK(CLK), .RN(n12575), .QN(
        n10439) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n6729), .CK(CLK), .RN(n12506), .QN(
        n10471) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n6730), .CK(CLK), .RN(n12434), .QN(
        n10503) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n6731), .CK(CLK), .RN(n12649), .QN(
        n10535) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n6732), .CK(CLK), .RN(n12656), .QN(
        n5734) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n6733), .CK(CLK), .RN(n12619), .QN(
        n5766) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n6734), .CK(CLK), .RN(n12605), .QN(
        n5798) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n6735), .CK(CLK), .RN(n12612), .QN(
        n5830) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n6736), .CK(CLK), .RN(n12583), .QN(
        n5862) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n6737), .CK(CLK), .RN(n12561), .QN(
        n5894) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n6738), .CK(CLK), .RN(n12539), .QN(
        n5926) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n6739), .CK(CLK), .RN(n12513), .QN(
        n5990) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n6740), .CK(CLK), .RN(n12627), .QN(
        n6307) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n6741), .CK(CLK), .RN(n12517), .QN(
        n9157) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n6742), .CK(CLK), .RN(n12524), .QN(
        n9189) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n6743), .CK(CLK), .RN(n12499), .QN(
        n9253) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n6744), .CK(CLK), .RN(n12590), .QN(
        n9587) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n6745), .CK(CLK), .RN(n12441), .QN(
        n9619) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n6746), .CK(CLK), .RN(n12448), .QN(
        n9651) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n6747), .CK(CLK), .RN(n12455), .QN(
        n10013) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n6748), .CK(CLK), .RN(n12634), .QN(
        n10045) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n6749), .CK(CLK), .RN(n12462), .QN(
        n10077) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n6750), .CK(CLK), .RN(n12469), .QN(
        n10109) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n6751), .CK(CLK), .RN(n12477), .QN(
        n10141) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n6752), .CK(CLK), .RN(n12568), .QN(
        n10173) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n6753), .CK(CLK), .RN(n12546), .QN(
        n10205) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n6754), .CK(CLK), .RN(n12553), .QN(
        n10239) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n6755), .CK(CLK), .RN(n12531), .QN(
        n10271) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n6756), .CK(CLK), .RN(n12641), .QN(
        n10306) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n6757), .CK(CLK), .RN(n12597), .QN(
        n10338) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n6758), .CK(CLK), .RN(n12484), .QN(
        n10370) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n6759), .CK(CLK), .RN(n12491), .QN(
        n10405) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n6760), .CK(CLK), .RN(n12575), .QN(
        n10437) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n6761), .CK(CLK), .RN(n12506), .QN(
        n10469) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n6762), .CK(CLK), .RN(n12434), .QN(
        n10501) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n6763), .CK(CLK), .RN(n12649), .QN(
        n10533) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n6764), .CK(CLK), .RN(n12656), .QN(
        n5735) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n6765), .CK(CLK), .RN(n12619), .QN(
        n5767) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n6766), .CK(CLK), .RN(n12605), .QN(
        n5799) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n6767), .CK(CLK), .RN(n12612), .QN(
        n5831) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n6768), .CK(CLK), .RN(n12583), .QN(
        n5863) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n6769), .CK(CLK), .RN(n12561), .QN(
        n5895) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n6770), .CK(CLK), .RN(n12539), .QN(
        n5927) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n6771), .CK(CLK), .RN(n12513), .QN(
        n5991) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n6772), .CK(CLK), .RN(n12627), .QN(
        n6308) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n6773), .CK(CLK), .RN(n12517), .QN(
        n9158) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n6774), .CK(CLK), .RN(n12524), .QN(
        n9190) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n6775), .CK(CLK), .RN(n12499), .QN(
        n9254) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n6776), .CK(CLK), .RN(n12590), .QN(
        n9588) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n6777), .CK(CLK), .RN(n12441), .QN(
        n9620) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n6778), .CK(CLK), .RN(n12448), .QN(
        n9652) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n6779), .CK(CLK), .RN(n12455), .QN(
        n10014) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n6780), .CK(CLK), .RN(n12634), .QN(
        n10046) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n6781), .CK(CLK), .RN(n12462), .QN(
        n10078) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n6782), .CK(CLK), .RN(n12469), .QN(
        n10110) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n6783), .CK(CLK), .RN(n12477), .QN(
        n10142) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n6784), .CK(CLK), .RN(n12568), .QN(
        n10174) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n6785), .CK(CLK), .RN(n12546), .QN(
        n10208) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n6786), .CK(CLK), .RN(n12553), .QN(
        n10240) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n6787), .CK(CLK), .RN(n12531), .QN(
        n10272) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n6788), .CK(CLK), .RN(n12641), .QN(
        n10307) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n6789), .CK(CLK), .RN(n12597), .QN(
        n10339) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n6790), .CK(CLK), .RN(n12484), .QN(
        n10371) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n6791), .CK(CLK), .RN(n12491), .QN(
        n10406) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n6792), .CK(CLK), .RN(n12575), .QN(
        n10438) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n6793), .CK(CLK), .RN(n12506), .QN(
        n10470) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n6794), .CK(CLK), .RN(n12434), .QN(
        n10502) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n6795), .CK(CLK), .RN(n12649), .QN(
        n10534) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n7036), .CK(CLK), .RN(n12635), .Q(n9999), .QN(n13060) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n7037), .CK(CLK), .RN(n12463), .Q(n9998), .QN(n13061) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n7038), .CK(CLK), .RN(n12470), .Q(n9997), .QN(n13062) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n7039), .CK(CLK), .RN(n12477), .Q(n9996), .QN(n13063) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n7040), .CK(CLK), .RN(n12569), .Q(n9995), .QN(n13064) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n7041), .CK(CLK), .RN(n12547), .Q(n9994), .QN(n13065) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n7042), .CK(CLK), .RN(n12554), .Q(n9993), 
        .QN(n13066) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n7043), .CK(CLK), .RN(n12532), .Q(n9992), 
        .QN(n13067) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n7044), .CK(CLK), .RN(n12642), .Q(n9991), 
        .QN(n13068) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n7045), .CK(CLK), .RN(n12598), .Q(n9990), 
        .QN(n13069) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n7046), .CK(CLK), .RN(n12485), .Q(n9989), 
        .QN(n13070) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n7047), .CK(CLK), .RN(n12492), .Q(n9988), 
        .QN(n13071) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n7048), .CK(CLK), .RN(n12576), .Q(n9987), 
        .QN(n13072) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n7049), .CK(CLK), .RN(n12507), .Q(n9986), 
        .QN(n13073) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n7050), .CK(CLK), .RN(n12434), .Q(n9985), 
        .QN(n13074) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n7051), .CK(CLK), .RN(n12649), .Q(n9984), 
        .QN(n13075) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n7052), .CK(CLK), .RN(n12657), .Q(n9983), .QN(n13076) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n7053), .CK(CLK), .RN(n12620), .Q(n9982), .QN(n13077) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n7054), .CK(CLK), .RN(n12605), .Q(n9981), .QN(n13078) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n7055), .CK(CLK), .RN(n12613), .Q(n9980), .QN(n13079) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n7056), .CK(CLK), .RN(n12583), .Q(n9979), .QN(n13080) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n7057), .CK(CLK), .RN(n12561), .Q(n9978), .QN(n13081) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n7058), .CK(CLK), .RN(n12539), .Q(n9977), .QN(n13082) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n7059), .CK(CLK), .RN(n12514), .Q(n9976), .QN(n13083) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n7060), .CK(CLK), .RN(n12627), .Q(n9975), .QN(n13084) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n7061), .CK(CLK), .RN(n12517), .Q(n9974), .QN(n13085) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n7062), .CK(CLK), .RN(n12525), .Q(n9973), .QN(n13086) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n7063), .CK(CLK), .RN(n12499), .Q(n9972), .QN(n13087) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n7064), .CK(CLK), .RN(n12591), .Q(n9971), .QN(n13088) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n7065), .CK(CLK), .RN(n12442), .Q(n9970), .QN(n13089) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n7066), .CK(CLK), .RN(n12449), .Q(n9969), .QN(n13090) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n7067), .CK(CLK), .RN(n12455), .Q(n9968), .QN(n13091) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n7068), .CK(CLK), .RN(n12635), .Q(n9967), .QN(n13092) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n7069), .CK(CLK), .RN(n12463), .Q(n9966), .QN(n13093) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n7070), .CK(CLK), .RN(n12470), .Q(n9965), .QN(n13094) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n7071), .CK(CLK), .RN(n12477), .Q(n9964), .QN(n13095) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n7072), .CK(CLK), .RN(n12569), .Q(n9963), .QN(n13096) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n7073), .CK(CLK), .RN(n12547), .Q(n9962), .QN(n13097) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n7074), .CK(CLK), .RN(n12554), .Q(n9961), 
        .QN(n13098) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n7075), .CK(CLK), .RN(n12532), .Q(n9960), 
        .QN(n13099) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n7076), .CK(CLK), .RN(n12642), .Q(n9959), 
        .QN(n13100) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n7077), .CK(CLK), .RN(n12598), .Q(n9958), 
        .QN(n13101) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n7078), .CK(CLK), .RN(n12485), .Q(n9957), 
        .QN(n13102) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n7079), .CK(CLK), .RN(n12492), .Q(n9956), 
        .QN(n13103) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n7080), .CK(CLK), .RN(n12576), .Q(n9955), 
        .QN(n13104) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n7081), .CK(CLK), .RN(n12507), .Q(n9954), 
        .QN(n13105) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n7082), .CK(CLK), .RN(n12434), .Q(n9953), 
        .QN(n13106) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n7083), .CK(CLK), .RN(n12649), .Q(n9952), 
        .QN(n13107) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n7084), .CK(CLK), .RN(n12657), .QN(
        n13108) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n7085), .CK(CLK), .RN(n12620), .QN(
        n13109) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n7086), .CK(CLK), .RN(n12606), .QN(
        n13110) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n7087), .CK(CLK), .RN(n12613), .QN(
        n13111) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n7088), .CK(CLK), .RN(n12584), .QN(
        n13112) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n7089), .CK(CLK), .RN(n12562), .QN(
        n13113) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n7090), .CK(CLK), .RN(n12540), .QN(
        n13114) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n7091), .CK(CLK), .RN(n12514), .QN(
        n13115) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n7092), .CK(CLK), .RN(n12628), .QN(
        n13116) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n7093), .CK(CLK), .RN(n12518), .QN(
        n13117) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n7094), .CK(CLK), .RN(n12525), .QN(
        n13118) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n7095), .CK(CLK), .RN(n12500), .QN(
        n13119) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n7096), .CK(CLK), .RN(n12591), .QN(
        n13120) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n7097), .CK(CLK), .RN(n12442), .QN(
        n13121) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n7098), .CK(CLK), .RN(n12449), .QN(
        n13122) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n7099), .CK(CLK), .RN(n12456), .QN(
        n13123) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n7100), .CK(CLK), .RN(n12635), .QN(
        n13124) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n7101), .CK(CLK), .RN(n12463), .QN(
        n13125) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n7102), .CK(CLK), .RN(n12470), .QN(
        n13126) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n7103), .CK(CLK), .RN(n12478), .QN(
        n13127) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n7104), .CK(CLK), .RN(n12569), .QN(
        n13128) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n7105), .CK(CLK), .RN(n12547), .QN(
        n13129) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n7106), .CK(CLK), .RN(n12554), .QN(
        n13130) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n7107), .CK(CLK), .RN(n12532), .QN(
        n13131) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n7108), .CK(CLK), .RN(n12642), .QN(
        n13132) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n7109), .CK(CLK), .RN(n12598), .QN(
        n13133) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n7110), .CK(CLK), .RN(n12485), .QN(
        n13134) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n7111), .CK(CLK), .RN(n12492), .QN(
        n13135) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n7112), .CK(CLK), .RN(n12576), .QN(
        n13136) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n7113), .CK(CLK), .RN(n12507), .QN(
        n13137) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n7114), .CK(CLK), .RN(n12435), .QN(
        n13138) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n7115), .CK(CLK), .RN(n12650), .QN(
        n13139) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n7116), .CK(CLK), .RN(n12657), .QN(
        n13140) );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n7117), .CK(CLK), .RN(n12620), .QN(
        n13141) );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n7118), .CK(CLK), .RN(n12606), .QN(
        n13142) );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n7119), .CK(CLK), .RN(n12613), .QN(
        n13143) );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n7120), .CK(CLK), .RN(n12584), .QN(
        n13144) );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n7121), .CK(CLK), .RN(n12562), .QN(
        n13145) );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n7122), .CK(CLK), .RN(n12540), .QN(
        n13146) );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n7123), .CK(CLK), .RN(n12514), .QN(
        n13147) );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n7124), .CK(CLK), .RN(n12628), .QN(
        n13148) );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n7125), .CK(CLK), .RN(n12518), .QN(
        n13149) );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n7126), .CK(CLK), .RN(n12525), .QN(
        n13150) );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n7127), .CK(CLK), .RN(n12500), .QN(
        n13151) );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n7128), .CK(CLK), .RN(n12591), .QN(
        n13152) );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n7129), .CK(CLK), .RN(n12442), .QN(
        n13153) );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n7130), .CK(CLK), .RN(n12449), .QN(
        n13154) );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n7131), .CK(CLK), .RN(n12456), .QN(
        n13155) );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n7132), .CK(CLK), .RN(n12635), .QN(
        n13156) );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n7133), .CK(CLK), .RN(n12463), .QN(
        n13157) );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n7134), .CK(CLK), .RN(n12470), .QN(
        n13158) );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n7135), .CK(CLK), .RN(n12478), .QN(
        n13159) );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n7136), .CK(CLK), .RN(n12569), .QN(
        n13160) );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n7137), .CK(CLK), .RN(n12547), .QN(
        n13161) );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n7138), .CK(CLK), .RN(n12554), .QN(
        n13162) );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n7139), .CK(CLK), .RN(n12532), .QN(
        n13163) );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n7140), .CK(CLK), .RN(n12642), .QN(
        n13164) );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n7141), .CK(CLK), .RN(n12598), .QN(
        n13165) );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n7142), .CK(CLK), .RN(n12485), .QN(
        n13166) );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n7143), .CK(CLK), .RN(n12492), .QN(
        n13167) );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n7144), .CK(CLK), .RN(n12576), .QN(
        n13168) );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n7145), .CK(CLK), .RN(n12507), .QN(
        n13169) );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n7146), .CK(CLK), .RN(n12435), .QN(
        n13170) );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n7147), .CK(CLK), .RN(n12650), .QN(
        n13171) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n7148), .CK(CLK), .RN(n12657), .QN(
        n13172) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n7149), .CK(CLK), .RN(n12620), .QN(
        n13173) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n7150), .CK(CLK), .RN(n12606), .QN(
        n13174) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n7151), .CK(CLK), .RN(n12613), .QN(
        n13175) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n7152), .CK(CLK), .RN(n12584), .QN(
        n13176) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n7153), .CK(CLK), .RN(n12562), .QN(
        n13177) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n7154), .CK(CLK), .RN(n12540), .QN(
        n13178) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n7155), .CK(CLK), .RN(n12514), .QN(
        n13179) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n7156), .CK(CLK), .RN(n12628), .QN(
        n13180) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n7157), .CK(CLK), .RN(n12518), .QN(
        n13181) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n7158), .CK(CLK), .RN(n12525), .QN(
        n13182) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n7159), .CK(CLK), .RN(n12500), .QN(
        n13183) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n7160), .CK(CLK), .RN(n12591), .QN(
        n13184) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n7161), .CK(CLK), .RN(n12442), .QN(
        n13185) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n7162), .CK(CLK), .RN(n12449), .QN(
        n13186) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n7163), .CK(CLK), .RN(n12456), .QN(
        n13187) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n7164), .CK(CLK), .RN(n12635), .QN(
        n13188) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n7165), .CK(CLK), .RN(n12463), .QN(
        n13189) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n7166), .CK(CLK), .RN(n12470), .QN(
        n13190) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n7167), .CK(CLK), .RN(n12478), .QN(
        n13191) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n7168), .CK(CLK), .RN(n12569), .QN(
        n13192) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n7169), .CK(CLK), .RN(n12547), .QN(
        n13193) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n7170), .CK(CLK), .RN(n12554), .QN(
        n13194) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n7171), .CK(CLK), .RN(n12532), .QN(
        n13195) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n7172), .CK(CLK), .RN(n12642), .QN(
        n13196) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n7173), .CK(CLK), .RN(n12598), .QN(
        n13197) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n7174), .CK(CLK), .RN(n12485), .QN(
        n13198) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n7175), .CK(CLK), .RN(n12492), .QN(
        n13199) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n7176), .CK(CLK), .RN(n12576), .QN(
        n13200) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n7177), .CK(CLK), .RN(n12507), .QN(
        n13201) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n7178), .CK(CLK), .RN(n12435), .QN(
        n13202) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n7179), .CK(CLK), .RN(n12650), .QN(
        n13203) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n7180), .CK(CLK), .RN(n12657), .Q(n9855), .QN(n13204) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n7181), .CK(CLK), .RN(n12620), .Q(n9854), .QN(n13205) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n7182), .CK(CLK), .RN(n12606), .Q(n9853), .QN(n13206) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n7183), .CK(CLK), .RN(n12613), .Q(n9852), .QN(n13207) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n7184), .CK(CLK), .RN(n12584), .Q(n9851), .QN(n13208) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n7185), .CK(CLK), .RN(n12562), .Q(n9850), .QN(n13209) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n7186), .CK(CLK), .RN(n12540), .Q(n9849), .QN(n13210) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n7187), .CK(CLK), .RN(n12514), .Q(n9848), .QN(n13211) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n7188), .CK(CLK), .RN(n12628), .Q(n9847), .QN(n13212) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n7189), .CK(CLK), .RN(n12518), .Q(n9846), .QN(n13213) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n7190), .CK(CLK), .RN(n12525), .Q(n9845), .QN(n13214) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n7191), .CK(CLK), .RN(n12500), .Q(n9844), .QN(n13215) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n7192), .CK(CLK), .RN(n12591), .Q(n9843), .QN(n13216) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n7193), .CK(CLK), .RN(n12442), .Q(n9842), .QN(n13217) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n7194), .CK(CLK), .RN(n12449), .Q(n9841), .QN(n13218) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n7195), .CK(CLK), .RN(n12456), .Q(n9840), .QN(n13219) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n7196), .CK(CLK), .RN(n12635), .Q(n9839), .QN(n13220) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n7197), .CK(CLK), .RN(n12463), .Q(n9838), .QN(n13221) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n7198), .CK(CLK), .RN(n12470), .Q(n9837), .QN(n13222) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n7199), .CK(CLK), .RN(n12478), .Q(n9836), .QN(n13223) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n7200), .CK(CLK), .RN(n12569), .Q(n9835), .QN(n13224) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n7201), .CK(CLK), .RN(n12547), .Q(n9834), .QN(n13225) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n7202), .CK(CLK), .RN(n12554), .Q(n9833), 
        .QN(n13226) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n7203), .CK(CLK), .RN(n12532), .Q(n9832), 
        .QN(n13227) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n7204), .CK(CLK), .RN(n12642), .Q(n9831), 
        .QN(n13228) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n7205), .CK(CLK), .RN(n12598), .Q(n9830), 
        .QN(n13229) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n7206), .CK(CLK), .RN(n12485), .Q(n9829), 
        .QN(n13230) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n7207), .CK(CLK), .RN(n12492), .Q(n9828), 
        .QN(n13231) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n7208), .CK(CLK), .RN(n12576), .Q(n9827), 
        .QN(n13232) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n7209), .CK(CLK), .RN(n12507), .Q(n9826), 
        .QN(n13233) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n7210), .CK(CLK), .RN(n12435), .Q(n9825), 
        .QN(n13234) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n7211), .CK(CLK), .RN(n12650), .Q(n9824), 
        .QN(n13235) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n7212), .CK(CLK), .RN(n12657), .Q(n9823), .QN(n13236) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n7213), .CK(CLK), .RN(n12621), .Q(n9822), .QN(n13237) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n7214), .CK(CLK), .RN(n12606), .Q(n9821), .QN(n13238) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n7215), .CK(CLK), .RN(n12613), .Q(n9820), .QN(n13239) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n7216), .CK(CLK), .RN(n12584), .Q(n9819), .QN(n13240) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n7217), .CK(CLK), .RN(n12562), .Q(n9818), .QN(n13241) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n7218), .CK(CLK), .RN(n12540), .Q(n9817), .QN(n13242) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n7219), .CK(CLK), .RN(n12515), .Q(n9816), .QN(n13243) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n7220), .CK(CLK), .RN(n12628), .Q(n9815), .QN(n13244) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n7221), .CK(CLK), .RN(n12518), .Q(n9814), .QN(n13245) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n7222), .CK(CLK), .RN(n12525), .Q(n9813), .QN(n13246) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n7223), .CK(CLK), .RN(n12500), .Q(n9812), .QN(n13247) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n7224), .CK(CLK), .RN(n12591), .Q(n9811), .QN(n13248) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n7225), .CK(CLK), .RN(n12442), .Q(n9810), .QN(n13249) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n7226), .CK(CLK), .RN(n12450), .Q(n9809), .QN(n13250) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n7227), .CK(CLK), .RN(n12456), .Q(n9808), .QN(n13251) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n7228), .CK(CLK), .RN(n12635), .Q(n9807), .QN(n13252) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n7229), .CK(CLK), .RN(n12463), .Q(n9806), .QN(n13253) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n7230), .CK(CLK), .RN(n12471), .Q(n9805), .QN(n13254) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n7231), .CK(CLK), .RN(n12478), .Q(n9804), .QN(n13255) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n7232), .CK(CLK), .RN(n12569), .Q(n9803), .QN(n13256) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n7233), .CK(CLK), .RN(n12547), .Q(n9802), .QN(n13257) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n7234), .CK(CLK), .RN(n12555), .Q(n9801), 
        .QN(n13258) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n7235), .CK(CLK), .RN(n12533), .Q(n9800), 
        .QN(n13259) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n7236), .CK(CLK), .RN(n12643), .Q(n9799), 
        .QN(n13260) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n7237), .CK(CLK), .RN(n12599), .Q(n9798), 
        .QN(n13261) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n7238), .CK(CLK), .RN(n12485), .Q(n9797), 
        .QN(n13262) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n7239), .CK(CLK), .RN(n12493), .Q(n9796), 
        .QN(n13263) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n7240), .CK(CLK), .RN(n12577), .Q(n9795), 
        .QN(n13264) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n7241), .CK(CLK), .RN(n12507), .Q(n9794), 
        .QN(n13265) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n7242), .CK(CLK), .RN(n12435), .Q(n9793), 
        .QN(n13266) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n7243), .CK(CLK), .RN(n12650), .Q(n9792), 
        .QN(n13267) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n7244), .CK(CLK), .RN(n12657), .Q(n9791), .QN(n13268) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n7245), .CK(CLK), .RN(n12621), .Q(n9790), .QN(n13269) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n7246), .CK(CLK), .RN(n12606), .Q(n9789), .QN(n13270) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n7247), .CK(CLK), .RN(n12613), .Q(n9788), .QN(n13271) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n7248), .CK(CLK), .RN(n12584), .Q(n9787), .QN(n13272) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n7249), .CK(CLK), .RN(n12562), .Q(n9786), .QN(n13273) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n7250), .CK(CLK), .RN(n12540), .Q(n9785), .QN(n13274) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n7251), .CK(CLK), .RN(n12515), .Q(n9784), .QN(n13275) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n7252), .CK(CLK), .RN(n12628), .Q(n9783), .QN(n13276) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n7253), .CK(CLK), .RN(n12518), .Q(n9782), .QN(n13277) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n7254), .CK(CLK), .RN(n12525), .Q(n9781), .QN(n13278) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n7255), .CK(CLK), .RN(n12500), .Q(n9780), .QN(n13279) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n7256), .CK(CLK), .RN(n12591), .Q(n9779), .QN(n13280) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n7257), .CK(CLK), .RN(n12442), .Q(n9778), .QN(n13281) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n7258), .CK(CLK), .RN(n12450), .Q(n9777), .QN(n13282) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n7259), .CK(CLK), .RN(n12456), .Q(n9776), .QN(n13283) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n7260), .CK(CLK), .RN(n12635), .Q(n9775), .QN(n13284) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n7261), .CK(CLK), .RN(n12463), .Q(n9774), .QN(n13285) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n7262), .CK(CLK), .RN(n12471), .Q(n9773), .QN(n13286) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n7263), .CK(CLK), .RN(n12478), .Q(n9772), .QN(n13287) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n7264), .CK(CLK), .RN(n12569), .Q(n9771), .QN(n13288) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n7265), .CK(CLK), .RN(n12547), .Q(n9770), .QN(n13289) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n7266), .CK(CLK), .RN(n12555), .Q(n9769), 
        .QN(n13290) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n7267), .CK(CLK), .RN(n12533), .Q(n9768), 
        .QN(n13291) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n7268), .CK(CLK), .RN(n12643), .Q(n9767), 
        .QN(n13292) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n7269), .CK(CLK), .RN(n12599), .Q(n9766), 
        .QN(n13293) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n7270), .CK(CLK), .RN(n12485), .Q(n9765), 
        .QN(n13294) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n7271), .CK(CLK), .RN(n12493), .Q(n9764), 
        .QN(n13295) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n7272), .CK(CLK), .RN(n12577), .Q(n9763), 
        .QN(n13296) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n7273), .CK(CLK), .RN(n12507), .Q(n9762), 
        .QN(n13297) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n7274), .CK(CLK), .RN(n12435), .Q(n9761), 
        .QN(n13298) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n7275), .CK(CLK), .RN(n12650), .Q(n9760), 
        .QN(n13299) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n7276), .CK(CLK), .RN(n12657), .Q(n9759), .QN(n13300) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n7277), .CK(CLK), .RN(n12621), .Q(n9758), .QN(n13301) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n7278), .CK(CLK), .RN(n12606), .Q(n9757), .QN(n13302) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n7279), .CK(CLK), .RN(n12613), .Q(n9756), .QN(n13303) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n7280), .CK(CLK), .RN(n12584), .Q(n9755), .QN(n13304) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n7281), .CK(CLK), .RN(n12562), .Q(n9754), .QN(n13305) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n7282), .CK(CLK), .RN(n12540), .Q(n9753), .QN(n13306) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n7283), .CK(CLK), .RN(n12515), .Q(n9752), .QN(n13307) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n7284), .CK(CLK), .RN(n12628), .Q(n9751), .QN(n13308) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n7285), .CK(CLK), .RN(n12518), .Q(n9750), .QN(n13309) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n7286), .CK(CLK), .RN(n12525), .Q(n9749), .QN(n13310) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n7287), .CK(CLK), .RN(n12500), .Q(n9748), .QN(n13311) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n7288), .CK(CLK), .RN(n12591), .Q(n9747), .QN(n13312) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n7289), .CK(CLK), .RN(n12442), .Q(n9746), .QN(n13313) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n7290), .CK(CLK), .RN(n12450), .Q(n9745), .QN(n13314) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n7291), .CK(CLK), .RN(n12456), .Q(n9744), .QN(n13315) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n7292), .CK(CLK), .RN(n12635), .Q(n9743), .QN(n13316) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n7293), .CK(CLK), .RN(n12463), .Q(n9742), .QN(n13317) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n7294), .CK(CLK), .RN(n12471), .Q(n9741), .QN(n13318) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n7295), .CK(CLK), .RN(n12478), .Q(n9740), .QN(n13319) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n7296), .CK(CLK), .RN(n12569), .Q(n9739), .QN(n13320) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n7297), .CK(CLK), .RN(n12547), .Q(n9738), .QN(n13321) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n7298), .CK(CLK), .RN(n12555), .Q(n9737), 
        .QN(n13322) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n7299), .CK(CLK), .RN(n12533), .Q(n9736), 
        .QN(n13323) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n7300), .CK(CLK), .RN(n12643), .Q(n9735), 
        .QN(n13324) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n7301), .CK(CLK), .RN(n12599), .Q(n9734), 
        .QN(n13325) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n7302), .CK(CLK), .RN(n12485), .Q(n9733), 
        .QN(n13326) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n7303), .CK(CLK), .RN(n12493), .Q(n9732), 
        .QN(n13327) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n7304), .CK(CLK), .RN(n12577), .Q(n9731), 
        .QN(n13328) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n7305), .CK(CLK), .RN(n12507), .Q(n9730), 
        .QN(n13329) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n7306), .CK(CLK), .RN(n12435), .Q(n9729), 
        .QN(n13330) );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n7307), .CK(CLK), .RN(n12650), .Q(n9728), 
        .QN(n13331) );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n7308), .CK(CLK), .RN(n12657), .Q(n9727), .QN(n13332) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n7309), .CK(CLK), .RN(n12621), .Q(n9726), .QN(n13333) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n7310), .CK(CLK), .RN(n12606), .Q(n9725), .QN(n13334) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n7311), .CK(CLK), .RN(n12613), .Q(n9724), .QN(n13335) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n7312), .CK(CLK), .RN(n12584), .Q(n9723), .QN(n13336) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n7313), .CK(CLK), .RN(n12562), .Q(n9722), .QN(n13337) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n7314), .CK(CLK), .RN(n12540), .Q(n9721), .QN(n13338) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n7315), .CK(CLK), .RN(n12515), .Q(n9720), .QN(n13339) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n7316), .CK(CLK), .RN(n12628), .Q(n9719), .QN(n13340) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n7317), .CK(CLK), .RN(n12518), .Q(n9718), .QN(n13341) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n7318), .CK(CLK), .RN(n12525), .Q(n9717), .QN(n13342) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n7319), .CK(CLK), .RN(n12500), .Q(n9716), .QN(n13343) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n7320), .CK(CLK), .RN(n12591), .Q(n9715), .QN(n13344) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n7321), .CK(CLK), .RN(n12442), .Q(n9714), .QN(n13345) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n7322), .CK(CLK), .RN(n12450), .Q(n9713), .QN(n13346) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n7323), .CK(CLK), .RN(n12456), .Q(n9712), .QN(n13347) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n7324), .CK(CLK), .RN(n12635), .Q(n9711), .QN(n13348) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n7325), .CK(CLK), .RN(n12463), .Q(n9710), .QN(n13349) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n7326), .CK(CLK), .RN(n12471), .Q(n9709), .QN(n13350) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n7327), .CK(CLK), .RN(n12478), .Q(n9708), .QN(n13351) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n7328), .CK(CLK), .RN(n12569), .Q(n9707), .QN(n13352) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n7329), .CK(CLK), .RN(n12547), .Q(n9706), .QN(n13353) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n7330), .CK(CLK), .RN(n12555), .Q(n9705), 
        .QN(n13354) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n7331), .CK(CLK), .RN(n12533), .Q(n9704), 
        .QN(n13355) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n7332), .CK(CLK), .RN(n12643), .Q(n9703), 
        .QN(n13356) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n7333), .CK(CLK), .RN(n12599), .Q(n9702), 
        .QN(n13357) );
  DFFR_X1 \REGISTERS_reg[32][31]  ( .D(n7340), .CK(CLK), .RN(n12658), .Q(n9695), .QN(n13364) );
  DFFR_X1 \REGISTERS_reg[32][30]  ( .D(n7341), .CK(CLK), .RN(n12621), .Q(n9694), .QN(n13365) );
  DFFR_X1 \REGISTERS_reg[32][29]  ( .D(n7342), .CK(CLK), .RN(n12606), .Q(n9693), .QN(n13366) );
  DFFR_X1 \REGISTERS_reg[32][28]  ( .D(n7343), .CK(CLK), .RN(n12614), .Q(n9692), .QN(n13367) );
  DFFR_X1 \REGISTERS_reg[32][27]  ( .D(n7344), .CK(CLK), .RN(n12584), .Q(n9691), .QN(n13368) );
  DFFR_X1 \REGISTERS_reg[32][26]  ( .D(n7345), .CK(CLK), .RN(n12562), .Q(n9690), .QN(n13369) );
  DFFR_X1 \REGISTERS_reg[32][25]  ( .D(n7346), .CK(CLK), .RN(n12540), .Q(n9689), .QN(n13370) );
  DFFR_X1 \REGISTERS_reg[32][24]  ( .D(n7347), .CK(CLK), .RN(n12515), .Q(n9688), .QN(n13371) );
  DFFR_X1 \REGISTERS_reg[32][23]  ( .D(n7348), .CK(CLK), .RN(n12628), .Q(n9687), .QN(n13372) );
  DFFR_X1 \REGISTERS_reg[32][22]  ( .D(n7349), .CK(CLK), .RN(n12518), .Q(n9686), .QN(n13373) );
  DFFR_X1 \REGISTERS_reg[32][21]  ( .D(n7350), .CK(CLK), .RN(n12526), .Q(n9685), .QN(n13374) );
  DFFR_X1 \REGISTERS_reg[32][20]  ( .D(n7351), .CK(CLK), .RN(n12500), .Q(n9684), .QN(n13375) );
  DFFR_X1 \REGISTERS_reg[32][19]  ( .D(n7352), .CK(CLK), .RN(n12592), .Q(n9683), .QN(n13376) );
  DFFR_X1 \REGISTERS_reg[32][18]  ( .D(n7353), .CK(CLK), .RN(n12443), .Q(n9682), .QN(n13377) );
  DFFR_X1 \REGISTERS_reg[32][17]  ( .D(n7354), .CK(CLK), .RN(n12450), .Q(n9681), .QN(n13378) );
  DFFR_X1 \REGISTERS_reg[32][16]  ( .D(n7355), .CK(CLK), .RN(n12456), .Q(n9680), .QN(n13379) );
  DFFR_X1 \REGISTERS_reg[32][15]  ( .D(n7356), .CK(CLK), .RN(n12636), .Q(n9679), .QN(n13380) );
  DFFR_X1 \REGISTERS_reg[32][14]  ( .D(n7357), .CK(CLK), .RN(n12464), .Q(n9678), .QN(n13381) );
  DFFR_X1 \REGISTERS_reg[32][13]  ( .D(n7358), .CK(CLK), .RN(n12471), .Q(n9677), .QN(n13382) );
  DFFR_X1 \REGISTERS_reg[32][12]  ( .D(n7359), .CK(CLK), .RN(n12478), .Q(n9676), .QN(n13383) );
  DFFR_X1 \REGISTERS_reg[32][11]  ( .D(n7360), .CK(CLK), .RN(n12570), .Q(n9675), .QN(n13384) );
  DFFR_X1 \REGISTERS_reg[32][10]  ( .D(n7361), .CK(CLK), .RN(n12548), .Q(n9674), .QN(n13385) );
  DFFR_X1 \REGISTERS_reg[32][9]  ( .D(n7362), .CK(CLK), .RN(n12555), .Q(n9673), 
        .QN(n13386) );
  DFFR_X1 \REGISTERS_reg[32][8]  ( .D(n7363), .CK(CLK), .RN(n12533), .Q(n9672), 
        .QN(n13387) );
  DFFR_X1 \REGISTERS_reg[32][7]  ( .D(n7364), .CK(CLK), .RN(n12643), .Q(n9671), 
        .QN(n13388) );
  DFFR_X1 \REGISTERS_reg[32][6]  ( .D(n7365), .CK(CLK), .RN(n12599), .Q(n9670), 
        .QN(n13389) );
  DFFR_X1 \REGISTERS_reg[32][5]  ( .D(n7366), .CK(CLK), .RN(n12486), .Q(n9669), 
        .QN(n13390) );
  DFFR_X1 \REGISTERS_reg[32][4]  ( .D(n7367), .CK(CLK), .RN(n12493), .Q(n9668), 
        .QN(n13391) );
  DFFR_X1 \REGISTERS_reg[32][3]  ( .D(n7368), .CK(CLK), .RN(n12577), .Q(n9667), 
        .QN(n13392) );
  DFFR_X1 \REGISTERS_reg[32][2]  ( .D(n7369), .CK(CLK), .RN(n12508), .Q(n9666), 
        .QN(n13393) );
  DFFR_X1 \REGISTERS_reg[32][1]  ( .D(n7370), .CK(CLK), .RN(n12435), .Q(n9665), 
        .QN(n13394) );
  DFFR_X1 \REGISTERS_reg[32][0]  ( .D(n7371), .CK(CLK), .RN(n12650), .Q(n9664), 
        .QN(n13395) );
  DFFR_X1 \REGISTERS_reg[33][31]  ( .D(n7372), .CK(CLK), .RN(n12658), .QN(
        n5729) );
  DFFR_X1 \REGISTERS_reg[33][30]  ( .D(n7373), .CK(CLK), .RN(n12621), .QN(
        n5761) );
  DFFR_X1 \REGISTERS_reg[33][29]  ( .D(n7374), .CK(CLK), .RN(n12606), .QN(
        n5793) );
  DFFR_X1 \REGISTERS_reg[33][28]  ( .D(n7375), .CK(CLK), .RN(n12614), .QN(
        n5825) );
  DFFR_X1 \REGISTERS_reg[33][27]  ( .D(n7376), .CK(CLK), .RN(n12584), .QN(
        n5857) );
  DFFR_X1 \REGISTERS_reg[33][26]  ( .D(n7377), .CK(CLK), .RN(n12562), .QN(
        n5889) );
  DFFR_X1 \REGISTERS_reg[33][25]  ( .D(n7378), .CK(CLK), .RN(n12540), .QN(
        n5921) );
  DFFR_X1 \REGISTERS_reg[33][24]  ( .D(n7379), .CK(CLK), .RN(n12515), .QN(
        n5985) );
  DFFR_X1 \REGISTERS_reg[33][23]  ( .D(n7380), .CK(CLK), .RN(n12628), .QN(
        n6302) );
  DFFR_X1 \REGISTERS_reg[33][22]  ( .D(n7381), .CK(CLK), .RN(n12518), .QN(
        n9152) );
  DFFR_X1 \REGISTERS_reg[33][21]  ( .D(n7382), .CK(CLK), .RN(n12526), .QN(
        n9184) );
  DFFR_X1 \REGISTERS_reg[33][20]  ( .D(n7383), .CK(CLK), .RN(n12500), .QN(
        n9248) );
  DFFR_X1 \REGISTERS_reg[33][19]  ( .D(n7384), .CK(CLK), .RN(n12592), .QN(
        n9582) );
  DFFR_X1 \REGISTERS_reg[33][18]  ( .D(n7385), .CK(CLK), .RN(n12443), .QN(
        n9614) );
  DFFR_X1 \REGISTERS_reg[33][17]  ( .D(n7386), .CK(CLK), .RN(n12450), .QN(
        n9646) );
  DFFR_X1 \REGISTERS_reg[33][16]  ( .D(n7387), .CK(CLK), .RN(n12456), .QN(
        n10008) );
  DFFR_X1 \REGISTERS_reg[33][15]  ( .D(n7388), .CK(CLK), .RN(n12636), .QN(
        n10040) );
  DFFR_X1 \REGISTERS_reg[33][14]  ( .D(n7389), .CK(CLK), .RN(n12464), .QN(
        n10072) );
  DFFR_X1 \REGISTERS_reg[33][13]  ( .D(n7390), .CK(CLK), .RN(n12471), .QN(
        n10104) );
  DFFR_X1 \REGISTERS_reg[33][12]  ( .D(n7391), .CK(CLK), .RN(n12478), .QN(
        n10136) );
  DFFR_X1 \REGISTERS_reg[33][11]  ( .D(n7392), .CK(CLK), .RN(n12570), .QN(
        n10168) );
  DFFR_X1 \REGISTERS_reg[33][10]  ( .D(n7393), .CK(CLK), .RN(n12548), .QN(
        n10200) );
  DFFR_X1 \REGISTERS_reg[33][9]  ( .D(n7394), .CK(CLK), .RN(n12555), .QN(
        n10234) );
  DFFR_X1 \REGISTERS_reg[33][8]  ( .D(n7395), .CK(CLK), .RN(n12533), .QN(
        n10266) );
  DFFR_X1 \REGISTERS_reg[33][7]  ( .D(n7396), .CK(CLK), .RN(n12643), .QN(
        n10298) );
  DFFR_X1 \REGISTERS_reg[33][6]  ( .D(n7397), .CK(CLK), .RN(n12599), .QN(
        n10333) );
  DFFR_X1 \REGISTERS_reg[33][5]  ( .D(n7398), .CK(CLK), .RN(n12486), .QN(
        n10365) );
  DFFR_X1 \REGISTERS_reg[33][4]  ( .D(n7399), .CK(CLK), .RN(n12493), .QN(
        n10400) );
  DFFR_X1 \REGISTERS_reg[33][3]  ( .D(n7400), .CK(CLK), .RN(n12577), .QN(
        n10432) );
  DFFR_X1 \REGISTERS_reg[33][2]  ( .D(n7401), .CK(CLK), .RN(n12508), .QN(
        n10464) );
  DFFR_X1 \REGISTERS_reg[33][1]  ( .D(n7402), .CK(CLK), .RN(n12435), .QN(
        n10496) );
  DFFR_X1 \REGISTERS_reg[33][0]  ( .D(n7403), .CK(CLK), .RN(n12650), .QN(
        n10528) );
  DFFR_X1 \REGISTERS_reg[34][31]  ( .D(n7404), .CK(CLK), .RN(n12658), .QN(
        n5728) );
  DFFR_X1 \REGISTERS_reg[34][30]  ( .D(n7405), .CK(CLK), .RN(n12621), .QN(
        n5760) );
  DFFR_X1 \REGISTERS_reg[34][29]  ( .D(n7406), .CK(CLK), .RN(n12606), .QN(
        n5792) );
  DFFR_X1 \REGISTERS_reg[34][28]  ( .D(n7407), .CK(CLK), .RN(n12614), .QN(
        n5824) );
  DFFR_X1 \REGISTERS_reg[34][27]  ( .D(n7408), .CK(CLK), .RN(n12584), .QN(
        n5856) );
  DFFR_X1 \REGISTERS_reg[34][26]  ( .D(n7409), .CK(CLK), .RN(n12562), .QN(
        n5888) );
  DFFR_X1 \REGISTERS_reg[34][25]  ( .D(n7410), .CK(CLK), .RN(n12540), .QN(
        n5920) );
  DFFR_X1 \REGISTERS_reg[34][24]  ( .D(n7411), .CK(CLK), .RN(n12515), .QN(
        n5984) );
  DFFR_X1 \REGISTERS_reg[34][23]  ( .D(n7412), .CK(CLK), .RN(n12628), .QN(
        n6301) );
  DFFR_X1 \REGISTERS_reg[34][22]  ( .D(n7413), .CK(CLK), .RN(n12518), .QN(
        n9151) );
  DFFR_X1 \REGISTERS_reg[34][21]  ( .D(n7414), .CK(CLK), .RN(n12526), .QN(
        n9183) );
  DFFR_X1 \REGISTERS_reg[34][20]  ( .D(n7415), .CK(CLK), .RN(n12500), .QN(
        n9215) );
  DFFR_X1 \REGISTERS_reg[34][19]  ( .D(n7416), .CK(CLK), .RN(n12592), .QN(
        n9581) );
  DFFR_X1 \REGISTERS_reg[34][18]  ( .D(n7417), .CK(CLK), .RN(n12443), .QN(
        n9613) );
  DFFR_X1 \REGISTERS_reg[34][17]  ( .D(n7418), .CK(CLK), .RN(n12450), .QN(
        n9645) );
  DFFR_X1 \REGISTERS_reg[34][16]  ( .D(n7419), .CK(CLK), .RN(n12456), .QN(
        n10007) );
  DFFR_X1 \REGISTERS_reg[34][15]  ( .D(n7420), .CK(CLK), .RN(n12636), .QN(
        n10039) );
  DFFR_X1 \REGISTERS_reg[34][14]  ( .D(n7421), .CK(CLK), .RN(n12464), .QN(
        n10071) );
  DFFR_X1 \REGISTERS_reg[34][13]  ( .D(n7422), .CK(CLK), .RN(n12471), .QN(
        n10103) );
  DFFR_X1 \REGISTERS_reg[34][12]  ( .D(n7423), .CK(CLK), .RN(n12478), .QN(
        n10135) );
  DFFR_X1 \REGISTERS_reg[34][11]  ( .D(n7424), .CK(CLK), .RN(n12570), .QN(
        n10167) );
  DFFR_X1 \REGISTERS_reg[34][10]  ( .D(n7425), .CK(CLK), .RN(n12548), .QN(
        n10199) );
  DFFR_X1 \REGISTERS_reg[34][9]  ( .D(n7426), .CK(CLK), .RN(n12555), .QN(
        n10233) );
  DFFR_X1 \REGISTERS_reg[34][8]  ( .D(n7427), .CK(CLK), .RN(n12533), .QN(
        n10265) );
  DFFR_X1 \REGISTERS_reg[34][7]  ( .D(n7428), .CK(CLK), .RN(n12643), .QN(
        n10297) );
  DFFR_X1 \REGISTERS_reg[34][6]  ( .D(n7429), .CK(CLK), .RN(n12599), .QN(
        n10332) );
  DFFR_X1 \REGISTERS_reg[34][5]  ( .D(n7430), .CK(CLK), .RN(n12486), .QN(
        n10364) );
  DFFR_X1 \REGISTERS_reg[34][4]  ( .D(n7431), .CK(CLK), .RN(n12493), .QN(
        n10396) );
  DFFR_X1 \REGISTERS_reg[34][3]  ( .D(n7432), .CK(CLK), .RN(n12577), .QN(
        n10431) );
  DFFR_X1 \REGISTERS_reg[34][2]  ( .D(n7433), .CK(CLK), .RN(n12508), .QN(
        n10463) );
  DFFR_X1 \REGISTERS_reg[34][1]  ( .D(n7434), .CK(CLK), .RN(n12435), .QN(
        n10495) );
  DFFR_X1 \REGISTERS_reg[34][0]  ( .D(n7435), .CK(CLK), .RN(n12650), .QN(
        n10527) );
  DFFR_X1 \REGISTERS_reg[35][31]  ( .D(n7436), .CK(CLK), .RN(n12658), .QN(
        n5726) );
  DFFR_X1 \REGISTERS_reg[35][30]  ( .D(n7437), .CK(CLK), .RN(n12621), .QN(
        n5758) );
  DFFR_X1 \REGISTERS_reg[35][29]  ( .D(n7438), .CK(CLK), .RN(n12606), .QN(
        n5790) );
  DFFR_X1 \REGISTERS_reg[35][28]  ( .D(n7439), .CK(CLK), .RN(n12614), .QN(
        n5822) );
  DFFR_X1 \REGISTERS_reg[35][27]  ( .D(n7440), .CK(CLK), .RN(n12584), .QN(
        n5854) );
  DFFR_X1 \REGISTERS_reg[35][26]  ( .D(n7441), .CK(CLK), .RN(n12562), .QN(
        n5886) );
  DFFR_X1 \REGISTERS_reg[35][25]  ( .D(n7442), .CK(CLK), .RN(n12540), .QN(
        n5918) );
  DFFR_X1 \REGISTERS_reg[35][24]  ( .D(n7443), .CK(CLK), .RN(n12515), .QN(
        n5982) );
  DFFR_X1 \REGISTERS_reg[35][23]  ( .D(n7444), .CK(CLK), .RN(n12628), .QN(
        n6140) );
  DFFR_X1 \REGISTERS_reg[35][22]  ( .D(n7445), .CK(CLK), .RN(n12518), .QN(
        n9149) );
  DFFR_X1 \REGISTERS_reg[35][21]  ( .D(n7446), .CK(CLK), .RN(n12526), .QN(
        n9181) );
  DFFR_X1 \REGISTERS_reg[35][20]  ( .D(n7447), .CK(CLK), .RN(n12500), .QN(
        n9213) );
  DFFR_X1 \REGISTERS_reg[35][19]  ( .D(n7448), .CK(CLK), .RN(n12592), .QN(
        n9579) );
  DFFR_X1 \REGISTERS_reg[35][18]  ( .D(n7449), .CK(CLK), .RN(n12443), .QN(
        n9611) );
  DFFR_X1 \REGISTERS_reg[35][17]  ( .D(n7450), .CK(CLK), .RN(n12450), .QN(
        n9643) );
  DFFR_X1 \REGISTERS_reg[35][16]  ( .D(n7451), .CK(CLK), .RN(n12456), .QN(
        n10005) );
  DFFR_X1 \REGISTERS_reg[35][15]  ( .D(n7452), .CK(CLK), .RN(n12636), .QN(
        n10037) );
  DFFR_X1 \REGISTERS_reg[35][14]  ( .D(n7453), .CK(CLK), .RN(n12464), .QN(
        n10069) );
  DFFR_X1 \REGISTERS_reg[35][13]  ( .D(n7454), .CK(CLK), .RN(n12471), .QN(
        n10101) );
  DFFR_X1 \REGISTERS_reg[35][12]  ( .D(n7455), .CK(CLK), .RN(n12478), .QN(
        n10133) );
  DFFR_X1 \REGISTERS_reg[35][11]  ( .D(n7456), .CK(CLK), .RN(n12570), .QN(
        n10165) );
  DFFR_X1 \REGISTERS_reg[35][10]  ( .D(n7457), .CK(CLK), .RN(n12548), .QN(
        n10197) );
  DFFR_X1 \REGISTERS_reg[35][9]  ( .D(n7458), .CK(CLK), .RN(n12555), .QN(
        n10231) );
  DFFR_X1 \REGISTERS_reg[35][8]  ( .D(n7459), .CK(CLK), .RN(n12533), .QN(
        n10263) );
  DFFR_X1 \REGISTERS_reg[35][7]  ( .D(n7460), .CK(CLK), .RN(n12643), .QN(
        n10295) );
  DFFR_X1 \REGISTERS_reg[35][6]  ( .D(n7461), .CK(CLK), .RN(n12599), .QN(
        n10330) );
  DFFR_X1 \REGISTERS_reg[35][5]  ( .D(n7462), .CK(CLK), .RN(n12486), .QN(
        n10362) );
  DFFR_X1 \REGISTERS_reg[35][4]  ( .D(n7463), .CK(CLK), .RN(n12493), .QN(
        n10394) );
  DFFR_X1 \REGISTERS_reg[35][3]  ( .D(n7464), .CK(CLK), .RN(n12577), .QN(
        n10429) );
  DFFR_X1 \REGISTERS_reg[35][2]  ( .D(n7465), .CK(CLK), .RN(n12508), .QN(
        n10461) );
  DFFR_X1 \REGISTERS_reg[35][1]  ( .D(n7466), .CK(CLK), .RN(n12435), .QN(
        n10493) );
  DFFR_X1 \REGISTERS_reg[35][0]  ( .D(n7467), .CK(CLK), .RN(n12650), .QN(
        n10525) );
  DFFR_X1 \REGISTERS_reg[36][31]  ( .D(n7468), .CK(CLK), .RN(n12658), .QN(
        n5727) );
  DFFR_X1 \REGISTERS_reg[36][30]  ( .D(n7469), .CK(CLK), .RN(n12621), .QN(
        n5759) );
  DFFR_X1 \REGISTERS_reg[36][29]  ( .D(n7470), .CK(CLK), .RN(n12607), .QN(
        n5791) );
  DFFR_X1 \REGISTERS_reg[36][28]  ( .D(n7471), .CK(CLK), .RN(n12614), .QN(
        n5823) );
  DFFR_X1 \REGISTERS_reg[36][27]  ( .D(n7472), .CK(CLK), .RN(n12585), .QN(
        n5855) );
  DFFR_X1 \REGISTERS_reg[36][26]  ( .D(n7473), .CK(CLK), .RN(n12563), .QN(
        n5887) );
  DFFR_X1 \REGISTERS_reg[36][25]  ( .D(n7474), .CK(CLK), .RN(n12541), .QN(
        n5919) );
  DFFR_X1 \REGISTERS_reg[36][24]  ( .D(n7475), .CK(CLK), .RN(n12515), .QN(
        n5983) );
  DFFR_X1 \REGISTERS_reg[36][23]  ( .D(n7476), .CK(CLK), .RN(n12629), .QN(
        n6236) );
  DFFR_X1 \REGISTERS_reg[36][22]  ( .D(n7477), .CK(CLK), .RN(n12519), .QN(
        n9150) );
  DFFR_X1 \REGISTERS_reg[36][21]  ( .D(n7478), .CK(CLK), .RN(n12526), .QN(
        n9182) );
  DFFR_X1 \REGISTERS_reg[36][20]  ( .D(n7479), .CK(CLK), .RN(n12501), .QN(
        n9214) );
  DFFR_X1 \REGISTERS_reg[36][19]  ( .D(n7480), .CK(CLK), .RN(n12592), .QN(
        n9580) );
  DFFR_X1 \REGISTERS_reg[36][18]  ( .D(n7481), .CK(CLK), .RN(n12443), .QN(
        n9612) );
  DFFR_X1 \REGISTERS_reg[36][17]  ( .D(n7482), .CK(CLK), .RN(n12450), .QN(
        n9644) );
  DFFR_X1 \REGISTERS_reg[36][16]  ( .D(n7483), .CK(CLK), .RN(n12457), .QN(
        n10006) );
  DFFR_X1 \REGISTERS_reg[36][15]  ( .D(n7484), .CK(CLK), .RN(n12636), .QN(
        n10038) );
  DFFR_X1 \REGISTERS_reg[36][14]  ( .D(n7485), .CK(CLK), .RN(n12464), .QN(
        n10070) );
  DFFR_X1 \REGISTERS_reg[36][13]  ( .D(n7486), .CK(CLK), .RN(n12471), .QN(
        n10102) );
  DFFR_X1 \REGISTERS_reg[36][12]  ( .D(n7487), .CK(CLK), .RN(n12479), .QN(
        n10134) );
  DFFR_X1 \REGISTERS_reg[36][11]  ( .D(n7488), .CK(CLK), .RN(n12570), .QN(
        n10166) );
  DFFR_X1 \REGISTERS_reg[36][10]  ( .D(n7489), .CK(CLK), .RN(n12548), .QN(
        n10198) );
  DFFR_X1 \REGISTERS_reg[36][9]  ( .D(n7490), .CK(CLK), .RN(n12555), .QN(
        n10232) );
  DFFR_X1 \REGISTERS_reg[36][8]  ( .D(n7491), .CK(CLK), .RN(n12533), .QN(
        n10264) );
  DFFR_X1 \REGISTERS_reg[36][7]  ( .D(n7492), .CK(CLK), .RN(n12643), .QN(
        n10296) );
  DFFR_X1 \REGISTERS_reg[36][6]  ( .D(n7493), .CK(CLK), .RN(n12599), .QN(
        n10331) );
  DFFR_X1 \REGISTERS_reg[36][5]  ( .D(n7494), .CK(CLK), .RN(n12486), .QN(
        n10363) );
  DFFR_X1 \REGISTERS_reg[36][4]  ( .D(n7495), .CK(CLK), .RN(n12493), .QN(
        n10395) );
  DFFR_X1 \REGISTERS_reg[36][3]  ( .D(n7496), .CK(CLK), .RN(n12577), .QN(
        n10430) );
  DFFR_X1 \REGISTERS_reg[36][2]  ( .D(n7497), .CK(CLK), .RN(n12508), .QN(
        n10462) );
  DFFR_X1 \REGISTERS_reg[36][1]  ( .D(n7498), .CK(CLK), .RN(n12436), .QN(
        n10494) );
  DFFR_X1 \REGISTERS_reg[36][0]  ( .D(n7499), .CK(CLK), .RN(n12651), .QN(
        n10526) );
  DFFR_X1 \REGISTERS_reg[37][31]  ( .D(n7500), .CK(CLK), .RN(n12658), .QN(
        n5725) );
  DFFR_X1 \REGISTERS_reg[37][30]  ( .D(n7501), .CK(CLK), .RN(n12621), .QN(
        n5757) );
  DFFR_X1 \REGISTERS_reg[37][29]  ( .D(n7502), .CK(CLK), .RN(n12607), .QN(
        n5789) );
  DFFR_X1 \REGISTERS_reg[37][28]  ( .D(n7503), .CK(CLK), .RN(n12614), .QN(
        n5821) );
  DFFR_X1 \REGISTERS_reg[37][27]  ( .D(n7504), .CK(CLK), .RN(n12585), .QN(
        n5853) );
  DFFR_X1 \REGISTERS_reg[37][26]  ( .D(n7505), .CK(CLK), .RN(n12563), .QN(
        n5885) );
  DFFR_X1 \REGISTERS_reg[37][25]  ( .D(n7506), .CK(CLK), .RN(n12541), .QN(
        n5917) );
  DFFR_X1 \REGISTERS_reg[37][24]  ( .D(n7507), .CK(CLK), .RN(n12515), .QN(
        n5981) );
  DFFR_X1 \REGISTERS_reg[37][23]  ( .D(n7508), .CK(CLK), .RN(n12629), .QN(
        n6044) );
  DFFR_X1 \REGISTERS_reg[37][22]  ( .D(n7509), .CK(CLK), .RN(n12519), .QN(
        n9148) );
  DFFR_X1 \REGISTERS_reg[37][21]  ( .D(n7510), .CK(CLK), .RN(n12526), .QN(
        n9180) );
  DFFR_X1 \REGISTERS_reg[37][20]  ( .D(n7511), .CK(CLK), .RN(n12501), .QN(
        n9212) );
  DFFR_X1 \REGISTERS_reg[37][19]  ( .D(n7512), .CK(CLK), .RN(n12592), .QN(
        n9578) );
  DFFR_X1 \REGISTERS_reg[37][18]  ( .D(n7513), .CK(CLK), .RN(n12443), .QN(
        n9610) );
  DFFR_X1 \REGISTERS_reg[37][17]  ( .D(n7514), .CK(CLK), .RN(n12450), .QN(
        n9642) );
  DFFR_X1 \REGISTERS_reg[37][16]  ( .D(n7515), .CK(CLK), .RN(n12457), .QN(
        n10004) );
  DFFR_X1 \REGISTERS_reg[37][15]  ( .D(n7516), .CK(CLK), .RN(n12636), .QN(
        n10036) );
  DFFR_X1 \REGISTERS_reg[37][14]  ( .D(n7517), .CK(CLK), .RN(n12464), .QN(
        n10068) );
  DFFR_X1 \REGISTERS_reg[37][13]  ( .D(n7518), .CK(CLK), .RN(n12471), .QN(
        n10100) );
  DFFR_X1 \REGISTERS_reg[37][12]  ( .D(n7519), .CK(CLK), .RN(n12479), .QN(
        n10132) );
  DFFR_X1 \REGISTERS_reg[37][11]  ( .D(n7520), .CK(CLK), .RN(n12570), .QN(
        n10164) );
  DFFR_X1 \REGISTERS_reg[37][10]  ( .D(n7521), .CK(CLK), .RN(n12548), .QN(
        n10196) );
  DFFR_X1 \REGISTERS_reg[37][9]  ( .D(n7522), .CK(CLK), .RN(n12555), .QN(
        n10230) );
  DFFR_X1 \REGISTERS_reg[37][8]  ( .D(n7523), .CK(CLK), .RN(n12533), .QN(
        n10262) );
  DFFR_X1 \REGISTERS_reg[37][7]  ( .D(n7524), .CK(CLK), .RN(n12643), .QN(
        n10294) );
  DFFR_X1 \REGISTERS_reg[37][6]  ( .D(n7525), .CK(CLK), .RN(n12599), .QN(
        n10329) );
  DFFR_X1 \REGISTERS_reg[37][5]  ( .D(n7526), .CK(CLK), .RN(n12486), .QN(
        n10361) );
  DFFR_X1 \REGISTERS_reg[37][4]  ( .D(n7527), .CK(CLK), .RN(n12493), .QN(
        n10393) );
  DFFR_X1 \REGISTERS_reg[37][3]  ( .D(n7528), .CK(CLK), .RN(n12577), .QN(
        n10428) );
  DFFR_X1 \REGISTERS_reg[37][2]  ( .D(n7529), .CK(CLK), .RN(n12508), .QN(
        n10460) );
  DFFR_X1 \REGISTERS_reg[37][1]  ( .D(n7530), .CK(CLK), .RN(n12436), .QN(
        n10492) );
  DFFR_X1 \REGISTERS_reg[37][0]  ( .D(n7531), .CK(CLK), .RN(n12651), .QN(
        n10524) );
  DFFR_X1 \REGISTERS_reg[38][31]  ( .D(n7532), .CK(CLK), .RN(n12658), .QN(
        n5723) );
  DFFR_X1 \REGISTERS_reg[38][30]  ( .D(n7533), .CK(CLK), .RN(n12621), .QN(
        n5755) );
  DFFR_X1 \REGISTERS_reg[38][29]  ( .D(n7534), .CK(CLK), .RN(n12607), .QN(
        n5787) );
  DFFR_X1 \REGISTERS_reg[38][28]  ( .D(n7535), .CK(CLK), .RN(n12614), .QN(
        n5819) );
  DFFR_X1 \REGISTERS_reg[38][27]  ( .D(n7536), .CK(CLK), .RN(n12585), .QN(
        n5851) );
  DFFR_X1 \REGISTERS_reg[38][26]  ( .D(n7537), .CK(CLK), .RN(n12563), .QN(
        n5883) );
  DFFR_X1 \REGISTERS_reg[38][25]  ( .D(n7538), .CK(CLK), .RN(n12541), .QN(
        n5915) );
  DFFR_X1 \REGISTERS_reg[38][24]  ( .D(n7539), .CK(CLK), .RN(n12515), .QN(
        n5947) );
  DFFR_X1 \REGISTERS_reg[38][23]  ( .D(n7540), .CK(CLK), .RN(n12629), .QN(
        n6011) );
  DFFR_X1 \REGISTERS_reg[38][22]  ( .D(n7541), .CK(CLK), .RN(n12519), .QN(
        n9146) );
  DFFR_X1 \REGISTERS_reg[38][21]  ( .D(n7542), .CK(CLK), .RN(n12526), .QN(
        n9178) );
  DFFR_X1 \REGISTERS_reg[38][20]  ( .D(n7543), .CK(CLK), .RN(n12501), .QN(
        n9210) );
  DFFR_X1 \REGISTERS_reg[38][19]  ( .D(n7544), .CK(CLK), .RN(n12592), .QN(
        n9576) );
  DFFR_X1 \REGISTERS_reg[38][18]  ( .D(n7545), .CK(CLK), .RN(n12443), .QN(
        n9608) );
  DFFR_X1 \REGISTERS_reg[38][17]  ( .D(n7546), .CK(CLK), .RN(n12450), .QN(
        n9640) );
  DFFR_X1 \REGISTERS_reg[38][16]  ( .D(n7547), .CK(CLK), .RN(n12457), .QN(
        n10002) );
  DFFR_X1 \REGISTERS_reg[38][15]  ( .D(n7548), .CK(CLK), .RN(n12636), .QN(
        n10034) );
  DFFR_X1 \REGISTERS_reg[38][14]  ( .D(n7549), .CK(CLK), .RN(n12464), .QN(
        n10066) );
  DFFR_X1 \REGISTERS_reg[38][13]  ( .D(n7550), .CK(CLK), .RN(n12471), .QN(
        n10098) );
  DFFR_X1 \REGISTERS_reg[38][12]  ( .D(n7551), .CK(CLK), .RN(n12479), .QN(
        n10130) );
  DFFR_X1 \REGISTERS_reg[38][11]  ( .D(n7552), .CK(CLK), .RN(n12570), .QN(
        n10162) );
  DFFR_X1 \REGISTERS_reg[38][10]  ( .D(n7553), .CK(CLK), .RN(n12548), .QN(
        n10194) );
  DFFR_X1 \REGISTERS_reg[38][9]  ( .D(n7554), .CK(CLK), .RN(n12555), .QN(
        n10228) );
  DFFR_X1 \REGISTERS_reg[38][8]  ( .D(n7555), .CK(CLK), .RN(n12533), .QN(
        n10260) );
  DFFR_X1 \REGISTERS_reg[38][7]  ( .D(n7556), .CK(CLK), .RN(n12643), .QN(
        n10292) );
  DFFR_X1 \REGISTERS_reg[38][6]  ( .D(n7557), .CK(CLK), .RN(n12599), .QN(
        n10327) );
  DFFR_X1 \REGISTERS_reg[38][5]  ( .D(n7558), .CK(CLK), .RN(n12486), .QN(
        n10359) );
  DFFR_X1 \REGISTERS_reg[38][4]  ( .D(n7559), .CK(CLK), .RN(n12493), .QN(
        n10391) );
  DFFR_X1 \REGISTERS_reg[38][3]  ( .D(n7560), .CK(CLK), .RN(n12577), .QN(
        n10426) );
  DFFR_X1 \REGISTERS_reg[38][2]  ( .D(n7561), .CK(CLK), .RN(n12508), .QN(
        n10458) );
  DFFR_X1 \REGISTERS_reg[38][1]  ( .D(n7562), .CK(CLK), .RN(n12436), .QN(
        n10490) );
  DFFR_X1 \REGISTERS_reg[38][0]  ( .D(n7563), .CK(CLK), .RN(n12651), .QN(
        n10522) );
  DFFR_X1 \REGISTERS_reg[39][31]  ( .D(n7564), .CK(CLK), .RN(n12658), .QN(
        n13396) );
  DFFR_X1 \REGISTERS_reg[39][30]  ( .D(n7565), .CK(CLK), .RN(n12621), .QN(
        n13397) );
  DFFR_X1 \REGISTERS_reg[39][29]  ( .D(n7566), .CK(CLK), .RN(n12607), .QN(
        n13398) );
  DFFR_X1 \REGISTERS_reg[39][28]  ( .D(n7567), .CK(CLK), .RN(n12614), .QN(
        n13399) );
  DFFR_X1 \REGISTERS_reg[39][27]  ( .D(n7568), .CK(CLK), .RN(n12585), .QN(
        n13400) );
  DFFR_X1 \REGISTERS_reg[39][26]  ( .D(n7569), .CK(CLK), .RN(n12563), .QN(
        n13401) );
  DFFR_X1 \REGISTERS_reg[39][25]  ( .D(n7570), .CK(CLK), .RN(n12541), .QN(
        n13402) );
  DFFR_X1 \REGISTERS_reg[39][24]  ( .D(n7571), .CK(CLK), .RN(n12515), .QN(
        n13403) );
  DFFR_X1 \REGISTERS_reg[39][23]  ( .D(n7572), .CK(CLK), .RN(n12629), .QN(
        n13404) );
  DFFR_X1 \REGISTERS_reg[39][22]  ( .D(n7573), .CK(CLK), .RN(n12519), .QN(
        n13405) );
  DFFR_X1 \REGISTERS_reg[39][21]  ( .D(n7574), .CK(CLK), .RN(n12526), .QN(
        n13406) );
  DFFR_X1 \REGISTERS_reg[39][20]  ( .D(n7575), .CK(CLK), .RN(n12501), .QN(
        n13407) );
  DFFR_X1 \REGISTERS_reg[39][19]  ( .D(n7576), .CK(CLK), .RN(n12592), .QN(
        n13408) );
  DFFR_X1 \REGISTERS_reg[39][18]  ( .D(n7577), .CK(CLK), .RN(n12443), .QN(
        n13409) );
  DFFR_X1 \REGISTERS_reg[39][17]  ( .D(n7578), .CK(CLK), .RN(n12450), .QN(
        n13410) );
  DFFR_X1 \REGISTERS_reg[39][16]  ( .D(n7579), .CK(CLK), .RN(n12457), .QN(
        n13411) );
  DFFR_X1 \REGISTERS_reg[39][15]  ( .D(n7580), .CK(CLK), .RN(n12636), .QN(
        n13412) );
  DFFR_X1 \REGISTERS_reg[39][14]  ( .D(n7581), .CK(CLK), .RN(n12464), .QN(
        n13413) );
  DFFR_X1 \REGISTERS_reg[39][13]  ( .D(n7582), .CK(CLK), .RN(n12471), .QN(
        n13414) );
  DFFR_X1 \REGISTERS_reg[39][12]  ( .D(n7583), .CK(CLK), .RN(n12479), .QN(
        n13415) );
  DFFR_X1 \REGISTERS_reg[39][11]  ( .D(n7584), .CK(CLK), .RN(n12570), .QN(
        n13416) );
  DFFR_X1 \REGISTERS_reg[39][10]  ( .D(n7585), .CK(CLK), .RN(n12548), .QN(
        n13417) );
  DFFR_X1 \REGISTERS_reg[39][9]  ( .D(n7586), .CK(CLK), .RN(n12555), .QN(
        n13418) );
  DFFR_X1 \REGISTERS_reg[39][8]  ( .D(n7587), .CK(CLK), .RN(n12533), .QN(
        n13419) );
  DFFR_X1 \REGISTERS_reg[39][7]  ( .D(n7588), .CK(CLK), .RN(n12643), .QN(
        n13420) );
  DFFR_X1 \REGISTERS_reg[39][6]  ( .D(n7589), .CK(CLK), .RN(n12599), .QN(
        n13421) );
  DFFR_X1 \REGISTERS_reg[39][5]  ( .D(n7590), .CK(CLK), .RN(n12486), .QN(
        n13422) );
  DFFR_X1 \REGISTERS_reg[39][4]  ( .D(n7591), .CK(CLK), .RN(n12493), .QN(
        n13423) );
  DFFR_X1 \REGISTERS_reg[39][3]  ( .D(n7592), .CK(CLK), .RN(n12577), .QN(
        n13424) );
  DFFR_X1 \REGISTERS_reg[39][2]  ( .D(n7593), .CK(CLK), .RN(n12508), .QN(
        n13425) );
  DFFR_X1 \REGISTERS_reg[39][1]  ( .D(n7594), .CK(CLK), .RN(n12436), .QN(
        n13426) );
  DFFR_X1 \REGISTERS_reg[39][0]  ( .D(n7595), .CK(CLK), .RN(n12651), .QN(
        n13427) );
  DFFR_X1 \REGISTERS_reg[40][31]  ( .D(n7596), .CK(CLK), .RN(n12658), .QN(
        n5724) );
  DFFR_X1 \REGISTERS_reg[40][30]  ( .D(n7597), .CK(CLK), .RN(n12622), .QN(
        n5756) );
  DFFR_X1 \REGISTERS_reg[40][29]  ( .D(n7598), .CK(CLK), .RN(n12607), .QN(
        n5788) );
  DFFR_X1 \REGISTERS_reg[40][28]  ( .D(n7599), .CK(CLK), .RN(n12614), .QN(
        n5820) );
  DFFR_X1 \REGISTERS_reg[40][27]  ( .D(n7600), .CK(CLK), .RN(n12585), .QN(
        n5852) );
  DFFR_X1 \REGISTERS_reg[40][26]  ( .D(n7601), .CK(CLK), .RN(n12563), .QN(
        n5884) );
  DFFR_X1 \REGISTERS_reg[40][25]  ( .D(n7602), .CK(CLK), .RN(n12541), .QN(
        n5916) );
  DFFR_X1 \REGISTERS_reg[40][24]  ( .D(n7603), .CK(CLK), .RN(n12516), .QN(
        n5948) );
  DFFR_X1 \REGISTERS_reg[40][23]  ( .D(n7604), .CK(CLK), .RN(n12629), .QN(
        n6012) );
  DFFR_X1 \REGISTERS_reg[40][22]  ( .D(n7605), .CK(CLK), .RN(n12519), .QN(
        n9147) );
  DFFR_X1 \REGISTERS_reg[40][21]  ( .D(n7606), .CK(CLK), .RN(n12526), .QN(
        n9179) );
  DFFR_X1 \REGISTERS_reg[40][20]  ( .D(n7607), .CK(CLK), .RN(n12501), .QN(
        n9211) );
  DFFR_X1 \REGISTERS_reg[40][19]  ( .D(n7608), .CK(CLK), .RN(n12592), .QN(
        n9577) );
  DFFR_X1 \REGISTERS_reg[40][18]  ( .D(n7609), .CK(CLK), .RN(n12443), .QN(
        n9609) );
  DFFR_X1 \REGISTERS_reg[40][17]  ( .D(n7610), .CK(CLK), .RN(n12451), .QN(
        n9641) );
  DFFR_X1 \REGISTERS_reg[40][16]  ( .D(n7611), .CK(CLK), .RN(n12457), .QN(
        n10003) );
  DFFR_X1 \REGISTERS_reg[40][15]  ( .D(n7612), .CK(CLK), .RN(n12636), .QN(
        n10035) );
  DFFR_X1 \REGISTERS_reg[40][14]  ( .D(n7613), .CK(CLK), .RN(n12464), .QN(
        n10067) );
  DFFR_X1 \REGISTERS_reg[40][13]  ( .D(n7614), .CK(CLK), .RN(n12472), .QN(
        n10099) );
  DFFR_X1 \REGISTERS_reg[40][12]  ( .D(n7615), .CK(CLK), .RN(n12479), .QN(
        n10131) );
  DFFR_X1 \REGISTERS_reg[40][11]  ( .D(n7616), .CK(CLK), .RN(n12570), .QN(
        n10163) );
  DFFR_X1 \REGISTERS_reg[40][10]  ( .D(n7617), .CK(CLK), .RN(n12548), .QN(
        n10195) );
  DFFR_X1 \REGISTERS_reg[40][9]  ( .D(n7618), .CK(CLK), .RN(n12556), .QN(
        n10229) );
  DFFR_X1 \REGISTERS_reg[40][8]  ( .D(n7619), .CK(CLK), .RN(n12534), .QN(
        n10261) );
  DFFR_X1 \REGISTERS_reg[40][7]  ( .D(n7620), .CK(CLK), .RN(n12644), .QN(
        n10293) );
  DFFR_X1 \REGISTERS_reg[40][6]  ( .D(n7621), .CK(CLK), .RN(n12600), .QN(
        n10328) );
  DFFR_X1 \REGISTERS_reg[40][5]  ( .D(n7622), .CK(CLK), .RN(n12486), .QN(
        n10360) );
  DFFR_X1 \REGISTERS_reg[40][4]  ( .D(n7623), .CK(CLK), .RN(n12494), .QN(
        n10392) );
  DFFR_X1 \REGISTERS_reg[40][3]  ( .D(n7624), .CK(CLK), .RN(n12578), .QN(
        n10427) );
  DFFR_X1 \REGISTERS_reg[40][2]  ( .D(n7625), .CK(CLK), .RN(n12508), .QN(
        n10459) );
  DFFR_X1 \REGISTERS_reg[40][1]  ( .D(n7626), .CK(CLK), .RN(n12436), .QN(
        n10491) );
  DFFR_X1 \REGISTERS_reg[40][0]  ( .D(n7627), .CK(CLK), .RN(n12651), .QN(
        n10523) );
  DFFR_X1 \REGISTERS_reg[41][31]  ( .D(n7628), .CK(CLK), .RN(n12658), .QN(
        n13428) );
  DFFR_X1 \REGISTERS_reg[41][30]  ( .D(n7629), .CK(CLK), .RN(n12622), .QN(
        n13429) );
  DFFR_X1 \REGISTERS_reg[41][29]  ( .D(n7630), .CK(CLK), .RN(n12607), .QN(
        n13430) );
  DFFR_X1 \REGISTERS_reg[41][28]  ( .D(n7631), .CK(CLK), .RN(n12614), .QN(
        n13431) );
  DFFR_X1 \REGISTERS_reg[41][27]  ( .D(n7632), .CK(CLK), .RN(n12585), .QN(
        n13432) );
  DFFR_X1 \REGISTERS_reg[41][26]  ( .D(n7633), .CK(CLK), .RN(n12563), .QN(
        n13433) );
  DFFR_X1 \REGISTERS_reg[41][25]  ( .D(n7634), .CK(CLK), .RN(n12541), .QN(
        n13434) );
  DFFR_X1 \REGISTERS_reg[41][24]  ( .D(n7635), .CK(CLK), .RN(n12516), .QN(
        n13435) );
  DFFR_X1 \REGISTERS_reg[41][23]  ( .D(n7636), .CK(CLK), .RN(n12629), .QN(
        n13436) );
  DFFR_X1 \REGISTERS_reg[41][22]  ( .D(n7637), .CK(CLK), .RN(n12519), .QN(
        n13437) );
  DFFR_X1 \REGISTERS_reg[41][21]  ( .D(n7638), .CK(CLK), .RN(n12526), .QN(
        n13438) );
  DFFR_X1 \REGISTERS_reg[41][20]  ( .D(n7639), .CK(CLK), .RN(n12501), .QN(
        n13439) );
  DFFR_X1 \REGISTERS_reg[41][19]  ( .D(n7640), .CK(CLK), .RN(n12592), .QN(
        n13440) );
  DFFR_X1 \REGISTERS_reg[41][18]  ( .D(n7641), .CK(CLK), .RN(n12443), .QN(
        n13441) );
  DFFR_X1 \REGISTERS_reg[41][17]  ( .D(n7642), .CK(CLK), .RN(n12451), .QN(
        n13442) );
  DFFR_X1 \REGISTERS_reg[41][16]  ( .D(n7643), .CK(CLK), .RN(n12457), .QN(
        n13443) );
  DFFR_X1 \REGISTERS_reg[41][15]  ( .D(n7644), .CK(CLK), .RN(n12636), .QN(
        n13444) );
  DFFR_X1 \REGISTERS_reg[41][14]  ( .D(n7645), .CK(CLK), .RN(n12464), .QN(
        n13445) );
  DFFR_X1 \REGISTERS_reg[41][13]  ( .D(n7646), .CK(CLK), .RN(n12472), .QN(
        n13446) );
  DFFR_X1 \REGISTERS_reg[41][12]  ( .D(n7647), .CK(CLK), .RN(n12479), .QN(
        n13447) );
  DFFR_X1 \REGISTERS_reg[41][11]  ( .D(n7648), .CK(CLK), .RN(n12570), .QN(
        n13448) );
  DFFR_X1 \REGISTERS_reg[41][10]  ( .D(n7649), .CK(CLK), .RN(n12548), .QN(
        n13449) );
  DFFR_X1 \REGISTERS_reg[41][9]  ( .D(n7650), .CK(CLK), .RN(n12556), .QN(
        n13450) );
  DFFR_X1 \REGISTERS_reg[41][8]  ( .D(n7651), .CK(CLK), .RN(n12534), .QN(
        n13451) );
  DFFR_X1 \REGISTERS_reg[41][7]  ( .D(n7652), .CK(CLK), .RN(n12644), .QN(
        n13452) );
  DFFR_X1 \REGISTERS_reg[41][6]  ( .D(n7653), .CK(CLK), .RN(n12600), .QN(
        n13453) );
  DFFR_X1 \REGISTERS_reg[41][5]  ( .D(n7654), .CK(CLK), .RN(n12486), .QN(
        n13454) );
  DFFR_X1 \REGISTERS_reg[41][4]  ( .D(n7655), .CK(CLK), .RN(n12494), .QN(
        n13455) );
  DFFR_X1 \REGISTERS_reg[41][3]  ( .D(n7656), .CK(CLK), .RN(n12578), .QN(
        n13456) );
  DFFR_X1 \REGISTERS_reg[41][2]  ( .D(n7657), .CK(CLK), .RN(n12508), .QN(
        n13457) );
  DFFR_X1 \REGISTERS_reg[41][1]  ( .D(n7658), .CK(CLK), .RN(n12436), .QN(
        n13458) );
  DFFR_X1 \REGISTERS_reg[41][0]  ( .D(n7659), .CK(CLK), .RN(n12651), .QN(
        n13459) );
  DFFR_X1 \REGISTERS_reg[42][31]  ( .D(n7660), .CK(CLK), .RN(n12658), .QN(
        n5730) );
  DFFR_X1 \REGISTERS_reg[42][30]  ( .D(n7661), .CK(CLK), .RN(n12622), .QN(
        n5762) );
  DFFR_X1 \REGISTERS_reg[42][29]  ( .D(n7662), .CK(CLK), .RN(n12607), .QN(
        n5794) );
  DFFR_X1 \REGISTERS_reg[42][28]  ( .D(n7663), .CK(CLK), .RN(n12614), .QN(
        n5826) );
  DFFR_X1 \REGISTERS_reg[42][27]  ( .D(n7664), .CK(CLK), .RN(n12585), .QN(
        n5858) );
  DFFR_X1 \REGISTERS_reg[42][26]  ( .D(n7665), .CK(CLK), .RN(n12563), .QN(
        n5890) );
  DFFR_X1 \REGISTERS_reg[42][25]  ( .D(n7666), .CK(CLK), .RN(n12541), .QN(
        n5922) );
  DFFR_X1 \REGISTERS_reg[42][24]  ( .D(n7667), .CK(CLK), .RN(n12516), .QN(
        n5986) );
  DFFR_X1 \REGISTERS_reg[42][23]  ( .D(n7668), .CK(CLK), .RN(n12629), .QN(
        n6303) );
  DFFR_X1 \REGISTERS_reg[42][22]  ( .D(n7669), .CK(CLK), .RN(n12519), .QN(
        n9153) );
  DFFR_X1 \REGISTERS_reg[42][21]  ( .D(n7670), .CK(CLK), .RN(n12526), .QN(
        n9185) );
  DFFR_X1 \REGISTERS_reg[42][20]  ( .D(n7671), .CK(CLK), .RN(n12501), .QN(
        n9249) );
  DFFR_X1 \REGISTERS_reg[42][19]  ( .D(n7672), .CK(CLK), .RN(n12592), .QN(
        n9583) );
  DFFR_X1 \REGISTERS_reg[42][18]  ( .D(n7673), .CK(CLK), .RN(n12443), .QN(
        n9615) );
  DFFR_X1 \REGISTERS_reg[42][17]  ( .D(n7674), .CK(CLK), .RN(n12451), .QN(
        n9647) );
  DFFR_X1 \REGISTERS_reg[42][16]  ( .D(n7675), .CK(CLK), .RN(n12457), .QN(
        n10009) );
  DFFR_X1 \REGISTERS_reg[42][15]  ( .D(n7676), .CK(CLK), .RN(n12636), .QN(
        n10041) );
  DFFR_X1 \REGISTERS_reg[42][14]  ( .D(n7677), .CK(CLK), .RN(n12464), .QN(
        n10073) );
  DFFR_X1 \REGISTERS_reg[42][13]  ( .D(n7678), .CK(CLK), .RN(n12472), .QN(
        n10105) );
  DFFR_X1 \REGISTERS_reg[42][12]  ( .D(n7679), .CK(CLK), .RN(n12479), .QN(
        n10137) );
  DFFR_X1 \REGISTERS_reg[42][11]  ( .D(n7680), .CK(CLK), .RN(n12570), .QN(
        n10169) );
  DFFR_X1 \REGISTERS_reg[42][10]  ( .D(n7681), .CK(CLK), .RN(n12548), .QN(
        n10201) );
  DFFR_X1 \REGISTERS_reg[42][9]  ( .D(n7682), .CK(CLK), .RN(n12556), .QN(
        n10235) );
  DFFR_X1 \REGISTERS_reg[42][8]  ( .D(n7683), .CK(CLK), .RN(n12534), .QN(
        n10267) );
  DFFR_X1 \REGISTERS_reg[42][7]  ( .D(n7684), .CK(CLK), .RN(n12644), .QN(
        n10299) );
  DFFR_X1 \REGISTERS_reg[42][6]  ( .D(n7685), .CK(CLK), .RN(n12600), .QN(
        n10334) );
  DFFR_X1 \REGISTERS_reg[42][5]  ( .D(n7686), .CK(CLK), .RN(n12486), .QN(
        n10366) );
  DFFR_X1 \REGISTERS_reg[42][4]  ( .D(n7687), .CK(CLK), .RN(n12494), .QN(
        n10401) );
  DFFR_X1 \REGISTERS_reg[42][3]  ( .D(n7688), .CK(CLK), .RN(n12578), .QN(
        n10433) );
  DFFR_X1 \REGISTERS_reg[42][2]  ( .D(n7689), .CK(CLK), .RN(n12508), .QN(
        n10465) );
  DFFR_X1 \REGISTERS_reg[42][1]  ( .D(n7690), .CK(CLK), .RN(n12436), .QN(
        n10497) );
  DFFR_X1 \REGISTERS_reg[42][0]  ( .D(n7691), .CK(CLK), .RN(n12651), .QN(
        n10529) );
  DFFR_X1 \REGISTERS_reg[43][31]  ( .D(n7692), .CK(CLK), .RN(n12658), .QN(
        n13460) );
  DFFR_X1 \REGISTERS_reg[43][30]  ( .D(n7693), .CK(CLK), .RN(n12622), .QN(
        n13461) );
  DFFR_X1 \REGISTERS_reg[43][29]  ( .D(n7694), .CK(CLK), .RN(n12607), .QN(
        n13462) );
  DFFR_X1 \REGISTERS_reg[43][28]  ( .D(n7695), .CK(CLK), .RN(n12614), .QN(
        n13463) );
  DFFR_X1 \REGISTERS_reg[43][27]  ( .D(n7696), .CK(CLK), .RN(n12585), .QN(
        n13464) );
  DFFR_X1 \REGISTERS_reg[43][26]  ( .D(n7697), .CK(CLK), .RN(n12563), .QN(
        n13465) );
  DFFR_X1 \REGISTERS_reg[43][25]  ( .D(n7698), .CK(CLK), .RN(n12541), .QN(
        n13466) );
  DFFR_X1 \REGISTERS_reg[43][24]  ( .D(n7699), .CK(CLK), .RN(n12516), .QN(
        n13467) );
  DFFR_X1 \REGISTERS_reg[43][23]  ( .D(n7700), .CK(CLK), .RN(n12629), .QN(
        n13468) );
  DFFR_X1 \REGISTERS_reg[43][22]  ( .D(n7701), .CK(CLK), .RN(n12519), .QN(
        n13469) );
  DFFR_X1 \REGISTERS_reg[43][21]  ( .D(n7702), .CK(CLK), .RN(n12526), .QN(
        n13470) );
  DFFR_X1 \REGISTERS_reg[43][20]  ( .D(n7703), .CK(CLK), .RN(n12501), .QN(
        n13471) );
  DFFR_X1 \REGISTERS_reg[43][19]  ( .D(n7704), .CK(CLK), .RN(n12592), .QN(
        n13472) );
  DFFR_X1 \REGISTERS_reg[43][18]  ( .D(n7705), .CK(CLK), .RN(n12443), .QN(
        n13473) );
  DFFR_X1 \REGISTERS_reg[43][17]  ( .D(n7706), .CK(CLK), .RN(n12451), .QN(
        n13474) );
  DFFR_X1 \REGISTERS_reg[43][16]  ( .D(n7707), .CK(CLK), .RN(n12457), .QN(
        n13475) );
  DFFR_X1 \REGISTERS_reg[43][15]  ( .D(n7708), .CK(CLK), .RN(n12636), .QN(
        n13476) );
  DFFR_X1 \REGISTERS_reg[43][14]  ( .D(n7709), .CK(CLK), .RN(n12464), .QN(
        n13477) );
  DFFR_X1 \REGISTERS_reg[43][13]  ( .D(n7710), .CK(CLK), .RN(n12472), .QN(
        n13478) );
  DFFR_X1 \REGISTERS_reg[43][12]  ( .D(n7711), .CK(CLK), .RN(n12479), .QN(
        n13479) );
  DFFR_X1 \REGISTERS_reg[43][11]  ( .D(n7712), .CK(CLK), .RN(n12570), .QN(
        n13480) );
  DFFR_X1 \REGISTERS_reg[43][10]  ( .D(n7713), .CK(CLK), .RN(n12548), .QN(
        n13481) );
  DFFR_X1 \REGISTERS_reg[43][9]  ( .D(n7714), .CK(CLK), .RN(n12556), .QN(
        n13482) );
  DFFR_X1 \REGISTERS_reg[43][8]  ( .D(n7715), .CK(CLK), .RN(n12534), .QN(
        n13483) );
  DFFR_X1 \REGISTERS_reg[43][7]  ( .D(n7716), .CK(CLK), .RN(n12644), .QN(
        n13484) );
  DFFR_X1 \REGISTERS_reg[43][6]  ( .D(n7717), .CK(CLK), .RN(n12600), .QN(
        n13485) );
  DFFR_X1 \REGISTERS_reg[43][5]  ( .D(n7718), .CK(CLK), .RN(n12486), .QN(
        n13486) );
  DFFR_X1 \REGISTERS_reg[43][4]  ( .D(n7719), .CK(CLK), .RN(n12494), .QN(
        n13487) );
  DFFR_X1 \REGISTERS_reg[43][3]  ( .D(n7720), .CK(CLK), .RN(n12578), .QN(
        n13488) );
  DFFR_X1 \REGISTERS_reg[43][2]  ( .D(n7721), .CK(CLK), .RN(n12508), .QN(
        n13489) );
  DFFR_X1 \REGISTERS_reg[43][1]  ( .D(n7722), .CK(CLK), .RN(n12436), .QN(
        n13490) );
  DFFR_X1 \REGISTERS_reg[43][0]  ( .D(n7723), .CK(CLK), .RN(n12651), .QN(
        n13491) );
  DFFR_X1 \REGISTERS_reg[44][31]  ( .D(n7724), .CK(CLK), .RN(n12659), .Q(n9567), .QN(n13492) );
  DFFR_X1 \REGISTERS_reg[44][30]  ( .D(n7725), .CK(CLK), .RN(n12622), .Q(n9566), .QN(n13493) );
  DFFR_X1 \REGISTERS_reg[44][29]  ( .D(n7726), .CK(CLK), .RN(n12607), .Q(n9565), .QN(n13494) );
  DFFR_X1 \REGISTERS_reg[44][28]  ( .D(n7727), .CK(CLK), .RN(n12615), .Q(n9564), .QN(n13495) );
  DFFR_X1 \REGISTERS_reg[44][27]  ( .D(n7728), .CK(CLK), .RN(n12585), .Q(n9563), .QN(n13496) );
  DFFR_X1 \REGISTERS_reg[44][26]  ( .D(n7729), .CK(CLK), .RN(n12563), .Q(n9562), .QN(n13497) );
  DFFR_X1 \REGISTERS_reg[44][25]  ( .D(n7730), .CK(CLK), .RN(n12541), .Q(n9561), .QN(n13498) );
  DFFR_X1 \REGISTERS_reg[44][24]  ( .D(n7731), .CK(CLK), .RN(n12516), .Q(n9560), .QN(n13499) );
  DFFR_X1 \REGISTERS_reg[44][23]  ( .D(n7732), .CK(CLK), .RN(n12629), .Q(n9559), .QN(n13500) );
  DFFR_X1 \REGISTERS_reg[44][22]  ( .D(n7733), .CK(CLK), .RN(n12519), .Q(n9558), .QN(n13501) );
  DFFR_X1 \REGISTERS_reg[44][21]  ( .D(n7734), .CK(CLK), .RN(n12527), .Q(n9557), .QN(n13502) );
  DFFR_X1 \REGISTERS_reg[44][20]  ( .D(n7735), .CK(CLK), .RN(n12501), .Q(n9556), .QN(n13503) );
  DFFR_X1 \REGISTERS_reg[44][19]  ( .D(n7736), .CK(CLK), .RN(n12593), .Q(n9555), .QN(n13504) );
  DFFR_X1 \REGISTERS_reg[44][18]  ( .D(n7737), .CK(CLK), .RN(n12444), .Q(n9554), .QN(n13505) );
  DFFR_X1 \REGISTERS_reg[44][17]  ( .D(n7738), .CK(CLK), .RN(n12451), .Q(n9553), .QN(n13506) );
  DFFR_X1 \REGISTERS_reg[44][16]  ( .D(n7739), .CK(CLK), .RN(n12457), .Q(n9552), .QN(n13507) );
  DFFR_X1 \REGISTERS_reg[44][15]  ( .D(n7740), .CK(CLK), .RN(n12637), .Q(n9551), .QN(n13508) );
  DFFR_X1 \REGISTERS_reg[44][14]  ( .D(n7741), .CK(CLK), .RN(n12465), .Q(n9550), .QN(n13509) );
  DFFR_X1 \REGISTERS_reg[44][13]  ( .D(n7742), .CK(CLK), .RN(n12472), .Q(n9549), .QN(n13510) );
  DFFR_X1 \REGISTERS_reg[44][12]  ( .D(n7743), .CK(CLK), .RN(n12479), .Q(n9548), .QN(n13511) );
  DFFR_X1 \REGISTERS_reg[44][11]  ( .D(n7744), .CK(CLK), .RN(n12571), .Q(n9547), .QN(n13512) );
  DFFR_X1 \REGISTERS_reg[44][10]  ( .D(n7745), .CK(CLK), .RN(n12549), .Q(n9546), .QN(n13513) );
  DFFR_X1 \REGISTERS_reg[44][9]  ( .D(n7746), .CK(CLK), .RN(n12556), .Q(n9545), 
        .QN(n13514) );
  DFFR_X1 \REGISTERS_reg[44][8]  ( .D(n7747), .CK(CLK), .RN(n12534), .Q(n9544), 
        .QN(n13515) );
  DFFR_X1 \REGISTERS_reg[44][7]  ( .D(n7748), .CK(CLK), .RN(n12644), .Q(n9543), 
        .QN(n13516) );
  DFFR_X1 \REGISTERS_reg[44][6]  ( .D(n7749), .CK(CLK), .RN(n12600), .Q(n9542), 
        .QN(n13517) );
  DFFR_X1 \REGISTERS_reg[44][5]  ( .D(n7750), .CK(CLK), .RN(n12487), .Q(n9541), 
        .QN(n13518) );
  DFFR_X1 \REGISTERS_reg[44][4]  ( .D(n7751), .CK(CLK), .RN(n12494), .Q(n9540), 
        .QN(n13519) );
  DFFR_X1 \REGISTERS_reg[44][3]  ( .D(n7752), .CK(CLK), .RN(n12578), .Q(n9539), 
        .QN(n13520) );
  DFFR_X1 \REGISTERS_reg[44][2]  ( .D(n7753), .CK(CLK), .RN(n12509), .Q(n9538), 
        .QN(n13521) );
  DFFR_X1 \REGISTERS_reg[44][1]  ( .D(n7754), .CK(CLK), .RN(n12436), .Q(n9537), 
        .QN(n13522) );
  DFFR_X1 \REGISTERS_reg[44][0]  ( .D(n7755), .CK(CLK), .RN(n12651), .Q(n9536), 
        .QN(n13523) );
  DFFR_X1 \REGISTERS_reg[45][31]  ( .D(n7756), .CK(CLK), .RN(n12659), .Q(n9535), .QN(n13524) );
  DFFR_X1 \REGISTERS_reg[45][30]  ( .D(n7757), .CK(CLK), .RN(n12622), .Q(n9534), .QN(n13525) );
  DFFR_X1 \REGISTERS_reg[45][29]  ( .D(n7758), .CK(CLK), .RN(n12607), .Q(n9533), .QN(n13526) );
  DFFR_X1 \REGISTERS_reg[45][28]  ( .D(n7759), .CK(CLK), .RN(n12615), .Q(n9532), .QN(n13527) );
  DFFR_X1 \REGISTERS_reg[45][27]  ( .D(n7760), .CK(CLK), .RN(n12585), .Q(n9531), .QN(n13528) );
  DFFR_X1 \REGISTERS_reg[45][26]  ( .D(n7761), .CK(CLK), .RN(n12563), .Q(n9530), .QN(n13529) );
  DFFR_X1 \REGISTERS_reg[45][25]  ( .D(n7762), .CK(CLK), .RN(n12541), .Q(n9529), .QN(n13530) );
  DFFR_X1 \REGISTERS_reg[45][24]  ( .D(n7763), .CK(CLK), .RN(n12516), .Q(n9528), .QN(n13531) );
  DFFR_X1 \REGISTERS_reg[45][23]  ( .D(n7764), .CK(CLK), .RN(n12629), .Q(n9527), .QN(n13532) );
  DFFR_X1 \REGISTERS_reg[45][22]  ( .D(n7765), .CK(CLK), .RN(n12519), .Q(n9526), .QN(n13533) );
  DFFR_X1 \REGISTERS_reg[45][21]  ( .D(n7766), .CK(CLK), .RN(n12527), .Q(n9525), .QN(n13534) );
  DFFR_X1 \REGISTERS_reg[45][20]  ( .D(n7767), .CK(CLK), .RN(n12501), .Q(n9524), .QN(n13535) );
  DFFR_X1 \REGISTERS_reg[45][19]  ( .D(n7768), .CK(CLK), .RN(n12593), .Q(n9523), .QN(n13536) );
  DFFR_X1 \REGISTERS_reg[45][18]  ( .D(n7769), .CK(CLK), .RN(n12444), .Q(n9522), .QN(n13537) );
  DFFR_X1 \REGISTERS_reg[45][17]  ( .D(n7770), .CK(CLK), .RN(n12451), .Q(n9521), .QN(n13538) );
  DFFR_X1 \REGISTERS_reg[45][16]  ( .D(n7771), .CK(CLK), .RN(n12457), .Q(n9520), .QN(n13539) );
  DFFR_X1 \REGISTERS_reg[45][15]  ( .D(n7772), .CK(CLK), .RN(n12637), .Q(n9519), .QN(n13540) );
  DFFR_X1 \REGISTERS_reg[45][14]  ( .D(n7773), .CK(CLK), .RN(n12465), .Q(n9518), .QN(n13541) );
  DFFR_X1 \REGISTERS_reg[45][13]  ( .D(n7774), .CK(CLK), .RN(n12472), .Q(n9517), .QN(n13542) );
  DFFR_X1 \REGISTERS_reg[45][12]  ( .D(n7775), .CK(CLK), .RN(n12479), .Q(n9516), .QN(n13543) );
  DFFR_X1 \REGISTERS_reg[45][11]  ( .D(n7776), .CK(CLK), .RN(n12571), .Q(n9515), .QN(n13544) );
  DFFR_X1 \REGISTERS_reg[45][10]  ( .D(n7777), .CK(CLK), .RN(n12549), .Q(n9514), .QN(n13545) );
  DFFR_X1 \REGISTERS_reg[45][9]  ( .D(n7778), .CK(CLK), .RN(n12556), .Q(n9513), 
        .QN(n13546) );
  DFFR_X1 \REGISTERS_reg[45][8]  ( .D(n7779), .CK(CLK), .RN(n12534), .Q(n9512), 
        .QN(n13547) );
  DFFR_X1 \REGISTERS_reg[45][7]  ( .D(n7780), .CK(CLK), .RN(n12644), .Q(n9511), 
        .QN(n13548) );
  DFFR_X1 \REGISTERS_reg[45][6]  ( .D(n7781), .CK(CLK), .RN(n12600), .Q(n9510), 
        .QN(n13549) );
  DFFR_X1 \REGISTERS_reg[45][5]  ( .D(n7782), .CK(CLK), .RN(n12487), .Q(n9509), 
        .QN(n13550) );
  DFFR_X1 \REGISTERS_reg[45][4]  ( .D(n7783), .CK(CLK), .RN(n12494), .Q(n9508), 
        .QN(n13551) );
  DFFR_X1 \REGISTERS_reg[45][3]  ( .D(n7784), .CK(CLK), .RN(n12578), .Q(n9507), 
        .QN(n13552) );
  DFFR_X1 \REGISTERS_reg[45][2]  ( .D(n7785), .CK(CLK), .RN(n12509), .Q(n9506), 
        .QN(n13553) );
  DFFR_X1 \REGISTERS_reg[45][1]  ( .D(n7786), .CK(CLK), .RN(n12436), .Q(n9505), 
        .QN(n13554) );
  DFFR_X1 \REGISTERS_reg[45][0]  ( .D(n7787), .CK(CLK), .RN(n12651), .Q(n9504), 
        .QN(n13555) );
  DFFR_X1 \REGISTERS_reg[46][31]  ( .D(n7788), .CK(CLK), .RN(n12659), .QN(
        n13556) );
  DFFR_X1 \REGISTERS_reg[46][30]  ( .D(n7789), .CK(CLK), .RN(n12622), .QN(
        n13557) );
  DFFR_X1 \REGISTERS_reg[46][29]  ( .D(n7790), .CK(CLK), .RN(n12607), .QN(
        n13558) );
  DFFR_X1 \REGISTERS_reg[46][28]  ( .D(n7791), .CK(CLK), .RN(n12615), .QN(
        n13559) );
  DFFR_X1 \REGISTERS_reg[46][27]  ( .D(n7792), .CK(CLK), .RN(n12585), .QN(
        n13560) );
  DFFR_X1 \REGISTERS_reg[46][26]  ( .D(n7793), .CK(CLK), .RN(n12563), .QN(
        n13561) );
  DFFR_X1 \REGISTERS_reg[46][25]  ( .D(n7794), .CK(CLK), .RN(n12541), .QN(
        n13562) );
  DFFR_X1 \REGISTERS_reg[46][24]  ( .D(n7795), .CK(CLK), .RN(n12516), .QN(
        n13563) );
  DFFR_X1 \REGISTERS_reg[46][23]  ( .D(n7796), .CK(CLK), .RN(n12629), .QN(
        n13564) );
  DFFR_X1 \REGISTERS_reg[46][22]  ( .D(n7797), .CK(CLK), .RN(n12519), .QN(
        n13565) );
  DFFR_X1 \REGISTERS_reg[46][21]  ( .D(n7798), .CK(CLK), .RN(n12527), .QN(
        n13566) );
  DFFR_X1 \REGISTERS_reg[46][20]  ( .D(n7799), .CK(CLK), .RN(n12501), .QN(
        n13567) );
  DFFR_X1 \REGISTERS_reg[46][19]  ( .D(n7800), .CK(CLK), .RN(n12593), .QN(
        n13568) );
  DFFR_X1 \REGISTERS_reg[46][18]  ( .D(n7801), .CK(CLK), .RN(n12444), .QN(
        n13569) );
  DFFR_X1 \REGISTERS_reg[46][17]  ( .D(n7802), .CK(CLK), .RN(n12451), .QN(
        n13570) );
  DFFR_X1 \REGISTERS_reg[46][16]  ( .D(n7803), .CK(CLK), .RN(n12457), .QN(
        n13571) );
  DFFR_X1 \REGISTERS_reg[46][15]  ( .D(n7804), .CK(CLK), .RN(n12637), .QN(
        n13572) );
  DFFR_X1 \REGISTERS_reg[46][14]  ( .D(n7805), .CK(CLK), .RN(n12465), .QN(
        n13573) );
  DFFR_X1 \REGISTERS_reg[46][13]  ( .D(n7806), .CK(CLK), .RN(n12472), .QN(
        n13574) );
  DFFR_X1 \REGISTERS_reg[46][12]  ( .D(n7807), .CK(CLK), .RN(n12479), .QN(
        n13575) );
  DFFR_X1 \REGISTERS_reg[46][11]  ( .D(n7808), .CK(CLK), .RN(n12571), .QN(
        n13576) );
  DFFR_X1 \REGISTERS_reg[46][10]  ( .D(n7809), .CK(CLK), .RN(n12549), .QN(
        n13577) );
  DFFR_X1 \REGISTERS_reg[46][9]  ( .D(n7810), .CK(CLK), .RN(n12556), .QN(
        n13578) );
  DFFR_X1 \REGISTERS_reg[46][8]  ( .D(n7811), .CK(CLK), .RN(n12534), .QN(
        n13579) );
  DFFR_X1 \REGISTERS_reg[46][7]  ( .D(n7812), .CK(CLK), .RN(n12644), .QN(
        n13580) );
  DFFR_X1 \REGISTERS_reg[46][6]  ( .D(n7813), .CK(CLK), .RN(n12600), .QN(
        n13581) );
  DFFR_X1 \REGISTERS_reg[46][5]  ( .D(n7814), .CK(CLK), .RN(n12487), .QN(
        n13582) );
  DFFR_X1 \REGISTERS_reg[46][4]  ( .D(n7815), .CK(CLK), .RN(n12494), .QN(
        n13583) );
  DFFR_X1 \REGISTERS_reg[46][3]  ( .D(n7816), .CK(CLK), .RN(n12578), .QN(
        n13584) );
  DFFR_X1 \REGISTERS_reg[46][2]  ( .D(n7817), .CK(CLK), .RN(n12509), .QN(
        n13585) );
  DFFR_X1 \REGISTERS_reg[46][1]  ( .D(n7818), .CK(CLK), .RN(n12436), .QN(
        n13586) );
  DFFR_X1 \REGISTERS_reg[46][0]  ( .D(n7819), .CK(CLK), .RN(n12651), .QN(
        n13587) );
  DFFR_X1 \REGISTERS_reg[47][31]  ( .D(n7820), .CK(CLK), .RN(n12659), .QN(
        n13588) );
  DFFR_X1 \REGISTERS_reg[47][30]  ( .D(n7821), .CK(CLK), .RN(n12622), .QN(
        n13589) );
  DFFR_X1 \REGISTERS_reg[47][29]  ( .D(n7822), .CK(CLK), .RN(n12607), .QN(
        n13590) );
  DFFR_X1 \REGISTERS_reg[47][28]  ( .D(n7823), .CK(CLK), .RN(n12615), .QN(
        n13591) );
  DFFR_X1 \REGISTERS_reg[47][27]  ( .D(n7824), .CK(CLK), .RN(n12585), .QN(
        n13592) );
  DFFR_X1 \REGISTERS_reg[47][26]  ( .D(n7825), .CK(CLK), .RN(n12563), .QN(
        n13593) );
  DFFR_X1 \REGISTERS_reg[47][25]  ( .D(n7826), .CK(CLK), .RN(n12541), .QN(
        n13594) );
  DFFR_X1 \REGISTERS_reg[47][24]  ( .D(n7827), .CK(CLK), .RN(n12516), .QN(
        n13595) );
  DFFR_X1 \REGISTERS_reg[47][23]  ( .D(n7828), .CK(CLK), .RN(n12629), .QN(
        n13596) );
  DFFR_X1 \REGISTERS_reg[47][22]  ( .D(n7829), .CK(CLK), .RN(n12519), .QN(
        n13597) );
  DFFR_X1 \REGISTERS_reg[47][21]  ( .D(n7830), .CK(CLK), .RN(n12527), .QN(
        n13598) );
  DFFR_X1 \REGISTERS_reg[47][20]  ( .D(n7831), .CK(CLK), .RN(n12501), .QN(
        n13599) );
  DFFR_X1 \REGISTERS_reg[47][19]  ( .D(n7832), .CK(CLK), .RN(n12593), .QN(
        n13600) );
  DFFR_X1 \REGISTERS_reg[47][18]  ( .D(n7833), .CK(CLK), .RN(n12444), .QN(
        n13601) );
  DFFR_X1 \REGISTERS_reg[47][17]  ( .D(n7834), .CK(CLK), .RN(n12451), .QN(
        n13602) );
  DFFR_X1 \REGISTERS_reg[47][16]  ( .D(n7835), .CK(CLK), .RN(n12457), .QN(
        n13603) );
  DFFR_X1 \REGISTERS_reg[47][15]  ( .D(n7836), .CK(CLK), .RN(n12637), .QN(
        n13604) );
  DFFR_X1 \REGISTERS_reg[47][14]  ( .D(n7837), .CK(CLK), .RN(n12465), .QN(
        n13605) );
  DFFR_X1 \REGISTERS_reg[47][13]  ( .D(n7838), .CK(CLK), .RN(n12472), .QN(
        n13606) );
  DFFR_X1 \REGISTERS_reg[47][12]  ( .D(n7839), .CK(CLK), .RN(n12479), .QN(
        n13607) );
  DFFR_X1 \REGISTERS_reg[47][11]  ( .D(n7840), .CK(CLK), .RN(n12571), .QN(
        n13608) );
  DFFR_X1 \REGISTERS_reg[47][10]  ( .D(n7841), .CK(CLK), .RN(n12549), .QN(
        n13609) );
  DFFR_X1 \REGISTERS_reg[47][9]  ( .D(n7842), .CK(CLK), .RN(n12556), .QN(
        n13610) );
  DFFR_X1 \REGISTERS_reg[47][8]  ( .D(n7843), .CK(CLK), .RN(n12534), .QN(
        n13611) );
  DFFR_X1 \REGISTERS_reg[47][7]  ( .D(n7844), .CK(CLK), .RN(n12644), .QN(
        n13612) );
  DFFR_X1 \REGISTERS_reg[47][6]  ( .D(n7845), .CK(CLK), .RN(n12600), .QN(
        n13613) );
  DFFR_X1 \REGISTERS_reg[47][5]  ( .D(n7846), .CK(CLK), .RN(n12487), .QN(
        n13614) );
  DFFR_X1 \REGISTERS_reg[47][4]  ( .D(n7847), .CK(CLK), .RN(n12494), .QN(
        n13615) );
  DFFR_X1 \REGISTERS_reg[47][3]  ( .D(n7848), .CK(CLK), .RN(n12578), .QN(
        n13616) );
  DFFR_X1 \REGISTERS_reg[47][2]  ( .D(n7849), .CK(CLK), .RN(n12509), .QN(
        n13617) );
  DFFR_X1 \REGISTERS_reg[47][1]  ( .D(n7850), .CK(CLK), .RN(n12436), .QN(
        n13618) );
  DFFR_X1 \REGISTERS_reg[47][0]  ( .D(n7851), .CK(CLK), .RN(n12651), .QN(
        n13619) );
  DFFR_X1 \REGISTERS_reg[48][31]  ( .D(n7852), .CK(CLK), .RN(n12659), .QN(
        n13620) );
  DFFR_X1 \REGISTERS_reg[48][30]  ( .D(n7853), .CK(CLK), .RN(n12622), .QN(
        n13621) );
  DFFR_X1 \REGISTERS_reg[48][29]  ( .D(n7854), .CK(CLK), .RN(n12608), .QN(
        n13622) );
  DFFR_X1 \REGISTERS_reg[48][28]  ( .D(n7855), .CK(CLK), .RN(n12615), .QN(
        n13623) );
  DFFR_X1 \REGISTERS_reg[48][27]  ( .D(n7856), .CK(CLK), .RN(n12586), .QN(
        n13624) );
  DFFR_X1 \REGISTERS_reg[48][26]  ( .D(n7857), .CK(CLK), .RN(n12564), .QN(
        n13625) );
  DFFR_X1 \REGISTERS_reg[48][25]  ( .D(n7858), .CK(CLK), .RN(n12542), .QN(
        n13626) );
  DFFR_X1 \REGISTERS_reg[48][24]  ( .D(n7859), .CK(CLK), .RN(n12516), .QN(
        n13627) );
  DFFR_X1 \REGISTERS_reg[48][23]  ( .D(n7860), .CK(CLK), .RN(n12630), .QN(
        n13628) );
  DFFR_X1 \REGISTERS_reg[48][22]  ( .D(n7861), .CK(CLK), .RN(n12520), .QN(
        n13629) );
  DFFR_X1 \REGISTERS_reg[48][21]  ( .D(n7862), .CK(CLK), .RN(n12527), .QN(
        n13630) );
  DFFR_X1 \REGISTERS_reg[48][20]  ( .D(n7863), .CK(CLK), .RN(n12502), .QN(
        n13631) );
  DFFR_X1 \REGISTERS_reg[48][19]  ( .D(n7864), .CK(CLK), .RN(n12593), .QN(
        n13632) );
  DFFR_X1 \REGISTERS_reg[48][18]  ( .D(n7865), .CK(CLK), .RN(n12444), .QN(
        n13633) );
  DFFR_X1 \REGISTERS_reg[48][17]  ( .D(n7866), .CK(CLK), .RN(n12451), .QN(
        n13634) );
  DFFR_X1 \REGISTERS_reg[48][16]  ( .D(n7867), .CK(CLK), .RN(n12458), .QN(
        n13635) );
  DFFR_X1 \REGISTERS_reg[48][15]  ( .D(n7868), .CK(CLK), .RN(n12637), .QN(
        n13636) );
  DFFR_X1 \REGISTERS_reg[48][14]  ( .D(n7869), .CK(CLK), .RN(n12465), .QN(
        n13637) );
  DFFR_X1 \REGISTERS_reg[48][13]  ( .D(n7870), .CK(CLK), .RN(n12472), .QN(
        n13638) );
  DFFR_X1 \REGISTERS_reg[48][12]  ( .D(n7871), .CK(CLK), .RN(n12480), .QN(
        n13639) );
  DFFR_X1 \REGISTERS_reg[48][11]  ( .D(n7872), .CK(CLK), .RN(n12571), .QN(
        n13640) );
  DFFR_X1 \REGISTERS_reg[48][10]  ( .D(n7873), .CK(CLK), .RN(n12549), .QN(
        n13641) );
  DFFR_X1 \REGISTERS_reg[48][9]  ( .D(n7874), .CK(CLK), .RN(n12556), .QN(
        n13642) );
  DFFR_X1 \REGISTERS_reg[48][8]  ( .D(n7875), .CK(CLK), .RN(n12534), .QN(
        n13643) );
  DFFR_X1 \REGISTERS_reg[48][7]  ( .D(n7876), .CK(CLK), .RN(n12644), .QN(
        n13644) );
  DFFR_X1 \REGISTERS_reg[48][6]  ( .D(n7877), .CK(CLK), .RN(n12600), .QN(
        n13645) );
  DFFR_X1 \REGISTERS_reg[48][5]  ( .D(n7878), .CK(CLK), .RN(n12487), .QN(
        n13646) );
  DFFR_X1 \REGISTERS_reg[48][4]  ( .D(n7879), .CK(CLK), .RN(n12494), .QN(
        n13647) );
  DFFR_X1 \REGISTERS_reg[48][3]  ( .D(n7880), .CK(CLK), .RN(n12578), .QN(
        n13648) );
  DFFR_X1 \REGISTERS_reg[48][2]  ( .D(n7881), .CK(CLK), .RN(n12509), .QN(
        n13649) );
  DFFR_X1 \REGISTERS_reg[48][1]  ( .D(n7882), .CK(CLK), .RN(n12437), .QN(
        n13650) );
  DFFR_X1 \REGISTERS_reg[48][0]  ( .D(n7883), .CK(CLK), .RN(n12652), .QN(
        n13651) );
  DFFR_X1 \REGISTERS_reg[49][31]  ( .D(n7884), .CK(CLK), .RN(n12659), .Q(n9407), .QN(n13652) );
  DFFR_X1 \REGISTERS_reg[49][30]  ( .D(n7885), .CK(CLK), .RN(n12622), .Q(n9406), .QN(n13653) );
  DFFR_X1 \REGISTERS_reg[49][29]  ( .D(n7886), .CK(CLK), .RN(n12608), .Q(n9405), .QN(n13654) );
  DFFR_X1 \REGISTERS_reg[49][28]  ( .D(n7887), .CK(CLK), .RN(n12615), .Q(n9404), .QN(n13655) );
  DFFR_X1 \REGISTERS_reg[49][27]  ( .D(n7888), .CK(CLK), .RN(n12586), .Q(n9403), .QN(n13656) );
  DFFR_X1 \REGISTERS_reg[49][26]  ( .D(n7889), .CK(CLK), .RN(n12564), .Q(n9402), .QN(n13657) );
  DFFR_X1 \REGISTERS_reg[49][25]  ( .D(n7890), .CK(CLK), .RN(n12542), .Q(n9401), .QN(n13658) );
  DFFR_X1 \REGISTERS_reg[49][24]  ( .D(n7891), .CK(CLK), .RN(n12516), .Q(n9400), .QN(n13659) );
  DFFR_X1 \REGISTERS_reg[49][23]  ( .D(n7892), .CK(CLK), .RN(n12630), .Q(n9399), .QN(n13660) );
  DFFR_X1 \REGISTERS_reg[49][22]  ( .D(n7893), .CK(CLK), .RN(n12520), .Q(n9398), .QN(n13661) );
  DFFR_X1 \REGISTERS_reg[49][21]  ( .D(n7894), .CK(CLK), .RN(n12527), .Q(n9397), .QN(n13662) );
  DFFR_X1 \REGISTERS_reg[49][20]  ( .D(n7895), .CK(CLK), .RN(n12502), .Q(n9396), .QN(n13663) );
  DFFR_X1 \REGISTERS_reg[49][19]  ( .D(n7896), .CK(CLK), .RN(n12593), .Q(n9395), .QN(n13664) );
  DFFR_X1 \REGISTERS_reg[49][18]  ( .D(n7897), .CK(CLK), .RN(n12444), .Q(n9394), .QN(n13665) );
  DFFR_X1 \REGISTERS_reg[49][17]  ( .D(n7898), .CK(CLK), .RN(n12451), .Q(n9393), .QN(n13666) );
  DFFR_X1 \REGISTERS_reg[49][16]  ( .D(n7899), .CK(CLK), .RN(n12458), .Q(n9392), .QN(n13667) );
  DFFR_X1 \REGISTERS_reg[49][15]  ( .D(n7900), .CK(CLK), .RN(n12637), .Q(n9391), .QN(n13668) );
  DFFR_X1 \REGISTERS_reg[49][14]  ( .D(n7901), .CK(CLK), .RN(n12465), .Q(n9390), .QN(n13669) );
  DFFR_X1 \REGISTERS_reg[49][13]  ( .D(n7902), .CK(CLK), .RN(n12472), .Q(n9389), .QN(n13670) );
  DFFR_X1 \REGISTERS_reg[49][12]  ( .D(n7903), .CK(CLK), .RN(n12480), .Q(n9388), .QN(n13671) );
  DFFR_X1 \REGISTERS_reg[49][11]  ( .D(n7904), .CK(CLK), .RN(n12571), .Q(n9387), .QN(n13672) );
  DFFR_X1 \REGISTERS_reg[49][10]  ( .D(n7905), .CK(CLK), .RN(n12549), .Q(n9386), .QN(n13673) );
  DFFR_X1 \REGISTERS_reg[49][9]  ( .D(n7906), .CK(CLK), .RN(n12556), .Q(n9385), 
        .QN(n13674) );
  DFFR_X1 \REGISTERS_reg[49][8]  ( .D(n7907), .CK(CLK), .RN(n12534), .Q(n9384), 
        .QN(n13675) );
  DFFR_X1 \REGISTERS_reg[49][7]  ( .D(n7908), .CK(CLK), .RN(n12644), .Q(n9383), 
        .QN(n13676) );
  DFFR_X1 \REGISTERS_reg[49][6]  ( .D(n7909), .CK(CLK), .RN(n12600), .Q(n9382), 
        .QN(n13677) );
  DFFR_X1 \REGISTERS_reg[49][5]  ( .D(n7910), .CK(CLK), .RN(n12487), .Q(n9381), 
        .QN(n13678) );
  DFFR_X1 \REGISTERS_reg[49][4]  ( .D(n7911), .CK(CLK), .RN(n12494), .Q(n9380), 
        .QN(n13679) );
  DFFR_X1 \REGISTERS_reg[49][3]  ( .D(n7912), .CK(CLK), .RN(n12578), .Q(n9379), 
        .QN(n13680) );
  DFFR_X1 \REGISTERS_reg[49][2]  ( .D(n7913), .CK(CLK), .RN(n12509), .Q(n9378), 
        .QN(n13681) );
  DFFR_X1 \REGISTERS_reg[49][1]  ( .D(n7914), .CK(CLK), .RN(n12437), .Q(n9377), 
        .QN(n13682) );
  DFFR_X1 \REGISTERS_reg[49][0]  ( .D(n7915), .CK(CLK), .RN(n12652), .Q(n9376), 
        .QN(n13683) );
  DFFR_X1 \REGISTERS_reg[50][31]  ( .D(n7916), .CK(CLK), .RN(n12659), .Q(n9375), .QN(n13684) );
  DFFR_X1 \REGISTERS_reg[50][30]  ( .D(n7917), .CK(CLK), .RN(n12622), .Q(n9374), .QN(n13685) );
  DFFR_X1 \REGISTERS_reg[50][29]  ( .D(n7918), .CK(CLK), .RN(n12608), .Q(n9373), .QN(n13686) );
  DFFR_X1 \REGISTERS_reg[50][28]  ( .D(n7919), .CK(CLK), .RN(n12615), .Q(n9372), .QN(n13687) );
  DFFR_X1 \REGISTERS_reg[50][27]  ( .D(n7920), .CK(CLK), .RN(n12586), .Q(n9371), .QN(n13688) );
  DFFR_X1 \REGISTERS_reg[50][26]  ( .D(n7921), .CK(CLK), .RN(n12564), .Q(n9370), .QN(n13689) );
  DFFR_X1 \REGISTERS_reg[50][25]  ( .D(n7922), .CK(CLK), .RN(n12542), .Q(n9369), .QN(n13690) );
  DFFR_X1 \REGISTERS_reg[50][24]  ( .D(n7923), .CK(CLK), .RN(n12516), .Q(n9368), .QN(n13691) );
  DFFR_X1 \REGISTERS_reg[50][23]  ( .D(n7924), .CK(CLK), .RN(n12630), .Q(n9367), .QN(n13692) );
  DFFR_X1 \REGISTERS_reg[50][22]  ( .D(n7925), .CK(CLK), .RN(n12520), .Q(n9366), .QN(n13693) );
  DFFR_X1 \REGISTERS_reg[50][21]  ( .D(n7926), .CK(CLK), .RN(n12527), .Q(n9365), .QN(n13694) );
  DFFR_X1 \REGISTERS_reg[50][20]  ( .D(n7927), .CK(CLK), .RN(n12502), .Q(n9364), .QN(n13695) );
  DFFR_X1 \REGISTERS_reg[50][19]  ( .D(n7928), .CK(CLK), .RN(n12593), .Q(n9363), .QN(n13696) );
  DFFR_X1 \REGISTERS_reg[50][18]  ( .D(n7929), .CK(CLK), .RN(n12444), .Q(n9362), .QN(n13697) );
  DFFR_X1 \REGISTERS_reg[50][17]  ( .D(n7930), .CK(CLK), .RN(n12451), .Q(n9361), .QN(n13698) );
  DFFR_X1 \REGISTERS_reg[50][16]  ( .D(n7931), .CK(CLK), .RN(n12458), .Q(n9360), .QN(n13699) );
  DFFR_X1 \REGISTERS_reg[50][15]  ( .D(n7932), .CK(CLK), .RN(n12637), .Q(n9359), .QN(n13700) );
  DFFR_X1 \REGISTERS_reg[50][14]  ( .D(n7933), .CK(CLK), .RN(n12465), .Q(n9358), .QN(n13701) );
  DFFR_X1 \REGISTERS_reg[50][13]  ( .D(n7934), .CK(CLK), .RN(n12472), .Q(n9357), .QN(n13702) );
  DFFR_X1 \REGISTERS_reg[50][12]  ( .D(n7935), .CK(CLK), .RN(n12480), .Q(n9356), .QN(n13703) );
  DFFR_X1 \REGISTERS_reg[50][11]  ( .D(n7936), .CK(CLK), .RN(n12571), .Q(n9355), .QN(n13704) );
  DFFR_X1 \REGISTERS_reg[50][10]  ( .D(n7937), .CK(CLK), .RN(n12549), .Q(n9354), .QN(n13705) );
  DFFR_X1 \REGISTERS_reg[50][9]  ( .D(n7938), .CK(CLK), .RN(n12556), .Q(n9353), 
        .QN(n13706) );
  DFFR_X1 \REGISTERS_reg[50][8]  ( .D(n7939), .CK(CLK), .RN(n12534), .Q(n9352), 
        .QN(n13707) );
  DFFR_X1 \REGISTERS_reg[50][7]  ( .D(n7940), .CK(CLK), .RN(n12644), .Q(n9351), 
        .QN(n13708) );
  DFFR_X1 \REGISTERS_reg[50][6]  ( .D(n7941), .CK(CLK), .RN(n12600), .Q(n9350), 
        .QN(n13709) );
  DFFR_X1 \REGISTERS_reg[50][5]  ( .D(n7942), .CK(CLK), .RN(n12487), .Q(n9349), 
        .QN(n13710) );
  DFFR_X1 \REGISTERS_reg[50][4]  ( .D(n7943), .CK(CLK), .RN(n12494), .Q(n9348), 
        .QN(n13711) );
  DFFR_X1 \REGISTERS_reg[50][3]  ( .D(n7944), .CK(CLK), .RN(n12578), .Q(n9347), 
        .QN(n13712) );
  DFFR_X1 \REGISTERS_reg[50][2]  ( .D(n7945), .CK(CLK), .RN(n12509), .Q(n9346), 
        .QN(n13713) );
  DFFR_X1 \REGISTERS_reg[50][1]  ( .D(n7946), .CK(CLK), .RN(n12437), .Q(n9345), 
        .QN(n13714) );
  DFFR_X1 \REGISTERS_reg[50][0]  ( .D(n7947), .CK(CLK), .RN(n12652), .Q(n9344), 
        .QN(n13715) );
  DFFR_X1 \REGISTERS_reg[51][31]  ( .D(n7948), .CK(CLK), .RN(n12659), .Q(n9343), .QN(n13716) );
  DFFR_X1 \REGISTERS_reg[51][30]  ( .D(n7949), .CK(CLK), .RN(n12622), .Q(n9342), .QN(n13717) );
  DFFR_X1 \REGISTERS_reg[51][29]  ( .D(n7950), .CK(CLK), .RN(n12608), .Q(n9341), .QN(n13718) );
  DFFR_X1 \REGISTERS_reg[51][28]  ( .D(n7951), .CK(CLK), .RN(n12615), .Q(n9340), .QN(n13719) );
  DFFR_X1 \REGISTERS_reg[51][27]  ( .D(n7952), .CK(CLK), .RN(n12586), .Q(n9339), .QN(n13720) );
  DFFR_X1 \REGISTERS_reg[51][26]  ( .D(n7953), .CK(CLK), .RN(n12564), .Q(n9338), .QN(n13721) );
  DFFR_X1 \REGISTERS_reg[51][25]  ( .D(n7954), .CK(CLK), .RN(n12542), .Q(n9337), .QN(n13722) );
  DFFR_X1 \REGISTERS_reg[51][24]  ( .D(n7955), .CK(CLK), .RN(n12516), .Q(n9336), .QN(n13723) );
  DFFR_X1 \REGISTERS_reg[51][23]  ( .D(n7956), .CK(CLK), .RN(n12630), .Q(n9335), .QN(n13724) );
  DFFR_X1 \REGISTERS_reg[51][22]  ( .D(n7957), .CK(CLK), .RN(n12520), .Q(n9334), .QN(n13725) );
  DFFR_X1 \REGISTERS_reg[51][21]  ( .D(n7958), .CK(CLK), .RN(n12527), .Q(n9333), .QN(n13726) );
  DFFR_X1 \REGISTERS_reg[51][20]  ( .D(n7959), .CK(CLK), .RN(n12502), .Q(n9332), .QN(n13727) );
  DFFR_X1 \REGISTERS_reg[51][19]  ( .D(n7960), .CK(CLK), .RN(n12593), .Q(n9331), .QN(n13728) );
  DFFR_X1 \REGISTERS_reg[51][18]  ( .D(n7961), .CK(CLK), .RN(n12444), .Q(n9330), .QN(n13729) );
  DFFR_X1 \REGISTERS_reg[51][17]  ( .D(n7962), .CK(CLK), .RN(n12451), .Q(n9329), .QN(n13730) );
  DFFR_X1 \REGISTERS_reg[51][16]  ( .D(n7963), .CK(CLK), .RN(n12458), .Q(n9328), .QN(n13731) );
  DFFR_X1 \REGISTERS_reg[51][15]  ( .D(n7964), .CK(CLK), .RN(n12637), .Q(n9327), .QN(n13732) );
  DFFR_X1 \REGISTERS_reg[51][14]  ( .D(n7965), .CK(CLK), .RN(n12465), .Q(n9326), .QN(n13733) );
  DFFR_X1 \REGISTERS_reg[51][13]  ( .D(n7966), .CK(CLK), .RN(n12472), .Q(n9325), .QN(n13734) );
  DFFR_X1 \REGISTERS_reg[51][12]  ( .D(n7967), .CK(CLK), .RN(n12480), .Q(n9324), .QN(n13735) );
  DFFR_X1 \REGISTERS_reg[51][11]  ( .D(n7968), .CK(CLK), .RN(n12571), .Q(n9323), .QN(n13736) );
  DFFR_X1 \REGISTERS_reg[51][10]  ( .D(n7969), .CK(CLK), .RN(n12549), .Q(n9322), .QN(n13737) );
  DFFR_X1 \REGISTERS_reg[51][9]  ( .D(n7970), .CK(CLK), .RN(n12556), .Q(n9321), 
        .QN(n13738) );
  DFFR_X1 \REGISTERS_reg[51][8]  ( .D(n7971), .CK(CLK), .RN(n12534), .Q(n9320), 
        .QN(n13739) );
  DFFR_X1 \REGISTERS_reg[51][7]  ( .D(n7972), .CK(CLK), .RN(n12644), .Q(n9319), 
        .QN(n13740) );
  DFFR_X1 \REGISTERS_reg[51][6]  ( .D(n7973), .CK(CLK), .RN(n12600), .Q(n9318), 
        .QN(n13741) );
  DFFR_X1 \REGISTERS_reg[51][5]  ( .D(n7974), .CK(CLK), .RN(n12487), .Q(n9317), 
        .QN(n13742) );
  DFFR_X1 \REGISTERS_reg[51][4]  ( .D(n7975), .CK(CLK), .RN(n12494), .Q(n9316), 
        .QN(n13743) );
  DFFR_X1 \REGISTERS_reg[51][3]  ( .D(n7976), .CK(CLK), .RN(n12578), .Q(n9315), 
        .QN(n13744) );
  DFFR_X1 \REGISTERS_reg[51][2]  ( .D(n7977), .CK(CLK), .RN(n12509), .Q(n9314), 
        .QN(n13745) );
  DFFR_X1 \REGISTERS_reg[51][1]  ( .D(n7978), .CK(CLK), .RN(n12437), .Q(n9313), 
        .QN(n13746) );
  DFFR_X1 \REGISTERS_reg[51][0]  ( .D(n7979), .CK(CLK), .RN(n12652), .Q(n9312), 
        .QN(n13747) );
  DFFR_X1 \REGISTERS_reg[52][30]  ( .D(n7981), .CK(CLK), .RN(n12623), .Q(n9310), .QN(n13749) );
  DFFR_X1 \REGISTERS_reg[52][29]  ( .D(n7982), .CK(CLK), .RN(n12608), .Q(n9309), .QN(n13750) );
  DFFR_X1 \REGISTERS_reg[52][28]  ( .D(n7983), .CK(CLK), .RN(n12615), .Q(n9308), .QN(n13751) );
  DFFR_X1 \REGISTERS_reg[52][27]  ( .D(n7984), .CK(CLK), .RN(n12586), .Q(n9307), .QN(n13752) );
  DFFR_X1 \REGISTERS_reg[52][26]  ( .D(n7985), .CK(CLK), .RN(n12564), .Q(n9306), .QN(n13753) );
  DFFR_X1 \REGISTERS_reg[52][25]  ( .D(n7986), .CK(CLK), .RN(n12542), .Q(n9305), .QN(n13754) );
  DFFR_X1 \REGISTERS_reg[52][24]  ( .D(n7987), .CK(CLK), .RN(n12463), .Q(n9304), .QN(n13755) );
  DFFR_X1 \REGISTERS_reg[52][23]  ( .D(n7988), .CK(CLK), .RN(n12630), .Q(n9303), .QN(n13756) );
  DFFR_X1 \REGISTERS_reg[52][22]  ( .D(n7989), .CK(CLK), .RN(n12520), .Q(n9302), .QN(n13757) );
  DFFR_X1 \REGISTERS_reg[52][21]  ( .D(n7990), .CK(CLK), .RN(n12527), .Q(n9301), .QN(n13758) );
  DFFR_X1 \REGISTERS_reg[52][20]  ( .D(n7991), .CK(CLK), .RN(n12502), .Q(n9300), .QN(n13759) );
  DFFR_X1 \REGISTERS_reg[52][19]  ( .D(n7992), .CK(CLK), .RN(n12593), .Q(n9299), .QN(n13760) );
  DFFR_X1 \REGISTERS_reg[52][18]  ( .D(n7993), .CK(CLK), .RN(n12444), .Q(n9298), .QN(n13761) );
  DFFR_X1 \REGISTERS_reg[52][17]  ( .D(n7994), .CK(CLK), .RN(n12452), .Q(n9297), .QN(n13762) );
  DFFR_X1 \REGISTERS_reg[52][16]  ( .D(n7995), .CK(CLK), .RN(n12458), .Q(n9296), .QN(n13763) );
  DFFR_X1 \REGISTERS_reg[52][15]  ( .D(n7996), .CK(CLK), .RN(n12637), .Q(n9295), .QN(n13764) );
  DFFR_X1 \REGISTERS_reg[52][14]  ( .D(n7997), .CK(CLK), .RN(n12465), .Q(n9294), .QN(n13765) );
  DFFR_X1 \REGISTERS_reg[52][13]  ( .D(n7998), .CK(CLK), .RN(n12473), .Q(n9293), .QN(n13766) );
  DFFR_X1 \REGISTERS_reg[52][12]  ( .D(n7999), .CK(CLK), .RN(n12480), .Q(n9292), .QN(n13767) );
  DFFR_X1 \REGISTERS_reg[52][11]  ( .D(n8000), .CK(CLK), .RN(n12571), .Q(n9291), .QN(n13768) );
  DFFR_X1 \REGISTERS_reg[52][10]  ( .D(n8001), .CK(CLK), .RN(n12549), .Q(n9290), .QN(n13769) );
  DFFR_X1 \REGISTERS_reg[52][9]  ( .D(n8002), .CK(CLK), .RN(n12557), .Q(n9289), 
        .QN(n13770) );
  DFFR_X1 \REGISTERS_reg[52][8]  ( .D(n8003), .CK(CLK), .RN(n12535), .Q(n9288), 
        .QN(n13771) );
  DFFR_X1 \REGISTERS_reg[52][7]  ( .D(n8004), .CK(CLK), .RN(n12645), .Q(n9287), 
        .QN(n13772) );
  DFFR_X1 \REGISTERS_reg[52][6]  ( .D(n8005), .CK(CLK), .RN(n12601), .Q(n9286), 
        .QN(n13773) );
  DFFR_X1 \REGISTERS_reg[52][5]  ( .D(n8006), .CK(CLK), .RN(n12487), .Q(n9285), 
        .QN(n13774) );
  DFFR_X1 \REGISTERS_reg[52][4]  ( .D(n8007), .CK(CLK), .RN(n12495), .Q(n9284), 
        .QN(n13775) );
  DFFR_X1 \REGISTERS_reg[52][3]  ( .D(n8008), .CK(CLK), .RN(n12579), .Q(n9283), 
        .QN(n13776) );
  DFFR_X1 \REGISTERS_reg[52][2]  ( .D(n8009), .CK(CLK), .RN(n12509), .Q(n9282), 
        .QN(n13777) );
  DFFR_X1 \REGISTERS_reg[52][1]  ( .D(n8010), .CK(CLK), .RN(n12437), .Q(n9281), 
        .QN(n13778) );
  DFFR_X1 \REGISTERS_reg[52][0]  ( .D(n8011), .CK(CLK), .RN(n12652), .Q(n9280), 
        .QN(n13779) );
  DFFR_X1 \REGISTERS_reg[53][31]  ( .D(n8012), .CK(CLK), .RN(n12659), .Q(n9279), .QN(n13780) );
  DFFR_X1 \REGISTERS_reg[53][30]  ( .D(n8013), .CK(CLK), .RN(n12623), .Q(n9278), .QN(n13781) );
  DFFR_X1 \REGISTERS_reg[53][29]  ( .D(n8014), .CK(CLK), .RN(n12608), .Q(n9277), .QN(n13782) );
  DFFR_X1 \REGISTERS_reg[53][28]  ( .D(n8015), .CK(CLK), .RN(n12615), .Q(n9276), .QN(n13783) );
  DFFR_X1 \REGISTERS_reg[53][27]  ( .D(n8016), .CK(CLK), .RN(n12586), .Q(n9275), .QN(n13784) );
  DFFR_X1 \REGISTERS_reg[53][26]  ( .D(n8017), .CK(CLK), .RN(n12564), .Q(n9274), .QN(n13785) );
  DFFR_X1 \REGISTERS_reg[53][25]  ( .D(n8018), .CK(CLK), .RN(n12542), .Q(n9273), .QN(n13786) );
  DFFR_X1 \REGISTERS_reg[53][24]  ( .D(n8019), .CK(CLK), .RN(n12462), .Q(n9272), .QN(n13787) );
  DFFR_X1 \REGISTERS_reg[53][23]  ( .D(n8020), .CK(CLK), .RN(n12630), .Q(n9271), .QN(n13788) );
  DFFR_X1 \REGISTERS_reg[53][22]  ( .D(n8021), .CK(CLK), .RN(n12520), .Q(n9270), .QN(n13789) );
  DFFR_X1 \REGISTERS_reg[53][21]  ( .D(n8022), .CK(CLK), .RN(n12527), .Q(n9269), .QN(n13790) );
  DFFR_X1 \REGISTERS_reg[53][20]  ( .D(n8023), .CK(CLK), .RN(n12502), .Q(n9268), .QN(n13791) );
  DFFR_X1 \REGISTERS_reg[53][19]  ( .D(n8024), .CK(CLK), .RN(n12593), .Q(n9267), .QN(n13792) );
  DFFR_X1 \REGISTERS_reg[53][18]  ( .D(n8025), .CK(CLK), .RN(n12444), .Q(n9266), .QN(n13793) );
  DFFR_X1 \REGISTERS_reg[53][17]  ( .D(n8026), .CK(CLK), .RN(n12452), .Q(n9265), .QN(n13794) );
  DFFR_X1 \REGISTERS_reg[54][31]  ( .D(n8044), .CK(CLK), .RN(n12659), .Q(n9247), .QN(n13812) );
  DFFR_X1 \REGISTERS_reg[54][30]  ( .D(n8045), .CK(CLK), .RN(n12623), .Q(n9246), .QN(n13813) );
  DFFR_X1 \REGISTERS_reg[54][29]  ( .D(n8046), .CK(CLK), .RN(n12608), .Q(n9245), .QN(n13814) );
  DFFR_X1 \REGISTERS_reg[54][28]  ( .D(n8047), .CK(CLK), .RN(n12615), .Q(n9244), .QN(n13815) );
  DFFR_X1 \REGISTERS_reg[54][27]  ( .D(n8048), .CK(CLK), .RN(n12586), .Q(n9243), .QN(n13816) );
  DFFR_X1 \REGISTERS_reg[54][26]  ( .D(n8049), .CK(CLK), .RN(n12564), .Q(n9242), .QN(n13817) );
  DFFR_X1 \REGISTERS_reg[54][25]  ( .D(n8050), .CK(CLK), .RN(n12542), .Q(n9241), .QN(n13818) );
  DFFR_X1 \REGISTERS_reg[54][24]  ( .D(n8051), .CK(CLK), .RN(n12481), .Q(n9240), .QN(n13819) );
  DFFR_X1 \REGISTERS_reg[54][23]  ( .D(n8052), .CK(CLK), .RN(n12630), .Q(n9239), .QN(n13820) );
  DFFR_X1 \REGISTERS_reg[54][22]  ( .D(n8053), .CK(CLK), .RN(n12520), .Q(n9238), .QN(n13821) );
  DFFR_X1 \REGISTERS_reg[54][21]  ( .D(n8054), .CK(CLK), .RN(n12527), .Q(n9237), .QN(n13822) );
  DFFR_X1 \REGISTERS_reg[54][20]  ( .D(n8055), .CK(CLK), .RN(n12502), .Q(n9236), .QN(n13823) );
  DFFR_X1 \REGISTERS_reg[54][19]  ( .D(n8056), .CK(CLK), .RN(n12593), .Q(n9235), .QN(n13824) );
  DFFR_X1 \REGISTERS_reg[54][18]  ( .D(n8057), .CK(CLK), .RN(n12444), .Q(n9234), .QN(n13825) );
  DFFR_X1 \REGISTERS_reg[54][17]  ( .D(n8058), .CK(CLK), .RN(n12452), .Q(n9233), .QN(n13826) );
  DFFR_X1 \REGISTERS_reg[54][16]  ( .D(n8059), .CK(CLK), .RN(n12458), .Q(n9232), .QN(n13827) );
  DFFR_X1 \REGISTERS_reg[54][15]  ( .D(n8060), .CK(CLK), .RN(n12637), .Q(n9231), .QN(n13828) );
  DFFR_X1 \REGISTERS_reg[54][14]  ( .D(n8061), .CK(CLK), .RN(n12465), .Q(n9230), .QN(n13829) );
  DFFR_X1 \REGISTERS_reg[54][13]  ( .D(n8062), .CK(CLK), .RN(n12473), .Q(n9229), .QN(n13830) );
  DFFR_X1 \REGISTERS_reg[54][12]  ( .D(n8063), .CK(CLK), .RN(n12480), .Q(n9228), .QN(n13831) );
  DFFR_X1 \REGISTERS_reg[54][11]  ( .D(n8064), .CK(CLK), .RN(n12571), .Q(n9227), .QN(n13832) );
  DFFR_X1 \REGISTERS_reg[54][10]  ( .D(n8065), .CK(CLK), .RN(n12549), .Q(n9226), .QN(n13833) );
  DFFR_X1 \REGISTERS_reg[54][9]  ( .D(n8066), .CK(CLK), .RN(n12557), .Q(n9225), 
        .QN(n13834) );
  DFFR_X1 \REGISTERS_reg[54][8]  ( .D(n8067), .CK(CLK), .RN(n12535), .Q(n9224), 
        .QN(n13835) );
  DFFR_X1 \REGISTERS_reg[54][7]  ( .D(n8068), .CK(CLK), .RN(n12645), .Q(n9223), 
        .QN(n13836) );
  DFFR_X1 \REGISTERS_reg[54][6]  ( .D(n8069), .CK(CLK), .RN(n12601), .Q(n9222), 
        .QN(n13837) );
  DFFR_X1 \REGISTERS_reg[54][5]  ( .D(n8070), .CK(CLK), .RN(n12487), .Q(n9221), 
        .QN(n13838) );
  DFFR_X1 \REGISTERS_reg[54][4]  ( .D(n8071), .CK(CLK), .RN(n12495), .Q(n9220), 
        .QN(n13839) );
  DFFR_X1 \REGISTERS_reg[54][3]  ( .D(n8072), .CK(CLK), .RN(n12579), .Q(n9219), 
        .QN(n13840) );
  DFFR_X1 \REGISTERS_reg[54][2]  ( .D(n8073), .CK(CLK), .RN(n12509), .Q(n9218), 
        .QN(n13841) );
  DFFR_X1 \REGISTERS_reg[54][1]  ( .D(n8074), .CK(CLK), .RN(n12437), .Q(n9217), 
        .QN(n13842) );
  DFFR_X1 \REGISTERS_reg[54][0]  ( .D(n8075), .CK(CLK), .RN(n12652), .Q(n9216), 
        .QN(n13843) );
  DFFR_X1 \REGISTERS_reg[55][31]  ( .D(n8076), .CK(CLK), .RN(n12659), .QN(
        n5721) );
  DFFR_X1 \REGISTERS_reg[55][30]  ( .D(n8077), .CK(CLK), .RN(n12623), .QN(
        n5753) );
  DFFR_X1 \REGISTERS_reg[55][29]  ( .D(n8078), .CK(CLK), .RN(n12608), .QN(
        n5785) );
  DFFR_X1 \REGISTERS_reg[55][28]  ( .D(n8079), .CK(CLK), .RN(n12615), .QN(
        n5817) );
  DFFR_X1 \REGISTERS_reg[55][27]  ( .D(n8080), .CK(CLK), .RN(n12586), .QN(
        n5849) );
  DFFR_X1 \REGISTERS_reg[55][26]  ( .D(n8081), .CK(CLK), .RN(n12564), .QN(
        n5881) );
  DFFR_X1 \REGISTERS_reg[55][25]  ( .D(n8082), .CK(CLK), .RN(n12542), .QN(
        n5913) );
  DFFR_X1 \REGISTERS_reg[55][24]  ( .D(n8083), .CK(CLK), .RN(n12480), .QN(
        n5945) );
  DFFR_X1 \REGISTERS_reg[55][23]  ( .D(n8084), .CK(CLK), .RN(n12630), .QN(
        n6009) );
  DFFR_X1 \REGISTERS_reg[55][22]  ( .D(n8085), .CK(CLK), .RN(n12520), .QN(
        n9144) );
  DFFR_X1 \REGISTERS_reg[55][21]  ( .D(n8086), .CK(CLK), .RN(n12527), .QN(
        n9176) );
  DFFR_X1 \REGISTERS_reg[55][20]  ( .D(n8087), .CK(CLK), .RN(n12502), .QN(
        n9208) );
  DFFR_X1 \REGISTERS_reg[55][19]  ( .D(n8088), .CK(CLK), .RN(n12593), .QN(
        n9574) );
  DFFR_X1 \REGISTERS_reg[55][18]  ( .D(n8089), .CK(CLK), .RN(n12444), .QN(
        n9606) );
  DFFR_X1 \REGISTERS_reg[55][17]  ( .D(n8090), .CK(CLK), .RN(n12452), .QN(
        n9638) );
  DFFR_X1 \REGISTERS_reg[55][16]  ( .D(n8091), .CK(CLK), .RN(n12458), .QN(
        n10000) );
  DFFR_X1 \REGISTERS_reg[55][15]  ( .D(n8092), .CK(CLK), .RN(n12637), .QN(
        n10032) );
  DFFR_X1 \REGISTERS_reg[55][14]  ( .D(n8093), .CK(CLK), .RN(n12465), .QN(
        n10064) );
  DFFR_X1 \REGISTERS_reg[55][13]  ( .D(n8094), .CK(CLK), .RN(n12473), .QN(
        n10096) );
  DFFR_X1 \REGISTERS_reg[55][12]  ( .D(n8095), .CK(CLK), .RN(n12480), .QN(
        n10128) );
  DFFR_X1 \REGISTERS_reg[55][11]  ( .D(n8096), .CK(CLK), .RN(n12571), .QN(
        n10160) );
  DFFR_X1 \REGISTERS_reg[55][10]  ( .D(n8097), .CK(CLK), .RN(n12549), .QN(
        n10192) );
  DFFR_X1 \REGISTERS_reg[55][9]  ( .D(n8098), .CK(CLK), .RN(n12557), .QN(
        n10226) );
  DFFR_X1 \REGISTERS_reg[55][8]  ( .D(n8099), .CK(CLK), .RN(n12535), .QN(
        n10258) );
  DFFR_X1 \REGISTERS_reg[55][7]  ( .D(n8100), .CK(CLK), .RN(n12645), .QN(
        n10290) );
  DFFR_X1 \REGISTERS_reg[55][6]  ( .D(n8101), .CK(CLK), .RN(n12601), .QN(
        n10325) );
  DFFR_X1 \REGISTERS_reg[55][5]  ( .D(n8102), .CK(CLK), .RN(n12487), .QN(
        n10357) );
  DFFR_X1 \REGISTERS_reg[55][4]  ( .D(n8103), .CK(CLK), .RN(n12495), .QN(
        n10389) );
  DFFR_X1 \REGISTERS_reg[55][3]  ( .D(n8104), .CK(CLK), .RN(n12579), .QN(
        n10424) );
  DFFR_X1 \REGISTERS_reg[55][2]  ( .D(n8105), .CK(CLK), .RN(n12509), .QN(
        n10456) );
  DFFR_X1 \REGISTERS_reg[55][1]  ( .D(n8106), .CK(CLK), .RN(n12437), .QN(
        n10488) );
  DFFR_X1 \REGISTERS_reg[55][0]  ( .D(n8107), .CK(CLK), .RN(n12652), .QN(
        n10520) );
  DFFR_X1 \REGISTERS_reg[56][31]  ( .D(n8108), .CK(CLK), .RN(n12660), .QN(
        n5720) );
  DFFR_X1 \REGISTERS_reg[56][30]  ( .D(n8109), .CK(CLK), .RN(n12623), .QN(
        n5752) );
  DFFR_X1 \REGISTERS_reg[56][29]  ( .D(n8110), .CK(CLK), .RN(n12608), .QN(
        n5784) );
  DFFR_X1 \REGISTERS_reg[56][28]  ( .D(n8111), .CK(CLK), .RN(n12616), .QN(
        n5816) );
  DFFR_X1 \REGISTERS_reg[56][27]  ( .D(n8112), .CK(CLK), .RN(n12586), .QN(
        n5848) );
  DFFR_X1 \REGISTERS_reg[56][26]  ( .D(n8113), .CK(CLK), .RN(n12564), .QN(
        n5880) );
  DFFR_X1 \REGISTERS_reg[56][25]  ( .D(n8114), .CK(CLK), .RN(n12542), .QN(
        n5912) );
  DFFR_X1 \REGISTERS_reg[56][24]  ( .D(n8115), .CK(CLK), .RN(n12479), .QN(
        n5944) );
  DFFR_X1 \REGISTERS_reg[56][23]  ( .D(n8116), .CK(CLK), .RN(n12630), .QN(
        n6008) );
  DFFR_X1 \REGISTERS_reg[56][22]  ( .D(n8117), .CK(CLK), .RN(n12520), .QN(
        n9143) );
  DFFR_X1 \REGISTERS_reg[56][21]  ( .D(n8118), .CK(CLK), .RN(n12528), .QN(
        n9175) );
  DFFR_X1 \REGISTERS_reg[56][20]  ( .D(n8119), .CK(CLK), .RN(n12502), .QN(
        n9207) );
  DFFR_X1 \REGISTERS_reg[56][19]  ( .D(n8120), .CK(CLK), .RN(n12594), .QN(
        n9573) );
  DFFR_X1 \REGISTERS_reg[56][18]  ( .D(n8121), .CK(CLK), .RN(n12445), .QN(
        n9605) );
  DFFR_X1 \REGISTERS_reg[56][17]  ( .D(n8122), .CK(CLK), .RN(n12452), .QN(
        n9637) );
  DFFR_X1 \REGISTERS_reg[56][16]  ( .D(n8123), .CK(CLK), .RN(n12458), .QN(
        n9701) );
  DFFR_X1 \REGISTERS_reg[56][15]  ( .D(n8124), .CK(CLK), .RN(n12638), .QN(
        n10031) );
  DFFR_X1 \REGISTERS_reg[56][14]  ( .D(n8125), .CK(CLK), .RN(n12466), .QN(
        n10063) );
  DFFR_X1 \REGISTERS_reg[56][13]  ( .D(n8126), .CK(CLK), .RN(n12473), .QN(
        n10095) );
  DFFR_X1 \REGISTERS_reg[56][12]  ( .D(n8127), .CK(CLK), .RN(n12480), .QN(
        n10127) );
  DFFR_X1 \REGISTERS_reg[56][11]  ( .D(n8128), .CK(CLK), .RN(n12572), .QN(
        n10159) );
  DFFR_X1 \REGISTERS_reg[56][10]  ( .D(n8129), .CK(CLK), .RN(n12550), .QN(
        n10191) );
  DFFR_X1 \REGISTERS_reg[56][9]  ( .D(n8130), .CK(CLK), .RN(n12557), .QN(
        n10225) );
  DFFR_X1 \REGISTERS_reg[56][8]  ( .D(n8131), .CK(CLK), .RN(n12535), .QN(
        n10257) );
  DFFR_X1 \REGISTERS_reg[56][7]  ( .D(n8132), .CK(CLK), .RN(n12645), .QN(
        n10289) );
  DFFR_X1 \REGISTERS_reg[56][6]  ( .D(n8133), .CK(CLK), .RN(n12601), .QN(
        n10324) );
  DFFR_X1 \REGISTERS_reg[56][5]  ( .D(n8134), .CK(CLK), .RN(n12488), .QN(
        n10356) );
  DFFR_X1 \REGISTERS_reg[56][4]  ( .D(n8135), .CK(CLK), .RN(n12495), .QN(
        n10388) );
  DFFR_X1 \REGISTERS_reg[56][3]  ( .D(n8136), .CK(CLK), .RN(n12579), .QN(
        n10423) );
  DFFR_X1 \REGISTERS_reg[56][2]  ( .D(n8137), .CK(CLK), .RN(n12510), .QN(
        n10455) );
  DFFR_X1 \REGISTERS_reg[56][1]  ( .D(n8138), .CK(CLK), .RN(n12437), .QN(
        n10487) );
  DFFR_X1 \REGISTERS_reg[56][0]  ( .D(n8139), .CK(CLK), .RN(n12652), .QN(
        n10519) );
  DFFR_X1 \REGISTERS_reg[57][31]  ( .D(n8140), .CK(CLK), .RN(n12660), .QN(
        n5718) );
  DFFR_X1 \REGISTERS_reg[57][30]  ( .D(n8141), .CK(CLK), .RN(n12623), .QN(
        n5750) );
  DFFR_X1 \REGISTERS_reg[57][29]  ( .D(n8142), .CK(CLK), .RN(n12608), .QN(
        n5782) );
  DFFR_X1 \REGISTERS_reg[57][28]  ( .D(n8143), .CK(CLK), .RN(n12616), .QN(
        n5814) );
  DFFR_X1 \REGISTERS_reg[57][27]  ( .D(n8144), .CK(CLK), .RN(n12586), .QN(
        n5846) );
  DFFR_X1 \REGISTERS_reg[57][26]  ( .D(n8145), .CK(CLK), .RN(n12564), .QN(
        n5878) );
  DFFR_X1 \REGISTERS_reg[57][25]  ( .D(n8146), .CK(CLK), .RN(n12542), .QN(
        n5910) );
  DFFR_X1 \REGISTERS_reg[57][24]  ( .D(n8147), .CK(CLK), .RN(n12478), .QN(
        n5942) );
  DFFR_X1 \REGISTERS_reg[57][23]  ( .D(n8148), .CK(CLK), .RN(n12630), .QN(
        n6006) );
  DFFR_X1 \REGISTERS_reg[57][22]  ( .D(n8149), .CK(CLK), .RN(n12520), .QN(
        n9141) );
  DFFR_X1 \REGISTERS_reg[57][21]  ( .D(n8150), .CK(CLK), .RN(n12528), .QN(
        n9173) );
  DFFR_X1 \REGISTERS_reg[57][20]  ( .D(n8151), .CK(CLK), .RN(n12502), .QN(
        n9205) );
  DFFR_X1 \REGISTERS_reg[57][19]  ( .D(n8152), .CK(CLK), .RN(n12594), .QN(
        n9571) );
  DFFR_X1 \REGISTERS_reg[57][18]  ( .D(n8153), .CK(CLK), .RN(n12445), .QN(
        n9603) );
  DFFR_X1 \REGISTERS_reg[57][17]  ( .D(n8154), .CK(CLK), .RN(n12452), .QN(
        n9635) );
  DFFR_X1 \REGISTERS_reg[57][16]  ( .D(n8155), .CK(CLK), .RN(n12458), .QN(
        n9699) );
  DFFR_X1 \REGISTERS_reg[57][15]  ( .D(n8156), .CK(CLK), .RN(n12638), .QN(
        n10029) );
  DFFR_X1 \REGISTERS_reg[57][14]  ( .D(n8157), .CK(CLK), .RN(n12466), .QN(
        n10061) );
  DFFR_X1 \REGISTERS_reg[57][13]  ( .D(n8158), .CK(CLK), .RN(n12473), .QN(
        n10093) );
  DFFR_X1 \REGISTERS_reg[57][12]  ( .D(n8159), .CK(CLK), .RN(n12480), .QN(
        n10125) );
  DFFR_X1 \REGISTERS_reg[57][11]  ( .D(n8160), .CK(CLK), .RN(n12572), .QN(
        n10157) );
  DFFR_X1 \REGISTERS_reg[57][10]  ( .D(n8161), .CK(CLK), .RN(n12550), .QN(
        n10189) );
  DFFR_X1 \REGISTERS_reg[57][9]  ( .D(n8162), .CK(CLK), .RN(n12557), .QN(
        n10223) );
  DFFR_X1 \REGISTERS_reg[57][8]  ( .D(n8163), .CK(CLK), .RN(n12535), .QN(
        n10255) );
  DFFR_X1 \REGISTERS_reg[57][7]  ( .D(n8164), .CK(CLK), .RN(n12645), .QN(
        n10287) );
  DFFR_X1 \REGISTERS_reg[57][6]  ( .D(n8165), .CK(CLK), .RN(n12601), .QN(
        n10322) );
  DFFR_X1 \REGISTERS_reg[57][5]  ( .D(n8166), .CK(CLK), .RN(n12488), .QN(
        n10354) );
  DFFR_X1 \REGISTERS_reg[57][4]  ( .D(n8167), .CK(CLK), .RN(n12495), .QN(
        n10386) );
  DFFR_X1 \REGISTERS_reg[57][3]  ( .D(n8168), .CK(CLK), .RN(n12579), .QN(
        n10421) );
  DFFR_X1 \REGISTERS_reg[57][2]  ( .D(n8169), .CK(CLK), .RN(n12510), .QN(
        n10453) );
  DFFR_X1 \REGISTERS_reg[57][1]  ( .D(n8170), .CK(CLK), .RN(n12437), .QN(
        n10485) );
  DFFR_X1 \REGISTERS_reg[57][0]  ( .D(n8171), .CK(CLK), .RN(n12652), .QN(
        n10517) );
  DFFR_X1 \REGISTERS_reg[58][31]  ( .D(n8172), .CK(CLK), .RN(n12660), .QN(
        n5719) );
  DFFR_X1 \REGISTERS_reg[58][30]  ( .D(n8173), .CK(CLK), .RN(n12623), .QN(
        n5751) );
  DFFR_X1 \REGISTERS_reg[58][29]  ( .D(n8174), .CK(CLK), .RN(n12608), .QN(
        n5783) );
  DFFR_X1 \REGISTERS_reg[58][28]  ( .D(n8175), .CK(CLK), .RN(n12616), .QN(
        n5815) );
  DFFR_X1 \REGISTERS_reg[58][27]  ( .D(n8176), .CK(CLK), .RN(n12586), .QN(
        n5847) );
  DFFR_X1 \REGISTERS_reg[58][26]  ( .D(n8177), .CK(CLK), .RN(n12564), .QN(
        n5879) );
  DFFR_X1 \REGISTERS_reg[58][25]  ( .D(n8178), .CK(CLK), .RN(n12542), .QN(
        n5911) );
  DFFR_X1 \REGISTERS_reg[58][24]  ( .D(n8179), .CK(CLK), .RN(n12477), .QN(
        n5943) );
  DFFR_X1 \REGISTERS_reg[58][23]  ( .D(n8180), .CK(CLK), .RN(n12630), .QN(
        n6007) );
  DFFR_X1 \REGISTERS_reg[58][22]  ( .D(n8181), .CK(CLK), .RN(n12520), .QN(
        n9142) );
  DFFR_X1 \REGISTERS_reg[58][21]  ( .D(n8182), .CK(CLK), .RN(n12528), .QN(
        n9174) );
  DFFR_X1 \REGISTERS_reg[58][20]  ( .D(n8183), .CK(CLK), .RN(n12502), .QN(
        n9206) );
  DFFR_X1 \REGISTERS_reg[58][19]  ( .D(n8184), .CK(CLK), .RN(n12594), .QN(
        n9572) );
  DFFR_X1 \REGISTERS_reg[58][18]  ( .D(n8185), .CK(CLK), .RN(n12445), .QN(
        n9604) );
  DFFR_X1 \REGISTERS_reg[58][17]  ( .D(n8186), .CK(CLK), .RN(n12452), .QN(
        n9636) );
  DFFR_X1 \REGISTERS_reg[58][16]  ( .D(n8187), .CK(CLK), .RN(n12458), .QN(
        n9700) );
  DFFR_X1 \REGISTERS_reg[58][15]  ( .D(n8188), .CK(CLK), .RN(n12638), .QN(
        n10030) );
  DFFR_X1 \REGISTERS_reg[58][14]  ( .D(n8189), .CK(CLK), .RN(n12466), .QN(
        n10062) );
  DFFR_X1 \REGISTERS_reg[58][13]  ( .D(n8190), .CK(CLK), .RN(n12473), .QN(
        n10094) );
  DFFR_X1 \REGISTERS_reg[58][12]  ( .D(n8191), .CK(CLK), .RN(n12480), .QN(
        n10126) );
  DFFR_X1 \REGISTERS_reg[58][11]  ( .D(n8192), .CK(CLK), .RN(n12572), .QN(
        n10158) );
  DFFR_X1 \REGISTERS_reg[58][10]  ( .D(n8193), .CK(CLK), .RN(n12550), .QN(
        n10190) );
  DFFR_X1 \REGISTERS_reg[58][9]  ( .D(n8194), .CK(CLK), .RN(n12557), .QN(
        n10224) );
  DFFR_X1 \REGISTERS_reg[58][8]  ( .D(n8195), .CK(CLK), .RN(n12535), .QN(
        n10256) );
  DFFR_X1 \REGISTERS_reg[58][7]  ( .D(n8196), .CK(CLK), .RN(n12645), .QN(
        n10288) );
  DFFR_X1 \REGISTERS_reg[58][6]  ( .D(n8197), .CK(CLK), .RN(n12601), .QN(
        n10323) );
  DFFR_X1 \REGISTERS_reg[58][5]  ( .D(n8198), .CK(CLK), .RN(n12488), .QN(
        n10355) );
  DFFR_X1 \REGISTERS_reg[58][4]  ( .D(n8199), .CK(CLK), .RN(n12495), .QN(
        n10387) );
  DFFR_X1 \REGISTERS_reg[58][3]  ( .D(n8200), .CK(CLK), .RN(n12579), .QN(
        n10422) );
  DFFR_X1 \REGISTERS_reg[58][2]  ( .D(n8201), .CK(CLK), .RN(n12510), .QN(
        n10454) );
  DFFR_X1 \REGISTERS_reg[58][1]  ( .D(n8202), .CK(CLK), .RN(n12437), .QN(
        n10486) );
  DFFR_X1 \REGISTERS_reg[58][0]  ( .D(n8203), .CK(CLK), .RN(n12652), .QN(
        n10518) );
  DFFR_X1 \REGISTERS_reg[59][31]  ( .D(n8204), .CK(CLK), .RN(n12660), .QN(
        n5717) );
  DFFR_X1 \REGISTERS_reg[59][30]  ( .D(n8205), .CK(CLK), .RN(n12623), .QN(
        n5749) );
  DFFR_X1 \REGISTERS_reg[59][29]  ( .D(n8206), .CK(CLK), .RN(n12608), .QN(
        n5781) );
  DFFR_X1 \REGISTERS_reg[59][28]  ( .D(n8207), .CK(CLK), .RN(n12616), .QN(
        n5813) );
  DFFR_X1 \REGISTERS_reg[59][27]  ( .D(n8208), .CK(CLK), .RN(n12586), .QN(
        n5845) );
  DFFR_X1 \REGISTERS_reg[59][26]  ( .D(n8209), .CK(CLK), .RN(n12564), .QN(
        n5877) );
  DFFR_X1 \REGISTERS_reg[59][25]  ( .D(n8210), .CK(CLK), .RN(n12542), .QN(
        n5909) );
  DFFR_X1 \REGISTERS_reg[59][24]  ( .D(n8211), .CK(CLK), .RN(n12476), .QN(
        n5941) );
  DFFR_X1 \REGISTERS_reg[59][23]  ( .D(n8212), .CK(CLK), .RN(n12630), .QN(
        n6005) );
  DFFR_X1 \REGISTERS_reg[59][22]  ( .D(n8213), .CK(CLK), .RN(n12520), .QN(
        n9140) );
  DFFR_X1 \REGISTERS_reg[59][21]  ( .D(n8214), .CK(CLK), .RN(n12528), .QN(
        n9172) );
  DFFR_X1 \REGISTERS_reg[59][20]  ( .D(n8215), .CK(CLK), .RN(n12502), .QN(
        n9204) );
  DFFR_X1 \REGISTERS_reg[59][19]  ( .D(n8216), .CK(CLK), .RN(n12594), .QN(
        n9570) );
  DFFR_X1 \REGISTERS_reg[59][18]  ( .D(n8217), .CK(CLK), .RN(n12445), .QN(
        n9602) );
  DFFR_X1 \REGISTERS_reg[59][17]  ( .D(n8218), .CK(CLK), .RN(n12452), .QN(
        n9634) );
  DFFR_X1 \REGISTERS_reg[59][16]  ( .D(n8219), .CK(CLK), .RN(n12458), .QN(
        n9698) );
  DFFR_X1 \REGISTERS_reg[59][15]  ( .D(n8220), .CK(CLK), .RN(n12638), .QN(
        n10028) );
  DFFR_X1 \REGISTERS_reg[59][14]  ( .D(n8221), .CK(CLK), .RN(n12466), .QN(
        n10060) );
  DFFR_X1 \REGISTERS_reg[59][13]  ( .D(n8222), .CK(CLK), .RN(n12473), .QN(
        n10092) );
  DFFR_X1 \REGISTERS_reg[59][12]  ( .D(n8223), .CK(CLK), .RN(n12480), .QN(
        n10124) );
  DFFR_X1 \REGISTERS_reg[59][11]  ( .D(n8224), .CK(CLK), .RN(n12572), .QN(
        n10156) );
  DFFR_X1 \REGISTERS_reg[59][10]  ( .D(n8225), .CK(CLK), .RN(n12550), .QN(
        n10188) );
  DFFR_X1 \REGISTERS_reg[59][9]  ( .D(n8226), .CK(CLK), .RN(n12557), .QN(
        n10222) );
  DFFR_X1 \REGISTERS_reg[59][8]  ( .D(n8227), .CK(CLK), .RN(n12535), .QN(
        n10254) );
  DFFR_X1 \REGISTERS_reg[59][7]  ( .D(n8228), .CK(CLK), .RN(n12645), .QN(
        n10286) );
  DFFR_X1 \REGISTERS_reg[59][6]  ( .D(n8229), .CK(CLK), .RN(n12601), .QN(
        n10321) );
  DFFR_X1 \REGISTERS_reg[59][5]  ( .D(n8230), .CK(CLK), .RN(n12488), .QN(
        n10353) );
  DFFR_X1 \REGISTERS_reg[59][4]  ( .D(n8231), .CK(CLK), .RN(n12495), .QN(
        n10385) );
  DFFR_X1 \REGISTERS_reg[59][3]  ( .D(n8232), .CK(CLK), .RN(n12579), .QN(
        n10420) );
  DFFR_X1 \REGISTERS_reg[59][2]  ( .D(n8233), .CK(CLK), .RN(n12510), .QN(
        n10452) );
  DFFR_X1 \REGISTERS_reg[59][1]  ( .D(n8234), .CK(CLK), .RN(n12437), .QN(
        n10484) );
  DFFR_X1 \REGISTERS_reg[59][0]  ( .D(n8235), .CK(CLK), .RN(n12652), .QN(
        n10516) );
  DFFR_X1 \REGISTERS_reg[60][31]  ( .D(n8236), .CK(CLK), .RN(n12660), .QN(
        n5715) );
  DFFR_X1 \REGISTERS_reg[60][30]  ( .D(n8237), .CK(CLK), .RN(n12623), .QN(
        n5747) );
  DFFR_X1 \REGISTERS_reg[60][29]  ( .D(n8238), .CK(CLK), .RN(n12609), .QN(
        n5779) );
  DFFR_X1 \REGISTERS_reg[60][28]  ( .D(n8239), .CK(CLK), .RN(n12616), .QN(
        n5811) );
  DFFR_X1 \REGISTERS_reg[60][27]  ( .D(n8240), .CK(CLK), .RN(n12587), .QN(
        n5843) );
  DFFR_X1 \REGISTERS_reg[60][26]  ( .D(n8241), .CK(CLK), .RN(n12565), .QN(
        n5875) );
  DFFR_X1 \REGISTERS_reg[60][25]  ( .D(n8242), .CK(CLK), .RN(n12543), .QN(
        n5907) );
  DFFR_X1 \REGISTERS_reg[60][24]  ( .D(n8243), .CK(CLK), .RN(n12475), .QN(
        n5939) );
  DFFR_X1 \REGISTERS_reg[60][23]  ( .D(n8244), .CK(CLK), .RN(n12631), .QN(
        n6003) );
  DFFR_X1 \REGISTERS_reg[60][22]  ( .D(n8245), .CK(CLK), .RN(n12521), .QN(
        n9138) );
  DFFR_X1 \REGISTERS_reg[60][21]  ( .D(n8246), .CK(CLK), .RN(n12528), .QN(
        n9170) );
  DFFR_X1 \REGISTERS_reg[60][20]  ( .D(n8247), .CK(CLK), .RN(n12503), .QN(
        n9202) );
  DFFR_X1 \REGISTERS_reg[60][19]  ( .D(n8248), .CK(CLK), .RN(n12594), .QN(
        n9568) );
  DFFR_X1 \REGISTERS_reg[60][18]  ( .D(n8249), .CK(CLK), .RN(n12445), .QN(
        n9600) );
  DFFR_X1 \REGISTERS_reg[60][17]  ( .D(n8250), .CK(CLK), .RN(n12452), .QN(
        n9632) );
  DFFR_X1 \REGISTERS_reg[60][16]  ( .D(n8251), .CK(CLK), .RN(n12459), .QN(
        n9696) );
  DFFR_X1 \REGISTERS_reg[60][15]  ( .D(n8252), .CK(CLK), .RN(n12638), .QN(
        n10026) );
  DFFR_X1 \REGISTERS_reg[60][14]  ( .D(n8253), .CK(CLK), .RN(n12466), .QN(
        n10058) );
  DFFR_X1 \REGISTERS_reg[60][13]  ( .D(n8254), .CK(CLK), .RN(n12473), .QN(
        n10090) );
  DFFR_X1 \REGISTERS_reg[60][12]  ( .D(n8255), .CK(CLK), .RN(n12481), .QN(
        n10122) );
  DFFR_X1 \REGISTERS_reg[60][11]  ( .D(n8256), .CK(CLK), .RN(n12572), .QN(
        n10154) );
  DFFR_X1 \REGISTERS_reg[60][10]  ( .D(n8257), .CK(CLK), .RN(n12550), .QN(
        n10186) );
  DFFR_X1 \REGISTERS_reg[60][9]  ( .D(n8258), .CK(CLK), .RN(n12557), .QN(
        n10220) );
  DFFR_X1 \REGISTERS_reg[60][8]  ( .D(n8259), .CK(CLK), .RN(n12535), .QN(
        n10252) );
  DFFR_X1 \REGISTERS_reg[60][7]  ( .D(n8260), .CK(CLK), .RN(n12645), .QN(
        n10284) );
  DFFR_X1 \REGISTERS_reg[60][6]  ( .D(n8261), .CK(CLK), .RN(n12601), .QN(
        n10319) );
  DFFR_X1 \REGISTERS_reg[60][5]  ( .D(n8262), .CK(CLK), .RN(n12488), .QN(
        n10351) );
  DFFR_X1 \REGISTERS_reg[60][4]  ( .D(n8263), .CK(CLK), .RN(n12495), .QN(
        n10383) );
  DFFR_X1 \REGISTERS_reg[60][3]  ( .D(n8264), .CK(CLK), .RN(n12579), .QN(
        n10418) );
  DFFR_X1 \REGISTERS_reg[60][2]  ( .D(n8265), .CK(CLK), .RN(n12510), .QN(
        n10450) );
  DFFR_X1 \REGISTERS_reg[60][1]  ( .D(n8266), .CK(CLK), .RN(n12438), .QN(
        n10482) );
  DFFR_X1 \REGISTERS_reg[60][0]  ( .D(n8267), .CK(CLK), .RN(n12653), .QN(
        n10514) );
  DFFR_X1 \REGISTERS_reg[61][31]  ( .D(n8268), .CK(CLK), .RN(n12660), .QN(
        n13844) );
  DFFR_X1 \REGISTERS_reg[61][30]  ( .D(n8269), .CK(CLK), .RN(n12623), .QN(
        n13845) );
  DFFR_X1 \REGISTERS_reg[61][29]  ( .D(n8270), .CK(CLK), .RN(n12609), .QN(
        n13846) );
  DFFR_X1 \REGISTERS_reg[61][28]  ( .D(n8271), .CK(CLK), .RN(n12616), .QN(
        n13847) );
  DFFR_X1 \REGISTERS_reg[61][27]  ( .D(n8272), .CK(CLK), .RN(n12587), .QN(
        n13848) );
  DFFR_X1 \REGISTERS_reg[61][26]  ( .D(n8273), .CK(CLK), .RN(n12565), .QN(
        n13849) );
  DFFR_X1 \REGISTERS_reg[61][25]  ( .D(n8274), .CK(CLK), .RN(n12543), .QN(
        n13850) );
  DFFR_X1 \REGISTERS_reg[61][24]  ( .D(n8275), .CK(CLK), .RN(n12488), .QN(
        n13851) );
  DFFR_X1 \REGISTERS_reg[61][23]  ( .D(n8276), .CK(CLK), .RN(n12631), .QN(
        n13852) );
  DFFR_X1 \REGISTERS_reg[61][22]  ( .D(n8277), .CK(CLK), .RN(n12521), .QN(
        n13853) );
  DFFR_X1 \REGISTERS_reg[61][21]  ( .D(n8278), .CK(CLK), .RN(n12528), .QN(
        n13854) );
  DFFR_X1 \REGISTERS_reg[61][20]  ( .D(n8279), .CK(CLK), .RN(n12503), .QN(
        n13855) );
  DFFR_X1 \REGISTERS_reg[61][19]  ( .D(n8280), .CK(CLK), .RN(n12594), .QN(
        n13856) );
  DFFR_X1 \REGISTERS_reg[61][18]  ( .D(n8281), .CK(CLK), .RN(n12445), .QN(
        n13857) );
  DFFR_X1 \REGISTERS_reg[61][17]  ( .D(n8282), .CK(CLK), .RN(n12452), .QN(
        n13858) );
  DFFR_X1 \REGISTERS_reg[61][16]  ( .D(n8283), .CK(CLK), .RN(n12459), .QN(
        n13859) );
  DFFR_X1 \REGISTERS_reg[61][15]  ( .D(n8284), .CK(CLK), .RN(n12638), .QN(
        n13860) );
  DFFR_X1 \REGISTERS_reg[61][14]  ( .D(n8285), .CK(CLK), .RN(n12466), .QN(
        n13861) );
  DFFR_X1 \REGISTERS_reg[61][13]  ( .D(n8286), .CK(CLK), .RN(n12473), .QN(
        n13862) );
  DFFR_X1 \REGISTERS_reg[61][12]  ( .D(n8287), .CK(CLK), .RN(n12481), .QN(
        n13863) );
  DFFR_X1 \REGISTERS_reg[61][11]  ( .D(n8288), .CK(CLK), .RN(n12572), .QN(
        n13864) );
  DFFR_X1 \REGISTERS_reg[61][10]  ( .D(n8289), .CK(CLK), .RN(n12550), .QN(
        n13865) );
  DFFR_X1 \REGISTERS_reg[61][9]  ( .D(n8290), .CK(CLK), .RN(n12557), .QN(
        n13866) );
  DFFR_X1 \REGISTERS_reg[61][8]  ( .D(n8291), .CK(CLK), .RN(n12535), .QN(
        n13867) );
  DFFR_X1 \REGISTERS_reg[61][7]  ( .D(n8292), .CK(CLK), .RN(n12645), .QN(
        n13868) );
  DFFR_X1 \REGISTERS_reg[61][6]  ( .D(n8293), .CK(CLK), .RN(n12601), .QN(
        n13869) );
  DFFR_X1 \REGISTERS_reg[61][5]  ( .D(n8294), .CK(CLK), .RN(n12488), .QN(
        n13870) );
  DFFR_X1 \REGISTERS_reg[61][4]  ( .D(n8295), .CK(CLK), .RN(n12495), .QN(
        n13871) );
  DFFR_X1 \REGISTERS_reg[61][3]  ( .D(n8296), .CK(CLK), .RN(n12579), .QN(
        n13872) );
  DFFR_X1 \REGISTERS_reg[61][2]  ( .D(n8297), .CK(CLK), .RN(n12510), .QN(
        n13873) );
  DFFR_X1 \REGISTERS_reg[61][1]  ( .D(n8298), .CK(CLK), .RN(n12438), .QN(
        n13874) );
  DFFR_X1 \REGISTERS_reg[61][0]  ( .D(n8299), .CK(CLK), .RN(n12653), .QN(
        n13875) );
  DFFR_X1 \REGISTERS_reg[62][31]  ( .D(n8300), .CK(CLK), .RN(n12660), .QN(
        n5716) );
  DFFR_X1 \REGISTERS_reg[62][30]  ( .D(n8301), .CK(CLK), .RN(n12623), .QN(
        n5748) );
  DFFR_X1 \REGISTERS_reg[62][29]  ( .D(n8302), .CK(CLK), .RN(n12609), .QN(
        n5780) );
  DFFR_X1 \REGISTERS_reg[62][28]  ( .D(n8303), .CK(CLK), .RN(n12616), .QN(
        n5812) );
  DFFR_X1 \REGISTERS_reg[62][27]  ( .D(n8304), .CK(CLK), .RN(n12587), .QN(
        n5844) );
  DFFR_X1 \REGISTERS_reg[62][26]  ( .D(n8305), .CK(CLK), .RN(n12565), .QN(
        n5876) );
  DFFR_X1 \REGISTERS_reg[62][25]  ( .D(n8306), .CK(CLK), .RN(n12543), .QN(
        n5908) );
  DFFR_X1 \REGISTERS_reg[62][24]  ( .D(n8307), .CK(CLK), .RN(n12487), .QN(
        n5940) );
  DFFR_X1 \REGISTERS_reg[62][23]  ( .D(n8308), .CK(CLK), .RN(n12631), .QN(
        n6004) );
  DFFR_X1 \REGISTERS_reg[62][22]  ( .D(n8309), .CK(CLK), .RN(n12521), .QN(
        n9139) );
  DFFR_X1 \REGISTERS_reg[62][21]  ( .D(n8310), .CK(CLK), .RN(n12528), .QN(
        n9171) );
  DFFR_X1 \REGISTERS_reg[62][20]  ( .D(n8311), .CK(CLK), .RN(n12503), .QN(
        n9203) );
  DFFR_X1 \REGISTERS_reg[62][19]  ( .D(n8312), .CK(CLK), .RN(n12594), .QN(
        n9569) );
  DFFR_X1 \REGISTERS_reg[62][18]  ( .D(n8313), .CK(CLK), .RN(n12445), .QN(
        n9601) );
  DFFR_X1 \REGISTERS_reg[62][17]  ( .D(n8314), .CK(CLK), .RN(n12452), .QN(
        n9633) );
  DFFR_X1 \REGISTERS_reg[62][16]  ( .D(n8315), .CK(CLK), .RN(n12459), .QN(
        n9697) );
  DFFR_X1 \REGISTERS_reg[62][15]  ( .D(n8316), .CK(CLK), .RN(n12638), .QN(
        n10027) );
  DFFR_X1 \REGISTERS_reg[62][14]  ( .D(n8317), .CK(CLK), .RN(n12466), .QN(
        n10059) );
  DFFR_X1 \REGISTERS_reg[62][13]  ( .D(n8318), .CK(CLK), .RN(n12473), .QN(
        n10091) );
  DFFR_X1 \REGISTERS_reg[62][12]  ( .D(n8319), .CK(CLK), .RN(n12481), .QN(
        n10123) );
  DFFR_X1 \REGISTERS_reg[62][11]  ( .D(n8320), .CK(CLK), .RN(n12572), .QN(
        n10155) );
  DFFR_X1 \REGISTERS_reg[62][10]  ( .D(n8321), .CK(CLK), .RN(n12550), .QN(
        n10187) );
  DFFR_X1 \REGISTERS_reg[62][9]  ( .D(n8322), .CK(CLK), .RN(n12557), .QN(
        n10221) );
  DFFR_X1 \REGISTERS_reg[62][8]  ( .D(n8323), .CK(CLK), .RN(n12535), .QN(
        n10253) );
  DFFR_X1 \REGISTERS_reg[62][7]  ( .D(n8324), .CK(CLK), .RN(n12645), .QN(
        n10285) );
  DFFR_X1 \REGISTERS_reg[62][6]  ( .D(n8325), .CK(CLK), .RN(n12601), .QN(
        n10320) );
  DFFR_X1 \REGISTERS_reg[62][5]  ( .D(n8326), .CK(CLK), .RN(n12488), .QN(
        n10352) );
  DFFR_X1 \REGISTERS_reg[62][4]  ( .D(n8327), .CK(CLK), .RN(n12495), .QN(
        n10384) );
  DFFR_X1 \REGISTERS_reg[62][3]  ( .D(n8328), .CK(CLK), .RN(n12579), .QN(
        n10419) );
  DFFR_X1 \REGISTERS_reg[62][2]  ( .D(n8329), .CK(CLK), .RN(n12510), .QN(
        n10451) );
  DFFR_X1 \REGISTERS_reg[62][1]  ( .D(n8330), .CK(CLK), .RN(n12438), .QN(
        n10483) );
  DFFR_X1 \REGISTERS_reg[62][0]  ( .D(n8331), .CK(CLK), .RN(n12653), .QN(
        n10515) );
  DFFR_X1 \REGISTERS_reg[63][31]  ( .D(n8332), .CK(CLK), .RN(n12660), .QN(
        n13876) );
  DFFR_X1 \REGISTERS_reg[63][30]  ( .D(n8333), .CK(CLK), .RN(n12623), .QN(
        n13877) );
  DFFR_X1 \REGISTERS_reg[63][29]  ( .D(n8334), .CK(CLK), .RN(n12609), .QN(
        n13878) );
  DFFR_X1 \REGISTERS_reg[63][28]  ( .D(n8335), .CK(CLK), .RN(n12616), .QN(
        n13879) );
  DFFR_X1 \REGISTERS_reg[63][27]  ( .D(n8336), .CK(CLK), .RN(n12587), .QN(
        n13880) );
  DFFR_X1 \REGISTERS_reg[63][26]  ( .D(n8337), .CK(CLK), .RN(n12565), .QN(
        n13881) );
  DFFR_X1 \REGISTERS_reg[63][25]  ( .D(n8338), .CK(CLK), .RN(n12543), .QN(
        n13882) );
  DFFR_X1 \REGISTERS_reg[63][24]  ( .D(n8339), .CK(CLK), .RN(n12464), .QN(
        n13883) );
  DFFR_X1 \REGISTERS_reg[63][23]  ( .D(n8340), .CK(CLK), .RN(n12631), .QN(
        n13884) );
  DFFR_X1 \REGISTERS_reg[63][22]  ( .D(n8341), .CK(CLK), .RN(n12521), .QN(
        n13885) );
  DFFR_X1 \REGISTERS_reg[63][21]  ( .D(n8342), .CK(CLK), .RN(n12528), .QN(
        n13886) );
  DFFR_X1 \REGISTERS_reg[63][20]  ( .D(n8343), .CK(CLK), .RN(n12503), .QN(
        n13887) );
  DFFR_X1 \REGISTERS_reg[63][19]  ( .D(n8344), .CK(CLK), .RN(n12594), .QN(
        n13888) );
  DFFR_X1 \REGISTERS_reg[63][18]  ( .D(n8345), .CK(CLK), .RN(n12445), .QN(
        n13889) );
  DFFR_X1 \REGISTERS_reg[63][17]  ( .D(n8346), .CK(CLK), .RN(n12452), .QN(
        n13890) );
  DFFR_X1 \REGISTERS_reg[63][16]  ( .D(n8347), .CK(CLK), .RN(n12459), .QN(
        n13891) );
  DFFR_X1 \REGISTERS_reg[63][15]  ( .D(n8348), .CK(CLK), .RN(n12638), .QN(
        n13892) );
  DFFR_X1 \REGISTERS_reg[63][14]  ( .D(n8349), .CK(CLK), .RN(n12466), .QN(
        n13893) );
  DFFR_X1 \REGISTERS_reg[63][13]  ( .D(n8350), .CK(CLK), .RN(n12473), .QN(
        n13894) );
  DFFR_X1 \REGISTERS_reg[63][12]  ( .D(n8351), .CK(CLK), .RN(n12481), .QN(
        n13895) );
  DFFR_X1 \REGISTERS_reg[63][11]  ( .D(n8352), .CK(CLK), .RN(n12572), .QN(
        n13896) );
  DFFR_X1 \REGISTERS_reg[63][10]  ( .D(n8353), .CK(CLK), .RN(n12550), .QN(
        n13897) );
  DFFR_X1 \REGISTERS_reg[63][9]  ( .D(n8354), .CK(CLK), .RN(n12557), .QN(
        n13898) );
  DFFR_X1 \REGISTERS_reg[63][8]  ( .D(n8355), .CK(CLK), .RN(n12535), .QN(
        n13899) );
  DFFR_X1 \REGISTERS_reg[63][7]  ( .D(n8356), .CK(CLK), .RN(n12645), .QN(
        n13900) );
  DFFR_X1 \REGISTERS_reg[63][6]  ( .D(n8357), .CK(CLK), .RN(n12601), .QN(
        n13901) );
  DFFR_X1 \REGISTERS_reg[63][5]  ( .D(n8358), .CK(CLK), .RN(n12488), .QN(
        n13902) );
  DFFR_X1 \REGISTERS_reg[63][4]  ( .D(n8359), .CK(CLK), .RN(n12495), .QN(
        n13903) );
  DFFR_X1 \REGISTERS_reg[63][3]  ( .D(n8360), .CK(CLK), .RN(n12579), .QN(
        n13904) );
  DFFR_X1 \REGISTERS_reg[63][2]  ( .D(n8361), .CK(CLK), .RN(n12510), .QN(
        n13905) );
  DFFR_X1 \REGISTERS_reg[63][1]  ( .D(n8362), .CK(CLK), .RN(n12438), .QN(
        n13906) );
  DFFR_X1 \REGISTERS_reg[63][0]  ( .D(n8363), .CK(CLK), .RN(n12653), .QN(
        n13907) );
  DFFR_X1 \REGISTERS_reg[64][31]  ( .D(n8364), .CK(CLK), .RN(n12660), .QN(
        n5722) );
  DFFR_X1 \REGISTERS_reg[64][30]  ( .D(n8365), .CK(CLK), .RN(n12624), .QN(
        n5754) );
  DFFR_X1 \REGISTERS_reg[64][29]  ( .D(n8366), .CK(CLK), .RN(n12609), .QN(
        n5786) );
  DFFR_X1 \REGISTERS_reg[64][28]  ( .D(n8367), .CK(CLK), .RN(n12616), .QN(
        n5818) );
  DFFR_X1 \REGISTERS_reg[64][27]  ( .D(n8368), .CK(CLK), .RN(n12587), .QN(
        n5850) );
  DFFR_X1 \REGISTERS_reg[64][26]  ( .D(n8369), .CK(CLK), .RN(n12565), .QN(
        n5882) );
  DFFR_X1 \REGISTERS_reg[64][25]  ( .D(n8370), .CK(CLK), .RN(n12543), .QN(
        n5914) );
  DFFR_X1 \REGISTERS_reg[64][24]  ( .D(n8371), .CK(CLK), .RN(n12449), .QN(
        n5946) );
  DFFR_X1 \REGISTERS_reg[64][23]  ( .D(n8372), .CK(CLK), .RN(n12631), .QN(
        n6010) );
  DFFR_X1 \REGISTERS_reg[64][22]  ( .D(n8373), .CK(CLK), .RN(n12521), .QN(
        n9145) );
  DFFR_X1 \REGISTERS_reg[64][21]  ( .D(n8374), .CK(CLK), .RN(n12528), .QN(
        n9177) );
  DFFR_X1 \REGISTERS_reg[64][20]  ( .D(n8375), .CK(CLK), .RN(n12503), .QN(
        n9209) );
  DFFR_X1 \REGISTERS_reg[64][19]  ( .D(n8376), .CK(CLK), .RN(n12594), .QN(
        n9575) );
  DFFR_X1 \REGISTERS_reg[64][18]  ( .D(n8377), .CK(CLK), .RN(n12445), .QN(
        n9607) );
  DFFR_X1 \REGISTERS_reg[64][17]  ( .D(n8378), .CK(CLK), .RN(n12453), .QN(
        n9639) );
  DFFR_X1 \REGISTERS_reg[64][16]  ( .D(n8379), .CK(CLK), .RN(n12459), .QN(
        n10001) );
  DFFR_X1 \REGISTERS_reg[64][15]  ( .D(n8380), .CK(CLK), .RN(n12638), .QN(
        n10033) );
  DFFR_X1 \REGISTERS_reg[64][14]  ( .D(n8381), .CK(CLK), .RN(n12466), .QN(
        n10065) );
  DFFR_X1 \REGISTERS_reg[64][13]  ( .D(n8382), .CK(CLK), .RN(n12474), .QN(
        n10097) );
  DFFR_X1 \REGISTERS_reg[64][12]  ( .D(n8383), .CK(CLK), .RN(n12481), .QN(
        n10129) );
  DFFR_X1 \REGISTERS_reg[64][11]  ( .D(n8384), .CK(CLK), .RN(n12572), .QN(
        n10161) );
  DFFR_X1 \REGISTERS_reg[64][10]  ( .D(n8385), .CK(CLK), .RN(n12550), .QN(
        n10193) );
  DFFR_X1 \REGISTERS_reg[64][9]  ( .D(n8386), .CK(CLK), .RN(n12558), .QN(
        n10227) );
  DFFR_X1 \REGISTERS_reg[64][8]  ( .D(n8387), .CK(CLK), .RN(n12536), .QN(
        n10259) );
  DFFR_X1 \REGISTERS_reg[64][7]  ( .D(n8388), .CK(CLK), .RN(n12646), .QN(
        n10291) );
  DFFR_X1 \REGISTERS_reg[64][6]  ( .D(n8389), .CK(CLK), .RN(n12602), .QN(
        n10326) );
  DFFR_X1 \REGISTERS_reg[64][5]  ( .D(n8390), .CK(CLK), .RN(n12488), .QN(
        n10358) );
  DFFR_X1 \REGISTERS_reg[64][4]  ( .D(n8391), .CK(CLK), .RN(n12496), .QN(
        n10390) );
  DFFR_X1 \REGISTERS_reg[64][3]  ( .D(n8392), .CK(CLK), .RN(n12580), .QN(
        n10425) );
  DFFR_X1 \REGISTERS_reg[64][2]  ( .D(n8393), .CK(CLK), .RN(n12510), .QN(
        n10457) );
  DFFR_X1 \REGISTERS_reg[64][1]  ( .D(n8394), .CK(CLK), .RN(n12438), .QN(
        n10489) );
  DFFR_X1 \REGISTERS_reg[64][0]  ( .D(n8395), .CK(CLK), .RN(n12653), .QN(
        n10521) );
  DFFR_X1 \REGISTERS_reg[65][31]  ( .D(n8396), .CK(CLK), .RN(n12660), .QN(
        n13908) );
  DFFR_X1 \REGISTERS_reg[65][30]  ( .D(n8397), .CK(CLK), .RN(n12624), .QN(
        n13909) );
  DFFR_X1 \REGISTERS_reg[65][29]  ( .D(n8398), .CK(CLK), .RN(n12609), .QN(
        n13910) );
  DFFR_X1 \REGISTERS_reg[65][28]  ( .D(n8399), .CK(CLK), .RN(n12616), .QN(
        n13911) );
  DFFR_X1 \REGISTERS_reg[65][27]  ( .D(n8400), .CK(CLK), .RN(n12587), .QN(
        n13912) );
  DFFR_X1 \REGISTERS_reg[65][26]  ( .D(n8401), .CK(CLK), .RN(n12565), .QN(
        n13913) );
  DFFR_X1 \REGISTERS_reg[65][25]  ( .D(n8402), .CK(CLK), .RN(n12543), .QN(
        n13914) );
  DFFR_X1 \REGISTERS_reg[65][24]  ( .D(n8403), .CK(CLK), .RN(n12461), .QN(
        n13915) );
  DFFR_X1 \REGISTERS_reg[65][23]  ( .D(n8404), .CK(CLK), .RN(n12631), .QN(
        n13916) );
  DFFR_X1 \REGISTERS_reg[65][22]  ( .D(n8405), .CK(CLK), .RN(n12521), .QN(
        n13917) );
  DFFR_X1 \REGISTERS_reg[65][21]  ( .D(n8406), .CK(CLK), .RN(n12528), .QN(
        n13918) );
  DFFR_X1 \REGISTERS_reg[65][20]  ( .D(n8407), .CK(CLK), .RN(n12503), .QN(
        n13919) );
  DFFR_X1 \REGISTERS_reg[65][19]  ( .D(n8408), .CK(CLK), .RN(n12594), .QN(
        n13920) );
  DFFR_X1 \REGISTERS_reg[65][18]  ( .D(n8409), .CK(CLK), .RN(n12445), .QN(
        n13921) );
  DFFR_X1 \REGISTERS_reg[65][17]  ( .D(n8410), .CK(CLK), .RN(n12453), .QN(
        n13922) );
  DFFR_X1 \REGISTERS_reg[65][16]  ( .D(n8411), .CK(CLK), .RN(n12459), .QN(
        n13923) );
  DFFR_X1 \REGISTERS_reg[65][15]  ( .D(n8412), .CK(CLK), .RN(n12638), .QN(
        n13924) );
  DFFR_X1 \REGISTERS_reg[65][14]  ( .D(n8413), .CK(CLK), .RN(n12466), .QN(
        n13925) );
  DFFR_X1 \REGISTERS_reg[65][13]  ( .D(n8414), .CK(CLK), .RN(n12474), .QN(
        n13926) );
  DFFR_X1 \REGISTERS_reg[65][12]  ( .D(n8415), .CK(CLK), .RN(n12481), .QN(
        n13927) );
  DFFR_X1 \REGISTERS_reg[65][11]  ( .D(n8416), .CK(CLK), .RN(n12572), .QN(
        n13928) );
  DFFR_X1 \REGISTERS_reg[65][10]  ( .D(n8417), .CK(CLK), .RN(n12550), .QN(
        n13929) );
  DFFR_X1 \REGISTERS_reg[65][9]  ( .D(n8418), .CK(CLK), .RN(n12558), .QN(
        n13930) );
  DFFR_X1 \REGISTERS_reg[65][8]  ( .D(n8419), .CK(CLK), .RN(n12536), .QN(
        n13931) );
  DFFR_X1 \REGISTERS_reg[65][7]  ( .D(n8420), .CK(CLK), .RN(n12646), .QN(
        n13932) );
  DFFR_X1 \REGISTERS_reg[65][6]  ( .D(n8421), .CK(CLK), .RN(n12602), .QN(
        n13933) );
  DFFR_X1 \REGISTERS_reg[65][5]  ( .D(n8422), .CK(CLK), .RN(n12488), .QN(
        n13934) );
  DFFR_X1 \REGISTERS_reg[65][4]  ( .D(n8423), .CK(CLK), .RN(n12496), .QN(
        n13935) );
  DFFR_X1 \REGISTERS_reg[65][3]  ( .D(n8424), .CK(CLK), .RN(n12580), .QN(
        n13936) );
  DFFR_X1 \REGISTERS_reg[65][2]  ( .D(n8425), .CK(CLK), .RN(n12510), .QN(
        n13937) );
  DFFR_X1 \REGISTERS_reg[65][1]  ( .D(n8426), .CK(CLK), .RN(n12438), .QN(
        n13938) );
  DFFR_X1 \REGISTERS_reg[65][0]  ( .D(n8427), .CK(CLK), .RN(n12653), .QN(
        n13939) );
  DFFR_X1 \REGISTERS_reg[66][31]  ( .D(n8428), .CK(CLK), .RN(n12660), .QN(
        n13940) );
  DFFR_X1 \REGISTERS_reg[66][30]  ( .D(n8429), .CK(CLK), .RN(n12624), .QN(
        n13941) );
  DFFR_X1 \REGISTERS_reg[66][29]  ( .D(n8430), .CK(CLK), .RN(n12609), .QN(
        n13942) );
  DFFR_X1 \REGISTERS_reg[66][28]  ( .D(n8431), .CK(CLK), .RN(n12616), .QN(
        n13943) );
  DFFR_X1 \REGISTERS_reg[66][27]  ( .D(n8432), .CK(CLK), .RN(n12587), .QN(
        n13944) );
  DFFR_X1 \REGISTERS_reg[66][26]  ( .D(n8433), .CK(CLK), .RN(n12565), .QN(
        n13945) );
  DFFR_X1 \REGISTERS_reg[66][25]  ( .D(n8434), .CK(CLK), .RN(n12543), .QN(
        n13946) );
  DFFR_X1 \REGISTERS_reg[66][24]  ( .D(n8435), .CK(CLK), .RN(n12460), .QN(
        n13947) );
  DFFR_X1 \REGISTERS_reg[66][23]  ( .D(n8436), .CK(CLK), .RN(n12631), .QN(
        n13948) );
  DFFR_X1 \REGISTERS_reg[66][22]  ( .D(n8437), .CK(CLK), .RN(n12521), .QN(
        n13949) );
  DFFR_X1 \REGISTERS_reg[66][21]  ( .D(n8438), .CK(CLK), .RN(n12528), .QN(
        n13950) );
  DFFR_X1 \REGISTERS_reg[66][20]  ( .D(n8439), .CK(CLK), .RN(n12503), .QN(
        n13951) );
  DFFR_X1 \REGISTERS_reg[66][19]  ( .D(n8440), .CK(CLK), .RN(n12594), .QN(
        n13952) );
  DFFR_X1 \REGISTERS_reg[66][18]  ( .D(n8441), .CK(CLK), .RN(n12445), .QN(
        n13953) );
  DFFR_X1 \REGISTERS_reg[66][17]  ( .D(n8442), .CK(CLK), .RN(n12453), .QN(
        n13954) );
  DFFR_X1 \REGISTERS_reg[66][16]  ( .D(n8443), .CK(CLK), .RN(n12459), .QN(
        n13955) );
  DFFR_X1 \REGISTERS_reg[66][15]  ( .D(n8444), .CK(CLK), .RN(n12638), .QN(
        n13956) );
  DFFR_X1 \REGISTERS_reg[66][14]  ( .D(n8445), .CK(CLK), .RN(n12466), .QN(
        n13957) );
  DFFR_X1 \REGISTERS_reg[66][13]  ( .D(n8446), .CK(CLK), .RN(n12474), .QN(
        n13958) );
  DFFR_X1 \REGISTERS_reg[66][12]  ( .D(n8447), .CK(CLK), .RN(n12481), .QN(
        n13959) );
  DFFR_X1 \REGISTERS_reg[66][11]  ( .D(n8448), .CK(CLK), .RN(n12572), .QN(
        n13960) );
  DFFR_X1 \REGISTERS_reg[66][10]  ( .D(n8449), .CK(CLK), .RN(n12550), .QN(
        n13961) );
  DFFR_X1 \REGISTERS_reg[66][9]  ( .D(n8450), .CK(CLK), .RN(n12558), .QN(
        n13962) );
  DFFR_X1 \REGISTERS_reg[66][8]  ( .D(n8451), .CK(CLK), .RN(n12536), .QN(
        n13963) );
  DFFR_X1 \REGISTERS_reg[66][7]  ( .D(n8452), .CK(CLK), .RN(n12646), .QN(
        n13964) );
  DFFR_X1 \REGISTERS_reg[66][6]  ( .D(n8453), .CK(CLK), .RN(n12602), .QN(
        n13965) );
  DFFR_X1 \REGISTERS_reg[66][5]  ( .D(n8454), .CK(CLK), .RN(n12488), .QN(
        n13966) );
  DFFR_X1 \REGISTERS_reg[66][4]  ( .D(n8455), .CK(CLK), .RN(n12496), .QN(
        n13967) );
  DFFR_X1 \REGISTERS_reg[66][3]  ( .D(n8456), .CK(CLK), .RN(n12580), .QN(
        n13968) );
  DFFR_X1 \REGISTERS_reg[66][2]  ( .D(n8457), .CK(CLK), .RN(n12510), .QN(
        n13969) );
  DFFR_X1 \REGISTERS_reg[66][1]  ( .D(n8458), .CK(CLK), .RN(n12438), .QN(
        n13970) );
  DFFR_X1 \REGISTERS_reg[66][0]  ( .D(n8459), .CK(CLK), .RN(n12653), .QN(
        n13971) );
  DFFR_X1 \REGISTERS_reg[67][31]  ( .D(n8460), .CK(CLK), .RN(n12660), .QN(
        n13972) );
  DFFR_X1 \REGISTERS_reg[67][30]  ( .D(n8461), .CK(CLK), .RN(n12624), .QN(
        n13973) );
  DFFR_X1 \REGISTERS_reg[67][29]  ( .D(n8462), .CK(CLK), .RN(n12609), .QN(
        n13974) );
  DFFR_X1 \REGISTERS_reg[67][28]  ( .D(n8463), .CK(CLK), .RN(n12616), .QN(
        n13975) );
  DFFR_X1 \REGISTERS_reg[67][27]  ( .D(n8464), .CK(CLK), .RN(n12587), .QN(
        n13976) );
  DFFR_X1 \REGISTERS_reg[67][26]  ( .D(n8465), .CK(CLK), .RN(n12565), .QN(
        n13977) );
  DFFR_X1 \REGISTERS_reg[67][25]  ( .D(n8466), .CK(CLK), .RN(n12543), .QN(
        n13978) );
  DFFR_X1 \REGISTERS_reg[67][24]  ( .D(n8467), .CK(CLK), .RN(n12459), .QN(
        n13979) );
  DFFR_X1 \REGISTERS_reg[67][23]  ( .D(n8468), .CK(CLK), .RN(n12631), .QN(
        n13980) );
  DFFR_X1 \REGISTERS_reg[67][22]  ( .D(n8469), .CK(CLK), .RN(n12521), .QN(
        n13981) );
  DFFR_X1 \REGISTERS_reg[67][21]  ( .D(n8470), .CK(CLK), .RN(n12528), .QN(
        n13982) );
  DFFR_X1 \REGISTERS_reg[67][20]  ( .D(n8471), .CK(CLK), .RN(n12503), .QN(
        n13983) );
  DFFR_X1 \REGISTERS_reg[67][19]  ( .D(n8472), .CK(CLK), .RN(n12594), .QN(
        n13984) );
  DFFR_X1 \REGISTERS_reg[67][18]  ( .D(n8473), .CK(CLK), .RN(n12445), .QN(
        n13985) );
  DFFR_X1 \REGISTERS_reg[67][17]  ( .D(n8474), .CK(CLK), .RN(n12453), .QN(
        n13986) );
  DFFR_X1 \REGISTERS_reg[67][16]  ( .D(n8475), .CK(CLK), .RN(n12459), .QN(
        n13987) );
  DFFR_X1 \REGISTERS_reg[67][15]  ( .D(n8476), .CK(CLK), .RN(n12638), .QN(
        n13988) );
  DFFR_X1 \REGISTERS_reg[67][14]  ( .D(n8477), .CK(CLK), .RN(n12466), .QN(
        n13989) );
  DFFR_X1 \REGISTERS_reg[67][13]  ( .D(n8478), .CK(CLK), .RN(n12474), .QN(
        n13990) );
  DFFR_X1 \REGISTERS_reg[67][12]  ( .D(n8479), .CK(CLK), .RN(n12481), .QN(
        n13991) );
  DFFR_X1 \REGISTERS_reg[67][11]  ( .D(n8480), .CK(CLK), .RN(n12572), .QN(
        n13992) );
  DFFR_X1 \REGISTERS_reg[67][10]  ( .D(n8481), .CK(CLK), .RN(n12550), .QN(
        n13993) );
  DFFR_X1 \REGISTERS_reg[67][9]  ( .D(n8482), .CK(CLK), .RN(n12558), .QN(
        n13994) );
  DFFR_X1 \REGISTERS_reg[67][8]  ( .D(n8483), .CK(CLK), .RN(n12536), .QN(
        n13995) );
  DFFR_X1 \REGISTERS_reg[67][7]  ( .D(n8484), .CK(CLK), .RN(n12646), .QN(
        n13996) );
  DFFR_X1 \REGISTERS_reg[67][6]  ( .D(n8485), .CK(CLK), .RN(n12602), .QN(
        n13997) );
  DFFR_X1 \REGISTERS_reg[67][5]  ( .D(n8486), .CK(CLK), .RN(n12488), .QN(
        n13998) );
  DFFR_X1 \REGISTERS_reg[67][4]  ( .D(n8487), .CK(CLK), .RN(n12496), .QN(
        n13999) );
  DFFR_X1 \REGISTERS_reg[67][3]  ( .D(n8488), .CK(CLK), .RN(n12580), .QN(
        n14000) );
  DFFR_X1 \REGISTERS_reg[67][2]  ( .D(n8489), .CK(CLK), .RN(n12510), .QN(
        n14001) );
  DFFR_X1 \REGISTERS_reg[67][1]  ( .D(n8490), .CK(CLK), .RN(n12438), .QN(
        n14002) );
  DFFR_X1 \REGISTERS_reg[67][0]  ( .D(n8491), .CK(CLK), .RN(n12653), .QN(
        n14003) );
  DFFR_X1 \REGISTERS_reg[68][31]  ( .D(n8492), .CK(CLK), .RN(n12661), .QN(n998) );
  DFFR_X1 \REGISTERS_reg[68][30]  ( .D(n8493), .CK(CLK), .RN(n12624), .QN(
        n14004) );
  DFFR_X1 \REGISTERS_reg[68][29]  ( .D(n8494), .CK(CLK), .RN(n12609), .QN(
        n14005) );
  DFFR_X1 \REGISTERS_reg[68][28]  ( .D(n8495), .CK(CLK), .RN(n12617), .QN(
        n14006) );
  DFFR_X1 \REGISTERS_reg[68][27]  ( .D(n8496), .CK(CLK), .RN(n12587), .QN(
        n14007) );
  DFFR_X1 \REGISTERS_reg[68][26]  ( .D(n8497), .CK(CLK), .RN(n12565), .QN(
        n14008) );
  DFFR_X1 \REGISTERS_reg[68][25]  ( .D(n8498), .CK(CLK), .RN(n12543), .QN(
        n14009) );
  DFFR_X1 \REGISTERS_reg[68][24]  ( .D(n8499), .CK(CLK), .RN(n12458), .QN(
        n14010) );
  DFFR_X1 \REGISTERS_reg[68][23]  ( .D(n8500), .CK(CLK), .RN(n12631), .QN(
        n14011) );
  DFFR_X1 \REGISTERS_reg[68][22]  ( .D(n8501), .CK(CLK), .RN(n12521), .QN(
        n14012) );
  DFFR_X1 \REGISTERS_reg[68][21]  ( .D(n8502), .CK(CLK), .RN(n12529), .QN(
        n14013) );
  DFFR_X1 \REGISTERS_reg[68][20]  ( .D(n8503), .CK(CLK), .RN(n12503), .QN(
        n14014) );
  DFFR_X1 \REGISTERS_reg[68][19]  ( .D(n8504), .CK(CLK), .RN(n12595), .QN(
        n14015) );
  DFFR_X1 \REGISTERS_reg[68][18]  ( .D(n8505), .CK(CLK), .RN(n12446), .QN(
        n14016) );
  DFFR_X1 \REGISTERS_reg[68][17]  ( .D(n8506), .CK(CLK), .RN(n12453), .QN(
        n14017) );
  DFFR_X1 \REGISTERS_reg[68][16]  ( .D(n8507), .CK(CLK), .RN(n12459), .QN(
        n14018) );
  DFFR_X1 \REGISTERS_reg[68][15]  ( .D(n8508), .CK(CLK), .RN(n12639), .QN(
        n14019) );
  DFFR_X1 \REGISTERS_reg[68][14]  ( .D(n8509), .CK(CLK), .RN(n12467), .QN(
        n14020) );
  DFFR_X1 \REGISTERS_reg[68][13]  ( .D(n8510), .CK(CLK), .RN(n12474), .QN(
        n14021) );
  DFFR_X1 \REGISTERS_reg[68][12]  ( .D(n8511), .CK(CLK), .RN(n12481), .QN(
        n14022) );
  DFFR_X1 \REGISTERS_reg[68][11]  ( .D(n8512), .CK(CLK), .RN(n12573), .QN(
        n14023) );
  DFFR_X1 \REGISTERS_reg[68][10]  ( .D(n8513), .CK(CLK), .RN(n12551), .QN(
        n14024) );
  DFFR_X1 \REGISTERS_reg[68][9]  ( .D(n8514), .CK(CLK), .RN(n12558), .QN(
        n14025) );
  DFFR_X1 \REGISTERS_reg[68][8]  ( .D(n8515), .CK(CLK), .RN(n12536), .QN(
        n14026) );
  DFFR_X1 \REGISTERS_reg[68][7]  ( .D(n8516), .CK(CLK), .RN(n12646), .QN(
        n14027) );
  DFFR_X1 \REGISTERS_reg[68][6]  ( .D(n8517), .CK(CLK), .RN(n12602), .QN(
        n14028) );
  DFFR_X1 \REGISTERS_reg[68][5]  ( .D(n8518), .CK(CLK), .RN(n12489), .QN(
        n14029) );
  DFFR_X1 \REGISTERS_reg[68][4]  ( .D(n8519), .CK(CLK), .RN(n12496), .QN(
        n14030) );
  DFFR_X1 \REGISTERS_reg[68][3]  ( .D(n8520), .CK(CLK), .RN(n12580), .QN(
        n14031) );
  DFFR_X1 \REGISTERS_reg[68][2]  ( .D(n8521), .CK(CLK), .RN(n12511), .QN(
        n14032) );
  DFFR_X1 \REGISTERS_reg[68][1]  ( .D(n8522), .CK(CLK), .RN(n12438), .QN(
        n14033) );
  DFFR_X1 \REGISTERS_reg[68][0]  ( .D(n8523), .CK(CLK), .RN(n12653), .QN(
        n14034) );
  DFFR_X1 \REGISTERS_reg[69][31]  ( .D(n8524), .CK(CLK), .RN(n12661), .QN(
        n14035) );
  DFFR_X1 \REGISTERS_reg[69][30]  ( .D(n8525), .CK(CLK), .RN(n12624), .QN(
        n14036) );
  DFFR_X1 \REGISTERS_reg[69][29]  ( .D(n8526), .CK(CLK), .RN(n12609), .QN(
        n14037) );
  DFFR_X1 \REGISTERS_reg[69][28]  ( .D(n8527), .CK(CLK), .RN(n12617), .QN(
        n14038) );
  DFFR_X1 \REGISTERS_reg[69][27]  ( .D(n8528), .CK(CLK), .RN(n12587), .QN(
        n14039) );
  DFFR_X1 \REGISTERS_reg[69][26]  ( .D(n8529), .CK(CLK), .RN(n12565), .QN(
        n14040) );
  DFFR_X1 \REGISTERS_reg[69][25]  ( .D(n8530), .CK(CLK), .RN(n12543), .QN(
        n14041) );
  DFFR_X1 \REGISTERS_reg[69][24]  ( .D(n8531), .CK(CLK), .RN(n12467), .QN(
        n14042) );
  DFFR_X1 \REGISTERS_reg[69][23]  ( .D(n8532), .CK(CLK), .RN(n12631), .QN(
        n14043) );
  DFFR_X1 \REGISTERS_reg[69][22]  ( .D(n8533), .CK(CLK), .RN(n12521), .QN(
        n14044) );
  DFFR_X1 \REGISTERS_reg[69][21]  ( .D(n8534), .CK(CLK), .RN(n12529), .QN(
        n14045) );
  DFFR_X1 \REGISTERS_reg[69][20]  ( .D(n8535), .CK(CLK), .RN(n12503), .QN(
        n14046) );
  DFFR_X1 \REGISTERS_reg[69][19]  ( .D(n8536), .CK(CLK), .RN(n12595), .QN(
        n14047) );
  DFFR_X1 \REGISTERS_reg[69][18]  ( .D(n8537), .CK(CLK), .RN(n12446), .QN(
        n14048) );
  DFFR_X1 \REGISTERS_reg[69][17]  ( .D(n8538), .CK(CLK), .RN(n12453), .QN(
        n14049) );
  DFFR_X1 \REGISTERS_reg[69][16]  ( .D(n8539), .CK(CLK), .RN(n12459), .QN(
        n14050) );
  DFFR_X1 \REGISTERS_reg[69][15]  ( .D(n8540), .CK(CLK), .RN(n12639), .QN(
        n14051) );
  DFFR_X1 \REGISTERS_reg[69][14]  ( .D(n8541), .CK(CLK), .RN(n12467), .QN(
        n14052) );
  DFFR_X1 \REGISTERS_reg[69][13]  ( .D(n8542), .CK(CLK), .RN(n12474), .QN(
        n14053) );
  DFFR_X1 \REGISTERS_reg[69][12]  ( .D(n8543), .CK(CLK), .RN(n12481), .QN(
        n14054) );
  DFFR_X1 \REGISTERS_reg[69][11]  ( .D(n8544), .CK(CLK), .RN(n12573), .QN(
        n14055) );
  DFFR_X1 \REGISTERS_reg[69][10]  ( .D(n8545), .CK(CLK), .RN(n12551), .QN(
        n14056) );
  DFFR_X1 \REGISTERS_reg[69][9]  ( .D(n8546), .CK(CLK), .RN(n12558), .QN(
        n14057) );
  DFFR_X1 \REGISTERS_reg[69][8]  ( .D(n8547), .CK(CLK), .RN(n12536), .QN(
        n14058) );
  DFFR_X1 \REGISTERS_reg[69][7]  ( .D(n8548), .CK(CLK), .RN(n12646), .QN(
        n14059) );
  DFFR_X1 \REGISTERS_reg[69][6]  ( .D(n8549), .CK(CLK), .RN(n12602), .QN(
        n14060) );
  DFFR_X1 \REGISTERS_reg[69][5]  ( .D(n8550), .CK(CLK), .RN(n12489), .QN(
        n14061) );
  DFFR_X1 \REGISTERS_reg[69][4]  ( .D(n8551), .CK(CLK), .RN(n12496), .QN(
        n14062) );
  DFFR_X1 \REGISTERS_reg[69][3]  ( .D(n8552), .CK(CLK), .RN(n12580), .QN(
        n14063) );
  DFFR_X1 \REGISTERS_reg[69][2]  ( .D(n8553), .CK(CLK), .RN(n12511), .QN(
        n14064) );
  DFFR_X1 \REGISTERS_reg[69][1]  ( .D(n8554), .CK(CLK), .RN(n12438), .QN(
        n14065) );
  DFFR_X1 \REGISTERS_reg[69][0]  ( .D(n8555), .CK(CLK), .RN(n12653), .QN(
        n14066) );
  DFFR_X1 \REGISTERS_reg[70][31]  ( .D(n8556), .CK(CLK), .RN(n12661), .QN(
        n14067) );
  DFFR_X1 \REGISTERS_reg[70][30]  ( .D(n8557), .CK(CLK), .RN(n12624), .QN(
        n14068) );
  DFFR_X1 \REGISTERS_reg[70][29]  ( .D(n8558), .CK(CLK), .RN(n12609), .QN(
        n14069) );
  DFFR_X1 \REGISTERS_reg[70][28]  ( .D(n8559), .CK(CLK), .RN(n12617), .QN(
        n14070) );
  DFFR_X1 \REGISTERS_reg[70][27]  ( .D(n8560), .CK(CLK), .RN(n12587), .QN(
        n14071) );
  DFFR_X1 \REGISTERS_reg[70][26]  ( .D(n8561), .CK(CLK), .RN(n12565), .QN(
        n14072) );
  DFFR_X1 \REGISTERS_reg[70][25]  ( .D(n8562), .CK(CLK), .RN(n12543), .QN(
        n14073) );
  DFFR_X1 \REGISTERS_reg[70][24]  ( .D(n8563), .CK(CLK), .RN(n12457), .QN(
        n14074) );
  DFFR_X1 \REGISTERS_reg[70][23]  ( .D(n8564), .CK(CLK), .RN(n12631), .QN(
        n14075) );
  DFFR_X1 \REGISTERS_reg[70][22]  ( .D(n8565), .CK(CLK), .RN(n12521), .QN(
        n14076) );
  DFFR_X1 \REGISTERS_reg[70][21]  ( .D(n8566), .CK(CLK), .RN(n12529), .QN(
        n14077) );
  DFFR_X1 \REGISTERS_reg[70][20]  ( .D(n8567), .CK(CLK), .RN(n12503), .QN(
        n14078) );
  DFFR_X1 \REGISTERS_reg[70][19]  ( .D(n8568), .CK(CLK), .RN(n12595), .QN(
        n14079) );
  DFFR_X1 \REGISTERS_reg[70][18]  ( .D(n8569), .CK(CLK), .RN(n12446), .QN(
        n14080) );
  DFFR_X1 \REGISTERS_reg[70][17]  ( .D(n8570), .CK(CLK), .RN(n12453), .QN(
        n14081) );
  DFFR_X1 \REGISTERS_reg[70][16]  ( .D(n8571), .CK(CLK), .RN(n12459), .QN(
        n14082) );
  DFFR_X1 \REGISTERS_reg[70][15]  ( .D(n8572), .CK(CLK), .RN(n12639), .QN(
        n14083) );
  DFFR_X1 \REGISTERS_reg[70][14]  ( .D(n8573), .CK(CLK), .RN(n12467), .QN(
        n14084) );
  DFFR_X1 \REGISTERS_reg[70][13]  ( .D(n8574), .CK(CLK), .RN(n12474), .QN(
        n14085) );
  DFFR_X1 \REGISTERS_reg[70][12]  ( .D(n8575), .CK(CLK), .RN(n12481), .QN(
        n14086) );
  DFFR_X1 \REGISTERS_reg[70][11]  ( .D(n8576), .CK(CLK), .RN(n12573), .QN(
        n14087) );
  DFFR_X1 \REGISTERS_reg[70][10]  ( .D(n8577), .CK(CLK), .RN(n12551), .QN(
        n14088) );
  DFFR_X1 \REGISTERS_reg[70][9]  ( .D(n8578), .CK(CLK), .RN(n12558), .QN(
        n14089) );
  DFFR_X1 \REGISTERS_reg[70][8]  ( .D(n8579), .CK(CLK), .RN(n12536), .QN(
        n14090) );
  DFFR_X1 \REGISTERS_reg[70][7]  ( .D(n8580), .CK(CLK), .RN(n12646), .QN(
        n14091) );
  DFFR_X1 \REGISTERS_reg[70][6]  ( .D(n8581), .CK(CLK), .RN(n12602), .QN(
        n14092) );
  DFFR_X1 \REGISTERS_reg[70][5]  ( .D(n8582), .CK(CLK), .RN(n12489), .QN(
        n14093) );
  DFFR_X1 \REGISTERS_reg[70][4]  ( .D(n8583), .CK(CLK), .RN(n12496), .QN(
        n14094) );
  DFFR_X1 \REGISTERS_reg[70][3]  ( .D(n8584), .CK(CLK), .RN(n12580), .QN(
        n14095) );
  DFFR_X1 \REGISTERS_reg[70][2]  ( .D(n8585), .CK(CLK), .RN(n12511), .QN(
        n14096) );
  DFFR_X1 \REGISTERS_reg[70][1]  ( .D(n8586), .CK(CLK), .RN(n12438), .QN(
        n14097) );
  DFFR_X1 \REGISTERS_reg[70][0]  ( .D(n8587), .CK(CLK), .RN(n12653), .QN(
        n14098) );
  DFFR_X1 \REGISTERS_reg[71][31]  ( .D(n8588), .CK(CLK), .RN(n12661), .QN(n997) );
  DFFR_X1 \REGISTERS_reg[71][30]  ( .D(n8589), .CK(CLK), .RN(n12624), .QN(
        n14099) );
  DFFR_X1 \REGISTERS_reg[71][29]  ( .D(n8590), .CK(CLK), .RN(n12609), .QN(
        n14100) );
  DFFR_X1 \REGISTERS_reg[71][28]  ( .D(n8591), .CK(CLK), .RN(n12617), .QN(
        n14101) );
  DFFR_X1 \REGISTERS_reg[71][27]  ( .D(n8592), .CK(CLK), .RN(n12587), .QN(
        n14102) );
  DFFR_X1 \REGISTERS_reg[71][26]  ( .D(n8593), .CK(CLK), .RN(n12565), .QN(
        n14103) );
  DFFR_X1 \REGISTERS_reg[71][25]  ( .D(n8594), .CK(CLK), .RN(n12543), .QN(
        n14104) );
  DFFR_X1 \REGISTERS_reg[71][24]  ( .D(n8595), .CK(CLK), .RN(n12456), .QN(
        n14105) );
  DFFR_X1 \REGISTERS_reg[71][23]  ( .D(n8596), .CK(CLK), .RN(n12631), .QN(
        n14106) );
  DFFR_X1 \REGISTERS_reg[71][22]  ( .D(n8597), .CK(CLK), .RN(n12521), .QN(
        n14107) );
  DFFR_X1 \REGISTERS_reg[71][21]  ( .D(n8598), .CK(CLK), .RN(n12529), .QN(
        n14108) );
  DFFR_X1 \REGISTERS_reg[71][20]  ( .D(n8599), .CK(CLK), .RN(n12503), .QN(
        n14109) );
  DFFR_X1 \REGISTERS_reg[71][19]  ( .D(n8600), .CK(CLK), .RN(n12595), .QN(
        n14110) );
  DFFR_X1 \REGISTERS_reg[71][18]  ( .D(n8601), .CK(CLK), .RN(n12446), .QN(
        n14111) );
  DFFR_X1 \REGISTERS_reg[71][17]  ( .D(n8602), .CK(CLK), .RN(n12453), .QN(
        n14112) );
  DFFR_X1 \REGISTERS_reg[71][16]  ( .D(n8603), .CK(CLK), .RN(n12459), .QN(
        n14113) );
  DFFR_X1 \REGISTERS_reg[71][15]  ( .D(n8604), .CK(CLK), .RN(n12639), .QN(
        n14114) );
  DFFR_X1 \REGISTERS_reg[71][14]  ( .D(n8605), .CK(CLK), .RN(n12467), .QN(
        n14115) );
  DFFR_X1 \REGISTERS_reg[71][13]  ( .D(n8606), .CK(CLK), .RN(n12474), .QN(
        n14116) );
  DFFR_X1 \REGISTERS_reg[71][12]  ( .D(n8607), .CK(CLK), .RN(n12481), .QN(
        n14117) );
  DFFR_X1 \REGISTERS_reg[71][11]  ( .D(n8608), .CK(CLK), .RN(n12573), .QN(
        n14118) );
  DFFR_X1 \REGISTERS_reg[71][10]  ( .D(n8609), .CK(CLK), .RN(n12551), .QN(
        n14119) );
  DFFR_X1 \REGISTERS_reg[71][9]  ( .D(n8610), .CK(CLK), .RN(n12558), .QN(
        n14120) );
  DFFR_X1 \REGISTERS_reg[71][8]  ( .D(n8611), .CK(CLK), .RN(n12536), .QN(
        n14121) );
  DFFR_X1 \REGISTERS_reg[71][7]  ( .D(n8612), .CK(CLK), .RN(n12646), .QN(
        n14122) );
  DFFR_X1 \REGISTERS_reg[71][6]  ( .D(n8613), .CK(CLK), .RN(n12602), .QN(
        n14123) );
  DFFR_X1 \REGISTERS_reg[71][5]  ( .D(n8614), .CK(CLK), .RN(n12489), .QN(
        n14124) );
  DFFR_X1 \REGISTERS_reg[71][4]  ( .D(n8615), .CK(CLK), .RN(n12496), .QN(
        n14125) );
  DFFR_X1 \REGISTERS_reg[71][3]  ( .D(n8616), .CK(CLK), .RN(n12580), .QN(
        n14126) );
  DFFR_X1 \REGISTERS_reg[71][2]  ( .D(n8617), .CK(CLK), .RN(n12511), .QN(
        n14127) );
  DFFR_X1 \REGISTERS_reg[71][1]  ( .D(n8618), .CK(CLK), .RN(n12438), .QN(
        n14128) );
  DFFR_X1 \REGISTERS_reg[71][0]  ( .D(n8619), .CK(CLK), .RN(n12653), .QN(
        n14129) );
  DFFR_X1 \REGISTERS_reg[72][31]  ( .D(n8620), .CK(CLK), .RN(n12661), .QN(
        n14130) );
  DFFR_X1 \REGISTERS_reg[72][30]  ( .D(n8621), .CK(CLK), .RN(n12624), .QN(
        n14131) );
  DFFR_X1 \REGISTERS_reg[72][29]  ( .D(n8622), .CK(CLK), .RN(n12610), .QN(
        n14132) );
  DFFR_X1 \REGISTERS_reg[72][28]  ( .D(n8623), .CK(CLK), .RN(n12617), .QN(
        n14133) );
  DFFR_X1 \REGISTERS_reg[72][27]  ( .D(n8624), .CK(CLK), .RN(n12588), .QN(
        n14134) );
  DFFR_X1 \REGISTERS_reg[72][26]  ( .D(n8625), .CK(CLK), .RN(n12566), .QN(
        n14135) );
  DFFR_X1 \REGISTERS_reg[72][25]  ( .D(n8626), .CK(CLK), .RN(n12544), .QN(
        n14136) );
  DFFR_X1 \REGISTERS_reg[72][24]  ( .D(n8627), .CK(CLK), .RN(n12466), .QN(
        n14137) );
  DFFR_X1 \REGISTERS_reg[72][23]  ( .D(n8628), .CK(CLK), .RN(n12632), .QN(
        n14138) );
  DFFR_X1 \REGISTERS_reg[72][22]  ( .D(n8629), .CK(CLK), .RN(n12522), .QN(
        n14139) );
  DFFR_X1 \REGISTERS_reg[72][21]  ( .D(n8630), .CK(CLK), .RN(n12529), .QN(
        n14140) );
  DFFR_X1 \REGISTERS_reg[72][20]  ( .D(n8631), .CK(CLK), .RN(n12504), .QN(
        n14141) );
  DFFR_X1 \REGISTERS_reg[72][19]  ( .D(n8632), .CK(CLK), .RN(n12595), .QN(
        n14142) );
  DFFR_X1 \REGISTERS_reg[72][18]  ( .D(n8633), .CK(CLK), .RN(n12446), .QN(
        n14143) );
  DFFR_X1 \REGISTERS_reg[72][17]  ( .D(n8634), .CK(CLK), .RN(n12453), .QN(
        n14144) );
  DFFR_X1 \REGISTERS_reg[72][16]  ( .D(n8635), .CK(CLK), .RN(n12460), .QN(
        n14145) );
  DFFR_X1 \REGISTERS_reg[72][15]  ( .D(n8636), .CK(CLK), .RN(n12639), .QN(
        n14146) );
  DFFR_X1 \REGISTERS_reg[72][14]  ( .D(n8637), .CK(CLK), .RN(n12467), .QN(
        n14147) );
  DFFR_X1 \REGISTERS_reg[72][13]  ( .D(n8638), .CK(CLK), .RN(n12474), .QN(
        n14148) );
  DFFR_X1 \REGISTERS_reg[72][12]  ( .D(n8639), .CK(CLK), .RN(n12482), .QN(
        n14149) );
  DFFR_X1 \REGISTERS_reg[72][11]  ( .D(n8640), .CK(CLK), .RN(n12573), .QN(
        n14150) );
  DFFR_X1 \REGISTERS_reg[72][10]  ( .D(n8641), .CK(CLK), .RN(n12551), .QN(
        n14151) );
  DFFR_X1 \REGISTERS_reg[72][9]  ( .D(n8642), .CK(CLK), .RN(n12558), .QN(
        n14152) );
  DFFR_X1 \REGISTERS_reg[72][8]  ( .D(n8643), .CK(CLK), .RN(n12536), .QN(
        n14153) );
  DFFR_X1 \REGISTERS_reg[72][7]  ( .D(n8644), .CK(CLK), .RN(n12646), .QN(
        n14154) );
  DFFR_X1 \REGISTERS_reg[72][6]  ( .D(n8645), .CK(CLK), .RN(n12602), .QN(
        n14155) );
  DFFR_X1 \REGISTERS_reg[72][5]  ( .D(n8646), .CK(CLK), .RN(n12489), .QN(
        n14156) );
  DFFR_X1 \REGISTERS_reg[72][4]  ( .D(n8647), .CK(CLK), .RN(n12496), .QN(
        n14157) );
  DFFR_X1 \REGISTERS_reg[72][3]  ( .D(n8648), .CK(CLK), .RN(n12580), .QN(
        n14158) );
  DFFR_X1 \REGISTERS_reg[72][2]  ( .D(n8649), .CK(CLK), .RN(n12511), .QN(
        n14159) );
  DFFR_X1 \REGISTERS_reg[72][1]  ( .D(n8650), .CK(CLK), .RN(n12439), .QN(
        n14160) );
  DFFR_X1 \REGISTERS_reg[72][0]  ( .D(n8651), .CK(CLK), .RN(n12654), .QN(
        n14161) );
  DFFR_X1 \REGISTERS_reg[73][31]  ( .D(n8652), .CK(CLK), .RN(n12661), .QN(
        n14162) );
  DFFR_X1 \REGISTERS_reg[73][30]  ( .D(n8653), .CK(CLK), .RN(n12624), .QN(
        n14163) );
  DFFR_X1 \REGISTERS_reg[73][29]  ( .D(n8654), .CK(CLK), .RN(n12610), .QN(
        n14164) );
  DFFR_X1 \REGISTERS_reg[73][28]  ( .D(n8655), .CK(CLK), .RN(n12617), .QN(
        n14165) );
  DFFR_X1 \REGISTERS_reg[73][27]  ( .D(n8656), .CK(CLK), .RN(n12588), .QN(
        n14166) );
  DFFR_X1 \REGISTERS_reg[73][26]  ( .D(n8657), .CK(CLK), .RN(n12566), .QN(
        n14167) );
  DFFR_X1 \REGISTERS_reg[73][25]  ( .D(n8658), .CK(CLK), .RN(n12544), .QN(
        n14168) );
  DFFR_X1 \REGISTERS_reg[73][24]  ( .D(n8659), .CK(CLK), .RN(n12455), .QN(
        n14169) );
  DFFR_X1 \REGISTERS_reg[73][23]  ( .D(n8660), .CK(CLK), .RN(n12632), .QN(
        n14170) );
  DFFR_X1 \REGISTERS_reg[73][22]  ( .D(n8661), .CK(CLK), .RN(n12522), .QN(
        n14171) );
  DFFR_X1 \REGISTERS_reg[73][21]  ( .D(n8662), .CK(CLK), .RN(n12529), .QN(
        n14172) );
  DFFR_X1 \REGISTERS_reg[73][20]  ( .D(n8663), .CK(CLK), .RN(n12504), .QN(
        n14173) );
  DFFR_X1 \REGISTERS_reg[73][19]  ( .D(n8664), .CK(CLK), .RN(n12595), .QN(
        n14174) );
  DFFR_X1 \REGISTERS_reg[73][18]  ( .D(n8665), .CK(CLK), .RN(n12446), .QN(
        n14175) );
  DFFR_X1 \REGISTERS_reg[73][17]  ( .D(n8666), .CK(CLK), .RN(n12453), .QN(
        n14176) );
  DFFR_X1 \REGISTERS_reg[73][16]  ( .D(n8667), .CK(CLK), .RN(n12460), .QN(
        n14177) );
  DFFR_X1 \REGISTERS_reg[73][15]  ( .D(n8668), .CK(CLK), .RN(n12639), .QN(
        n14178) );
  DFFR_X1 \REGISTERS_reg[73][14]  ( .D(n8669), .CK(CLK), .RN(n12467), .QN(
        n14179) );
  DFFR_X1 \REGISTERS_reg[73][13]  ( .D(n8670), .CK(CLK), .RN(n12474), .QN(
        n14180) );
  DFFR_X1 \REGISTERS_reg[73][12]  ( .D(n8671), .CK(CLK), .RN(n12482), .QN(
        n14181) );
  DFFR_X1 \REGISTERS_reg[73][11]  ( .D(n8672), .CK(CLK), .RN(n12573), .QN(
        n14182) );
  DFFR_X1 \REGISTERS_reg[73][10]  ( .D(n8673), .CK(CLK), .RN(n12551), .QN(
        n14183) );
  DFFR_X1 \REGISTERS_reg[73][9]  ( .D(n8674), .CK(CLK), .RN(n12558), .QN(
        n14184) );
  DFFR_X1 \REGISTERS_reg[73][8]  ( .D(n8675), .CK(CLK), .RN(n12536), .QN(
        n14185) );
  DFFR_X1 \REGISTERS_reg[73][7]  ( .D(n8676), .CK(CLK), .RN(n12646), .QN(
        n14186) );
  DFFR_X1 \REGISTERS_reg[73][6]  ( .D(n8677), .CK(CLK), .RN(n12602), .QN(
        n14187) );
  DFFR_X1 \REGISTERS_reg[73][5]  ( .D(n8678), .CK(CLK), .RN(n12489), .QN(
        n14188) );
  DFFR_X1 \REGISTERS_reg[73][4]  ( .D(n8679), .CK(CLK), .RN(n12496), .QN(
        n14189) );
  DFFR_X1 \REGISTERS_reg[73][3]  ( .D(n8680), .CK(CLK), .RN(n12580), .QN(
        n14190) );
  DFFR_X1 \REGISTERS_reg[73][2]  ( .D(n8681), .CK(CLK), .RN(n12511), .QN(
        n14191) );
  DFFR_X1 \REGISTERS_reg[73][1]  ( .D(n8682), .CK(CLK), .RN(n12439), .QN(
        n14192) );
  DFFR_X1 \REGISTERS_reg[73][0]  ( .D(n8683), .CK(CLK), .RN(n12654), .QN(
        n14193) );
  DFFR_X1 \REGISTERS_reg[74][31]  ( .D(n8684), .CK(CLK), .RN(n12661), .QN(n996) );
  DFFR_X1 \REGISTERS_reg[74][30]  ( .D(n8685), .CK(CLK), .RN(n12624), .QN(
        n14194) );
  DFFR_X1 \REGISTERS_reg[74][29]  ( .D(n8686), .CK(CLK), .RN(n12610), .QN(
        n14195) );
  DFFR_X1 \REGISTERS_reg[74][28]  ( .D(n8687), .CK(CLK), .RN(n12617), .QN(
        n14196) );
  DFFR_X1 \REGISTERS_reg[74][27]  ( .D(n8688), .CK(CLK), .RN(n12588), .QN(
        n14197) );
  DFFR_X1 \REGISTERS_reg[74][26]  ( .D(n8689), .CK(CLK), .RN(n12566), .QN(
        n14198) );
  DFFR_X1 \REGISTERS_reg[74][25]  ( .D(n8690), .CK(CLK), .RN(n12544), .QN(
        n14199) );
  DFFR_X1 \REGISTERS_reg[74][24]  ( .D(n8691), .CK(CLK), .RN(n12468), .QN(
        n14200) );
  DFFR_X1 \REGISTERS_reg[74][23]  ( .D(n8692), .CK(CLK), .RN(n12632), .QN(
        n14201) );
  DFFR_X1 \REGISTERS_reg[74][22]  ( .D(n8693), .CK(CLK), .RN(n12522), .QN(
        n14202) );
  DFFR_X1 \REGISTERS_reg[74][21]  ( .D(n8694), .CK(CLK), .RN(n12529), .QN(
        n14203) );
  DFFR_X1 \REGISTERS_reg[74][20]  ( .D(n8695), .CK(CLK), .RN(n12504), .QN(
        n14204) );
  DFFR_X1 \REGISTERS_reg[74][19]  ( .D(n8696), .CK(CLK), .RN(n12595), .QN(
        n14205) );
  DFFR_X1 \REGISTERS_reg[74][18]  ( .D(n8697), .CK(CLK), .RN(n12446), .QN(
        n14206) );
  DFFR_X1 \REGISTERS_reg[74][17]  ( .D(n8698), .CK(CLK), .RN(n12453), .QN(
        n14207) );
  DFFR_X1 \REGISTERS_reg[74][16]  ( .D(n8699), .CK(CLK), .RN(n12460), .QN(
        n14208) );
  DFFR_X1 \REGISTERS_reg[74][15]  ( .D(n8700), .CK(CLK), .RN(n12639), .QN(
        n14209) );
  DFFR_X1 \REGISTERS_reg[74][14]  ( .D(n8701), .CK(CLK), .RN(n12467), .QN(
        n14210) );
  DFFR_X1 \REGISTERS_reg[74][13]  ( .D(n8702), .CK(CLK), .RN(n12474), .QN(
        n14211) );
  DFFR_X1 \REGISTERS_reg[74][12]  ( .D(n8703), .CK(CLK), .RN(n12482), .QN(
        n14212) );
  DFFR_X1 \REGISTERS_reg[74][11]  ( .D(n8704), .CK(CLK), .RN(n12573), .QN(
        n14213) );
  DFFR_X1 \REGISTERS_reg[74][10]  ( .D(n8705), .CK(CLK), .RN(n12551), .QN(
        n14214) );
  DFFR_X1 \REGISTERS_reg[74][9]  ( .D(n8706), .CK(CLK), .RN(n12558), .QN(
        n14215) );
  DFFR_X1 \REGISTERS_reg[74][8]  ( .D(n8707), .CK(CLK), .RN(n12536), .QN(
        n14216) );
  DFFR_X1 \REGISTERS_reg[74][7]  ( .D(n8708), .CK(CLK), .RN(n12646), .QN(
        n14217) );
  DFFR_X1 \REGISTERS_reg[74][6]  ( .D(n8709), .CK(CLK), .RN(n12602), .QN(
        n14218) );
  DFFR_X1 \REGISTERS_reg[74][5]  ( .D(n8710), .CK(CLK), .RN(n12489), .QN(
        n14219) );
  DFFR_X1 \REGISTERS_reg[74][4]  ( .D(n8711), .CK(CLK), .RN(n12496), .QN(
        n14220) );
  DFFR_X1 \REGISTERS_reg[74][3]  ( .D(n8712), .CK(CLK), .RN(n12580), .QN(
        n14221) );
  DFFR_X1 \REGISTERS_reg[74][2]  ( .D(n8713), .CK(CLK), .RN(n12511), .QN(
        n14222) );
  DFFR_X1 \REGISTERS_reg[74][1]  ( .D(n8714), .CK(CLK), .RN(n12439), .QN(
        n14223) );
  DFFR_X1 \REGISTERS_reg[74][0]  ( .D(n8715), .CK(CLK), .RN(n12654), .QN(
        n14224) );
  DFFR_X1 \REGISTERS_reg[75][31]  ( .D(n8716), .CK(CLK), .RN(n12661), .QN(n868) );
  DFFR_X1 \REGISTERS_reg[75][30]  ( .D(n8717), .CK(CLK), .RN(n12624), .QN(n872) );
  DFFR_X1 \REGISTERS_reg[75][29]  ( .D(n8718), .CK(CLK), .RN(n12610), .QN(n876) );
  DFFR_X1 \REGISTERS_reg[75][28]  ( .D(n8719), .CK(CLK), .RN(n12617), .QN(n880) );
  DFFR_X1 \REGISTERS_reg[75][27]  ( .D(n8720), .CK(CLK), .RN(n12588), .QN(n884) );
  DFFR_X1 \REGISTERS_reg[75][26]  ( .D(n8721), .CK(CLK), .RN(n12566), .QN(n888) );
  DFFR_X1 \REGISTERS_reg[75][25]  ( .D(n8722), .CK(CLK), .RN(n12544), .QN(n892) );
  DFFR_X1 \REGISTERS_reg[75][24]  ( .D(n8723), .CK(CLK), .RN(n12465), .QN(n896) );
  DFFR_X1 \REGISTERS_reg[75][23]  ( .D(n8724), .CK(CLK), .RN(n12632), .QN(n900) );
  DFFR_X1 \REGISTERS_reg[75][22]  ( .D(n8725), .CK(CLK), .RN(n12522), .QN(n904) );
  DFFR_X1 \REGISTERS_reg[75][21]  ( .D(n8726), .CK(CLK), .RN(n12529), .QN(n908) );
  DFFR_X1 \REGISTERS_reg[75][20]  ( .D(n8727), .CK(CLK), .RN(n12504), .QN(n912) );
  DFFR_X1 \REGISTERS_reg[75][19]  ( .D(n8728), .CK(CLK), .RN(n12595), .QN(n916) );
  DFFR_X1 \REGISTERS_reg[75][18]  ( .D(n8729), .CK(CLK), .RN(n12446), .QN(n920) );
  DFFR_X1 \REGISTERS_reg[75][17]  ( .D(n8730), .CK(CLK), .RN(n12453), .QN(n924) );
  DFFR_X1 \REGISTERS_reg[75][16]  ( .D(n8731), .CK(CLK), .RN(n12460), .QN(n928) );
  DFFR_X1 \REGISTERS_reg[75][15]  ( .D(n8732), .CK(CLK), .RN(n12639), .QN(n932) );
  DFFR_X1 \REGISTERS_reg[75][14]  ( .D(n8733), .CK(CLK), .RN(n12467), .QN(n936) );
  DFFR_X1 \REGISTERS_reg[75][13]  ( .D(n8734), .CK(CLK), .RN(n12474), .QN(n940) );
  DFFR_X1 \REGISTERS_reg[75][12]  ( .D(n8735), .CK(CLK), .RN(n12482), .QN(n944) );
  DFFR_X1 \REGISTERS_reg[75][11]  ( .D(n8736), .CK(CLK), .RN(n12573), .QN(n948) );
  DFFR_X1 \REGISTERS_reg[75][10]  ( .D(n8737), .CK(CLK), .RN(n12551), .QN(n952) );
  DFFR_X1 \REGISTERS_reg[75][9]  ( .D(n8738), .CK(CLK), .RN(n12558), .QN(n956)
         );
  DFFR_X1 \REGISTERS_reg[75][8]  ( .D(n8739), .CK(CLK), .RN(n12536), .QN(n960)
         );
  DFFR_X1 \REGISTERS_reg[75][7]  ( .D(n8740), .CK(CLK), .RN(n12646), .QN(n964)
         );
  DFFR_X1 \REGISTERS_reg[75][6]  ( .D(n8741), .CK(CLK), .RN(n12602), .QN(n968)
         );
  DFFR_X1 \REGISTERS_reg[75][5]  ( .D(n8742), .CK(CLK), .RN(n12489), .QN(n972)
         );
  DFFR_X1 \REGISTERS_reg[75][4]  ( .D(n8743), .CK(CLK), .RN(n12496), .QN(n976)
         );
  DFFR_X1 \REGISTERS_reg[75][3]  ( .D(n8744), .CK(CLK), .RN(n12580), .QN(n980)
         );
  DFFR_X1 \REGISTERS_reg[75][2]  ( .D(n8745), .CK(CLK), .RN(n12511), .QN(n984)
         );
  DFFR_X1 \REGISTERS_reg[75][1]  ( .D(n8746), .CK(CLK), .RN(n12439), .QN(n988)
         );
  DFFR_X1 \REGISTERS_reg[75][0]  ( .D(n8747), .CK(CLK), .RN(n12654), .QN(n992)
         );
  DFFR_X1 \REGISTERS_reg[76][31]  ( .D(n8748), .CK(CLK), .RN(n12661), .QN(
        n14225) );
  DFFR_X1 \REGISTERS_reg[76][30]  ( .D(n8749), .CK(CLK), .RN(n12625), .QN(
        n14226) );
  DFFR_X1 \REGISTERS_reg[76][29]  ( .D(n8750), .CK(CLK), .RN(n12610), .QN(
        n14227) );
  DFFR_X1 \REGISTERS_reg[76][28]  ( .D(n8751), .CK(CLK), .RN(n12617), .QN(
        n14228) );
  DFFR_X1 \REGISTERS_reg[76][27]  ( .D(n8752), .CK(CLK), .RN(n12588), .QN(
        n14229) );
  DFFR_X1 \REGISTERS_reg[76][26]  ( .D(n8753), .CK(CLK), .RN(n12566), .QN(
        n14230) );
  DFFR_X1 \REGISTERS_reg[76][25]  ( .D(n8754), .CK(CLK), .RN(n12544), .QN(
        n14231) );
  DFFR_X1 \REGISTERS_reg[76][24]  ( .D(n8755), .CK(CLK), .RN(n12508), .QN(
        n14232) );
  DFFR_X1 \REGISTERS_reg[76][23]  ( .D(n8756), .CK(CLK), .RN(n12632), .QN(
        n14233) );
  DFFR_X1 \REGISTERS_reg[76][22]  ( .D(n8757), .CK(CLK), .RN(n12522), .QN(
        n14234) );
  DFFR_X1 \REGISTERS_reg[76][21]  ( .D(n8758), .CK(CLK), .RN(n12529), .QN(
        n14235) );
  DFFR_X1 \REGISTERS_reg[76][20]  ( .D(n8759), .CK(CLK), .RN(n12504), .QN(
        n14236) );
  DFFR_X1 \REGISTERS_reg[76][19]  ( .D(n8760), .CK(CLK), .RN(n12595), .QN(
        n14237) );
  DFFR_X1 \REGISTERS_reg[76][18]  ( .D(n8761), .CK(CLK), .RN(n12446), .QN(
        n14238) );
  DFFR_X1 \REGISTERS_reg[76][17]  ( .D(n8762), .CK(CLK), .RN(n12454), .QN(
        n14239) );
  DFFR_X1 \REGISTERS_reg[76][16]  ( .D(n8763), .CK(CLK), .RN(n12460), .QN(
        n14240) );
  DFFR_X1 \REGISTERS_reg[76][15]  ( .D(n8764), .CK(CLK), .RN(n12639), .QN(
        n14241) );
  DFFR_X1 \REGISTERS_reg[76][14]  ( .D(n8765), .CK(CLK), .RN(n12467), .QN(
        n14242) );
  DFFR_X1 \REGISTERS_reg[76][13]  ( .D(n8766), .CK(CLK), .RN(n12475), .QN(
        n14243) );
  DFFR_X1 \REGISTERS_reg[76][12]  ( .D(n8767), .CK(CLK), .RN(n12482), .QN(
        n14244) );
  DFFR_X1 \REGISTERS_reg[76][11]  ( .D(n8768), .CK(CLK), .RN(n12573), .QN(
        n14245) );
  DFFR_X1 \REGISTERS_reg[76][10]  ( .D(n8769), .CK(CLK), .RN(n12551), .QN(
        n14246) );
  DFFR_X1 \REGISTERS_reg[76][9]  ( .D(n8770), .CK(CLK), .RN(n12559), .QN(
        n14247) );
  DFFR_X1 \REGISTERS_reg[76][8]  ( .D(n8771), .CK(CLK), .RN(n12537), .QN(
        n14248) );
  DFFR_X1 \REGISTERS_reg[76][7]  ( .D(n8772), .CK(CLK), .RN(n12647), .QN(
        n14249) );
  DFFR_X1 \REGISTERS_reg[76][6]  ( .D(n8773), .CK(CLK), .RN(n12603), .QN(
        n14250) );
  DFFR_X1 \REGISTERS_reg[76][5]  ( .D(n8774), .CK(CLK), .RN(n12489), .QN(
        n14251) );
  DFFR_X1 \REGISTERS_reg[76][4]  ( .D(n8775), .CK(CLK), .RN(n12497), .QN(
        n14252) );
  DFFR_X1 \REGISTERS_reg[76][3]  ( .D(n8776), .CK(CLK), .RN(n12581), .QN(
        n14253) );
  DFFR_X1 \REGISTERS_reg[76][2]  ( .D(n8777), .CK(CLK), .RN(n12511), .QN(
        n14254) );
  DFFR_X1 \REGISTERS_reg[76][1]  ( .D(n8778), .CK(CLK), .RN(n12439), .QN(
        n14255) );
  DFFR_X1 \REGISTERS_reg[76][0]  ( .D(n8779), .CK(CLK), .RN(n12654), .QN(
        n14256) );
  DFFR_X1 \REGISTERS_reg[78][31]  ( .D(n8812), .CK(CLK), .RN(n12661), .QN(
        n5712) );
  DFFR_X1 \REGISTERS_reg[78][30]  ( .D(n8813), .CK(CLK), .RN(n12625), .QN(
        n5744) );
  DFFR_X1 \REGISTERS_reg[78][29]  ( .D(n8814), .CK(CLK), .RN(n12610), .QN(
        n5776) );
  DFFR_X1 \REGISTERS_reg[78][28]  ( .D(n8815), .CK(CLK), .RN(n12617), .QN(
        n5808) );
  DFFR_X1 \REGISTERS_reg[78][27]  ( .D(n8816), .CK(CLK), .RN(n12588), .QN(
        n5840) );
  DFFR_X1 \REGISTERS_reg[78][26]  ( .D(n8817), .CK(CLK), .RN(n12566), .QN(
        n5872) );
  DFFR_X1 \REGISTERS_reg[78][25]  ( .D(n8818), .CK(CLK), .RN(n12544), .QN(
        n5904) );
  DFFR_X1 \REGISTERS_reg[78][24]  ( .D(n8819), .CK(CLK), .RN(n12507), .QN(
        n5936) );
  DFFR_X1 \REGISTERS_reg[78][23]  ( .D(n8820), .CK(CLK), .RN(n12632), .QN(
        n6000) );
  DFFR_X1 \REGISTERS_reg[78][22]  ( .D(n8821), .CK(CLK), .RN(n12522), .QN(
        n9135) );
  DFFR_X1 \REGISTERS_reg[78][21]  ( .D(n8822), .CK(CLK), .RN(n12529), .QN(
        n9167) );
  DFFR_X1 \REGISTERS_reg[78][20]  ( .D(n8823), .CK(CLK), .RN(n12504), .QN(
        n9199) );
  DFFR_X1 \REGISTERS_reg[78][19]  ( .D(n8824), .CK(CLK), .RN(n12595), .QN(
        n9263) );
  DFFR_X1 \REGISTERS_reg[78][18]  ( .D(n8825), .CK(CLK), .RN(n12446), .QN(
        n9597) );
  DFFR_X1 \REGISTERS_reg[78][17]  ( .D(n8826), .CK(CLK), .RN(n12454), .QN(
        n9629) );
  DFFR_X1 \REGISTERS_reg[78][16]  ( .D(n8827), .CK(CLK), .RN(n12460), .QN(
        n9661) );
  DFFR_X1 \REGISTERS_reg[78][15]  ( .D(n8828), .CK(CLK), .RN(n12639), .QN(
        n10023) );
  DFFR_X1 \REGISTERS_reg[78][14]  ( .D(n8829), .CK(CLK), .RN(n12467), .QN(
        n10055) );
  DFFR_X1 \REGISTERS_reg[78][13]  ( .D(n8830), .CK(CLK), .RN(n12475), .QN(
        n10087) );
  DFFR_X1 \REGISTERS_reg[78][12]  ( .D(n8831), .CK(CLK), .RN(n12482), .QN(
        n10119) );
  DFFR_X1 \REGISTERS_reg[78][11]  ( .D(n8832), .CK(CLK), .RN(n12573), .QN(
        n10151) );
  DFFR_X1 \REGISTERS_reg[78][10]  ( .D(n8833), .CK(CLK), .RN(n12551), .QN(
        n10183) );
  DFFR_X1 \REGISTERS_reg[78][9]  ( .D(n8834), .CK(CLK), .RN(n12559), .QN(
        n10217) );
  DFFR_X1 \REGISTERS_reg[78][8]  ( .D(n8835), .CK(CLK), .RN(n12537), .QN(
        n10249) );
  DFFR_X1 \REGISTERS_reg[78][7]  ( .D(n8836), .CK(CLK), .RN(n12647), .QN(
        n10281) );
  DFFR_X1 \REGISTERS_reg[78][6]  ( .D(n8837), .CK(CLK), .RN(n12603), .QN(
        n10316) );
  DFFR_X1 \REGISTERS_reg[78][5]  ( .D(n8838), .CK(CLK), .RN(n12489), .QN(
        n10348) );
  DFFR_X1 \REGISTERS_reg[78][4]  ( .D(n8839), .CK(CLK), .RN(n12497), .QN(
        n10380) );
  DFFR_X1 \REGISTERS_reg[78][3]  ( .D(n8840), .CK(CLK), .RN(n12581), .QN(
        n10415) );
  DFFR_X1 \REGISTERS_reg[78][2]  ( .D(n8841), .CK(CLK), .RN(n12511), .QN(
        n10447) );
  DFFR_X1 \REGISTERS_reg[78][1]  ( .D(n8842), .CK(CLK), .RN(n12439), .QN(
        n10479) );
  DFFR_X1 \REGISTERS_reg[78][0]  ( .D(n8843), .CK(CLK), .RN(n12654), .QN(
        n10511) );
  DFFR_X1 \REGISTERS_reg[79][31]  ( .D(n8844), .CK(CLK), .RN(n12661), .QN(
        n5710) );
  DFFR_X1 \REGISTERS_reg[79][30]  ( .D(n8845), .CK(CLK), .RN(n12625), .QN(
        n5742) );
  DFFR_X1 \REGISTERS_reg[79][29]  ( .D(n8846), .CK(CLK), .RN(n12610), .QN(
        n5774) );
  DFFR_X1 \REGISTERS_reg[79][28]  ( .D(n8847), .CK(CLK), .RN(n12617), .QN(
        n5806) );
  DFFR_X1 \REGISTERS_reg[79][27]  ( .D(n8848), .CK(CLK), .RN(n12588), .QN(
        n5838) );
  DFFR_X1 \REGISTERS_reg[79][26]  ( .D(n8849), .CK(CLK), .RN(n12566), .QN(
        n5870) );
  DFFR_X1 \REGISTERS_reg[79][25]  ( .D(n8850), .CK(CLK), .RN(n12544), .QN(
        n5902) );
  DFFR_X1 \REGISTERS_reg[79][24]  ( .D(n8851), .CK(CLK), .RN(n12506), .QN(
        n5934) );
  DFFR_X1 \REGISTERS_reg[79][23]  ( .D(n8852), .CK(CLK), .RN(n12632), .QN(
        n5998) );
  DFFR_X1 \REGISTERS_reg[79][22]  ( .D(n8853), .CK(CLK), .RN(n12522), .QN(
        n6315) );
  DFFR_X1 \REGISTERS_reg[79][21]  ( .D(n8854), .CK(CLK), .RN(n12529), .QN(
        n9165) );
  DFFR_X1 \REGISTERS_reg[79][20]  ( .D(n8855), .CK(CLK), .RN(n12504), .QN(
        n9197) );
  DFFR_X1 \REGISTERS_reg[79][19]  ( .D(n8856), .CK(CLK), .RN(n12595), .QN(
        n9261) );
  DFFR_X1 \REGISTERS_reg[79][18]  ( .D(n8857), .CK(CLK), .RN(n12446), .QN(
        n9595) );
  DFFR_X1 \REGISTERS_reg[79][17]  ( .D(n8858), .CK(CLK), .RN(n12454), .QN(
        n9627) );
  DFFR_X1 \REGISTERS_reg[79][16]  ( .D(n8859), .CK(CLK), .RN(n12460), .QN(
        n9659) );
  DFFR_X1 \REGISTERS_reg[79][15]  ( .D(n8860), .CK(CLK), .RN(n12639), .QN(
        n10021) );
  DFFR_X1 \REGISTERS_reg[79][14]  ( .D(n8861), .CK(CLK), .RN(n12467), .QN(
        n10053) );
  DFFR_X1 \REGISTERS_reg[79][13]  ( .D(n8862), .CK(CLK), .RN(n12475), .QN(
        n10085) );
  DFFR_X1 \REGISTERS_reg[79][12]  ( .D(n8863), .CK(CLK), .RN(n12482), .QN(
        n10117) );
  DFFR_X1 \REGISTERS_reg[79][11]  ( .D(n8864), .CK(CLK), .RN(n12573), .QN(
        n10149) );
  DFFR_X1 \REGISTERS_reg[79][10]  ( .D(n8865), .CK(CLK), .RN(n12551), .QN(
        n10181) );
  DFFR_X1 \REGISTERS_reg[79][9]  ( .D(n8866), .CK(CLK), .RN(n12559), .QN(
        n10215) );
  DFFR_X1 \REGISTERS_reg[79][8]  ( .D(n8867), .CK(CLK), .RN(n12537), .QN(
        n10247) );
  DFFR_X1 \REGISTERS_reg[79][7]  ( .D(n8868), .CK(CLK), .RN(n12647), .QN(
        n10279) );
  DFFR_X1 \REGISTERS_reg[79][6]  ( .D(n8869), .CK(CLK), .RN(n12603), .QN(
        n10314) );
  DFFR_X1 \REGISTERS_reg[79][5]  ( .D(n8870), .CK(CLK), .RN(n12489), .QN(
        n10346) );
  DFFR_X1 \REGISTERS_reg[79][4]  ( .D(n8871), .CK(CLK), .RN(n12497), .QN(
        n10378) );
  DFFR_X1 \REGISTERS_reg[79][3]  ( .D(n8872), .CK(CLK), .RN(n12581), .QN(
        n10413) );
  DFFR_X1 \REGISTERS_reg[79][2]  ( .D(n8873), .CK(CLK), .RN(n12511), .QN(
        n10445) );
  DFFR_X1 \REGISTERS_reg[79][1]  ( .D(n8874), .CK(CLK), .RN(n12439), .QN(
        n10477) );
  DFFR_X1 \REGISTERS_reg[79][0]  ( .D(n8875), .CK(CLK), .RN(n12654), .QN(
        n10509) );
  DFFR_X1 \REGISTERS_reg[80][6]  ( .D(n8901), .CK(CLK), .RN(n12603), .QN(
        n10315) );
  DFFR_X1 \REGISTERS_reg[80][5]  ( .D(n8902), .CK(CLK), .RN(n12490), .QN(
        n10347) );
  DFFR_X1 \REGISTERS_reg[80][4]  ( .D(n8903), .CK(CLK), .RN(n12497), .QN(
        n10379) );
  DFFR_X1 \REGISTERS_reg[80][3]  ( .D(n8904), .CK(CLK), .RN(n12581), .QN(
        n10414) );
  DFFR_X1 \REGISTERS_reg[80][2]  ( .D(n8905), .CK(CLK), .RN(n12512), .QN(
        n10446) );
  DFFR_X1 \REGISTERS_reg[80][1]  ( .D(n8906), .CK(CLK), .RN(n12439), .QN(
        n10478) );
  DFFR_X1 \REGISTERS_reg[80][0]  ( .D(n8907), .CK(CLK), .RN(n12654), .QN(
        n10510) );
  DLH_X1 \OUT2_reg[31]  ( .G(n12426), .D(N8767), .Q(OUT2[31]) );
  DLH_X1 \OUT1_reg[31]  ( .G(n12429), .D(N8734), .Q(OUT1[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(n12428), .D(N8766), .Q(OUT2[30]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n12429), .D(N8733), .Q(OUT1[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(n12428), .D(N8765), .Q(OUT2[29]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n12429), .D(N8732), .Q(OUT1[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(n12426), .D(N8764), .Q(OUT2[28]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n12429), .D(N8731), .Q(OUT1[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(n12428), .D(N8763), .Q(OUT2[27]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n12429), .D(N8730), .Q(OUT1[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(n12428), .D(N8762), .Q(OUT2[26]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n12430), .D(N8729), .Q(OUT1[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(n12428), .D(N8761), .Q(OUT2[25]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n12430), .D(N8728), .Q(OUT1[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(n12428), .D(N8760), .Q(OUT2[24]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n12430), .D(N8727), .Q(OUT1[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(n12426), .D(N8759), .Q(OUT2[23]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n12429), .D(N8726), .Q(OUT1[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(n12428), .D(N8758), .Q(OUT2[22]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n12430), .D(N8725), .Q(OUT1[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(n12426), .D(N8757), .Q(OUT2[21]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n12430), .D(N8724), .Q(OUT1[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(n12427), .D(N8756), .Q(OUT2[20]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n12431), .D(N8723), .Q(OUT1[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(n12426), .D(N8755), .Q(OUT2[19]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n12429), .D(N8722), .Q(OUT1[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(n12427), .D(N8754), .Q(OUT2[18]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n12431), .D(N8721), .Q(OUT1[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(n12427), .D(N8753), .Q(OUT2[17]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n12431), .D(N8720), .Q(OUT1[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(n12427), .D(N8752), .Q(OUT2[16]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n12431), .D(N8719), .Q(OUT1[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(n12426), .D(N8751), .Q(OUT2[15]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n12429), .D(N8718), .Q(OUT1[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(n12427), .D(N8750), .Q(OUT2[14]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n12431), .D(N8717), .Q(OUT1[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(n12427), .D(N8749), .Q(OUT2[13]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n12431), .D(N8716), .Q(OUT1[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(n12427), .D(N8748), .Q(OUT2[12]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n12431), .D(N8715), .Q(OUT1[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(n12428), .D(N8747), .Q(OUT2[11]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n12430), .D(N8714), .Q(OUT1[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(n12428), .D(N8746), .Q(OUT2[10]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n12430), .D(N8713), .Q(OUT1[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(n12426), .D(N8745), .Q(OUT2[9]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n12430), .D(N8712), .Q(OUT1[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(n12428), .D(N8744), .Q(OUT2[8]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n12430), .D(N8711), .Q(OUT1[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(n12426), .D(N8743), .Q(OUT2[7]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n12429), .D(N8710), .Q(OUT1[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(n12426), .D(N8742), .Q(OUT2[6]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n12429), .D(N8709), .Q(OUT1[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(n12427), .D(N8741), .Q(OUT2[5]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n12431), .D(N8708), .Q(OUT1[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(n12427), .D(N8740), .Q(OUT2[4]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n12431), .D(N8707), .Q(OUT1[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(n12426), .D(N8739), .Q(OUT2[3]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n12430), .D(N8706), .Q(OUT1[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(n12427), .D(N8738), .Q(OUT2[2]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n12430), .D(N8705), .Q(OUT1[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(n12427), .D(N8737), .Q(OUT2[1]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n12431), .D(N8704), .Q(OUT1[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(n12426), .D(N8736), .Q(OUT2[0]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n12429), .D(N8703), .Q(OUT1[0]) );
  NOR3_X2 U4359 ( .A1(N8580), .A2(N8581), .A3(N8579), .ZN(n4219) );
  NOR3_X2 U5825 ( .A1(N8436), .A2(N8437), .A3(N8435), .ZN(n5652) );
  NAND3_X1 U7835 ( .A1(n14517), .A2(n2483), .A3(RETRN), .ZN(n2480) );
  NAND3_X1 U7836 ( .A1(n2489), .A2(n14518), .A3(n14517), .ZN(n2481) );
  NAND3_X1 U7837 ( .A1(n2936), .A2(n2935), .A3(n2937), .ZN(n2483) );
  NAND3_X1 U7838 ( .A1(WR), .A2(ENABLE), .A3(wr_signal), .ZN(n2597) );
  XOR2_X1 \r486/U4  ( .A(\U3/U99/Z_5 ), .B(\r486/carry[5] ), .Z(N8580) );
  FA_X1 \r486/U1_4  ( .A(\U3/U99/Z_4 ), .B(ADD_RD2[4]), .CI(\r486/carry[4] ), 
        .CO(\r486/carry[5] ), .S(N8579) );
  XOR2_X1 \r480/U4  ( .A(\U3/U98/Z_5 ), .B(\r480/carry[5] ), .Z(N8436) );
  FA_X1 \r480/U1_4  ( .A(\U3/U98/Z_4 ), .B(ADD_RD1[4]), .CI(\r480/carry[4] ), 
        .CO(\r480/carry[5] ), .S(N8435) );
  XOR2_X1 \r472/U3  ( .A(\U3/U97/Z_5 ), .B(\r472/carry[5] ), .Z(N2172) );
  FA_X1 \r472/U1_4  ( .A(ADD_WR[4]), .B(\U3/U97/Z_4 ), .CI(\r472/carry[4] ), 
        .CO(\r472/carry[5] ), .S(N2171) );
  DFFR_X1 \REGISTERS_reg[87][31]  ( .D(n9100), .CK(CLK), .RN(RESET), .Q(n14481), .QN(n2882) );
  DFFR_X1 \REGISTERS_reg[87][30]  ( .D(n9101), .CK(CLK), .RN(n12625), .Q(
        n14482), .QN(n2883) );
  DFFR_X1 \REGISTERS_reg[87][29]  ( .D(n9102), .CK(CLK), .RN(n12611), .Q(
        n14483), .QN(n2884) );
  DFFR_X1 \REGISTERS_reg[87][28]  ( .D(n9103), .CK(CLK), .RN(n12618), .Q(
        n14484), .QN(n2885) );
  DFFR_X1 \REGISTERS_reg[87][27]  ( .D(n9104), .CK(CLK), .RN(n12589), .Q(
        n14485), .QN(n2886) );
  DFFR_X1 \REGISTERS_reg[87][26]  ( .D(n9105), .CK(CLK), .RN(n12567), .Q(
        n14486), .QN(n2887) );
  DFFR_X1 \REGISTERS_reg[87][25]  ( .D(n9106), .CK(CLK), .RN(n12545), .Q(
        n14487), .QN(n2888) );
  DFFR_X1 \REGISTERS_reg[87][24]  ( .D(n9107), .CK(CLK), .RN(n12505), .Q(
        n14488), .QN(n2889) );
  DFFR_X1 \REGISTERS_reg[87][23]  ( .D(n9108), .CK(CLK), .RN(n12633), .Q(
        n14489), .QN(n2890) );
  DFFR_X1 \REGISTERS_reg[87][22]  ( .D(n9109), .CK(CLK), .RN(n12523), .Q(
        n14490), .QN(n2891) );
  DFFR_X1 \REGISTERS_reg[87][21]  ( .D(n9110), .CK(CLK), .RN(n12530), .Q(
        n14491), .QN(n2892) );
  DFFR_X1 \REGISTERS_reg[87][20]  ( .D(n9111), .CK(CLK), .RN(n12505), .Q(
        n14492), .QN(n2893) );
  DFFR_X1 \REGISTERS_reg[87][19]  ( .D(n9112), .CK(CLK), .RN(n12596), .Q(
        n14493), .QN(n2894) );
  DFFR_X1 \REGISTERS_reg[87][18]  ( .D(n9113), .CK(CLK), .RN(n12447), .Q(
        n14494), .QN(n2895) );
  DFFR_X1 \REGISTERS_reg[87][17]  ( .D(n9114), .CK(CLK), .RN(n12454), .Q(
        n14495), .QN(n2896) );
  DFFR_X1 \REGISTERS_reg[87][16]  ( .D(n9115), .CK(CLK), .RN(n12461), .Q(
        n14496), .QN(n2897) );
  DFFR_X1 \REGISTERS_reg[87][15]  ( .D(n9116), .CK(CLK), .RN(n12640), .Q(
        n14497), .QN(n2898) );
  DFFR_X1 \REGISTERS_reg[87][14]  ( .D(n9117), .CK(CLK), .RN(n12468), .Q(
        n14498), .QN(n2899) );
  DFFR_X1 \REGISTERS_reg[87][13]  ( .D(n9118), .CK(CLK), .RN(n12475), .Q(
        n14499), .QN(n2900) );
  DFFR_X1 \REGISTERS_reg[87][12]  ( .D(n9119), .CK(CLK), .RN(n12483), .Q(
        n14500), .QN(n2901) );
  DFFR_X1 \REGISTERS_reg[87][11]  ( .D(n9120), .CK(CLK), .RN(n12574), .Q(
        n14501), .QN(n2902) );
  DFFR_X1 \REGISTERS_reg[87][10]  ( .D(n9121), .CK(CLK), .RN(n12552), .Q(
        n14502), .QN(n2903) );
  DFFR_X1 \REGISTERS_reg[87][9]  ( .D(n9122), .CK(CLK), .RN(n12559), .Q(n14503), .QN(n2904) );
  DFFR_X1 \REGISTERS_reg[87][8]  ( .D(n9123), .CK(CLK), .RN(n12537), .Q(n14504), .QN(n2905) );
  DFFR_X1 \REGISTERS_reg[87][7]  ( .D(n9124), .CK(CLK), .RN(n12647), .Q(n14505), .QN(n2906) );
  DFFR_X1 \REGISTERS_reg[87][6]  ( .D(n9125), .CK(CLK), .RN(n12603), .Q(n14506), .QN(n2907) );
  DFFR_X1 \REGISTERS_reg[87][5]  ( .D(n9126), .CK(CLK), .RN(n12490), .Q(n14507), .QN(n2908) );
  DFFR_X1 \REGISTERS_reg[87][4]  ( .D(n9127), .CK(CLK), .RN(n12497), .Q(n14508), .QN(n2909) );
  DFFR_X1 \REGISTERS_reg[87][3]  ( .D(n9128), .CK(CLK), .RN(n12581), .Q(n14509), .QN(n2910) );
  DFFR_X1 \REGISTERS_reg[87][2]  ( .D(n9129), .CK(CLK), .RN(n12512), .Q(n14510), .QN(n2911) );
  DFFR_X1 \REGISTERS_reg[87][1]  ( .D(n9130), .CK(CLK), .RN(n12440), .Q(n14511), .QN(n2912) );
  DFFR_X1 \REGISTERS_reg[87][0]  ( .D(n9131), .CK(CLK), .RN(n12655), .Q(n14512), .QN(n2913) );
  DFFR_X1 \REGISTERS_reg[86][31]  ( .D(n9068), .CK(CLK), .RN(n12662), .Q(
        n14449), .QN(n5714) );
  DFFR_X1 \REGISTERS_reg[86][30]  ( .D(n9069), .CK(CLK), .RN(n12625), .Q(
        n14450), .QN(n5746) );
  DFFR_X1 \REGISTERS_reg[86][29]  ( .D(n9070), .CK(CLK), .RN(n12611), .Q(
        n14451), .QN(n5778) );
  DFFR_X1 \REGISTERS_reg[86][28]  ( .D(n9071), .CK(CLK), .RN(n12618), .Q(
        n14452), .QN(n5810) );
  DFFR_X1 \REGISTERS_reg[86][27]  ( .D(n9072), .CK(CLK), .RN(n12589), .Q(
        n14453), .QN(n5842) );
  DFFR_X1 \REGISTERS_reg[86][26]  ( .D(n9073), .CK(CLK), .RN(n12567), .Q(
        n14454), .QN(n5874) );
  DFFR_X1 \REGISTERS_reg[86][25]  ( .D(n9074), .CK(CLK), .RN(n12545), .Q(
        n14455), .QN(n5906) );
  DFFR_X1 \REGISTERS_reg[86][24]  ( .D(n9075), .CK(CLK), .RN(n12504), .Q(
        n14456), .QN(n5938) );
  DFFR_X1 \REGISTERS_reg[86][23]  ( .D(n9076), .CK(CLK), .RN(n12633), .Q(
        n14457), .QN(n6002) );
  DFFR_X1 \REGISTERS_reg[86][22]  ( .D(n9077), .CK(CLK), .RN(n12523), .Q(
        n14458), .QN(n9137) );
  DFFR_X1 \REGISTERS_reg[86][21]  ( .D(n9078), .CK(CLK), .RN(n12530), .Q(
        n14459), .QN(n9169) );
  DFFR_X1 \REGISTERS_reg[86][20]  ( .D(n9079), .CK(CLK), .RN(n12505), .Q(
        n14460), .QN(n9201) );
  DFFR_X1 \REGISTERS_reg[86][19]  ( .D(n9080), .CK(CLK), .RN(n12596), .Q(
        n14461), .QN(n9311) );
  DFFR_X1 \REGISTERS_reg[86][18]  ( .D(n9081), .CK(CLK), .RN(n12447), .Q(
        n14462), .QN(n9599) );
  DFFR_X1 \REGISTERS_reg[86][17]  ( .D(n9082), .CK(CLK), .RN(n12454), .Q(
        n14463), .QN(n9631) );
  DFFR_X1 \REGISTERS_reg[86][16]  ( .D(n9083), .CK(CLK), .RN(n12461), .Q(
        n14464), .QN(n9663) );
  DFFR_X1 \REGISTERS_reg[86][15]  ( .D(n9084), .CK(CLK), .RN(n12640), .Q(
        n14465), .QN(n10025) );
  DFFR_X1 \REGISTERS_reg[86][14]  ( .D(n9085), .CK(CLK), .RN(n12468), .Q(
        n14466), .QN(n10057) );
  DFFR_X1 \REGISTERS_reg[86][13]  ( .D(n9086), .CK(CLK), .RN(n12475), .Q(
        n14467), .QN(n10089) );
  DFFR_X1 \REGISTERS_reg[86][12]  ( .D(n9087), .CK(CLK), .RN(n12483), .Q(
        n14468), .QN(n10121) );
  DFFR_X1 \REGISTERS_reg[86][11]  ( .D(n9088), .CK(CLK), .RN(n12574), .Q(
        n14469), .QN(n10153) );
  DFFR_X1 \REGISTERS_reg[86][10]  ( .D(n9089), .CK(CLK), .RN(n12552), .Q(
        n14470), .QN(n10185) );
  DFFR_X1 \REGISTERS_reg[86][9]  ( .D(n9090), .CK(CLK), .RN(n12559), .Q(n14471), .QN(n10219) );
  DFFR_X1 \REGISTERS_reg[86][8]  ( .D(n9091), .CK(CLK), .RN(n12537), .Q(n14472), .QN(n10251) );
  DFFR_X1 \REGISTERS_reg[86][7]  ( .D(n9092), .CK(CLK), .RN(n12647), .Q(n14473), .QN(n10283) );
  DFFR_X1 \REGISTERS_reg[86][6]  ( .D(n9093), .CK(CLK), .RN(n12603), .Q(n14474), .QN(n10318) );
  DFFR_X1 \REGISTERS_reg[86][5]  ( .D(n9094), .CK(CLK), .RN(n12490), .Q(n14475), .QN(n10350) );
  DFFR_X1 \REGISTERS_reg[86][4]  ( .D(n9095), .CK(CLK), .RN(n12497), .Q(n14476), .QN(n10382) );
  DFFR_X1 \REGISTERS_reg[86][3]  ( .D(n9096), .CK(CLK), .RN(n12581), .Q(n14477), .QN(n10417) );
  DFFR_X1 \REGISTERS_reg[86][2]  ( .D(n9097), .CK(CLK), .RN(n12512), .Q(n14478), .QN(n10449) );
  DFFR_X1 \REGISTERS_reg[86][1]  ( .D(n9098), .CK(CLK), .RN(n12440), .Q(n14479), .QN(n10481) );
  DFFR_X1 \REGISTERS_reg[86][0]  ( .D(n9099), .CK(CLK), .RN(n12655), .Q(n14480), .QN(n10513) );
  DFFR_X1 \REGISTERS_reg[85][31]  ( .D(n9036), .CK(CLK), .RN(n12662), .Q(
        n14417), .QN(n2818) );
  DFFR_X1 \REGISTERS_reg[85][30]  ( .D(n9037), .CK(CLK), .RN(n12625), .Q(
        n14418), .QN(n2819) );
  DFFR_X1 \REGISTERS_reg[85][29]  ( .D(n9038), .CK(CLK), .RN(n12611), .Q(
        n14419), .QN(n2820) );
  DFFR_X1 \REGISTERS_reg[85][28]  ( .D(n9039), .CK(CLK), .RN(n12618), .Q(
        n14420), .QN(n2821) );
  DFFR_X1 \REGISTERS_reg[85][27]  ( .D(n9040), .CK(CLK), .RN(n12589), .Q(
        n14421), .QN(n2822) );
  DFFR_X1 \REGISTERS_reg[85][26]  ( .D(n9041), .CK(CLK), .RN(n12567), .Q(
        n14422), .QN(n2823) );
  DFFR_X1 \REGISTERS_reg[85][25]  ( .D(n9042), .CK(CLK), .RN(n12545), .Q(
        n14423), .QN(n2824) );
  DFFR_X1 \REGISTERS_reg[85][24]  ( .D(n9043), .CK(CLK), .RN(n12503), .Q(
        n14424), .QN(n2825) );
  DFFR_X1 \REGISTERS_reg[85][23]  ( .D(n9044), .CK(CLK), .RN(n12633), .Q(
        n14425), .QN(n2826) );
  DFFR_X1 \REGISTERS_reg[85][22]  ( .D(n9045), .CK(CLK), .RN(n12523), .Q(
        n14426), .QN(n2827) );
  DFFR_X1 \REGISTERS_reg[85][21]  ( .D(n9046), .CK(CLK), .RN(n12530), .Q(
        n14427), .QN(n2828) );
  DFFR_X1 \REGISTERS_reg[85][20]  ( .D(n9047), .CK(CLK), .RN(n12505), .Q(
        n14428), .QN(n2829) );
  DFFR_X1 \REGISTERS_reg[85][19]  ( .D(n9048), .CK(CLK), .RN(n12596), .Q(
        n14429), .QN(n2830) );
  DFFR_X1 \REGISTERS_reg[85][18]  ( .D(n9049), .CK(CLK), .RN(n12447), .Q(
        n14430), .QN(n2831) );
  DFFR_X1 \REGISTERS_reg[85][17]  ( .D(n9050), .CK(CLK), .RN(n12454), .Q(
        n14431), .QN(n2832) );
  DFFR_X1 \REGISTERS_reg[85][16]  ( .D(n9051), .CK(CLK), .RN(n12461), .Q(
        n14432), .QN(n2833) );
  DFFR_X1 \REGISTERS_reg[85][15]  ( .D(n9052), .CK(CLK), .RN(n12640), .Q(
        n14433), .QN(n2834) );
  DFFR_X1 \REGISTERS_reg[85][14]  ( .D(n9053), .CK(CLK), .RN(n12468), .Q(
        n14434), .QN(n2835) );
  DFFR_X1 \REGISTERS_reg[85][13]  ( .D(n9054), .CK(CLK), .RN(n12475), .Q(
        n14435), .QN(n2836) );
  DFFR_X1 \REGISTERS_reg[85][12]  ( .D(n9055), .CK(CLK), .RN(n12483), .Q(
        n14436), .QN(n2837) );
  DFFR_X1 \REGISTERS_reg[85][11]  ( .D(n9056), .CK(CLK), .RN(n12574), .Q(
        n14437), .QN(n2838) );
  DFFR_X1 \REGISTERS_reg[85][10]  ( .D(n9057), .CK(CLK), .RN(n12552), .Q(
        n14438), .QN(n2839) );
  DFFR_X1 \REGISTERS_reg[85][9]  ( .D(n9058), .CK(CLK), .RN(n12559), .Q(n14439), .QN(n2840) );
  DFFR_X1 \REGISTERS_reg[85][8]  ( .D(n9059), .CK(CLK), .RN(n12537), .Q(n14440), .QN(n2841) );
  DFFR_X1 \REGISTERS_reg[85][7]  ( .D(n9060), .CK(CLK), .RN(n12647), .Q(n14441), .QN(n2842) );
  DFFR_X1 \REGISTERS_reg[85][6]  ( .D(n9061), .CK(CLK), .RN(n12603), .Q(n14442), .QN(n2843) );
  DFFR_X1 \REGISTERS_reg[85][5]  ( .D(n9062), .CK(CLK), .RN(n12490), .Q(n14443), .QN(n2844) );
  DFFR_X1 \REGISTERS_reg[85][4]  ( .D(n9063), .CK(CLK), .RN(n12497), .Q(n14444), .QN(n2845) );
  DFFR_X1 \REGISTERS_reg[85][3]  ( .D(n9064), .CK(CLK), .RN(n12581), .Q(n14445), .QN(n2846) );
  DFFR_X1 \REGISTERS_reg[85][2]  ( .D(n9065), .CK(CLK), .RN(n12512), .Q(n14446), .QN(n2847) );
  DFFR_X1 \REGISTERS_reg[85][1]  ( .D(n9066), .CK(CLK), .RN(n12440), .Q(n14447), .QN(n2848) );
  DFFR_X1 \REGISTERS_reg[85][0]  ( .D(n9067), .CK(CLK), .RN(n12655), .Q(n14448), .QN(n2849) );
  DFFR_X1 \REGISTERS_reg[84][31]  ( .D(n9004), .CK(CLK), .RN(n12662), .Q(
        n14385), .QN(n5708) );
  DFFR_X1 \REGISTERS_reg[84][30]  ( .D(n9005), .CK(CLK), .RN(n12625), .Q(
        n14386), .QN(n5740) );
  DFFR_X1 \REGISTERS_reg[84][29]  ( .D(n9006), .CK(CLK), .RN(n12611), .Q(
        n14387), .QN(n5772) );
  DFFR_X1 \REGISTERS_reg[84][28]  ( .D(n9007), .CK(CLK), .RN(n12618), .Q(
        n14388), .QN(n5804) );
  DFFR_X1 \REGISTERS_reg[84][27]  ( .D(n9008), .CK(CLK), .RN(n12589), .Q(
        n14389), .QN(n5836) );
  DFFR_X1 \REGISTERS_reg[84][26]  ( .D(n9009), .CK(CLK), .RN(n12567), .Q(
        n14390), .QN(n5868) );
  DFFR_X1 \REGISTERS_reg[84][25]  ( .D(n9010), .CK(CLK), .RN(n12545), .Q(
        n14391), .QN(n5900) );
  DFFR_X1 \REGISTERS_reg[84][24]  ( .D(n9011), .CK(CLK), .RN(n12509), .Q(
        n14392), .QN(n5932) );
  DFFR_X1 \REGISTERS_reg[84][23]  ( .D(n9012), .CK(CLK), .RN(n12633), .Q(
        n14393), .QN(n5996) );
  DFFR_X1 \REGISTERS_reg[84][22]  ( .D(n9013), .CK(CLK), .RN(n12523), .Q(
        n14394), .QN(n6313) );
  DFFR_X1 \REGISTERS_reg[84][21]  ( .D(n9014), .CK(CLK), .RN(n12530), .Q(
        n14395), .QN(n9163) );
  DFFR_X1 \REGISTERS_reg[84][20]  ( .D(n9015), .CK(CLK), .RN(n12505), .Q(
        n14396), .QN(n9195) );
  DFFR_X1 \REGISTERS_reg[84][19]  ( .D(n9016), .CK(CLK), .RN(n12596), .Q(
        n14397), .QN(n9259) );
  DFFR_X1 \REGISTERS_reg[84][18]  ( .D(n9017), .CK(CLK), .RN(n12447), .Q(
        n14398), .QN(n9593) );
  DFFR_X1 \REGISTERS_reg[84][17]  ( .D(n9018), .CK(CLK), .RN(n12454), .Q(
        n14399), .QN(n9625) );
  DFFR_X1 \REGISTERS_reg[84][16]  ( .D(n9019), .CK(CLK), .RN(n12461), .Q(
        n14400), .QN(n9657) );
  DFFR_X1 \REGISTERS_reg[84][15]  ( .D(n9020), .CK(CLK), .RN(n12640), .Q(
        n14401), .QN(n10019) );
  DFFR_X1 \REGISTERS_reg[84][14]  ( .D(n9021), .CK(CLK), .RN(n12468), .Q(
        n14402), .QN(n10051) );
  DFFR_X1 \REGISTERS_reg[84][13]  ( .D(n9022), .CK(CLK), .RN(n12475), .Q(
        n14403), .QN(n10083) );
  DFFR_X1 \REGISTERS_reg[84][12]  ( .D(n9023), .CK(CLK), .RN(n12483), .Q(
        n14404), .QN(n10115) );
  DFFR_X1 \REGISTERS_reg[84][11]  ( .D(n9024), .CK(CLK), .RN(n12574), .Q(
        n14405), .QN(n10147) );
  DFFR_X1 \REGISTERS_reg[84][10]  ( .D(n9025), .CK(CLK), .RN(n12552), .Q(
        n14406), .QN(n10179) );
  DFFR_X1 \REGISTERS_reg[84][9]  ( .D(n9026), .CK(CLK), .RN(n12559), .Q(n14407), .QN(n10213) );
  DFFR_X1 \REGISTERS_reg[84][8]  ( .D(n9027), .CK(CLK), .RN(n12537), .Q(n14408), .QN(n10245) );
  DFFR_X1 \REGISTERS_reg[84][7]  ( .D(n9028), .CK(CLK), .RN(n12647), .Q(n14409), .QN(n10277) );
  DFFR_X1 \REGISTERS_reg[84][6]  ( .D(n9029), .CK(CLK), .RN(n12603), .Q(n14410), .QN(n10312) );
  DFFR_X1 \REGISTERS_reg[84][5]  ( .D(n9030), .CK(CLK), .RN(n12490), .Q(n14411), .QN(n10344) );
  DFFR_X1 \REGISTERS_reg[84][4]  ( .D(n9031), .CK(CLK), .RN(n12497), .Q(n14412), .QN(n10376) );
  DFFR_X1 \REGISTERS_reg[84][3]  ( .D(n9032), .CK(CLK), .RN(n12581), .Q(n14413), .QN(n10411) );
  DFFR_X1 \REGISTERS_reg[84][2]  ( .D(n9033), .CK(CLK), .RN(n12512), .Q(n14414), .QN(n10443) );
  DFFR_X1 \REGISTERS_reg[84][1]  ( .D(n9034), .CK(CLK), .RN(n12440), .Q(n14415), .QN(n10475) );
  DFFR_X1 \REGISTERS_reg[84][0]  ( .D(n9035), .CK(CLK), .RN(n12655), .Q(n14416), .QN(n10507) );
  DFFR_X1 \REGISTERS_reg[83][31]  ( .D(n8972), .CK(CLK), .RN(n12662), .Q(
        n14353), .QN(n2754) );
  DFFR_X1 \REGISTERS_reg[83][30]  ( .D(n8973), .CK(CLK), .RN(n12625), .Q(
        n14354), .QN(n2755) );
  DFFR_X1 \REGISTERS_reg[83][29]  ( .D(n8974), .CK(CLK), .RN(n12610), .Q(
        n14355), .QN(n2756) );
  DFFR_X1 \REGISTERS_reg[83][28]  ( .D(n8975), .CK(CLK), .RN(n12618), .Q(
        n14356), .QN(n2757) );
  DFFR_X1 \REGISTERS_reg[83][27]  ( .D(n8976), .CK(CLK), .RN(n12588), .Q(
        n14357), .QN(n2758) );
  DFFR_X1 \REGISTERS_reg[83][26]  ( .D(n8977), .CK(CLK), .RN(n12566), .Q(
        n14358), .QN(n2759) );
  DFFR_X1 \REGISTERS_reg[83][25]  ( .D(n8978), .CK(CLK), .RN(n12544), .Q(
        n14359), .QN(n2760) );
  DFFR_X1 \REGISTERS_reg[83][24]  ( .D(n8979), .CK(CLK), .RN(n12454), .Q(
        n14360), .QN(n2761) );
  DFFR_X1 \REGISTERS_reg[83][23]  ( .D(n8980), .CK(CLK), .RN(n12632), .Q(
        n14361), .QN(n2762) );
  DFFR_X1 \REGISTERS_reg[83][22]  ( .D(n8981), .CK(CLK), .RN(n12522), .Q(
        n14362), .QN(n2763) );
  DFFR_X1 \REGISTERS_reg[83][21]  ( .D(n8982), .CK(CLK), .RN(n12530), .Q(
        n14363), .QN(n2764) );
  DFFR_X1 \REGISTERS_reg[83][20]  ( .D(n8983), .CK(CLK), .RN(n12504), .Q(
        n14364), .QN(n2765) );
  DFFR_X1 \REGISTERS_reg[83][19]  ( .D(n8984), .CK(CLK), .RN(n12596), .Q(
        n14365), .QN(n2766) );
  DFFR_X1 \REGISTERS_reg[83][18]  ( .D(n8985), .CK(CLK), .RN(n12447), .Q(
        n14366), .QN(n2767) );
  DFFR_X1 \REGISTERS_reg[83][17]  ( .D(n8986), .CK(CLK), .RN(n12454), .Q(
        n14367), .QN(n2768) );
  DFFR_X1 \REGISTERS_reg[83][16]  ( .D(n8987), .CK(CLK), .RN(n12460), .Q(
        n14368), .QN(n2769) );
  DFFR_X1 \REGISTERS_reg[83][15]  ( .D(n8988), .CK(CLK), .RN(n12640), .Q(
        n14369), .QN(n2770) );
  DFFR_X1 \REGISTERS_reg[83][14]  ( .D(n8989), .CK(CLK), .RN(n12468), .Q(
        n14370), .QN(n2771) );
  DFFR_X1 \REGISTERS_reg[83][13]  ( .D(n8990), .CK(CLK), .RN(n12475), .Q(
        n14371), .QN(n2772) );
  DFFR_X1 \REGISTERS_reg[83][12]  ( .D(n8991), .CK(CLK), .RN(n12482), .Q(
        n14372), .QN(n2773) );
  DFFR_X1 \REGISTERS_reg[83][11]  ( .D(n8992), .CK(CLK), .RN(n12574), .Q(
        n14373), .QN(n2774) );
  DFFR_X1 \REGISTERS_reg[83][10]  ( .D(n8993), .CK(CLK), .RN(n12552), .Q(
        n14374), .QN(n2775) );
  DFFR_X1 \REGISTERS_reg[83][9]  ( .D(n8994), .CK(CLK), .RN(n12559), .Q(n14375), .QN(n2776) );
  DFFR_X1 \REGISTERS_reg[83][8]  ( .D(n8995), .CK(CLK), .RN(n12537), .Q(n14376), .QN(n2777) );
  DFFR_X1 \REGISTERS_reg[83][7]  ( .D(n8996), .CK(CLK), .RN(n12647), .Q(n14377), .QN(n2778) );
  DFFR_X1 \REGISTERS_reg[83][6]  ( .D(n8997), .CK(CLK), .RN(n12603), .Q(n14378), .QN(n2779) );
  DFFR_X1 \REGISTERS_reg[83][5]  ( .D(n8998), .CK(CLK), .RN(n12490), .Q(n14379), .QN(n2780) );
  DFFR_X1 \REGISTERS_reg[83][4]  ( .D(n8999), .CK(CLK), .RN(n12497), .Q(n14380), .QN(n2781) );
  DFFR_X1 \REGISTERS_reg[83][3]  ( .D(n9000), .CK(CLK), .RN(n12581), .Q(n14381), .QN(n2782) );
  DFFR_X1 \REGISTERS_reg[83][2]  ( .D(n9001), .CK(CLK), .RN(n12512), .Q(n14382), .QN(n2783) );
  DFFR_X1 \REGISTERS_reg[83][1]  ( .D(n9002), .CK(CLK), .RN(n12439), .Q(n14383), .QN(n2784) );
  DFFR_X1 \REGISTERS_reg[83][0]  ( .D(n9003), .CK(CLK), .RN(n12654), .Q(n14384), .QN(n2785) );
  DFFR_X1 \REGISTERS_reg[82][31]  ( .D(n8940), .CK(CLK), .RN(n12662), .Q(
        n14321), .QN(n5707) );
  DFFR_X1 \REGISTERS_reg[82][30]  ( .D(n8941), .CK(CLK), .RN(n12625), .Q(
        n14322), .QN(n5739) );
  DFFR_X1 \REGISTERS_reg[82][29]  ( .D(n8942), .CK(CLK), .RN(n12610), .Q(
        n14323), .QN(n5771) );
  DFFR_X1 \REGISTERS_reg[82][28]  ( .D(n8943), .CK(CLK), .RN(n12618), .Q(
        n14324), .QN(n5803) );
  DFFR_X1 \REGISTERS_reg[82][27]  ( .D(n8944), .CK(CLK), .RN(n12588), .Q(
        n14325), .QN(n5835) );
  DFFR_X1 \REGISTERS_reg[82][26]  ( .D(n8945), .CK(CLK), .RN(n12566), .Q(
        n14326), .QN(n5867) );
  DFFR_X1 \REGISTERS_reg[82][25]  ( .D(n8946), .CK(CLK), .RN(n12544), .Q(
        n14327), .QN(n5899) );
  DFFR_X1 \REGISTERS_reg[82][24]  ( .D(n8947), .CK(CLK), .RN(n12453), .Q(
        n14328), .QN(n5931) );
  DFFR_X1 \REGISTERS_reg[82][23]  ( .D(n8948), .CK(CLK), .RN(n12632), .Q(
        n14329), .QN(n5995) );
  DFFR_X1 \REGISTERS_reg[82][22]  ( .D(n8949), .CK(CLK), .RN(n12522), .Q(
        n14330), .QN(n6312) );
  DFFR_X1 \REGISTERS_reg[82][21]  ( .D(n8950), .CK(CLK), .RN(n12530), .Q(
        n14331), .QN(n9162) );
  DFFR_X1 \REGISTERS_reg[82][20]  ( .D(n8951), .CK(CLK), .RN(n12504), .Q(
        n14332), .QN(n9194) );
  DFFR_X1 \REGISTERS_reg[82][19]  ( .D(n8952), .CK(CLK), .RN(n12596), .Q(
        n14333), .QN(n9258) );
  DFFR_X1 \REGISTERS_reg[82][18]  ( .D(n8953), .CK(CLK), .RN(n12447), .Q(
        n14334), .QN(n9592) );
  DFFR_X1 \REGISTERS_reg[82][17]  ( .D(n8954), .CK(CLK), .RN(n12454), .Q(
        n14335), .QN(n9624) );
  DFFR_X1 \REGISTERS_reg[82][16]  ( .D(n8955), .CK(CLK), .RN(n12460), .Q(
        n14336), .QN(n9656) );
  DFFR_X1 \REGISTERS_reg[82][15]  ( .D(n8956), .CK(CLK), .RN(n12640), .Q(
        n14337), .QN(n10018) );
  DFFR_X1 \REGISTERS_reg[82][14]  ( .D(n8957), .CK(CLK), .RN(n12468), .Q(
        n14338), .QN(n10050) );
  DFFR_X1 \REGISTERS_reg[82][13]  ( .D(n8958), .CK(CLK), .RN(n12475), .Q(
        n14339), .QN(n10082) );
  DFFR_X1 \REGISTERS_reg[82][12]  ( .D(n8959), .CK(CLK), .RN(n12482), .Q(
        n14340), .QN(n10114) );
  DFFR_X1 \REGISTERS_reg[82][11]  ( .D(n8960), .CK(CLK), .RN(n12574), .Q(
        n14341), .QN(n10146) );
  DFFR_X1 \REGISTERS_reg[82][10]  ( .D(n8961), .CK(CLK), .RN(n12552), .Q(
        n14342), .QN(n10178) );
  DFFR_X1 \REGISTERS_reg[82][9]  ( .D(n8962), .CK(CLK), .RN(n12559), .Q(n14343), .QN(n10212) );
  DFFR_X1 \REGISTERS_reg[82][8]  ( .D(n8963), .CK(CLK), .RN(n12537), .Q(n14344), .QN(n10244) );
  DFFR_X1 \REGISTERS_reg[82][7]  ( .D(n8964), .CK(CLK), .RN(n12647), .Q(n14345), .QN(n10276) );
  DFFR_X1 \REGISTERS_reg[82][6]  ( .D(n8965), .CK(CLK), .RN(n12603), .Q(n14346), .QN(n10311) );
  DFFR_X1 \REGISTERS_reg[82][5]  ( .D(n8966), .CK(CLK), .RN(n12490), .Q(n14347), .QN(n10343) );
  DFFR_X1 \REGISTERS_reg[82][4]  ( .D(n8967), .CK(CLK), .RN(n12497), .Q(n14348), .QN(n10375) );
  DFFR_X1 \REGISTERS_reg[82][3]  ( .D(n8968), .CK(CLK), .RN(n12581), .Q(n14349), .QN(n10410) );
  DFFR_X1 \REGISTERS_reg[82][2]  ( .D(n8969), .CK(CLK), .RN(n12512), .Q(n14350), .QN(n10442) );
  DFFR_X1 \REGISTERS_reg[82][1]  ( .D(n8970), .CK(CLK), .RN(n12439), .Q(n14351), .QN(n10474) );
  DFFR_X1 \REGISTERS_reg[82][0]  ( .D(n8971), .CK(CLK), .RN(n12654), .Q(n14352), .QN(n10506) );
  DFFR_X1 \REGISTERS_reg[81][31]  ( .D(n8908), .CK(CLK), .RN(n12662), .Q(
        n14289), .QN(n5709) );
  DFFR_X1 \REGISTERS_reg[81][30]  ( .D(n8909), .CK(CLK), .RN(n12625), .Q(
        n14290), .QN(n5741) );
  DFFR_X1 \REGISTERS_reg[81][29]  ( .D(n8910), .CK(CLK), .RN(n12610), .Q(
        n14291), .QN(n5773) );
  DFFR_X1 \REGISTERS_reg[81][28]  ( .D(n8911), .CK(CLK), .RN(n12618), .Q(
        n14292), .QN(n5805) );
  DFFR_X1 \REGISTERS_reg[81][27]  ( .D(n8912), .CK(CLK), .RN(n12588), .Q(
        n14293), .QN(n5837) );
  DFFR_X1 \REGISTERS_reg[81][26]  ( .D(n8913), .CK(CLK), .RN(n12566), .Q(
        n14294), .QN(n5869) );
  DFFR_X1 \REGISTERS_reg[81][25]  ( .D(n8914), .CK(CLK), .RN(n12544), .Q(
        n14295), .QN(n5901) );
  DFFR_X1 \REGISTERS_reg[81][24]  ( .D(n8915), .CK(CLK), .RN(n12452), .Q(
        n14296), .QN(n5933) );
  DFFR_X1 \REGISTERS_reg[81][23]  ( .D(n8916), .CK(CLK), .RN(n12632), .Q(
        n14297), .QN(n5997) );
  DFFR_X1 \REGISTERS_reg[81][22]  ( .D(n8917), .CK(CLK), .RN(n12522), .Q(
        n14298), .QN(n6314) );
  DFFR_X1 \REGISTERS_reg[81][21]  ( .D(n8918), .CK(CLK), .RN(n12530), .Q(
        n14299), .QN(n9164) );
  DFFR_X1 \REGISTERS_reg[81][20]  ( .D(n8919), .CK(CLK), .RN(n12504), .Q(
        n14300), .QN(n9196) );
  DFFR_X1 \REGISTERS_reg[81][19]  ( .D(n8920), .CK(CLK), .RN(n12596), .Q(
        n14301), .QN(n9260) );
  DFFR_X1 \REGISTERS_reg[81][18]  ( .D(n8921), .CK(CLK), .RN(n12447), .Q(
        n14302), .QN(n9594) );
  DFFR_X1 \REGISTERS_reg[81][17]  ( .D(n8922), .CK(CLK), .RN(n12454), .Q(
        n14303), .QN(n9626) );
  DFFR_X1 \REGISTERS_reg[81][16]  ( .D(n8923), .CK(CLK), .RN(n12460), .Q(
        n14304), .QN(n9658) );
  DFFR_X1 \REGISTERS_reg[81][15]  ( .D(n8924), .CK(CLK), .RN(n12640), .Q(
        n14305), .QN(n10020) );
  DFFR_X1 \REGISTERS_reg[81][14]  ( .D(n8925), .CK(CLK), .RN(n12468), .Q(
        n14306), .QN(n10052) );
  DFFR_X1 \REGISTERS_reg[81][13]  ( .D(n8926), .CK(CLK), .RN(n12475), .Q(
        n14307), .QN(n10084) );
  DFFR_X1 \REGISTERS_reg[81][12]  ( .D(n8927), .CK(CLK), .RN(n12482), .Q(
        n14308), .QN(n10116) );
  DFFR_X1 \REGISTERS_reg[81][11]  ( .D(n8928), .CK(CLK), .RN(n12574), .Q(
        n14309), .QN(n10148) );
  DFFR_X1 \REGISTERS_reg[81][10]  ( .D(n8929), .CK(CLK), .RN(n12552), .Q(
        n14310), .QN(n10180) );
  DFFR_X1 \REGISTERS_reg[81][9]  ( .D(n8930), .CK(CLK), .RN(n12559), .Q(n14311), .QN(n10214) );
  DFFR_X1 \REGISTERS_reg[81][8]  ( .D(n8931), .CK(CLK), .RN(n12537), .Q(n14312), .QN(n10246) );
  DFFR_X1 \REGISTERS_reg[81][7]  ( .D(n8932), .CK(CLK), .RN(n12647), .Q(n14313), .QN(n10278) );
  DFFR_X1 \REGISTERS_reg[81][6]  ( .D(n8933), .CK(CLK), .RN(n12603), .Q(n14314), .QN(n10313) );
  DFFR_X1 \REGISTERS_reg[81][5]  ( .D(n8934), .CK(CLK), .RN(n12490), .Q(n14315), .QN(n10345) );
  DFFR_X1 \REGISTERS_reg[81][4]  ( .D(n8935), .CK(CLK), .RN(n12497), .Q(n14316), .QN(n10377) );
  DFFR_X1 \REGISTERS_reg[81][3]  ( .D(n8936), .CK(CLK), .RN(n12581), .Q(n14317), .QN(n10412) );
  DFFR_X1 \REGISTERS_reg[81][2]  ( .D(n8937), .CK(CLK), .RN(n12512), .Q(n14318), .QN(n10444) );
  DFFR_X1 \REGISTERS_reg[81][1]  ( .D(n8938), .CK(CLK), .RN(n12439), .Q(n14319), .QN(n10476) );
  DFFR_X1 \REGISTERS_reg[81][0]  ( .D(n8939), .CK(CLK), .RN(n12654), .Q(n14320), .QN(n10508) );
  DFFR_X1 \REGISTERS_reg[77][31]  ( .D(n8780), .CK(CLK), .RN(n12661), .Q(
        n14257), .QN(n5713) );
  DFFR_X1 \REGISTERS_reg[77][30]  ( .D(n8781), .CK(CLK), .RN(n12625), .Q(
        n14258), .QN(n5745) );
  DFFR_X1 \REGISTERS_reg[77][29]  ( .D(n8782), .CK(CLK), .RN(n12610), .Q(
        n14259), .QN(n5777) );
  DFFR_X1 \REGISTERS_reg[77][28]  ( .D(n8783), .CK(CLK), .RN(n12617), .Q(
        n14260), .QN(n5809) );
  DFFR_X1 \REGISTERS_reg[77][27]  ( .D(n8784), .CK(CLK), .RN(n12588), .Q(
        n14261), .QN(n5841) );
  DFFR_X1 \REGISTERS_reg[77][26]  ( .D(n8785), .CK(CLK), .RN(n12566), .Q(
        n14262), .QN(n5873) );
  DFFR_X1 \REGISTERS_reg[77][25]  ( .D(n8786), .CK(CLK), .RN(n12544), .Q(
        n14263), .QN(n5905) );
  DFFR_X1 \REGISTERS_reg[77][24]  ( .D(n8787), .CK(CLK), .RN(n12451), .Q(
        n14264), .QN(n5937) );
  DFFR_X1 \REGISTERS_reg[77][23]  ( .D(n8788), .CK(CLK), .RN(n12632), .Q(
        n14265), .QN(n6001) );
  DFFR_X1 \REGISTERS_reg[77][22]  ( .D(n8789), .CK(CLK), .RN(n12522), .Q(
        n14266), .QN(n9136) );
  DFFR_X1 \REGISTERS_reg[77][21]  ( .D(n8790), .CK(CLK), .RN(n12529), .Q(
        n14267), .QN(n9168) );
  DFFR_X1 \REGISTERS_reg[77][20]  ( .D(n8791), .CK(CLK), .RN(n12504), .Q(
        n14268), .QN(n9200) );
  DFFR_X1 \REGISTERS_reg[77][19]  ( .D(n8792), .CK(CLK), .RN(n12595), .Q(
        n14269), .QN(n9264) );
  DFFR_X1 \REGISTERS_reg[77][18]  ( .D(n8793), .CK(CLK), .RN(n12446), .Q(
        n14270), .QN(n9598) );
  DFFR_X1 \REGISTERS_reg[77][17]  ( .D(n8794), .CK(CLK), .RN(n12454), .Q(
        n14271), .QN(n9630) );
  DFFR_X1 \REGISTERS_reg[77][16]  ( .D(n8795), .CK(CLK), .RN(n12460), .Q(
        n14272), .QN(n9662) );
  DFFR_X1 \REGISTERS_reg[77][15]  ( .D(n8796), .CK(CLK), .RN(n12639), .Q(
        n14273), .QN(n10024) );
  DFFR_X1 \REGISTERS_reg[77][14]  ( .D(n8797), .CK(CLK), .RN(n12467), .Q(
        n14274), .QN(n10056) );
  DFFR_X1 \REGISTERS_reg[77][13]  ( .D(n8798), .CK(CLK), .RN(n12475), .Q(
        n14275), .QN(n10088) );
  DFFR_X1 \REGISTERS_reg[77][12]  ( .D(n8799), .CK(CLK), .RN(n12482), .Q(
        n14276), .QN(n10120) );
  DFFR_X1 \REGISTERS_reg[77][11]  ( .D(n8800), .CK(CLK), .RN(n12573), .Q(
        n14277), .QN(n10152) );
  DFFR_X1 \REGISTERS_reg[77][10]  ( .D(n8801), .CK(CLK), .RN(n12551), .Q(
        n14278), .QN(n10184) );
  DFFR_X1 \REGISTERS_reg[77][9]  ( .D(n8802), .CK(CLK), .RN(n12559), .Q(n14279), .QN(n10218) );
  DFFR_X1 \REGISTERS_reg[77][8]  ( .D(n8803), .CK(CLK), .RN(n12537), .Q(n14280), .QN(n10250) );
  DFFR_X1 \REGISTERS_reg[77][7]  ( .D(n8804), .CK(CLK), .RN(n12647), .Q(n14281), .QN(n10282) );
  DFFR_X1 \REGISTERS_reg[77][6]  ( .D(n8805), .CK(CLK), .RN(n12603), .Q(n14282), .QN(n10317) );
  DFFR_X1 \REGISTERS_reg[77][5]  ( .D(n8806), .CK(CLK), .RN(n12489), .Q(n14283), .QN(n10349) );
  DFFR_X1 \REGISTERS_reg[77][4]  ( .D(n8807), .CK(CLK), .RN(n12497), .Q(n14284), .QN(n10381) );
  DFFR_X1 \REGISTERS_reg[77][3]  ( .D(n8808), .CK(CLK), .RN(n12581), .Q(n14285), .QN(n10416) );
  DFFR_X1 \REGISTERS_reg[77][2]  ( .D(n8809), .CK(CLK), .RN(n12511), .Q(n14286), .QN(n10448) );
  DFFR_X1 \REGISTERS_reg[77][1]  ( .D(n8810), .CK(CLK), .RN(n12439), .Q(n14287), .QN(n10480) );
  DFFR_X1 \REGISTERS_reg[77][0]  ( .D(n8811), .CK(CLK), .RN(n12654), .Q(n14288), .QN(n10512) );
  DFFR_X1 \REGISTERS_reg[53][16]  ( .D(n8027), .CK(CLK), .RN(n12458), .Q(
        n13795), .QN(n929) );
  DFFR_X1 \REGISTERS_reg[53][15]  ( .D(n8028), .CK(CLK), .RN(n12637), .Q(
        n13796), .QN(n933) );
  DFFR_X1 \REGISTERS_reg[53][14]  ( .D(n8029), .CK(CLK), .RN(n12465), .Q(
        n13797), .QN(n937) );
  DFFR_X1 \REGISTERS_reg[53][13]  ( .D(n8030), .CK(CLK), .RN(n12473), .Q(
        n13798), .QN(n941) );
  DFFR_X1 \REGISTERS_reg[53][12]  ( .D(n8031), .CK(CLK), .RN(n12480), .Q(
        n13799), .QN(n945) );
  DFFR_X1 \REGISTERS_reg[53][11]  ( .D(n8032), .CK(CLK), .RN(n12571), .Q(
        n13800), .QN(n949) );
  DFFR_X1 \REGISTERS_reg[53][10]  ( .D(n8033), .CK(CLK), .RN(n12549), .Q(
        n13801), .QN(n953) );
  DFFR_X1 \REGISTERS_reg[53][9]  ( .D(n8034), .CK(CLK), .RN(n12557), .Q(n13802), .QN(n957) );
  DFFR_X1 \REGISTERS_reg[53][8]  ( .D(n8035), .CK(CLK), .RN(n12535), .Q(n13803), .QN(n961) );
  DFFR_X1 \REGISTERS_reg[53][7]  ( .D(n8036), .CK(CLK), .RN(n12645), .Q(n13804), .QN(n965) );
  DFFR_X1 \REGISTERS_reg[53][6]  ( .D(n8037), .CK(CLK), .RN(n12601), .Q(n13805), .QN(n969) );
  DFFR_X1 \REGISTERS_reg[53][5]  ( .D(n8038), .CK(CLK), .RN(n12487), .Q(n13806), .QN(n973) );
  DFFR_X1 \REGISTERS_reg[53][4]  ( .D(n8039), .CK(CLK), .RN(n12495), .Q(n13807), .QN(n977) );
  DFFR_X1 \REGISTERS_reg[53][3]  ( .D(n8040), .CK(CLK), .RN(n12579), .Q(n13808), .QN(n981) );
  DFFR_X1 \REGISTERS_reg[53][2]  ( .D(n8041), .CK(CLK), .RN(n12509), .Q(n13809), .QN(n985) );
  DFFR_X1 \REGISTERS_reg[53][1]  ( .D(n8042), .CK(CLK), .RN(n12437), .Q(n13810), .QN(n989) );
  DFFR_X1 \REGISTERS_reg[53][0]  ( .D(n8043), .CK(CLK), .RN(n12652), .Q(n13811), .QN(n993) );
  DFFR_X1 \REGISTERS_reg[52][31]  ( .D(n7980), .CK(CLK), .RN(n12659), .Q(
        n13748), .QN(n999) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n7334), .CK(CLK), .RN(n12485), .Q(n13358), .QN(n974) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n7335), .CK(CLK), .RN(n12493), .Q(n13359), .QN(n978) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n7336), .CK(CLK), .RN(n12577), .Q(n13360), .QN(n982) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n7337), .CK(CLK), .RN(n12507), .Q(n13361), .QN(n986) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n7338), .CK(CLK), .RN(n12435), .Q(n13362), .QN(n990) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n7339), .CK(CLK), .RN(n12650), .Q(n13363), .QN(n994) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n7020), .CK(CLK), .RN(n12657), .Q(
        n13044), .QN(n1868) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n7021), .CK(CLK), .RN(n12620), .Q(
        n13045), .QN(n1880) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n7022), .CK(CLK), .RN(n12605), .Q(
        n13046), .QN(n1892) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n7023), .CK(CLK), .RN(n12613), .Q(
        n13047), .QN(n1904) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n7024), .CK(CLK), .RN(n12583), .Q(
        n13048), .QN(n1916) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n7025), .CK(CLK), .RN(n12561), .Q(
        n13049), .QN(n1928) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n7026), .CK(CLK), .RN(n12539), .Q(
        n13050), .QN(n1940) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n7027), .CK(CLK), .RN(n12514), .Q(
        n13051), .QN(n1952) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n7028), .CK(CLK), .RN(n12627), .Q(
        n13052), .QN(n1964) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n7029), .CK(CLK), .RN(n12517), .Q(
        n13053), .QN(n1976) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n7030), .CK(CLK), .RN(n12525), .Q(
        n13054), .QN(n1988) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n7031), .CK(CLK), .RN(n12499), .Q(
        n13055), .QN(n2000) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n7032), .CK(CLK), .RN(n12591), .Q(
        n13056), .QN(n2012) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n7033), .CK(CLK), .RN(n12442), .Q(
        n13057), .QN(n2024) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n7034), .CK(CLK), .RN(n12449), .Q(
        n13058), .QN(n2036) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n7035), .CK(CLK), .RN(n12455), .Q(
        n13059), .QN(n2048) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n6988), .CK(CLK), .RN(n12657), .Q(
        n13012), .QN(n770) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n6989), .CK(CLK), .RN(n12620), .Q(
        n13013), .QN(n771) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n6990), .CK(CLK), .RN(n12605), .Q(
        n13014), .QN(n772) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n6991), .CK(CLK), .RN(n12613), .Q(
        n13015), .QN(n773) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n6992), .CK(CLK), .RN(n12583), .Q(
        n13016), .QN(n774) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n6993), .CK(CLK), .RN(n12561), .Q(
        n13017), .QN(n775) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n6994), .CK(CLK), .RN(n12539), .Q(
        n13018), .QN(n776) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n6995), .CK(CLK), .RN(n12514), .Q(
        n13019), .QN(n777) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n6996), .CK(CLK), .RN(n12627), .Q(
        n13020), .QN(n778) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n6997), .CK(CLK), .RN(n12517), .Q(
        n13021), .QN(n779) );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n6998), .CK(CLK), .RN(n12525), .Q(
        n13022), .QN(n780) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n6999), .CK(CLK), .RN(n12499), .Q(
        n13023), .QN(n781) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n7000), .CK(CLK), .RN(n12591), .Q(
        n13024), .QN(n782) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n7001), .CK(CLK), .RN(n12442), .Q(
        n13025), .QN(n783) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n7002), .CK(CLK), .RN(n12449), .Q(
        n13026), .QN(n784) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n7003), .CK(CLK), .RN(n12455), .Q(
        n13027), .QN(n785) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n7004), .CK(CLK), .RN(n12635), .Q(
        n13028), .QN(n786) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n7005), .CK(CLK), .RN(n12463), .Q(
        n13029), .QN(n787) );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n7006), .CK(CLK), .RN(n12470), .Q(
        n13030), .QN(n788) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n7007), .CK(CLK), .RN(n12477), .Q(
        n13031), .QN(n789) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n7008), .CK(CLK), .RN(n12569), .Q(
        n13032), .QN(n790) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n7009), .CK(CLK), .RN(n12547), .Q(
        n13033), .QN(n791) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n7010), .CK(CLK), .RN(n12554), .Q(n13034), .QN(n792) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n7011), .CK(CLK), .RN(n12532), .Q(n13035), .QN(n793) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n7012), .CK(CLK), .RN(n12642), .Q(n13036), .QN(n794) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n7013), .CK(CLK), .RN(n12598), .Q(n13037), .QN(n795) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n7014), .CK(CLK), .RN(n12485), .Q(n13038), .QN(n796) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n7015), .CK(CLK), .RN(n12492), .Q(n13039), .QN(n797) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n7016), .CK(CLK), .RN(n12576), .Q(n13040), .QN(n798) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n7017), .CK(CLK), .RN(n12507), .Q(n13041), .QN(n799) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n7018), .CK(CLK), .RN(n12434), .Q(n13042), .QN(n800) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n7019), .CK(CLK), .RN(n12649), .Q(n13043), .QN(n801) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n6956), .CK(CLK), .RN(n12657), .Q(
        n12980), .QN(n5738) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n6957), .CK(CLK), .RN(n12620), .Q(
        n12981), .QN(n5770) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n6958), .CK(CLK), .RN(n12605), .Q(
        n12982), .QN(n5802) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n6959), .CK(CLK), .RN(n12613), .Q(
        n12983), .QN(n5834) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n6960), .CK(CLK), .RN(n12583), .Q(
        n12984), .QN(n5866) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n6961), .CK(CLK), .RN(n12561), .Q(
        n12985), .QN(n5898) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n6962), .CK(CLK), .RN(n12539), .Q(
        n12986), .QN(n5930) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n6963), .CK(CLK), .RN(n12514), .Q(
        n12987), .QN(n5994) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n6964), .CK(CLK), .RN(n12627), .Q(
        n12988), .QN(n6311) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n6965), .CK(CLK), .RN(n12517), .Q(
        n12989), .QN(n9161) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n6966), .CK(CLK), .RN(n12525), .Q(
        n12990), .QN(n9193) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n6967), .CK(CLK), .RN(n12499), .Q(
        n12991), .QN(n9257) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n6968), .CK(CLK), .RN(n12591), .Q(
        n12992), .QN(n9591) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n6969), .CK(CLK), .RN(n12442), .Q(
        n12993), .QN(n9623) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n6970), .CK(CLK), .RN(n12449), .Q(
        n12994), .QN(n9655) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n6971), .CK(CLK), .RN(n12455), .Q(
        n12995), .QN(n10017) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n6972), .CK(CLK), .RN(n12635), .Q(
        n12996), .QN(n10049) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n6973), .CK(CLK), .RN(n12463), .Q(
        n12997), .QN(n10081) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n6974), .CK(CLK), .RN(n12470), .Q(
        n12998), .QN(n10113) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n6975), .CK(CLK), .RN(n12477), .Q(
        n12999), .QN(n10145) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n6976), .CK(CLK), .RN(n12569), .Q(
        n13000), .QN(n10177) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n6977), .CK(CLK), .RN(n12547), .Q(
        n13001), .QN(n10211) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n6978), .CK(CLK), .RN(n12554), .Q(n13002), .QN(n10243) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n6979), .CK(CLK), .RN(n12532), .Q(n13003), .QN(n10275) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n6980), .CK(CLK), .RN(n12642), .Q(n13004), .QN(n10310) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n6981), .CK(CLK), .RN(n12598), .Q(n13005), .QN(n10342) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n6982), .CK(CLK), .RN(n12485), .Q(n13006), .QN(n10374) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n6983), .CK(CLK), .RN(n12492), .Q(n13007), .QN(n10409) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n6984), .CK(CLK), .RN(n12576), .Q(n13008), .QN(n10441) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n6985), .CK(CLK), .RN(n12507), .Q(n13009), .QN(n10473) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n6986), .CK(CLK), .RN(n12434), .Q(n13010), .QN(n10505) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n6987), .CK(CLK), .RN(n12649), .Q(n13011), .QN(n10537) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n6924), .CK(CLK), .RN(n12656), .Q(
        n12948), .QN(n706) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n6925), .CK(CLK), .RN(n12620), .Q(
        n12949), .QN(n707) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n6926), .CK(CLK), .RN(n12605), .Q(
        n12950), .QN(n708) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n6927), .CK(CLK), .RN(n12612), .Q(
        n12951), .QN(n709) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n6928), .CK(CLK), .RN(n12583), .Q(
        n12952), .QN(n710) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n6929), .CK(CLK), .RN(n12561), .Q(
        n12953), .QN(n711) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n6930), .CK(CLK), .RN(n12539), .Q(
        n12954), .QN(n712) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n6931), .CK(CLK), .RN(n12514), .Q(
        n12955), .QN(n713) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n6932), .CK(CLK), .RN(n12627), .Q(
        n12956), .QN(n714) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n6933), .CK(CLK), .RN(n12517), .Q(
        n12957), .QN(n715) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n6934), .CK(CLK), .RN(n12524), .Q(
        n12958), .QN(n716) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n6935), .CK(CLK), .RN(n12499), .Q(
        n12959), .QN(n717) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n6936), .CK(CLK), .RN(n12590), .Q(
        n12960), .QN(n718) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n6937), .CK(CLK), .RN(n12441), .Q(
        n12961), .QN(n719) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n6938), .CK(CLK), .RN(n12449), .Q(
        n12962), .QN(n720) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n6939), .CK(CLK), .RN(n12455), .Q(
        n12963), .QN(n721) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n6940), .CK(CLK), .RN(n12634), .Q(
        n12964), .QN(n722) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n6941), .CK(CLK), .RN(n12462), .Q(
        n12965), .QN(n723) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n6942), .CK(CLK), .RN(n12470), .Q(
        n12966), .QN(n724) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n6943), .CK(CLK), .RN(n12477), .Q(
        n12967), .QN(n725) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n6944), .CK(CLK), .RN(n12568), .Q(
        n12968), .QN(n726) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n6945), .CK(CLK), .RN(n12546), .Q(
        n12969), .QN(n727) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n6946), .CK(CLK), .RN(n12554), .Q(n12970), .QN(n728) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n6947), .CK(CLK), .RN(n12532), .Q(n12971), .QN(n729) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n6948), .CK(CLK), .RN(n12642), .Q(n12972), .QN(n730) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n6949), .CK(CLK), .RN(n12598), .Q(n12973), .QN(n731) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n6950), .CK(CLK), .RN(n12484), .Q(n12974), .QN(n732) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n6951), .CK(CLK), .RN(n12492), .Q(n12975), .QN(n733) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n6952), .CK(CLK), .RN(n12576), .Q(n12976), .QN(n734) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n6953), .CK(CLK), .RN(n12506), .Q(n12977), .QN(n735) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n6954), .CK(CLK), .RN(n12434), .Q(n12978), .QN(n736) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n6955), .CK(CLK), .RN(n12649), .Q(n12979), .QN(n737) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n6892), .CK(CLK), .RN(n12656), .Q(
        n12916), .QN(n5732) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n6893), .CK(CLK), .RN(n12620), .Q(
        n12917), .QN(n5764) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n6894), .CK(CLK), .RN(n12605), .Q(
        n12918), .QN(n5796) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n6895), .CK(CLK), .RN(n12612), .Q(
        n12919), .QN(n5828) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n6896), .CK(CLK), .RN(n12583), .Q(
        n12920), .QN(n5860) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n6897), .CK(CLK), .RN(n12561), .Q(
        n12921), .QN(n5892) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n6898), .CK(CLK), .RN(n12539), .Q(
        n12922), .QN(n5924) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n6899), .CK(CLK), .RN(n12514), .Q(
        n12923), .QN(n5988) );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n6900), .CK(CLK), .RN(n12627), .Q(
        n12924), .QN(n6305) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n6901), .CK(CLK), .RN(n12517), .Q(
        n12925), .QN(n9155) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n6902), .CK(CLK), .RN(n12524), .Q(
        n12926), .QN(n9187) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n6903), .CK(CLK), .RN(n12499), .Q(
        n12927), .QN(n9251) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n6904), .CK(CLK), .RN(n12590), .Q(
        n12928), .QN(n9585) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n6905), .CK(CLK), .RN(n12441), .Q(
        n12929), .QN(n9617) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n6906), .CK(CLK), .RN(n12449), .Q(
        n12930), .QN(n9649) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n6907), .CK(CLK), .RN(n12455), .Q(
        n12931), .QN(n10011) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n6908), .CK(CLK), .RN(n12634), .Q(
        n12932), .QN(n10043) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n6909), .CK(CLK), .RN(n12462), .Q(
        n12933), .QN(n10075) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n6910), .CK(CLK), .RN(n12470), .Q(
        n12934), .QN(n10107) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n6911), .CK(CLK), .RN(n12477), .Q(
        n12935), .QN(n10139) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n6912), .CK(CLK), .RN(n12568), .Q(
        n12936), .QN(n10171) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n6913), .CK(CLK), .RN(n12546), .Q(
        n12937), .QN(n10203) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n6914), .CK(CLK), .RN(n12554), .Q(n12938), .QN(n10237) );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n6915), .CK(CLK), .RN(n12532), .Q(n12939), .QN(n10269) );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n6916), .CK(CLK), .RN(n12642), .Q(n12940), .QN(n10304) );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n6917), .CK(CLK), .RN(n12598), .Q(n12941), .QN(n10336) );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n6918), .CK(CLK), .RN(n12484), .Q(n12942), .QN(n10368) );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n6919), .CK(CLK), .RN(n12492), .Q(n12943), .QN(n10403) );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n6920), .CK(CLK), .RN(n12576), .Q(n12944), .QN(n10435) );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n6921), .CK(CLK), .RN(n12506), .Q(n12945), .QN(n10467) );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n6922), .CK(CLK), .RN(n12434), .Q(n12946), .QN(n10499) );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n6923), .CK(CLK), .RN(n12649), .Q(n12947), .QN(n10531) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n6860), .CK(CLK), .RN(n12656), .Q(
        n12884), .QN(n642) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n6861), .CK(CLK), .RN(n12620), .Q(
        n12885), .QN(n643) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n6862), .CK(CLK), .RN(n12605), .Q(
        n12886), .QN(n644) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n6863), .CK(CLK), .RN(n12612), .Q(
        n12887), .QN(n645) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n6864), .CK(CLK), .RN(n12583), .Q(
        n12888), .QN(n646) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n6865), .CK(CLK), .RN(n12561), .Q(
        n12889), .QN(n647) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n6866), .CK(CLK), .RN(n12539), .Q(
        n12890), .QN(n648) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n6867), .CK(CLK), .RN(n12514), .Q(
        n12891), .QN(n649) );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n6868), .CK(CLK), .RN(n12627), .Q(
        n12892), .QN(n650) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n6869), .CK(CLK), .RN(n12517), .Q(
        n12893), .QN(n651) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n6870), .CK(CLK), .RN(n12524), .Q(
        n12894), .QN(n652) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n6871), .CK(CLK), .RN(n12499), .Q(
        n12895), .QN(n653) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n6872), .CK(CLK), .RN(n12590), .Q(
        n12896), .QN(n654) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n6873), .CK(CLK), .RN(n12441), .Q(
        n12897), .QN(n655) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n6874), .CK(CLK), .RN(n12449), .Q(
        n12898), .QN(n656) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n6875), .CK(CLK), .RN(n12455), .Q(
        n12899), .QN(n657) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n6876), .CK(CLK), .RN(n12634), .Q(
        n12900), .QN(n658) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n6877), .CK(CLK), .RN(n12462), .Q(
        n12901), .QN(n659) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n6878), .CK(CLK), .RN(n12470), .Q(
        n12902), .QN(n660) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n6879), .CK(CLK), .RN(n12477), .Q(
        n12903), .QN(n661) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n6880), .CK(CLK), .RN(n12568), .Q(
        n12904), .QN(n662) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n6881), .CK(CLK), .RN(n12546), .Q(
        n12905), .QN(n663) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n6882), .CK(CLK), .RN(n12554), .Q(n12906), .QN(n664) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n6883), .CK(CLK), .RN(n12532), .Q(n12907), .QN(n665) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n6884), .CK(CLK), .RN(n12642), .Q(n12908), .QN(n666) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n6885), .CK(CLK), .RN(n12598), .Q(n12909), .QN(n667) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n6886), .CK(CLK), .RN(n12484), .Q(n12910), .QN(n668) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n6887), .CK(CLK), .RN(n12492), .Q(n12911), .QN(n669) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n6888), .CK(CLK), .RN(n12576), .Q(n12912), .QN(n670) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n6889), .CK(CLK), .RN(n12506), .Q(n12913), .QN(n671) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n6890), .CK(CLK), .RN(n12434), .Q(n12914), .QN(n672) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n6891), .CK(CLK), .RN(n12649), .Q(n12915), .QN(n673) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n6828), .CK(CLK), .RN(n12656), .Q(
        n12852), .QN(n5731) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n6829), .CK(CLK), .RN(n12620), .Q(
        n12853), .QN(n5763) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n6830), .CK(CLK), .RN(n12605), .Q(
        n12854), .QN(n5795) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n6831), .CK(CLK), .RN(n12612), .Q(
        n12855), .QN(n5827) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n6832), .CK(CLK), .RN(n12583), .Q(
        n12856), .QN(n5859) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n6833), .CK(CLK), .RN(n12561), .Q(
        n12857), .QN(n5891) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n6834), .CK(CLK), .RN(n12539), .Q(
        n12858), .QN(n5923) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n6835), .CK(CLK), .RN(n12514), .Q(
        n12859), .QN(n5987) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n6836), .CK(CLK), .RN(n12627), .Q(
        n12860), .QN(n6304) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n6837), .CK(CLK), .RN(n12517), .Q(
        n12861), .QN(n9154) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n6838), .CK(CLK), .RN(n12524), .Q(
        n12862), .QN(n9186) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n6839), .CK(CLK), .RN(n12499), .Q(
        n12863), .QN(n9250) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n6840), .CK(CLK), .RN(n12590), .Q(
        n12864), .QN(n9584) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n6841), .CK(CLK), .RN(n12441), .Q(
        n12865), .QN(n9616) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n6842), .CK(CLK), .RN(n12449), .Q(
        n12866), .QN(n9648) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n6843), .CK(CLK), .RN(n12455), .Q(
        n12867), .QN(n10010) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n6844), .CK(CLK), .RN(n12634), .Q(
        n12868), .QN(n10042) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n6845), .CK(CLK), .RN(n12462), .Q(
        n12869), .QN(n10074) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n6846), .CK(CLK), .RN(n12470), .Q(
        n12870), .QN(n10106) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n6847), .CK(CLK), .RN(n12477), .Q(
        n12871), .QN(n10138) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n6848), .CK(CLK), .RN(n12568), .Q(
        n12872), .QN(n10170) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n6849), .CK(CLK), .RN(n12546), .Q(
        n12873), .QN(n10202) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n6850), .CK(CLK), .RN(n12554), .Q(n12874), .QN(n10236) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n6851), .CK(CLK), .RN(n12532), .Q(n12875), .QN(n10268) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n6852), .CK(CLK), .RN(n12642), .Q(n12876), .QN(n10300) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n6853), .CK(CLK), .RN(n12598), .Q(n12877), .QN(n10335) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n6854), .CK(CLK), .RN(n12484), .Q(n12878), .QN(n10367) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n6855), .CK(CLK), .RN(n12492), .Q(n12879), .QN(n10402) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n6856), .CK(CLK), .RN(n12576), .Q(n12880), .QN(n10434) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n6857), .CK(CLK), .RN(n12506), .Q(n12881), .QN(n10466) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n6858), .CK(CLK), .RN(n12434), .Q(n12882), .QN(n10498) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n6859), .CK(CLK), .RN(n12649), .Q(n12883), .QN(n10530) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n6796), .CK(CLK), .RN(n12656), .Q(
        n12820), .QN(n5733) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n6797), .CK(CLK), .RN(n12619), .Q(
        n12821), .QN(n5765) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n6798), .CK(CLK), .RN(n12605), .Q(
        n12822), .QN(n5797) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n6799), .CK(CLK), .RN(n12612), .Q(
        n12823), .QN(n5829) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n6800), .CK(CLK), .RN(n12583), .Q(
        n12824), .QN(n5861) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n6801), .CK(CLK), .RN(n12561), .Q(
        n12825), .QN(n5893) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n6802), .CK(CLK), .RN(n12539), .Q(
        n12826), .QN(n5925) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n6803), .CK(CLK), .RN(n12513), .Q(
        n12827), .QN(n5989) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n6804), .CK(CLK), .RN(n12627), .Q(
        n12828), .QN(n6306) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n6805), .CK(CLK), .RN(n12517), .Q(
        n12829), .QN(n9156) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n6806), .CK(CLK), .RN(n12524), .Q(
        n12830), .QN(n9188) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n6807), .CK(CLK), .RN(n12499), .Q(
        n12831), .QN(n9252) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n6808), .CK(CLK), .RN(n12590), .Q(
        n12832), .QN(n9586) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n6809), .CK(CLK), .RN(n12441), .Q(
        n12833), .QN(n9618) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n6810), .CK(CLK), .RN(n12448), .Q(
        n12834), .QN(n9650) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n6811), .CK(CLK), .RN(n12455), .Q(
        n12835), .QN(n10012) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n6812), .CK(CLK), .RN(n12634), .Q(
        n12836), .QN(n10044) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n6813), .CK(CLK), .RN(n12462), .Q(
        n12837), .QN(n10076) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n6814), .CK(CLK), .RN(n12469), .Q(
        n12838), .QN(n10108) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n6815), .CK(CLK), .RN(n12477), .Q(
        n12839), .QN(n10140) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n6816), .CK(CLK), .RN(n12568), .Q(
        n12840), .QN(n10172) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n6817), .CK(CLK), .RN(n12546), .Q(
        n12841), .QN(n10204) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n6818), .CK(CLK), .RN(n12553), .Q(n12842), .QN(n10238) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n6819), .CK(CLK), .RN(n12531), .Q(n12843), .QN(n10270) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n6820), .CK(CLK), .RN(n12641), .Q(n12844), .QN(n10305) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n6821), .CK(CLK), .RN(n12597), .Q(n12845), .QN(n10337) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n6822), .CK(CLK), .RN(n12484), .Q(n12846), .QN(n10369) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n6823), .CK(CLK), .RN(n12491), .Q(n12847), .QN(n10404) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n6824), .CK(CLK), .RN(n12575), .Q(n12848), .QN(n10436) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n6825), .CK(CLK), .RN(n12506), .Q(n12849), .QN(n10468) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n6826), .CK(CLK), .RN(n12434), .Q(n12850), .QN(n10500) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n6827), .CK(CLK), .RN(n12649), .Q(n12851), .QN(n10532) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n6668), .CK(CLK), .RN(n12656), .Q(
        n12788), .QN(n5737) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n6669), .CK(CLK), .RN(n12619), .Q(
        n12789), .QN(n5769) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n6670), .CK(CLK), .RN(n12604), .Q(
        n12790), .QN(n5801) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n6671), .CK(CLK), .RN(n12612), .Q(
        n12791), .QN(n5833) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n6672), .CK(CLK), .RN(n12582), .Q(
        n12792), .QN(n5865) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n6673), .CK(CLK), .RN(n12560), .Q(
        n12793), .QN(n5897) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n6674), .CK(CLK), .RN(n12538), .Q(
        n12794), .QN(n5929) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n6675), .CK(CLK), .RN(n12513), .Q(
        n12795), .QN(n5993) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n6676), .CK(CLK), .RN(n12626), .Q(
        n12796), .QN(n6310) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n6677), .CK(CLK), .RN(n12469), .Q(
        n12797), .QN(n9160) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n6678), .CK(CLK), .RN(n12524), .Q(
        n12798), .QN(n9192) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n6679), .CK(CLK), .RN(n12498), .Q(
        n12799), .QN(n9256) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n6680), .CK(CLK), .RN(n12590), .Q(
        n12800), .QN(n9590) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n6681), .CK(CLK), .RN(n12441), .Q(
        n12801), .QN(n9622) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n6682), .CK(CLK), .RN(n12448), .Q(
        n12802), .QN(n9654) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n6683), .CK(CLK), .RN(n12489), .Q(
        n12803), .QN(n10016) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n6684), .CK(CLK), .RN(n12634), .Q(
        n12804), .QN(n10048) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n6685), .CK(CLK), .RN(n12462), .Q(
        n12805), .QN(n10080) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n6686), .CK(CLK), .RN(n12469), .Q(
        n12806), .QN(n10112) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n6687), .CK(CLK), .RN(n12476), .Q(
        n12807), .QN(n10144) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n6688), .CK(CLK), .RN(n12568), .Q(
        n12808), .QN(n10176) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n6689), .CK(CLK), .RN(n12546), .Q(
        n12809), .QN(n10210) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n6690), .CK(CLK), .RN(n12553), .Q(n12810), .QN(n10242) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n6691), .CK(CLK), .RN(n12531), .Q(n12811), .QN(n10274) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n6692), .CK(CLK), .RN(n12641), .Q(n12812), .QN(n10309) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n6693), .CK(CLK), .RN(n12597), .Q(n12813), .QN(n10341) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n6694), .CK(CLK), .RN(n12484), .Q(n12814), .QN(n10373) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n6695), .CK(CLK), .RN(n12491), .Q(n12815), .QN(n10408) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n6696), .CK(CLK), .RN(n12575), .Q(n12816), .QN(n10440) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n6697), .CK(CLK), .RN(n12506), .Q(n12817), .QN(n10472) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n6698), .CK(CLK), .RN(n12433), .Q(n12818), .QN(n10504) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n6699), .CK(CLK), .RN(n12648), .Q(n12819), .QN(n10536) );
  DFFR_X1 \REGISTERS_reg[80][31]  ( .D(n8876), .CK(CLK), .RN(n12662), .QN(
        n5711) );
  DFFR_X1 \REGISTERS_reg[80][30]  ( .D(n8877), .CK(CLK), .RN(n12625), .QN(
        n5743) );
  DFFR_X1 \REGISTERS_reg[80][29]  ( .D(n8878), .CK(CLK), .RN(n12610), .QN(
        n5775) );
  DFFR_X1 \REGISTERS_reg[80][28]  ( .D(n8879), .CK(CLK), .RN(n12618), .QN(
        n5807) );
  DFFR_X1 \REGISTERS_reg[80][27]  ( .D(n8880), .CK(CLK), .RN(n12588), .QN(
        n5839) );
  DFFR_X1 \REGISTERS_reg[80][26]  ( .D(n8881), .CK(CLK), .RN(n12566), .QN(
        n5871) );
  DFFR_X1 \REGISTERS_reg[80][25]  ( .D(n8882), .CK(CLK), .RN(n12544), .QN(
        n5903) );
  DFFR_X1 \REGISTERS_reg[80][24]  ( .D(n8883), .CK(CLK), .RN(n12450), .QN(
        n5935) );
  DFFR_X1 \REGISTERS_reg[80][23]  ( .D(n8884), .CK(CLK), .RN(n12632), .QN(
        n5999) );
  DFFR_X1 \REGISTERS_reg[80][22]  ( .D(n8885), .CK(CLK), .RN(n12522), .QN(
        n9134) );
  DFFR_X1 \REGISTERS_reg[80][21]  ( .D(n8886), .CK(CLK), .RN(n12530), .QN(
        n9166) );
  DFFR_X1 \REGISTERS_reg[80][20]  ( .D(n8887), .CK(CLK), .RN(n12504), .QN(
        n9198) );
  DFFR_X1 \REGISTERS_reg[80][19]  ( .D(n8888), .CK(CLK), .RN(n12596), .QN(
        n9262) );
  DFFR_X1 \REGISTERS_reg[80][18]  ( .D(n8889), .CK(CLK), .RN(n12447), .QN(
        n9596) );
  DFFR_X1 \REGISTERS_reg[80][17]  ( .D(n8890), .CK(CLK), .RN(n12454), .QN(
        n9628) );
  DFFR_X1 \REGISTERS_reg[80][16]  ( .D(n8891), .CK(CLK), .RN(n12460), .QN(
        n9660) );
  DFFR_X1 \REGISTERS_reg[80][15]  ( .D(n8892), .CK(CLK), .RN(n12640), .QN(
        n10022) );
  DFFR_X1 \REGISTERS_reg[80][14]  ( .D(n8893), .CK(CLK), .RN(n12468), .QN(
        n10054) );
  DFFR_X1 \REGISTERS_reg[80][13]  ( .D(n8894), .CK(CLK), .RN(n12475), .QN(
        n10086) );
  DFFR_X1 \REGISTERS_reg[80][12]  ( .D(n8895), .CK(CLK), .RN(n12482), .QN(
        n10118) );
  DFFR_X1 \REGISTERS_reg[80][11]  ( .D(n8896), .CK(CLK), .RN(n12574), .QN(
        n10150) );
  DFFR_X1 \REGISTERS_reg[80][10]  ( .D(n8897), .CK(CLK), .RN(n12552), .QN(
        n10182) );
  DFFR_X1 \REGISTERS_reg[80][9]  ( .D(n8898), .CK(CLK), .RN(n12559), .QN(
        n10216) );
  DFFR_X1 \REGISTERS_reg[80][8]  ( .D(n8899), .CK(CLK), .RN(n12537), .QN(
        n10248) );
  DFFR_X1 \REGISTERS_reg[80][7]  ( .D(n8900), .CK(CLK), .RN(n12647), .QN(
        n10280) );
  XNOR2_X1 U3 ( .A(\U3/U98/Z_6 ), .B(\r480/n4 ), .ZN(N8437) );
  XNOR2_X1 U4 ( .A(\U3/U99/Z_6 ), .B(\r486/n4 ), .ZN(N8581) );
  AND2_X1 U5 ( .A1(n2574), .A2(n2491), .ZN(n10538) );
  AND2_X1 U6 ( .A1(n2574), .A2(n2494), .ZN(n10539) );
  AND2_X1 U7 ( .A1(n2574), .A2(n2496), .ZN(n10540) );
  AND2_X1 U8 ( .A1(n2574), .A2(n2498), .ZN(n10541) );
  AND2_X1 U9 ( .A1(n2574), .A2(n2500), .ZN(n10542) );
  AND2_X1 U10 ( .A1(n2574), .A2(n2566), .ZN(n10543) );
  AND2_X1 U11 ( .A1(n2574), .A2(n2568), .ZN(n10544) );
  AND2_X1 U12 ( .A1(n2574), .A2(n2570), .ZN(n10545) );
  AND2_X1 U13 ( .A1(n2599), .A2(n2573), .ZN(n10546) );
  AND2_X1 U14 ( .A1(n2599), .A2(n2578), .ZN(n10547) );
  AND2_X1 U15 ( .A1(n2599), .A2(n2570), .ZN(n10548) );
  AND2_X1 U16 ( .A1(n2617), .A2(n2573), .ZN(n10549) );
  AND2_X1 U17 ( .A1(n2617), .A2(n2576), .ZN(n10550) );
  AND2_X1 U18 ( .A1(n2617), .A2(n2582), .ZN(n10551) );
  AND2_X1 U19 ( .A1(n2617), .A2(n2586), .ZN(n10552) );
  AND2_X1 U20 ( .A1(n2617), .A2(n2491), .ZN(n10553) );
  AND2_X1 U21 ( .A1(n2698), .A2(n2584), .ZN(n10554) );
  AND2_X1 U22 ( .A1(n2698), .A2(n2586), .ZN(n10555) );
  AND2_X1 U23 ( .A1(n2698), .A2(n2588), .ZN(n10556) );
  AND2_X1 U24 ( .A1(n2599), .A2(n2582), .ZN(n10557) );
  AND2_X1 U25 ( .A1(n2599), .A2(n2588), .ZN(n10558) );
  AND2_X1 U26 ( .A1(n2617), .A2(n2496), .ZN(n10559) );
  AND2_X1 U27 ( .A1(n2617), .A2(n2566), .ZN(n10560) );
  AND2_X1 U28 ( .A1(n2715), .A2(n2580), .ZN(n10561) );
  AND2_X1 U29 ( .A1(n2715), .A2(n2588), .ZN(n10562) );
  AND2_X1 U30 ( .A1(n2715), .A2(n2496), .ZN(n10563) );
  AND2_X1 U31 ( .A1(n2715), .A2(n2566), .ZN(n10564) );
  AND2_X1 U32 ( .A1(n2599), .A2(n2580), .ZN(n10565) );
  AND2_X1 U33 ( .A1(n2599), .A2(n2586), .ZN(n10566) );
  AND2_X1 U34 ( .A1(n2617), .A2(n2494), .ZN(n10567) );
  AND2_X1 U35 ( .A1(n2617), .A2(n2500), .ZN(n10568) );
  AND2_X1 U36 ( .A1(n2715), .A2(n2578), .ZN(n10569) );
  AND2_X1 U37 ( .A1(n2715), .A2(n2584), .ZN(n10570) );
  AND2_X1 U38 ( .A1(n2715), .A2(n2491), .ZN(n10571) );
  AND2_X1 U39 ( .A1(n2715), .A2(n2498), .ZN(n10572) );
  AND2_X1 U40 ( .A1(n2599), .A2(n2576), .ZN(n10573) );
  AND2_X1 U41 ( .A1(n2599), .A2(n2584), .ZN(n10574) );
  AND2_X1 U42 ( .A1(n2617), .A2(n2588), .ZN(n10575) );
  AND2_X1 U43 ( .A1(n2617), .A2(n2498), .ZN(n10576) );
  AND2_X1 U44 ( .A1(n2715), .A2(n2576), .ZN(n10577) );
  AND2_X1 U45 ( .A1(n2715), .A2(n2586), .ZN(n10578) );
  AND2_X1 U46 ( .A1(n2715), .A2(n2494), .ZN(n10579) );
  AND2_X1 U47 ( .A1(n2715), .A2(n2500), .ZN(n10580) );
  AND2_X1 U48 ( .A1(n2599), .A2(n2491), .ZN(n10581) );
  AND2_X1 U49 ( .A1(n2617), .A2(n2568), .ZN(n10582) );
  AND2_X1 U50 ( .A1(n2715), .A2(n2568), .ZN(n10583) );
  AND2_X1 U51 ( .A1(n2617), .A2(n2584), .ZN(n10584) );
  AND2_X1 U52 ( .A1(n2715), .A2(n2570), .ZN(n10585) );
  AND2_X1 U53 ( .A1(n2599), .A2(n2496), .ZN(n10586) );
  AND2_X1 U54 ( .A1(n2698), .A2(n2496), .ZN(n10587) );
  AND2_X1 U55 ( .A1(n2698), .A2(n2498), .ZN(n10588) );
  AND2_X1 U56 ( .A1(n2698), .A2(n2500), .ZN(n10589) );
  AND2_X1 U57 ( .A1(n2698), .A2(n2566), .ZN(n10590) );
  AND2_X1 U58 ( .A1(n2698), .A2(n2568), .ZN(n10591) );
  AND2_X1 U59 ( .A1(n2698), .A2(n2570), .ZN(n10592) );
  AND2_X1 U60 ( .A1(n2715), .A2(n2573), .ZN(n10593) );
  AND2_X1 U61 ( .A1(n2715), .A2(n2582), .ZN(n10594) );
  AND2_X1 U62 ( .A1(n2599), .A2(n2494), .ZN(n10595) );
  AND2_X1 U63 ( .A1(n2599), .A2(n2498), .ZN(n10596) );
  AND2_X1 U64 ( .A1(n2599), .A2(n2500), .ZN(n10597) );
  AND2_X1 U65 ( .A1(n2599), .A2(n2566), .ZN(n10598) );
  AND2_X1 U66 ( .A1(n2599), .A2(n2568), .ZN(n10599) );
  AND2_X1 U67 ( .A1(n2617), .A2(n2578), .ZN(n10600) );
  AND2_X1 U68 ( .A1(n2617), .A2(n2580), .ZN(n10601) );
  AND2_X1 U69 ( .A1(n2617), .A2(n2570), .ZN(n10602) );
  AND2_X1 U70 ( .A1(n2698), .A2(n2573), .ZN(n10603) );
  AND2_X1 U71 ( .A1(n2698), .A2(n2576), .ZN(n10604) );
  AND2_X1 U72 ( .A1(n2698), .A2(n2578), .ZN(n10605) );
  AND2_X1 U73 ( .A1(n2698), .A2(n2580), .ZN(n10606) );
  AND2_X1 U74 ( .A1(n2698), .A2(n2582), .ZN(n10607) );
  AND2_X1 U75 ( .A1(n2698), .A2(n2491), .ZN(n10608) );
  AND2_X1 U76 ( .A1(n2698), .A2(n2494), .ZN(n10609) );
  AND2_X1 U77 ( .A1(n2580), .A2(n2574), .ZN(n10610) );
  AND2_X1 U78 ( .A1(n2584), .A2(n2574), .ZN(n10611) );
  AND2_X1 U79 ( .A1(n2586), .A2(n2574), .ZN(n10612) );
  AND2_X1 U80 ( .A1(n2588), .A2(n2574), .ZN(n10613) );
  AND2_X1 U81 ( .A1(n2576), .A2(n2574), .ZN(n10614) );
  AND2_X1 U82 ( .A1(n2573), .A2(n2574), .ZN(n10615) );
  AND2_X1 U83 ( .A1(n2582), .A2(n2574), .ZN(n10616) );
  AND2_X1 U84 ( .A1(n2578), .A2(n2574), .ZN(n10617) );
  AND2_X1 U85 ( .A1(n2570), .A2(n2492), .ZN(n10618) );
  AND2_X1 U86 ( .A1(n2494), .A2(n2492), .ZN(n10619) );
  AND2_X1 U87 ( .A1(n2496), .A2(n2492), .ZN(n10620) );
  AND2_X1 U88 ( .A1(n2498), .A2(n2492), .ZN(n10621) );
  AND2_X1 U89 ( .A1(n2500), .A2(n2492), .ZN(n10622) );
  AND2_X1 U90 ( .A1(n2566), .A2(n2492), .ZN(n10623) );
  AND2_X1 U91 ( .A1(n2568), .A2(n2492), .ZN(n10624) );
  NOR2_X1 U92 ( .A1(n12770), .A2(N8435), .ZN(n5675) );
  NOR2_X1 U93 ( .A1(n12774), .A2(N8579), .ZN(n4242) );
  AND3_X1 U94 ( .A1(n2615), .A2(N2171), .A3(N2172), .ZN(n2599) );
  AND3_X1 U95 ( .A1(N2171), .A2(n12732), .A3(n2615), .ZN(n2698) );
  INV_X1 U96 ( .A(n12290), .ZN(n12280) );
  INV_X1 U97 ( .A(n12290), .ZN(n12279) );
  INV_X1 U98 ( .A(n12242), .ZN(n12232) );
  INV_X1 U99 ( .A(n12242), .ZN(n12231) );
  INV_X1 U100 ( .A(n11906), .ZN(n11896) );
  INV_X1 U101 ( .A(n11906), .ZN(n11895) );
  INV_X1 U102 ( .A(n11858), .ZN(n11848) );
  INV_X1 U103 ( .A(n11858), .ZN(n11847) );
  INV_X1 U104 ( .A(n11522), .ZN(n11512) );
  INV_X1 U105 ( .A(n11522), .ZN(n11511) );
  INV_X1 U106 ( .A(n11474), .ZN(n11464) );
  INV_X1 U107 ( .A(n11474), .ZN(n11463) );
  INV_X1 U108 ( .A(n12415), .ZN(n12406) );
  INV_X1 U109 ( .A(n12415), .ZN(n12405) );
  INV_X1 U110 ( .A(n12404), .ZN(n12395) );
  INV_X1 U111 ( .A(n12404), .ZN(n12394) );
  INV_X1 U112 ( .A(n12393), .ZN(n12384) );
  INV_X1 U113 ( .A(n12393), .ZN(n12383) );
  INV_X1 U114 ( .A(n12382), .ZN(n12373) );
  INV_X1 U115 ( .A(n12382), .ZN(n12372) );
  INV_X1 U116 ( .A(n12371), .ZN(n12362) );
  INV_X1 U117 ( .A(n12371), .ZN(n12361) );
  INV_X1 U118 ( .A(n12360), .ZN(n12351) );
  INV_X1 U119 ( .A(n12360), .ZN(n12350) );
  INV_X1 U120 ( .A(n12349), .ZN(n12340) );
  INV_X1 U121 ( .A(n12349), .ZN(n12339) );
  INV_X1 U122 ( .A(n12338), .ZN(n12328) );
  INV_X1 U123 ( .A(n12338), .ZN(n12327) );
  INV_X1 U124 ( .A(n12326), .ZN(n12316) );
  INV_X1 U125 ( .A(n12326), .ZN(n12315) );
  INV_X1 U126 ( .A(n12314), .ZN(n12304) );
  INV_X1 U127 ( .A(n12314), .ZN(n12303) );
  INV_X1 U128 ( .A(n12302), .ZN(n12292) );
  INV_X1 U129 ( .A(n12302), .ZN(n12291) );
  INV_X1 U130 ( .A(n12278), .ZN(n12268) );
  INV_X1 U131 ( .A(n12278), .ZN(n12267) );
  INV_X1 U132 ( .A(n12266), .ZN(n12256) );
  INV_X1 U133 ( .A(n12266), .ZN(n12255) );
  INV_X1 U134 ( .A(n12254), .ZN(n12244) );
  INV_X1 U135 ( .A(n12254), .ZN(n12243) );
  INV_X1 U136 ( .A(n12230), .ZN(n12220) );
  INV_X1 U137 ( .A(n12230), .ZN(n12219) );
  INV_X1 U138 ( .A(n12218), .ZN(n12208) );
  INV_X1 U139 ( .A(n12218), .ZN(n12207) );
  INV_X1 U140 ( .A(n12206), .ZN(n12196) );
  INV_X1 U141 ( .A(n12206), .ZN(n12195) );
  INV_X1 U142 ( .A(n12194), .ZN(n12184) );
  INV_X1 U143 ( .A(n12194), .ZN(n12183) );
  INV_X1 U144 ( .A(n12182), .ZN(n12172) );
  INV_X1 U145 ( .A(n12182), .ZN(n12171) );
  INV_X1 U146 ( .A(n12170), .ZN(n12160) );
  INV_X1 U147 ( .A(n12170), .ZN(n12159) );
  INV_X1 U148 ( .A(n12158), .ZN(n12148) );
  INV_X1 U149 ( .A(n12158), .ZN(n12147) );
  INV_X1 U150 ( .A(n12146), .ZN(n12136) );
  INV_X1 U151 ( .A(n12146), .ZN(n12135) );
  INV_X1 U152 ( .A(n12134), .ZN(n12124) );
  INV_X1 U153 ( .A(n12134), .ZN(n12123) );
  INV_X1 U154 ( .A(n12122), .ZN(n12112) );
  INV_X1 U155 ( .A(n12122), .ZN(n12111) );
  INV_X1 U156 ( .A(n12110), .ZN(n12100) );
  INV_X1 U157 ( .A(n12110), .ZN(n12099) );
  INV_X1 U158 ( .A(n12098), .ZN(n12088) );
  INV_X1 U159 ( .A(n12098), .ZN(n12087) );
  INV_X1 U160 ( .A(n12086), .ZN(n12076) );
  INV_X1 U161 ( .A(n12086), .ZN(n12075) );
  INV_X1 U162 ( .A(n12074), .ZN(n12064) );
  INV_X1 U163 ( .A(n12074), .ZN(n12063) );
  INV_X1 U164 ( .A(n12062), .ZN(n12052) );
  INV_X1 U165 ( .A(n12062), .ZN(n12051) );
  INV_X1 U166 ( .A(n12050), .ZN(n12040) );
  INV_X1 U167 ( .A(n12050), .ZN(n12039) );
  INV_X1 U168 ( .A(n12038), .ZN(n12028) );
  INV_X1 U169 ( .A(n12038), .ZN(n12027) );
  INV_X1 U170 ( .A(n12026), .ZN(n12016) );
  INV_X1 U171 ( .A(n12026), .ZN(n12015) );
  INV_X1 U172 ( .A(n12014), .ZN(n12004) );
  INV_X1 U173 ( .A(n12014), .ZN(n12003) );
  INV_X1 U174 ( .A(n12002), .ZN(n11992) );
  INV_X1 U175 ( .A(n12002), .ZN(n11991) );
  INV_X1 U176 ( .A(n11990), .ZN(n11980) );
  INV_X1 U177 ( .A(n11990), .ZN(n11979) );
  INV_X1 U178 ( .A(n11978), .ZN(n11968) );
  INV_X1 U179 ( .A(n11978), .ZN(n11967) );
  INV_X1 U180 ( .A(n11966), .ZN(n11956) );
  INV_X1 U181 ( .A(n11966), .ZN(n11955) );
  INV_X1 U182 ( .A(n11954), .ZN(n11944) );
  INV_X1 U183 ( .A(n11954), .ZN(n11943) );
  INV_X1 U184 ( .A(n11942), .ZN(n11932) );
  INV_X1 U185 ( .A(n11942), .ZN(n11931) );
  INV_X1 U186 ( .A(n11930), .ZN(n11920) );
  INV_X1 U187 ( .A(n11930), .ZN(n11919) );
  INV_X1 U188 ( .A(n11918), .ZN(n11908) );
  INV_X1 U189 ( .A(n11918), .ZN(n11907) );
  INV_X1 U191 ( .A(n11894), .ZN(n11884) );
  INV_X1 U192 ( .A(n11894), .ZN(n11883) );
  INV_X1 U193 ( .A(n11882), .ZN(n11872) );
  INV_X1 U194 ( .A(n11882), .ZN(n11871) );
  INV_X1 U195 ( .A(n11870), .ZN(n11860) );
  INV_X1 U196 ( .A(n11870), .ZN(n11859) );
  INV_X1 U197 ( .A(n11846), .ZN(n11836) );
  INV_X1 U198 ( .A(n11846), .ZN(n11835) );
  INV_X1 U199 ( .A(n11834), .ZN(n11824) );
  INV_X1 U200 ( .A(n11834), .ZN(n11823) );
  INV_X1 U201 ( .A(n11822), .ZN(n11812) );
  INV_X1 U202 ( .A(n11822), .ZN(n11811) );
  INV_X1 U203 ( .A(n11810), .ZN(n11800) );
  INV_X1 U204 ( .A(n11810), .ZN(n11799) );
  INV_X1 U205 ( .A(n11798), .ZN(n11788) );
  INV_X1 U206 ( .A(n11798), .ZN(n11787) );
  INV_X1 U207 ( .A(n11786), .ZN(n11776) );
  INV_X1 U208 ( .A(n11786), .ZN(n11775) );
  INV_X1 U209 ( .A(n11774), .ZN(n11764) );
  INV_X1 U210 ( .A(n11774), .ZN(n11763) );
  INV_X1 U211 ( .A(n11762), .ZN(n11752) );
  INV_X1 U212 ( .A(n11762), .ZN(n11751) );
  INV_X1 U213 ( .A(n11750), .ZN(n11740) );
  INV_X1 U214 ( .A(n11750), .ZN(n11739) );
  INV_X1 U215 ( .A(n11738), .ZN(n11728) );
  INV_X1 U216 ( .A(n11738), .ZN(n11727) );
  INV_X1 U217 ( .A(n11726), .ZN(n11716) );
  INV_X1 U218 ( .A(n11726), .ZN(n11715) );
  INV_X1 U219 ( .A(n11714), .ZN(n11704) );
  INV_X1 U220 ( .A(n11714), .ZN(n11703) );
  INV_X1 U221 ( .A(n11702), .ZN(n11692) );
  INV_X1 U222 ( .A(n11702), .ZN(n11691) );
  INV_X1 U223 ( .A(n11690), .ZN(n11680) );
  INV_X1 U225 ( .A(n11690), .ZN(n11679) );
  INV_X1 U226 ( .A(n11678), .ZN(n11668) );
  INV_X1 U227 ( .A(n11678), .ZN(n11667) );
  INV_X1 U228 ( .A(n11666), .ZN(n11656) );
  INV_X1 U229 ( .A(n11666), .ZN(n11655) );
  INV_X1 U230 ( .A(n11654), .ZN(n11644) );
  INV_X1 U231 ( .A(n11654), .ZN(n11643) );
  INV_X1 U232 ( .A(n11642), .ZN(n11632) );
  INV_X1 U233 ( .A(n11642), .ZN(n11631) );
  INV_X1 U234 ( .A(n11630), .ZN(n11620) );
  INV_X1 U235 ( .A(n11630), .ZN(n11619) );
  INV_X1 U236 ( .A(n11618), .ZN(n11608) );
  INV_X1 U237 ( .A(n11618), .ZN(n11607) );
  INV_X1 U238 ( .A(n11606), .ZN(n11596) );
  INV_X1 U239 ( .A(n11606), .ZN(n11595) );
  INV_X1 U240 ( .A(n11594), .ZN(n11584) );
  INV_X1 U241 ( .A(n11594), .ZN(n11583) );
  INV_X1 U242 ( .A(n11582), .ZN(n11572) );
  INV_X1 U243 ( .A(n11582), .ZN(n11571) );
  INV_X1 U244 ( .A(n11570), .ZN(n11560) );
  INV_X1 U245 ( .A(n11570), .ZN(n11559) );
  INV_X1 U246 ( .A(n11558), .ZN(n11548) );
  INV_X1 U247 ( .A(n11558), .ZN(n11547) );
  INV_X1 U248 ( .A(n11546), .ZN(n11536) );
  INV_X1 U249 ( .A(n11546), .ZN(n11535) );
  INV_X1 U250 ( .A(n11534), .ZN(n11524) );
  INV_X1 U251 ( .A(n11534), .ZN(n11523) );
  INV_X1 U252 ( .A(n11510), .ZN(n11500) );
  INV_X1 U253 ( .A(n11510), .ZN(n11499) );
  INV_X1 U254 ( .A(n11498), .ZN(n11488) );
  INV_X1 U255 ( .A(n11498), .ZN(n11487) );
  INV_X1 U256 ( .A(n11486), .ZN(n11476) );
  INV_X1 U257 ( .A(n11486), .ZN(n11475) );
  INV_X1 U258 ( .A(n11462), .ZN(n11452) );
  INV_X1 U259 ( .A(n11462), .ZN(n11451) );
  INV_X1 U260 ( .A(n11450), .ZN(n11440) );
  INV_X1 U261 ( .A(n11450), .ZN(n11439) );
  INV_X1 U262 ( .A(n11438), .ZN(n11428) );
  INV_X1 U263 ( .A(n11438), .ZN(n11427) );
  INV_X1 U264 ( .A(n11426), .ZN(n11416) );
  INV_X1 U265 ( .A(n11426), .ZN(n11415) );
  INV_X1 U266 ( .A(n11414), .ZN(n11404) );
  INV_X1 U267 ( .A(n11414), .ZN(n11403) );
  INV_X1 U268 ( .A(n11402), .ZN(n11392) );
  INV_X1 U269 ( .A(n11402), .ZN(n11391) );
  INV_X1 U270 ( .A(n11390), .ZN(n11380) );
  INV_X1 U271 ( .A(n11390), .ZN(n11379) );
  BUF_X1 U272 ( .A(n10594), .Z(n11514) );
  BUF_X1 U273 ( .A(n10594), .Z(n11515) );
  BUF_X1 U274 ( .A(n10594), .Z(n11516) );
  BUF_X1 U275 ( .A(n10594), .Z(n11517) );
  BUF_X1 U276 ( .A(n11522), .Z(n11518) );
  BUF_X1 U277 ( .A(n11520), .Z(n11519) );
  BUF_X1 U278 ( .A(n10594), .Z(n11520) );
  BUF_X1 U279 ( .A(n11522), .Z(n11521) );
  BUF_X1 U280 ( .A(n10571), .Z(n11466) );
  BUF_X1 U281 ( .A(n10571), .Z(n11467) );
  BUF_X1 U282 ( .A(n10571), .Z(n11468) );
  BUF_X1 U283 ( .A(n10571), .Z(n11469) );
  BUF_X1 U284 ( .A(n11474), .Z(n11470) );
  BUF_X1 U285 ( .A(n11472), .Z(n11471) );
  BUF_X1 U286 ( .A(n10571), .Z(n11472) );
  BUF_X1 U287 ( .A(n11474), .Z(n11473) );
  BUF_X1 U288 ( .A(n10616), .Z(n12282) );
  BUF_X1 U289 ( .A(n10616), .Z(n12283) );
  BUF_X1 U290 ( .A(n10616), .Z(n12284) );
  BUF_X1 U291 ( .A(n10616), .Z(n12285) );
  BUF_X1 U292 ( .A(n12290), .Z(n12286) );
  BUF_X1 U293 ( .A(n12288), .Z(n12287) );
  BUF_X1 U294 ( .A(n10616), .Z(n12288) );
  BUF_X1 U295 ( .A(n12290), .Z(n12289) );
  BUF_X1 U296 ( .A(n10538), .Z(n12234) );
  BUF_X1 U297 ( .A(n10538), .Z(n12235) );
  BUF_X1 U298 ( .A(n10538), .Z(n12236) );
  BUF_X1 U299 ( .A(n10538), .Z(n12237) );
  BUF_X1 U300 ( .A(n10538), .Z(n12238) );
  BUF_X1 U301 ( .A(n10538), .Z(n12239) );
  BUF_X1 U302 ( .A(n12234), .Z(n12240) );
  BUF_X1 U303 ( .A(n12236), .Z(n12241) );
  BUF_X1 U304 ( .A(n10551), .Z(n11898) );
  BUF_X1 U305 ( .A(n10551), .Z(n11899) );
  BUF_X1 U338 ( .A(n10551), .Z(n11900) );
  BUF_X1 U339 ( .A(n10551), .Z(n11901) );
  BUF_X1 U340 ( .A(n11906), .Z(n11902) );
  BUF_X1 U341 ( .A(n11904), .Z(n11903) );
  BUF_X1 U342 ( .A(n10551), .Z(n11904) );
  BUF_X1 U343 ( .A(n11906), .Z(n11905) );
  BUF_X1 U344 ( .A(n10553), .Z(n11850) );
  BUF_X1 U345 ( .A(n10553), .Z(n11851) );
  BUF_X1 U346 ( .A(n10553), .Z(n11852) );
  BUF_X1 U347 ( .A(n10553), .Z(n11853) );
  BUF_X1 U348 ( .A(n11858), .Z(n11854) );
  BUF_X1 U349 ( .A(n11856), .Z(n11855) );
  BUF_X1 U350 ( .A(n10553), .Z(n11856) );
  BUF_X1 U351 ( .A(n11858), .Z(n11857) );
  BUF_X1 U352 ( .A(n12237), .Z(n12242) );
  BUF_X1 U353 ( .A(n10551), .Z(n11906) );
  BUF_X1 U354 ( .A(n10553), .Z(n11858) );
  BUF_X1 U355 ( .A(n10594), .Z(n11522) );
  BUF_X1 U356 ( .A(n10571), .Z(n11474) );
  BUF_X1 U357 ( .A(n10616), .Z(n12290) );
  INV_X1 U358 ( .A(n12425), .ZN(n12417) );
  INV_X1 U359 ( .A(n12425), .ZN(n12416) );
  BUF_X1 U360 ( .A(n12714), .Z(n12708) );
  BUF_X1 U361 ( .A(n12713), .Z(n12711) );
  BUF_X1 U362 ( .A(n12722), .Z(n12685) );
  BUF_X1 U363 ( .A(n12719), .Z(n12693) );
  BUF_X1 U364 ( .A(n12723), .Z(n12680) );
  BUF_X1 U365 ( .A(n12716), .Z(n12703) );
  BUF_X1 U366 ( .A(n12723), .Z(n12682) );
  BUF_X1 U367 ( .A(n12722), .Z(n12683) );
  BUF_X1 U368 ( .A(n12717), .Z(n12700) );
  BUF_X1 U369 ( .A(n12719), .Z(n12694) );
  BUF_X1 U370 ( .A(n12715), .Z(n12706) );
  BUF_X1 U371 ( .A(n12714), .Z(n12707) );
  BUF_X1 U372 ( .A(n12715), .Z(n12704) );
  BUF_X1 U373 ( .A(n12722), .Z(n12684) );
  BUF_X1 U374 ( .A(n12721), .Z(n12686) );
  BUF_X1 U375 ( .A(n12721), .Z(n12687) );
  BUF_X1 U376 ( .A(n12718), .Z(n12695) );
  BUF_X1 U377 ( .A(n12721), .Z(n12688) );
  BUF_X1 U378 ( .A(n12720), .Z(n12689) );
  BUF_X1 U379 ( .A(n12720), .Z(n12690) );
  BUF_X1 U380 ( .A(n12716), .Z(n12701) );
  BUF_X1 U381 ( .A(n12723), .Z(n12681) );
  BUF_X1 U382 ( .A(n12713), .Z(n12710) );
  BUF_X1 U383 ( .A(n12718), .Z(n12696) );
  BUF_X1 U384 ( .A(n12724), .Z(n12679) );
  BUF_X1 U385 ( .A(n12714), .Z(n12709) );
  BUF_X1 U386 ( .A(n12715), .Z(n12705) );
  BUF_X1 U387 ( .A(n12716), .Z(n12702) );
  BUF_X1 U388 ( .A(n12717), .Z(n12698) );
  BUF_X1 U389 ( .A(n12717), .Z(n12699) );
  BUF_X1 U390 ( .A(n12718), .Z(n12697) );
  BUF_X1 U391 ( .A(n12719), .Z(n12692) );
  BUF_X1 U392 ( .A(n12720), .Z(n12691) );
  BUF_X1 U393 ( .A(n12726), .Z(n12672) );
  BUF_X1 U394 ( .A(n12726), .Z(n12673) );
  BUF_X1 U395 ( .A(n12728), .Z(n12665) );
  BUF_X1 U396 ( .A(n12725), .Z(n12674) );
  BUF_X1 U397 ( .A(n12728), .Z(n12666) );
  BUF_X1 U398 ( .A(n12725), .Z(n12675) );
  BUF_X1 U399 ( .A(n12728), .Z(n12667) );
  BUF_X1 U400 ( .A(n12725), .Z(n12676) );
  BUF_X1 U401 ( .A(n12727), .Z(n12668) );
  BUF_X1 U402 ( .A(n12724), .Z(n12677) );
  BUF_X1 U403 ( .A(n12727), .Z(n12669) );
  BUF_X1 U404 ( .A(n12724), .Z(n12678) );
  BUF_X1 U405 ( .A(n12727), .Z(n12670) );
  BUF_X1 U406 ( .A(n12726), .Z(n12671) );
  BUF_X1 U407 ( .A(n12729), .Z(n12663) );
  BUF_X1 U408 ( .A(n12729), .Z(n12664) );
  BUF_X1 U409 ( .A(n10545), .Z(n12150) );
  BUF_X1 U410 ( .A(n10545), .Z(n12151) );
  BUF_X1 U411 ( .A(n10545), .Z(n12152) );
  BUF_X1 U412 ( .A(n10545), .Z(n12153) );
  BUF_X1 U413 ( .A(n12158), .Z(n12154) );
  BUF_X1 U414 ( .A(n12156), .Z(n12155) );
  BUF_X1 U415 ( .A(n10545), .Z(n12156) );
  BUF_X1 U416 ( .A(n12158), .Z(n12157) );
  BUF_X1 U417 ( .A(n10573), .Z(n12126) );
  BUF_X1 U418 ( .A(n10573), .Z(n12127) );
  BUF_X1 U419 ( .A(n10573), .Z(n12128) );
  BUF_X1 U420 ( .A(n10573), .Z(n12129) );
  BUF_X1 U421 ( .A(n12134), .Z(n12130) );
  BUF_X1 U422 ( .A(n12132), .Z(n12131) );
  BUF_X1 U423 ( .A(n10573), .Z(n12132) );
  BUF_X1 U424 ( .A(n12134), .Z(n12133) );
  BUF_X1 U425 ( .A(n10565), .Z(n12102) );
  BUF_X1 U426 ( .A(n10565), .Z(n12103) );
  BUF_X1 U427 ( .A(n10565), .Z(n12104) );
  BUF_X1 U428 ( .A(n10565), .Z(n12105) );
  BUF_X1 U429 ( .A(n12110), .Z(n12106) );
  BUF_X1 U430 ( .A(n12108), .Z(n12107) );
  BUF_X1 U431 ( .A(n10565), .Z(n12108) );
  BUF_X1 U432 ( .A(n12110), .Z(n12109) );
  BUF_X1 U433 ( .A(n10557), .Z(n12090) );
  BUF_X1 U434 ( .A(n10557), .Z(n12091) );
  BUF_X1 U435 ( .A(n10557), .Z(n12092) );
  BUF_X1 U436 ( .A(n10557), .Z(n12093) );
  BUF_X1 U437 ( .A(n12098), .Z(n12094) );
  BUF_X1 U438 ( .A(n12096), .Z(n12095) );
  BUF_X1 U439 ( .A(n10557), .Z(n12096) );
  BUF_X1 U440 ( .A(n12098), .Z(n12097) );
  BUF_X1 U441 ( .A(n10574), .Z(n12078) );
  BUF_X1 U442 ( .A(n10574), .Z(n12079) );
  BUF_X1 U443 ( .A(n10574), .Z(n12080) );
  BUF_X1 U444 ( .A(n10574), .Z(n12081) );
  BUF_X1 U445 ( .A(n12086), .Z(n12082) );
  BUF_X1 U446 ( .A(n12084), .Z(n12083) );
  BUF_X1 U447 ( .A(n10574), .Z(n12084) );
  BUF_X1 U448 ( .A(n12086), .Z(n12085) );
  BUF_X1 U449 ( .A(n10566), .Z(n12066) );
  BUF_X1 U450 ( .A(n10566), .Z(n12067) );
  BUF_X1 U451 ( .A(n10566), .Z(n12068) );
  BUF_X1 U452 ( .A(n10566), .Z(n12069) );
  BUF_X1 U453 ( .A(n12074), .Z(n12070) );
  BUF_X1 U454 ( .A(n12072), .Z(n12071) );
  BUF_X1 U455 ( .A(n10566), .Z(n12072) );
  BUF_X1 U456 ( .A(n12074), .Z(n12073) );
  BUF_X1 U457 ( .A(n10558), .Z(n12054) );
  BUF_X1 U458 ( .A(n10558), .Z(n12055) );
  BUF_X1 U459 ( .A(n10558), .Z(n12056) );
  BUF_X1 U460 ( .A(n10558), .Z(n12057) );
  BUF_X1 U461 ( .A(n12062), .Z(n12058) );
  BUF_X1 U462 ( .A(n12060), .Z(n12059) );
  BUF_X1 U463 ( .A(n10558), .Z(n12060) );
  BUF_X1 U464 ( .A(n12062), .Z(n12061) );
  BUF_X1 U465 ( .A(n10581), .Z(n12042) );
  BUF_X1 U466 ( .A(n10581), .Z(n12043) );
  BUF_X1 U467 ( .A(n10581), .Z(n12044) );
  BUF_X1 U468 ( .A(n10581), .Z(n12045) );
  BUF_X1 U469 ( .A(n12050), .Z(n12046) );
  BUF_X1 U470 ( .A(n12048), .Z(n12047) );
  BUF_X1 U471 ( .A(n10581), .Z(n12048) );
  BUF_X1 U472 ( .A(n12050), .Z(n12049) );
  BUF_X1 U473 ( .A(n10586), .Z(n12018) );
  BUF_X1 U474 ( .A(n10586), .Z(n12019) );
  BUF_X1 U475 ( .A(n10586), .Z(n12020) );
  BUF_X1 U476 ( .A(n10586), .Z(n12021) );
  BUF_X1 U477 ( .A(n10584), .Z(n11886) );
  BUF_X1 U478 ( .A(n10584), .Z(n11887) );
  BUF_X1 U479 ( .A(n10584), .Z(n11888) );
  BUF_X1 U480 ( .A(n10584), .Z(n11889) );
  BUF_X1 U481 ( .A(n11894), .Z(n11890) );
  BUF_X1 U482 ( .A(n11892), .Z(n11891) );
  BUF_X1 U483 ( .A(n10584), .Z(n11892) );
  BUF_X1 U484 ( .A(n11894), .Z(n11893) );
  BUF_X1 U485 ( .A(n10575), .Z(n11862) );
  BUF_X1 U486 ( .A(n10575), .Z(n11863) );
  BUF_X1 U487 ( .A(n10575), .Z(n11864) );
  BUF_X1 U488 ( .A(n10575), .Z(n11865) );
  BUF_X1 U489 ( .A(n11870), .Z(n11866) );
  BUF_X1 U490 ( .A(n11868), .Z(n11867) );
  BUF_X1 U491 ( .A(n10575), .Z(n11868) );
  BUF_X1 U492 ( .A(n11870), .Z(n11869) );
  BUF_X1 U493 ( .A(n10567), .Z(n11838) );
  BUF_X1 U494 ( .A(n10567), .Z(n11839) );
  BUF_X1 U495 ( .A(n10567), .Z(n11840) );
  BUF_X1 U496 ( .A(n10567), .Z(n11841) );
  BUF_X1 U497 ( .A(n11846), .Z(n11842) );
  BUF_X1 U498 ( .A(n11844), .Z(n11843) );
  BUF_X1 U499 ( .A(n10567), .Z(n11844) );
  BUF_X1 U500 ( .A(n11846), .Z(n11845) );
  BUF_X1 U501 ( .A(n10559), .Z(n11826) );
  BUF_X1 U502 ( .A(n10559), .Z(n11827) );
  BUF_X1 U503 ( .A(n10559), .Z(n11828) );
  BUF_X1 U504 ( .A(n10559), .Z(n11829) );
  BUF_X1 U505 ( .A(n11834), .Z(n11830) );
  BUF_X1 U506 ( .A(n11832), .Z(n11831) );
  BUF_X1 U507 ( .A(n10559), .Z(n11832) );
  BUF_X1 U508 ( .A(n11834), .Z(n11833) );
  BUF_X1 U509 ( .A(n10576), .Z(n11814) );
  BUF_X1 U510 ( .A(n10576), .Z(n11815) );
  BUF_X1 U511 ( .A(n10576), .Z(n11816) );
  BUF_X1 U512 ( .A(n10576), .Z(n11817) );
  BUF_X1 U513 ( .A(n11822), .Z(n11818) );
  BUF_X1 U514 ( .A(n11820), .Z(n11819) );
  BUF_X1 U515 ( .A(n10576), .Z(n11820) );
  BUF_X1 U516 ( .A(n11822), .Z(n11821) );
  BUF_X1 U517 ( .A(n10568), .Z(n11802) );
  BUF_X1 U518 ( .A(n10568), .Z(n11803) );
  BUF_X1 U519 ( .A(n10568), .Z(n11804) );
  BUF_X1 U520 ( .A(n10568), .Z(n11805) );
  BUF_X1 U521 ( .A(n11810), .Z(n11806) );
  BUF_X1 U522 ( .A(n11808), .Z(n11807) );
  BUF_X1 U523 ( .A(n10568), .Z(n11808) );
  BUF_X1 U524 ( .A(n11810), .Z(n11809) );
  BUF_X1 U525 ( .A(n10560), .Z(n11790) );
  BUF_X1 U526 ( .A(n10560), .Z(n11791) );
  BUF_X1 U527 ( .A(n10560), .Z(n11792) );
  BUF_X1 U528 ( .A(n10560), .Z(n11793) );
  BUF_X1 U529 ( .A(n11798), .Z(n11794) );
  BUF_X1 U530 ( .A(n11796), .Z(n11795) );
  BUF_X1 U531 ( .A(n10560), .Z(n11796) );
  BUF_X1 U532 ( .A(n11798), .Z(n11797) );
  BUF_X1 U533 ( .A(n10582), .Z(n11778) );
  BUF_X1 U534 ( .A(n10582), .Z(n11779) );
  BUF_X1 U535 ( .A(n10582), .Z(n11780) );
  BUF_X1 U536 ( .A(n10582), .Z(n11781) );
  BUF_X1 U537 ( .A(n11786), .Z(n11782) );
  BUF_X1 U538 ( .A(n11784), .Z(n11783) );
  BUF_X1 U539 ( .A(n10582), .Z(n11784) );
  BUF_X1 U540 ( .A(n11786), .Z(n11785) );
  BUF_X1 U541 ( .A(n10603), .Z(n11754) );
  BUF_X1 U542 ( .A(n10609), .Z(n11646) );
  BUF_X1 U543 ( .A(n11654), .Z(n11647) );
  BUF_X1 U544 ( .A(n11649), .Z(n11648) );
  BUF_X1 U545 ( .A(n10609), .Z(n11649) );
  BUF_X1 U546 ( .A(n10587), .Z(n11634) );
  BUF_X1 U547 ( .A(n10587), .Z(n11635) );
  BUF_X1 U548 ( .A(n10587), .Z(n11636) );
  BUF_X1 U549 ( .A(n10587), .Z(n11637) );
  BUF_X1 U550 ( .A(n11642), .Z(n11638) );
  BUF_X1 U551 ( .A(n11640), .Z(n11639) );
  BUF_X1 U552 ( .A(n10587), .Z(n11640) );
  BUF_X1 U553 ( .A(n11642), .Z(n11641) );
  BUF_X1 U554 ( .A(n10588), .Z(n11622) );
  BUF_X1 U555 ( .A(n10588), .Z(n11623) );
  BUF_X1 U556 ( .A(n10588), .Z(n11624) );
  BUF_X1 U557 ( .A(n10588), .Z(n11625) );
  BUF_X1 U558 ( .A(n11630), .Z(n11626) );
  BUF_X1 U559 ( .A(n11628), .Z(n11627) );
  BUF_X1 U560 ( .A(n10588), .Z(n11628) );
  BUF_X1 U561 ( .A(n11630), .Z(n11629) );
  BUF_X1 U562 ( .A(n10589), .Z(n11610) );
  BUF_X1 U563 ( .A(n10589), .Z(n11611) );
  BUF_X1 U564 ( .A(n10589), .Z(n11612) );
  BUF_X1 U565 ( .A(n10589), .Z(n11613) );
  BUF_X1 U566 ( .A(n11618), .Z(n11614) );
  BUF_X1 U567 ( .A(n11616), .Z(n11615) );
  BUF_X1 U568 ( .A(n10589), .Z(n11616) );
  BUF_X1 U569 ( .A(n11618), .Z(n11617) );
  BUF_X1 U570 ( .A(n10590), .Z(n11598) );
  BUF_X1 U571 ( .A(n10590), .Z(n11599) );
  BUF_X1 U572 ( .A(n10590), .Z(n11600) );
  BUF_X1 U573 ( .A(n10590), .Z(n11601) );
  BUF_X1 U574 ( .A(n11606), .Z(n11602) );
  BUF_X1 U575 ( .A(n11604), .Z(n11603) );
  BUF_X1 U576 ( .A(n10590), .Z(n11604) );
  BUF_X1 U577 ( .A(n11606), .Z(n11605) );
  BUF_X1 U578 ( .A(n10591), .Z(n11586) );
  BUF_X1 U579 ( .A(n10591), .Z(n11587) );
  BUF_X1 U580 ( .A(n10591), .Z(n11588) );
  BUF_X1 U581 ( .A(n10591), .Z(n11589) );
  BUF_X1 U582 ( .A(n11594), .Z(n11590) );
  BUF_X1 U583 ( .A(n11592), .Z(n11591) );
  BUF_X1 U584 ( .A(n10591), .Z(n11592) );
  BUF_X1 U585 ( .A(n11594), .Z(n11593) );
  BUF_X1 U586 ( .A(n10592), .Z(n11574) );
  BUF_X1 U587 ( .A(n10592), .Z(n11575) );
  BUF_X1 U588 ( .A(n10592), .Z(n11576) );
  BUF_X1 U589 ( .A(n10592), .Z(n11577) );
  BUF_X1 U590 ( .A(n11582), .Z(n11578) );
  BUF_X1 U591 ( .A(n11580), .Z(n11579) );
  BUF_X1 U592 ( .A(n10592), .Z(n11580) );
  BUF_X1 U593 ( .A(n11582), .Z(n11581) );
  BUF_X1 U594 ( .A(n10593), .Z(n11562) );
  BUF_X1 U595 ( .A(n10593), .Z(n11563) );
  BUF_X1 U596 ( .A(n10593), .Z(n11564) );
  BUF_X1 U597 ( .A(n10593), .Z(n11565) );
  BUF_X1 U598 ( .A(n11570), .Z(n11566) );
  BUF_X1 U599 ( .A(n11568), .Z(n11567) );
  BUF_X1 U600 ( .A(n10593), .Z(n11568) );
  BUF_X1 U601 ( .A(n11570), .Z(n11569) );
  BUF_X1 U602 ( .A(n10577), .Z(n11550) );
  BUF_X1 U603 ( .A(n10577), .Z(n11551) );
  BUF_X1 U604 ( .A(n10577), .Z(n11552) );
  BUF_X1 U605 ( .A(n10577), .Z(n11553) );
  BUF_X1 U606 ( .A(n11558), .Z(n11554) );
  BUF_X1 U607 ( .A(n11556), .Z(n11555) );
  BUF_X1 U608 ( .A(n10577), .Z(n11556) );
  BUF_X1 U609 ( .A(n11558), .Z(n11557) );
  BUF_X1 U610 ( .A(n10569), .Z(n11538) );
  BUF_X1 U611 ( .A(n10569), .Z(n11539) );
  BUF_X1 U612 ( .A(n10569), .Z(n11540) );
  BUF_X1 U613 ( .A(n10569), .Z(n11541) );
  BUF_X1 U614 ( .A(n11546), .Z(n11542) );
  BUF_X1 U615 ( .A(n11544), .Z(n11543) );
  BUF_X1 U616 ( .A(n10569), .Z(n11544) );
  BUF_X1 U617 ( .A(n11546), .Z(n11545) );
  BUF_X1 U618 ( .A(n10561), .Z(n11526) );
  BUF_X1 U619 ( .A(n10561), .Z(n11527) );
  BUF_X1 U620 ( .A(n10561), .Z(n11528) );
  BUF_X1 U621 ( .A(n10561), .Z(n11529) );
  BUF_X1 U622 ( .A(n11534), .Z(n11530) );
  BUF_X1 U623 ( .A(n11532), .Z(n11531) );
  BUF_X1 U624 ( .A(n10561), .Z(n11532) );
  BUF_X1 U625 ( .A(n11534), .Z(n11533) );
  BUF_X1 U626 ( .A(n10570), .Z(n11502) );
  BUF_X1 U627 ( .A(n10570), .Z(n11503) );
  BUF_X1 U628 ( .A(n10570), .Z(n11504) );
  BUF_X1 U629 ( .A(n10570), .Z(n11505) );
  BUF_X1 U630 ( .A(n11510), .Z(n11506) );
  BUF_X1 U631 ( .A(n11508), .Z(n11507) );
  BUF_X1 U632 ( .A(n10570), .Z(n11508) );
  BUF_X1 U633 ( .A(n11510), .Z(n11509) );
  BUF_X1 U634 ( .A(n10578), .Z(n11490) );
  BUF_X1 U635 ( .A(n10578), .Z(n11491) );
  BUF_X1 U636 ( .A(n10578), .Z(n11492) );
  BUF_X1 U637 ( .A(n10578), .Z(n11493) );
  BUF_X1 U638 ( .A(n11498), .Z(n11494) );
  BUF_X1 U639 ( .A(n11496), .Z(n11495) );
  BUF_X1 U640 ( .A(n10578), .Z(n11496) );
  BUF_X1 U641 ( .A(n11498), .Z(n11497) );
  BUF_X1 U642 ( .A(n10562), .Z(n11478) );
  BUF_X1 U643 ( .A(n10562), .Z(n11479) );
  BUF_X1 U644 ( .A(n10562), .Z(n11480) );
  BUF_X1 U645 ( .A(n10562), .Z(n11481) );
  BUF_X1 U646 ( .A(n11486), .Z(n11482) );
  BUF_X1 U647 ( .A(n11484), .Z(n11483) );
  BUF_X1 U648 ( .A(n10562), .Z(n11484) );
  BUF_X1 U649 ( .A(n10579), .Z(n11454) );
  BUF_X1 U650 ( .A(n10579), .Z(n11455) );
  BUF_X1 U651 ( .A(n10579), .Z(n11456) );
  BUF_X1 U652 ( .A(n10579), .Z(n11457) );
  BUF_X1 U653 ( .A(n11462), .Z(n11458) );
  BUF_X1 U654 ( .A(n11460), .Z(n11459) );
  BUF_X1 U655 ( .A(n10579), .Z(n11460) );
  BUF_X1 U656 ( .A(n11462), .Z(n11461) );
  BUF_X1 U657 ( .A(n10563), .Z(n11442) );
  BUF_X1 U658 ( .A(n10563), .Z(n11443) );
  BUF_X1 U659 ( .A(n10563), .Z(n11444) );
  BUF_X1 U660 ( .A(n10563), .Z(n11445) );
  BUF_X1 U661 ( .A(n11450), .Z(n11446) );
  BUF_X1 U662 ( .A(n11448), .Z(n11447) );
  BUF_X1 U663 ( .A(n10563), .Z(n11448) );
  BUF_X1 U664 ( .A(n10572), .Z(n11430) );
  BUF_X1 U665 ( .A(n10572), .Z(n11431) );
  BUF_X1 U666 ( .A(n10572), .Z(n11432) );
  BUF_X1 U667 ( .A(n10572), .Z(n11433) );
  BUF_X1 U668 ( .A(n11438), .Z(n11434) );
  BUF_X1 U669 ( .A(n11436), .Z(n11435) );
  BUF_X1 U670 ( .A(n10572), .Z(n11436) );
  BUF_X1 U671 ( .A(n11438), .Z(n11437) );
  BUF_X1 U672 ( .A(n10580), .Z(n11418) );
  BUF_X1 U673 ( .A(n10580), .Z(n11419) );
  BUF_X1 U674 ( .A(n10580), .Z(n11420) );
  BUF_X1 U675 ( .A(n10580), .Z(n11421) );
  BUF_X1 U676 ( .A(n11426), .Z(n11422) );
  BUF_X1 U677 ( .A(n11424), .Z(n11423) );
  BUF_X1 U678 ( .A(n10580), .Z(n11424) );
  BUF_X1 U679 ( .A(n11426), .Z(n11425) );
  BUF_X1 U680 ( .A(n10564), .Z(n11406) );
  BUF_X1 U681 ( .A(n10564), .Z(n11407) );
  BUF_X1 U682 ( .A(n10564), .Z(n11408) );
  BUF_X1 U683 ( .A(n10564), .Z(n11409) );
  BUF_X1 U684 ( .A(n11414), .Z(n11410) );
  BUF_X1 U685 ( .A(n11412), .Z(n11411) );
  BUF_X1 U686 ( .A(n10564), .Z(n11412) );
  BUF_X1 U687 ( .A(n10583), .Z(n11394) );
  BUF_X1 U688 ( .A(n10583), .Z(n11395) );
  BUF_X1 U689 ( .A(n10583), .Z(n11396) );
  BUF_X1 U690 ( .A(n10583), .Z(n11397) );
  BUF_X1 U691 ( .A(n11402), .Z(n11398) );
  BUF_X1 U692 ( .A(n11400), .Z(n11399) );
  BUF_X1 U693 ( .A(n10583), .Z(n11400) );
  BUF_X1 U694 ( .A(n11402), .Z(n11401) );
  BUF_X1 U695 ( .A(n10585), .Z(n11382) );
  BUF_X1 U696 ( .A(n10585), .Z(n11383) );
  BUF_X1 U697 ( .A(n10585), .Z(n11384) );
  BUF_X1 U698 ( .A(n10585), .Z(n11385) );
  BUF_X1 U699 ( .A(n11390), .Z(n11386) );
  BUF_X1 U700 ( .A(n11388), .Z(n11387) );
  BUF_X1 U701 ( .A(n10585), .Z(n11388) );
  BUF_X1 U702 ( .A(n11390), .Z(n11389) );
  BUF_X1 U703 ( .A(n10619), .Z(n12407) );
  BUF_X1 U704 ( .A(n10619), .Z(n12408) );
  BUF_X1 U705 ( .A(n10619), .Z(n12409) );
  BUF_X1 U706 ( .A(n10619), .Z(n12410) );
  BUF_X1 U707 ( .A(n12415), .Z(n12411) );
  BUF_X1 U708 ( .A(n12413), .Z(n12412) );
  BUF_X1 U709 ( .A(n10619), .Z(n12413) );
  BUF_X1 U710 ( .A(n12415), .Z(n12414) );
  BUF_X1 U711 ( .A(n10620), .Z(n12396) );
  BUF_X1 U712 ( .A(n10620), .Z(n12397) );
  BUF_X1 U713 ( .A(n10620), .Z(n12398) );
  BUF_X1 U714 ( .A(n10620), .Z(n12399) );
  BUF_X1 U715 ( .A(n12404), .Z(n12400) );
  BUF_X1 U716 ( .A(n12402), .Z(n12401) );
  BUF_X1 U717 ( .A(n10620), .Z(n12402) );
  BUF_X1 U718 ( .A(n12404), .Z(n12403) );
  BUF_X1 U719 ( .A(n10621), .Z(n12385) );
  BUF_X1 U720 ( .A(n10621), .Z(n12386) );
  BUF_X1 U721 ( .A(n10621), .Z(n12387) );
  BUF_X1 U722 ( .A(n10621), .Z(n12388) );
  BUF_X1 U723 ( .A(n12393), .Z(n12389) );
  BUF_X1 U724 ( .A(n12391), .Z(n12390) );
  BUF_X1 U725 ( .A(n10621), .Z(n12391) );
  BUF_X1 U726 ( .A(n12393), .Z(n12392) );
  BUF_X1 U727 ( .A(n10622), .Z(n12374) );
  BUF_X1 U728 ( .A(n10622), .Z(n12375) );
  BUF_X1 U729 ( .A(n10622), .Z(n12376) );
  BUF_X1 U730 ( .A(n10622), .Z(n12377) );
  BUF_X1 U731 ( .A(n12382), .Z(n12378) );
  BUF_X1 U732 ( .A(n12380), .Z(n12379) );
  BUF_X1 U733 ( .A(n10622), .Z(n12380) );
  BUF_X1 U734 ( .A(n12382), .Z(n12381) );
  BUF_X1 U735 ( .A(n10623), .Z(n12363) );
  BUF_X1 U736 ( .A(n10623), .Z(n12364) );
  BUF_X1 U737 ( .A(n10623), .Z(n12365) );
  BUF_X1 U738 ( .A(n10623), .Z(n12366) );
  BUF_X1 U739 ( .A(n12371), .Z(n12367) );
  BUF_X1 U740 ( .A(n12369), .Z(n12368) );
  BUF_X1 U741 ( .A(n10623), .Z(n12369) );
  BUF_X1 U742 ( .A(n12371), .Z(n12370) );
  BUF_X1 U743 ( .A(n10624), .Z(n12352) );
  BUF_X1 U744 ( .A(n10624), .Z(n12353) );
  BUF_X1 U745 ( .A(n10624), .Z(n12354) );
  BUF_X1 U746 ( .A(n10624), .Z(n12355) );
  BUF_X1 U747 ( .A(n12360), .Z(n12356) );
  BUF_X1 U748 ( .A(n12358), .Z(n12357) );
  BUF_X1 U749 ( .A(n10624), .Z(n12358) );
  BUF_X1 U750 ( .A(n12360), .Z(n12359) );
  BUF_X1 U751 ( .A(n10618), .Z(n12341) );
  BUF_X1 U752 ( .A(n10618), .Z(n12342) );
  BUF_X1 U753 ( .A(n10618), .Z(n12343) );
  BUF_X1 U754 ( .A(n10618), .Z(n12344) );
  BUF_X1 U755 ( .A(n12349), .Z(n12345) );
  BUF_X1 U756 ( .A(n12347), .Z(n12346) );
  BUF_X1 U757 ( .A(n10618), .Z(n12347) );
  BUF_X1 U758 ( .A(n12349), .Z(n12348) );
  BUF_X1 U759 ( .A(n10615), .Z(n12330) );
  BUF_X1 U760 ( .A(n10615), .Z(n12331) );
  BUF_X1 U761 ( .A(n10615), .Z(n12332) );
  BUF_X1 U762 ( .A(n10615), .Z(n12333) );
  BUF_X1 U763 ( .A(n12338), .Z(n12334) );
  BUF_X1 U764 ( .A(n12336), .Z(n12335) );
  BUF_X1 U765 ( .A(n10615), .Z(n12336) );
  BUF_X1 U766 ( .A(n12338), .Z(n12337) );
  BUF_X1 U767 ( .A(n10614), .Z(n12318) );
  BUF_X1 U768 ( .A(n10614), .Z(n12319) );
  BUF_X1 U769 ( .A(n10614), .Z(n12320) );
  BUF_X1 U770 ( .A(n10614), .Z(n12321) );
  BUF_X1 U771 ( .A(n12326), .Z(n12322) );
  BUF_X1 U772 ( .A(n12324), .Z(n12323) );
  BUF_X1 U773 ( .A(n10614), .Z(n12324) );
  BUF_X1 U774 ( .A(n12326), .Z(n12325) );
  BUF_X1 U775 ( .A(n10617), .Z(n12306) );
  BUF_X1 U776 ( .A(n10617), .Z(n12307) );
  BUF_X1 U777 ( .A(n10617), .Z(n12308) );
  BUF_X1 U778 ( .A(n10617), .Z(n12309) );
  BUF_X1 U779 ( .A(n12314), .Z(n12310) );
  BUF_X1 U780 ( .A(n12312), .Z(n12311) );
  BUF_X1 U781 ( .A(n10617), .Z(n12312) );
  BUF_X1 U782 ( .A(n12314), .Z(n12313) );
  BUF_X1 U783 ( .A(n10603), .Z(n11755) );
  BUF_X1 U784 ( .A(n11486), .Z(n11485) );
  BUF_X1 U785 ( .A(n10541), .Z(n12198) );
  BUF_X1 U786 ( .A(n12026), .Z(n12022) );
  BUF_X1 U787 ( .A(n10596), .Z(n12006) );
  BUF_X1 U788 ( .A(n11450), .Z(n11449) );
  BUF_X1 U789 ( .A(n11414), .Z(n11413) );
  BUF_X1 U790 ( .A(n10611), .Z(n12270) );
  BUF_X1 U791 ( .A(n10539), .Z(n12222) );
  BUF_X1 U792 ( .A(n10539), .Z(n12223) );
  BUF_X1 U793 ( .A(n10539), .Z(n12224) );
  BUF_X1 U794 ( .A(n10539), .Z(n12225) );
  BUF_X1 U795 ( .A(n12230), .Z(n12226) );
  BUF_X1 U796 ( .A(n12228), .Z(n12227) );
  BUF_X1 U797 ( .A(n10539), .Z(n12228) );
  BUF_X1 U798 ( .A(n12230), .Z(n12229) );
  BUF_X1 U799 ( .A(n10540), .Z(n12210) );
  BUF_X1 U800 ( .A(n10540), .Z(n12211) );
  BUF_X1 U801 ( .A(n10540), .Z(n12212) );
  BUF_X1 U802 ( .A(n10540), .Z(n12213) );
  BUF_X1 U803 ( .A(n12218), .Z(n12214) );
  BUF_X1 U804 ( .A(n12216), .Z(n12215) );
  BUF_X1 U805 ( .A(n10540), .Z(n12216) );
  BUF_X1 U806 ( .A(n12218), .Z(n12217) );
  BUF_X1 U807 ( .A(n10541), .Z(n12199) );
  BUF_X1 U808 ( .A(n10541), .Z(n12200) );
  BUF_X1 U809 ( .A(n10541), .Z(n12201) );
  BUF_X1 U810 ( .A(n10541), .Z(n12202) );
  BUF_X1 U811 ( .A(n10541), .Z(n12203) );
  BUF_X1 U812 ( .A(n12198), .Z(n12204) );
  BUF_X1 U813 ( .A(n12200), .Z(n12205) );
  BUF_X1 U814 ( .A(n10542), .Z(n12186) );
  BUF_X1 U815 ( .A(n10542), .Z(n12187) );
  BUF_X1 U816 ( .A(n10542), .Z(n12188) );
  BUF_X1 U817 ( .A(n10542), .Z(n12189) );
  BUF_X1 U818 ( .A(n12194), .Z(n12190) );
  BUF_X1 U819 ( .A(n12192), .Z(n12191) );
  BUF_X1 U820 ( .A(n10542), .Z(n12192) );
  BUF_X1 U821 ( .A(n12194), .Z(n12193) );
  BUF_X1 U822 ( .A(n10543), .Z(n12174) );
  BUF_X1 U823 ( .A(n10543), .Z(n12175) );
  BUF_X1 U824 ( .A(n10543), .Z(n12176) );
  BUF_X1 U825 ( .A(n10543), .Z(n12177) );
  BUF_X1 U826 ( .A(n12182), .Z(n12178) );
  BUF_X1 U827 ( .A(n12180), .Z(n12179) );
  BUF_X1 U828 ( .A(n10543), .Z(n12180) );
  BUF_X1 U829 ( .A(n12182), .Z(n12181) );
  BUF_X1 U830 ( .A(n10544), .Z(n12162) );
  BUF_X1 U831 ( .A(n10544), .Z(n12163) );
  BUF_X1 U832 ( .A(n10544), .Z(n12164) );
  BUF_X1 U833 ( .A(n10544), .Z(n12165) );
  BUF_X1 U834 ( .A(n12170), .Z(n12166) );
  BUF_X1 U835 ( .A(n12168), .Z(n12167) );
  BUF_X1 U836 ( .A(n10544), .Z(n12168) );
  BUF_X1 U837 ( .A(n12170), .Z(n12169) );
  BUF_X1 U838 ( .A(n10546), .Z(n12138) );
  BUF_X1 U839 ( .A(n10546), .Z(n12139) );
  BUF_X1 U840 ( .A(n10546), .Z(n12140) );
  BUF_X1 U841 ( .A(n10546), .Z(n12141) );
  BUF_X1 U842 ( .A(n12146), .Z(n12142) );
  BUF_X1 U843 ( .A(n12144), .Z(n12143) );
  BUF_X1 U844 ( .A(n10546), .Z(n12144) );
  BUF_X1 U845 ( .A(n12146), .Z(n12145) );
  BUF_X1 U846 ( .A(n10547), .Z(n12114) );
  BUF_X1 U847 ( .A(n10547), .Z(n12115) );
  BUF_X1 U848 ( .A(n10547), .Z(n12116) );
  BUF_X1 U849 ( .A(n10547), .Z(n12117) );
  BUF_X1 U850 ( .A(n12122), .Z(n12118) );
  BUF_X1 U851 ( .A(n12120), .Z(n12119) );
  BUF_X1 U852 ( .A(n10547), .Z(n12120) );
  BUF_X1 U853 ( .A(n12122), .Z(n12121) );
  BUF_X1 U854 ( .A(n10595), .Z(n12030) );
  BUF_X1 U855 ( .A(n10595), .Z(n12031) );
  BUF_X1 U856 ( .A(n10595), .Z(n12032) );
  BUF_X1 U857 ( .A(n10595), .Z(n12033) );
  BUF_X1 U858 ( .A(n12038), .Z(n12034) );
  BUF_X1 U859 ( .A(n12036), .Z(n12035) );
  BUF_X1 U860 ( .A(n10595), .Z(n12036) );
  BUF_X1 U861 ( .A(n12038), .Z(n12037) );
  BUF_X1 U862 ( .A(n12018), .Z(n12023) );
  BUF_X1 U863 ( .A(n10586), .Z(n12024) );
  BUF_X1 U864 ( .A(n12026), .Z(n12025) );
  BUF_X1 U865 ( .A(n12014), .Z(n12007) );
  BUF_X1 U866 ( .A(n12012), .Z(n12008) );
  BUF_X1 U867 ( .A(n10596), .Z(n12009) );
  BUF_X1 U868 ( .A(n10596), .Z(n12010) );
  BUF_X1 U869 ( .A(n10596), .Z(n12011) );
  BUF_X1 U870 ( .A(n10596), .Z(n12012) );
  BUF_X1 U871 ( .A(n12014), .Z(n12013) );
  BUF_X1 U872 ( .A(n10597), .Z(n11994) );
  BUF_X1 U873 ( .A(n10597), .Z(n11995) );
  BUF_X1 U874 ( .A(n10597), .Z(n11996) );
  BUF_X1 U875 ( .A(n10597), .Z(n11997) );
  BUF_X1 U876 ( .A(n12002), .Z(n11998) );
  BUF_X1 U877 ( .A(n12000), .Z(n11999) );
  BUF_X1 U878 ( .A(n10597), .Z(n12000) );
  BUF_X1 U879 ( .A(n12002), .Z(n12001) );
  BUF_X1 U880 ( .A(n10598), .Z(n11982) );
  BUF_X1 U881 ( .A(n10598), .Z(n11983) );
  BUF_X1 U882 ( .A(n10598), .Z(n11984) );
  BUF_X1 U883 ( .A(n10598), .Z(n11985) );
  BUF_X1 U884 ( .A(n11990), .Z(n11986) );
  BUF_X1 U885 ( .A(n11988), .Z(n11987) );
  BUF_X1 U886 ( .A(n10598), .Z(n11988) );
  BUF_X1 U887 ( .A(n11990), .Z(n11989) );
  BUF_X1 U888 ( .A(n10599), .Z(n11970) );
  BUF_X1 U889 ( .A(n10599), .Z(n11971) );
  BUF_X1 U890 ( .A(n10599), .Z(n11972) );
  BUF_X1 U891 ( .A(n10599), .Z(n11973) );
  BUF_X1 U892 ( .A(n11978), .Z(n11974) );
  BUF_X1 U893 ( .A(n11976), .Z(n11975) );
  BUF_X1 U894 ( .A(n10599), .Z(n11976) );
  BUF_X1 U895 ( .A(n11978), .Z(n11977) );
  BUF_X1 U896 ( .A(n10548), .Z(n11958) );
  BUF_X1 U897 ( .A(n10548), .Z(n11959) );
  BUF_X1 U898 ( .A(n10548), .Z(n11960) );
  BUF_X1 U899 ( .A(n10548), .Z(n11961) );
  BUF_X1 U900 ( .A(n11966), .Z(n11962) );
  BUF_X1 U901 ( .A(n11964), .Z(n11963) );
  BUF_X1 U902 ( .A(n10548), .Z(n11964) );
  BUF_X1 U903 ( .A(n11966), .Z(n11965) );
  BUF_X1 U904 ( .A(n10549), .Z(n11946) );
  BUF_X1 U905 ( .A(n10549), .Z(n11947) );
  BUF_X1 U906 ( .A(n10549), .Z(n11948) );
  BUF_X1 U907 ( .A(n10549), .Z(n11949) );
  BUF_X1 U908 ( .A(n11954), .Z(n11950) );
  BUF_X1 U909 ( .A(n11952), .Z(n11951) );
  BUF_X1 U910 ( .A(n10549), .Z(n11952) );
  BUF_X1 U911 ( .A(n11954), .Z(n11953) );
  BUF_X1 U912 ( .A(n10550), .Z(n11934) );
  BUF_X1 U913 ( .A(n10550), .Z(n11935) );
  BUF_X1 U914 ( .A(n10550), .Z(n11936) );
  BUF_X1 U915 ( .A(n10550), .Z(n11937) );
  BUF_X1 U916 ( .A(n11942), .Z(n11938) );
  BUF_X1 U917 ( .A(n11940), .Z(n11939) );
  BUF_X1 U918 ( .A(n10550), .Z(n11940) );
  BUF_X1 U919 ( .A(n11942), .Z(n11941) );
  BUF_X1 U920 ( .A(n10600), .Z(n11922) );
  BUF_X1 U921 ( .A(n10600), .Z(n11923) );
  BUF_X1 U922 ( .A(n10600), .Z(n11924) );
  BUF_X1 U923 ( .A(n10600), .Z(n11925) );
  BUF_X1 U924 ( .A(n11930), .Z(n11926) );
  BUF_X1 U925 ( .A(n11928), .Z(n11927) );
  BUF_X1 U926 ( .A(n10600), .Z(n11928) );
  BUF_X1 U927 ( .A(n11930), .Z(n11929) );
  BUF_X1 U928 ( .A(n10601), .Z(n11910) );
  BUF_X1 U929 ( .A(n10601), .Z(n11911) );
  BUF_X1 U930 ( .A(n10601), .Z(n11912) );
  BUF_X1 U931 ( .A(n10601), .Z(n11913) );
  BUF_X1 U932 ( .A(n11918), .Z(n11914) );
  BUF_X1 U933 ( .A(n11916), .Z(n11915) );
  BUF_X1 U934 ( .A(n10601), .Z(n11916) );
  BUF_X1 U935 ( .A(n11918), .Z(n11917) );
  BUF_X1 U936 ( .A(n10552), .Z(n11874) );
  BUF_X1 U937 ( .A(n10552), .Z(n11875) );
  BUF_X1 U938 ( .A(n10552), .Z(n11876) );
  BUF_X1 U939 ( .A(n10552), .Z(n11877) );
  BUF_X1 U940 ( .A(n11882), .Z(n11878) );
  BUF_X1 U941 ( .A(n11880), .Z(n11879) );
  BUF_X1 U942 ( .A(n10552), .Z(n11880) );
  BUF_X1 U943 ( .A(n11882), .Z(n11881) );
  BUF_X1 U944 ( .A(n10602), .Z(n11766) );
  BUF_X1 U945 ( .A(n10602), .Z(n11767) );
  BUF_X1 U946 ( .A(n10602), .Z(n11768) );
  BUF_X1 U947 ( .A(n10602), .Z(n11769) );
  BUF_X1 U948 ( .A(n11774), .Z(n11770) );
  BUF_X1 U949 ( .A(n11772), .Z(n11771) );
  BUF_X1 U950 ( .A(n10602), .Z(n11772) );
  BUF_X1 U951 ( .A(n11774), .Z(n11773) );
  BUF_X1 U952 ( .A(n10603), .Z(n11756) );
  BUF_X1 U953 ( .A(n10603), .Z(n11757) );
  BUF_X1 U954 ( .A(n11762), .Z(n11758) );
  BUF_X1 U955 ( .A(n11754), .Z(n11759) );
  BUF_X1 U956 ( .A(n10603), .Z(n11760) );
  BUF_X1 U957 ( .A(n11762), .Z(n11761) );
  BUF_X1 U958 ( .A(n10604), .Z(n11742) );
  BUF_X1 U959 ( .A(n10604), .Z(n11743) );
  BUF_X1 U960 ( .A(n10604), .Z(n11744) );
  BUF_X1 U961 ( .A(n10604), .Z(n11745) );
  BUF_X1 U962 ( .A(n11750), .Z(n11746) );
  BUF_X1 U963 ( .A(n11748), .Z(n11747) );
  BUF_X1 U964 ( .A(n10604), .Z(n11748) );
  BUF_X1 U965 ( .A(n11750), .Z(n11749) );
  BUF_X1 U966 ( .A(n10605), .Z(n11730) );
  BUF_X1 U967 ( .A(n10605), .Z(n11731) );
  BUF_X1 U968 ( .A(n10605), .Z(n11732) );
  BUF_X1 U969 ( .A(n10605), .Z(n11733) );
  BUF_X1 U970 ( .A(n11738), .Z(n11734) );
  BUF_X1 U971 ( .A(n11736), .Z(n11735) );
  BUF_X1 U972 ( .A(n10605), .Z(n11736) );
  BUF_X1 U973 ( .A(n11738), .Z(n11737) );
  BUF_X1 U974 ( .A(n10606), .Z(n11718) );
  BUF_X1 U975 ( .A(n10606), .Z(n11719) );
  BUF_X1 U976 ( .A(n10606), .Z(n11720) );
  BUF_X1 U977 ( .A(n10606), .Z(n11721) );
  BUF_X1 U978 ( .A(n11726), .Z(n11722) );
  BUF_X1 U979 ( .A(n11724), .Z(n11723) );
  BUF_X1 U980 ( .A(n10606), .Z(n11724) );
  BUF_X1 U981 ( .A(n11726), .Z(n11725) );
  BUF_X1 U982 ( .A(n10607), .Z(n11706) );
  BUF_X1 U983 ( .A(n10607), .Z(n11707) );
  BUF_X1 U984 ( .A(n10607), .Z(n11708) );
  BUF_X1 U985 ( .A(n10607), .Z(n11709) );
  BUF_X1 U986 ( .A(n11714), .Z(n11710) );
  BUF_X1 U987 ( .A(n11712), .Z(n11711) );
  BUF_X1 U988 ( .A(n10607), .Z(n11712) );
  BUF_X1 U989 ( .A(n11714), .Z(n11713) );
  BUF_X1 U990 ( .A(n10554), .Z(n11694) );
  BUF_X1 U991 ( .A(n10554), .Z(n11695) );
  BUF_X1 U992 ( .A(n10554), .Z(n11696) );
  BUF_X1 U993 ( .A(n10554), .Z(n11697) );
  BUF_X1 U994 ( .A(n11702), .Z(n11698) );
  BUF_X1 U995 ( .A(n11700), .Z(n11699) );
  BUF_X1 U996 ( .A(n10554), .Z(n11700) );
  BUF_X1 U997 ( .A(n11702), .Z(n11701) );
  BUF_X1 U998 ( .A(n10555), .Z(n11682) );
  BUF_X1 U999 ( .A(n10555), .Z(n11683) );
  BUF_X1 U1000 ( .A(n10555), .Z(n11684) );
  BUF_X1 U1001 ( .A(n10555), .Z(n11685) );
  BUF_X1 U1002 ( .A(n11690), .Z(n11686) );
  BUF_X1 U1003 ( .A(n11688), .Z(n11687) );
  BUF_X1 U1004 ( .A(n10555), .Z(n11688) );
  BUF_X1 U1005 ( .A(n11690), .Z(n11689) );
  BUF_X1 U1006 ( .A(n10556), .Z(n11670) );
  BUF_X1 U1007 ( .A(n10556), .Z(n11671) );
  BUF_X1 U1008 ( .A(n10556), .Z(n11672) );
  BUF_X1 U1009 ( .A(n10556), .Z(n11673) );
  BUF_X1 U1010 ( .A(n11678), .Z(n11674) );
  BUF_X1 U1011 ( .A(n11676), .Z(n11675) );
  BUF_X1 U1012 ( .A(n10556), .Z(n11676) );
  BUF_X1 U1013 ( .A(n11678), .Z(n11677) );
  BUF_X1 U1014 ( .A(n10608), .Z(n11658) );
  BUF_X1 U1015 ( .A(n10608), .Z(n11659) );
  BUF_X1 U1016 ( .A(n10608), .Z(n11660) );
  BUF_X1 U1017 ( .A(n10608), .Z(n11661) );
  BUF_X1 U1018 ( .A(n11666), .Z(n11662) );
  BUF_X1 U1019 ( .A(n11664), .Z(n11663) );
  BUF_X1 U1020 ( .A(n10608), .Z(n11664) );
  BUF_X1 U1021 ( .A(n11666), .Z(n11665) );
  BUF_X1 U1022 ( .A(n10609), .Z(n11653) );
  BUF_X1 U1023 ( .A(n10609), .Z(n11652) );
  BUF_X1 U1024 ( .A(n11654), .Z(n11651) );
  BUF_X1 U1025 ( .A(n10609), .Z(n11650) );
  BUF_X1 U1026 ( .A(n10610), .Z(n12294) );
  BUF_X1 U1027 ( .A(n10610), .Z(n12295) );
  BUF_X1 U1028 ( .A(n10610), .Z(n12296) );
  BUF_X1 U1029 ( .A(n10610), .Z(n12297) );
  BUF_X1 U1030 ( .A(n12302), .Z(n12298) );
  BUF_X1 U1031 ( .A(n12300), .Z(n12299) );
  BUF_X1 U1032 ( .A(n10610), .Z(n12300) );
  BUF_X1 U1033 ( .A(n12302), .Z(n12301) );
  BUF_X1 U1034 ( .A(n10611), .Z(n12271) );
  BUF_X1 U1035 ( .A(n10611), .Z(n12272) );
  BUF_X1 U1036 ( .A(n10611), .Z(n12273) );
  BUF_X1 U1037 ( .A(n10611), .Z(n12274) );
  BUF_X1 U1038 ( .A(n10611), .Z(n12275) );
  BUF_X1 U1039 ( .A(n12270), .Z(n12276) );
  BUF_X1 U1040 ( .A(n12272), .Z(n12277) );
  BUF_X1 U1041 ( .A(n10612), .Z(n12258) );
  BUF_X1 U1042 ( .A(n10612), .Z(n12259) );
  BUF_X1 U1043 ( .A(n10612), .Z(n12260) );
  BUF_X1 U1044 ( .A(n10612), .Z(n12261) );
  BUF_X1 U1045 ( .A(n12266), .Z(n12262) );
  BUF_X1 U1046 ( .A(n12264), .Z(n12263) );
  BUF_X1 U1047 ( .A(n10612), .Z(n12264) );
  BUF_X1 U1048 ( .A(n12266), .Z(n12265) );
  BUF_X1 U1049 ( .A(n10613), .Z(n12246) );
  BUF_X1 U1050 ( .A(n10613), .Z(n12247) );
  BUF_X1 U1051 ( .A(n10613), .Z(n12248) );
  BUF_X1 U1052 ( .A(n10613), .Z(n12249) );
  BUF_X1 U1053 ( .A(n12254), .Z(n12250) );
  BUF_X1 U1054 ( .A(n12252), .Z(n12251) );
  BUF_X1 U1055 ( .A(n10613), .Z(n12252) );
  BUF_X1 U1056 ( .A(n12254), .Z(n12253) );
  BUF_X1 U1057 ( .A(n12713), .Z(n12712) );
  BUF_X1 U1058 ( .A(n10539), .Z(n12230) );
  BUF_X1 U1059 ( .A(n10540), .Z(n12218) );
  BUF_X1 U1060 ( .A(n12201), .Z(n12206) );
  BUF_X1 U1061 ( .A(n10542), .Z(n12194) );
  BUF_X1 U1062 ( .A(n10543), .Z(n12182) );
  BUF_X1 U1063 ( .A(n10544), .Z(n12170) );
  BUF_X1 U1064 ( .A(n10545), .Z(n12158) );
  BUF_X1 U1065 ( .A(n10546), .Z(n12146) );
  BUF_X1 U1066 ( .A(n10573), .Z(n12134) );
  BUF_X1 U1067 ( .A(n10547), .Z(n12122) );
  BUF_X1 U1068 ( .A(n10565), .Z(n12110) );
  BUF_X1 U1069 ( .A(n10557), .Z(n12098) );
  BUF_X1 U1070 ( .A(n10574), .Z(n12086) );
  BUF_X1 U1071 ( .A(n10566), .Z(n12074) );
  BUF_X1 U1072 ( .A(n10558), .Z(n12062) );
  BUF_X1 U1073 ( .A(n10581), .Z(n12050) );
  BUF_X1 U1074 ( .A(n10595), .Z(n12038) );
  BUF_X1 U1075 ( .A(n10586), .Z(n12026) );
  BUF_X1 U1076 ( .A(n10596), .Z(n12014) );
  BUF_X1 U1077 ( .A(n10597), .Z(n12002) );
  BUF_X1 U1078 ( .A(n10598), .Z(n11990) );
  BUF_X1 U1079 ( .A(n10599), .Z(n11978) );
  BUF_X1 U1080 ( .A(n10548), .Z(n11966) );
  BUF_X1 U1081 ( .A(n10549), .Z(n11954) );
  BUF_X1 U1082 ( .A(n10550), .Z(n11942) );
  BUF_X1 U1083 ( .A(n10600), .Z(n11930) );
  BUF_X1 U1084 ( .A(n10601), .Z(n11918) );
  BUF_X1 U1085 ( .A(n10584), .Z(n11894) );
  BUF_X1 U1086 ( .A(n10552), .Z(n11882) );
  BUF_X1 U1087 ( .A(n10575), .Z(n11870) );
  BUF_X1 U1088 ( .A(n10567), .Z(n11846) );
  BUF_X1 U1089 ( .A(n10559), .Z(n11834) );
  BUF_X1 U1090 ( .A(n10576), .Z(n11822) );
  BUF_X1 U1091 ( .A(n10568), .Z(n11810) );
  BUF_X1 U1092 ( .A(n10560), .Z(n11798) );
  BUF_X1 U1093 ( .A(n10582), .Z(n11786) );
  BUF_X1 U1094 ( .A(n10602), .Z(n11774) );
  BUF_X1 U1095 ( .A(n10603), .Z(n11762) );
  BUF_X1 U1096 ( .A(n10604), .Z(n11750) );
  BUF_X1 U1097 ( .A(n10605), .Z(n11738) );
  BUF_X1 U1098 ( .A(n10606), .Z(n11726) );
  BUF_X1 U1099 ( .A(n10607), .Z(n11714) );
  BUF_X1 U1100 ( .A(n10554), .Z(n11702) );
  BUF_X1 U1101 ( .A(n10555), .Z(n11690) );
  BUF_X1 U1102 ( .A(n10556), .Z(n11678) );
  BUF_X1 U1103 ( .A(n10608), .Z(n11666) );
  BUF_X1 U1104 ( .A(n10609), .Z(n11654) );
  BUF_X1 U1105 ( .A(n10587), .Z(n11642) );
  BUF_X1 U1106 ( .A(n10588), .Z(n11630) );
  BUF_X1 U1107 ( .A(n10589), .Z(n11618) );
  BUF_X1 U1108 ( .A(n10590), .Z(n11606) );
  BUF_X1 U1109 ( .A(n10591), .Z(n11594) );
  BUF_X1 U1110 ( .A(n10592), .Z(n11582) );
  BUF_X1 U1111 ( .A(n10593), .Z(n11570) );
  BUF_X1 U1112 ( .A(n10577), .Z(n11558) );
  BUF_X1 U1113 ( .A(n10569), .Z(n11546) );
  BUF_X1 U1114 ( .A(n10561), .Z(n11534) );
  BUF_X1 U1115 ( .A(n10570), .Z(n11510) );
  BUF_X1 U1116 ( .A(n10578), .Z(n11498) );
  BUF_X1 U1117 ( .A(n10562), .Z(n11486) );
  BUF_X1 U1118 ( .A(n10579), .Z(n11462) );
  BUF_X1 U1119 ( .A(n10563), .Z(n11450) );
  BUF_X1 U1120 ( .A(n10572), .Z(n11438) );
  BUF_X1 U1121 ( .A(n10580), .Z(n11426) );
  BUF_X1 U1122 ( .A(n10564), .Z(n11414) );
  BUF_X1 U1123 ( .A(n10583), .Z(n11402) );
  BUF_X1 U1124 ( .A(n10585), .Z(n11390) );
  BUF_X1 U1125 ( .A(n10619), .Z(n12415) );
  BUF_X1 U1126 ( .A(n10620), .Z(n12404) );
  BUF_X1 U1127 ( .A(n10621), .Z(n12393) );
  BUF_X1 U1128 ( .A(n10622), .Z(n12382) );
  BUF_X1 U1129 ( .A(n10623), .Z(n12371) );
  BUF_X1 U1130 ( .A(n10624), .Z(n12360) );
  BUF_X1 U1131 ( .A(n10618), .Z(n12349) );
  BUF_X1 U1132 ( .A(n10615), .Z(n12338) );
  BUF_X1 U1133 ( .A(n10614), .Z(n12326) );
  BUF_X1 U1134 ( .A(n10617), .Z(n12314) );
  BUF_X1 U1135 ( .A(n10610), .Z(n12302) );
  BUF_X1 U1136 ( .A(n12273), .Z(n12278) );
  BUF_X1 U1137 ( .A(n10612), .Z(n12266) );
  BUF_X1 U1138 ( .A(n10613), .Z(n12254) );
  BUF_X1 U1139 ( .A(n4339), .Z(n10986) );
  BUF_X1 U1140 ( .A(n2871), .Z(n11250) );
  BUF_X1 U1141 ( .A(n4339), .Z(n10987) );
  BUF_X1 U1142 ( .A(n2871), .Z(n11251) );
  BUF_X1 U1143 ( .A(n4337), .Z(n10992) );
  BUF_X1 U1144 ( .A(n4340), .Z(n10983) );
  BUF_X1 U1145 ( .A(n2869), .Z(n11256) );
  BUF_X1 U1146 ( .A(n2872), .Z(n11247) );
  BUF_X1 U1147 ( .A(n4337), .Z(n10993) );
  BUF_X1 U1148 ( .A(n4340), .Z(n10984) );
  BUF_X1 U1149 ( .A(n2869), .Z(n11257) );
  BUF_X1 U1150 ( .A(n2872), .Z(n11248) );
  BUF_X1 U1151 ( .A(n4318), .Z(n11046) );
  BUF_X1 U1152 ( .A(n2850), .Z(n11310) );
  BUF_X1 U1153 ( .A(n4318), .Z(n11047) );
  BUF_X1 U1154 ( .A(n2850), .Z(n11311) );
  BUF_X1 U1155 ( .A(n4298), .Z(n11079) );
  BUF_X1 U1156 ( .A(n2798), .Z(n11343) );
  BUF_X1 U1157 ( .A(n4298), .Z(n11080) );
  BUF_X1 U1158 ( .A(n2798), .Z(n11344) );
  BUF_X1 U1159 ( .A(n4360), .Z(n10947) );
  BUF_X1 U1160 ( .A(n2924), .Z(n11211) );
  BUF_X1 U1161 ( .A(n4360), .Z(n10948) );
  BUF_X1 U1162 ( .A(n2924), .Z(n11212) );
  BUF_X1 U1163 ( .A(n4307), .Z(n11055) );
  BUF_X1 U1164 ( .A(n2807), .Z(n11319) );
  BUF_X1 U1165 ( .A(n4307), .Z(n11056) );
  BUF_X1 U1166 ( .A(n2807), .Z(n11320) );
  BUF_X1 U1167 ( .A(n4335), .Z(n10998) );
  BUF_X1 U1168 ( .A(n4338), .Z(n10989) );
  BUF_X1 U1169 ( .A(n2867), .Z(n11262) );
  BUF_X1 U1170 ( .A(n2870), .Z(n11253) );
  BUF_X1 U1171 ( .A(n4335), .Z(n10999) );
  BUF_X1 U1172 ( .A(n4338), .Z(n10990) );
  BUF_X1 U1173 ( .A(n2867), .Z(n11263) );
  BUF_X1 U1174 ( .A(n2870), .Z(n11254) );
  BUF_X1 U1175 ( .A(n4361), .Z(n10944) );
  BUF_X1 U1176 ( .A(n2925), .Z(n11208) );
  BUF_X1 U1177 ( .A(n4361), .Z(n10945) );
  BUF_X1 U1178 ( .A(n2925), .Z(n11209) );
  BUF_X1 U1179 ( .A(n4297), .Z(n11082) );
  BUF_X1 U1180 ( .A(n4303), .Z(n11067) );
  BUF_X1 U1181 ( .A(n2797), .Z(n11346) );
  BUF_X1 U1182 ( .A(n2803), .Z(n11331) );
  BUF_X1 U1183 ( .A(n4297), .Z(n11083) );
  BUF_X1 U1184 ( .A(n4303), .Z(n11068) );
  BUF_X1 U1185 ( .A(n2797), .Z(n11347) );
  BUF_X1 U1186 ( .A(n2803), .Z(n11332) );
  BUF_X1 U1187 ( .A(n4334), .Z(n11001) );
  BUF_X1 U1188 ( .A(n2866), .Z(n11265) );
  BUF_X1 U1189 ( .A(n4334), .Z(n11002) );
  BUF_X1 U1190 ( .A(n2866), .Z(n11266) );
  BUF_X1 U1191 ( .A(n4328), .Z(n11016) );
  BUF_X1 U1192 ( .A(n4353), .Z(n10968) );
  BUF_X1 U1193 ( .A(n4356), .Z(n10959) );
  BUF_X1 U1194 ( .A(n4359), .Z(n10950) );
  BUF_X1 U1195 ( .A(n4365), .Z(n10935) );
  BUF_X1 U1196 ( .A(n2860), .Z(n11280) );
  BUF_X1 U1197 ( .A(n2917), .Z(n11232) );
  BUF_X1 U1198 ( .A(n2920), .Z(n11223) );
  BUF_X1 U1199 ( .A(n2923), .Z(n11214) );
  BUF_X1 U1200 ( .A(n2929), .Z(n11199) );
  BUF_X1 U1201 ( .A(n4328), .Z(n11017) );
  BUF_X1 U1202 ( .A(n4353), .Z(n10969) );
  BUF_X1 U1203 ( .A(n4356), .Z(n10960) );
  BUF_X1 U1204 ( .A(n4359), .Z(n10951) );
  BUF_X1 U1205 ( .A(n4365), .Z(n10936) );
  BUF_X1 U1206 ( .A(n2860), .Z(n11281) );
  BUF_X1 U1207 ( .A(n2917), .Z(n11233) );
  BUF_X1 U1208 ( .A(n2920), .Z(n11224) );
  BUF_X1 U1209 ( .A(n2923), .Z(n11215) );
  BUF_X1 U1210 ( .A(n2929), .Z(n11200) );
  BUF_X1 U1211 ( .A(n4295), .Z(n11088) );
  BUF_X1 U1212 ( .A(n4301), .Z(n11073) );
  BUF_X1 U1213 ( .A(n2795), .Z(n11352) );
  BUF_X1 U1214 ( .A(n2801), .Z(n11337) );
  BUF_X1 U1215 ( .A(n4295), .Z(n11089) );
  BUF_X1 U1216 ( .A(n4301), .Z(n11074) );
  BUF_X1 U1217 ( .A(n2795), .Z(n11353) );
  BUF_X1 U1218 ( .A(n2801), .Z(n11338) );
  BUF_X1 U1219 ( .A(n4296), .Z(n11085) );
  BUF_X1 U1220 ( .A(n4302), .Z(n11070) );
  BUF_X1 U1221 ( .A(n2796), .Z(n11349) );
  BUF_X1 U1222 ( .A(n2802), .Z(n11334) );
  BUF_X1 U1223 ( .A(n4296), .Z(n11086) );
  BUF_X1 U1224 ( .A(n4302), .Z(n11071) );
  BUF_X1 U1225 ( .A(n2796), .Z(n11350) );
  BUF_X1 U1226 ( .A(n2802), .Z(n11335) );
  BUF_X1 U1227 ( .A(n4332), .Z(n11007) );
  BUF_X1 U1228 ( .A(n2864), .Z(n11271) );
  BUF_X1 U1229 ( .A(n4332), .Z(n11008) );
  BUF_X1 U1230 ( .A(n2864), .Z(n11272) );
  BUF_X1 U1231 ( .A(n4323), .Z(n11031) );
  BUF_X1 U1232 ( .A(n4326), .Z(n11022) );
  BUF_X1 U1233 ( .A(n4351), .Z(n10974) );
  BUF_X1 U1234 ( .A(n4354), .Z(n10965) );
  BUF_X1 U1235 ( .A(n4363), .Z(n10941) );
  BUF_X1 U1236 ( .A(n2855), .Z(n11295) );
  BUF_X1 U1237 ( .A(n2858), .Z(n11286) );
  BUF_X1 U1238 ( .A(n2915), .Z(n11238) );
  BUF_X1 U1239 ( .A(n2918), .Z(n11229) );
  BUF_X1 U1240 ( .A(n2927), .Z(n11205) );
  BUF_X1 U1241 ( .A(n4323), .Z(n11032) );
  BUF_X1 U1242 ( .A(n4326), .Z(n11023) );
  BUF_X1 U1243 ( .A(n4351), .Z(n10975) );
  BUF_X1 U1244 ( .A(n4354), .Z(n10966) );
  BUF_X1 U1245 ( .A(n4363), .Z(n10942) );
  BUF_X1 U1246 ( .A(n2855), .Z(n11296) );
  BUF_X1 U1247 ( .A(n2858), .Z(n11287) );
  BUF_X1 U1248 ( .A(n2915), .Z(n11239) );
  BUF_X1 U1249 ( .A(n2918), .Z(n11230) );
  BUF_X1 U1250 ( .A(n2927), .Z(n11206) );
  BUF_X1 U1251 ( .A(n4333), .Z(n11004) );
  BUF_X1 U1252 ( .A(n2865), .Z(n11268) );
  BUF_X1 U1253 ( .A(n4333), .Z(n11005) );
  BUF_X1 U1254 ( .A(n2865), .Z(n11269) );
  BUF_X1 U1255 ( .A(n4352), .Z(n10971) );
  BUF_X1 U1256 ( .A(n4355), .Z(n10962) );
  BUF_X1 U1257 ( .A(n4358), .Z(n10953) );
  BUF_X1 U1258 ( .A(n2916), .Z(n11235) );
  BUF_X1 U1259 ( .A(n2919), .Z(n11226) );
  BUF_X1 U1260 ( .A(n2922), .Z(n11217) );
  BUF_X1 U1261 ( .A(n4352), .Z(n10972) );
  BUF_X1 U1262 ( .A(n4355), .Z(n10963) );
  BUF_X1 U1263 ( .A(n4358), .Z(n10954) );
  BUF_X1 U1264 ( .A(n2916), .Z(n11236) );
  BUF_X1 U1265 ( .A(n2919), .Z(n11227) );
  BUF_X1 U1266 ( .A(n2922), .Z(n11218) );
  BUF_X1 U1267 ( .A(n4318), .Z(n11048) );
  BUF_X1 U1268 ( .A(n2850), .Z(n11312) );
  BUF_X1 U1269 ( .A(n4298), .Z(n11081) );
  BUF_X1 U1270 ( .A(n2798), .Z(n11345) );
  BUF_X1 U1271 ( .A(n4360), .Z(n10949) );
  BUF_X1 U1272 ( .A(n2924), .Z(n11213) );
  BUF_X1 U1273 ( .A(n4307), .Z(n11057) );
  BUF_X1 U1274 ( .A(n2807), .Z(n11321) );
  BUF_X1 U1275 ( .A(n4335), .Z(n11000) );
  BUF_X1 U1276 ( .A(n4338), .Z(n10991) );
  BUF_X1 U1277 ( .A(n2867), .Z(n11264) );
  BUF_X1 U1278 ( .A(n2870), .Z(n11255) );
  BUF_X1 U1279 ( .A(n4361), .Z(n10946) );
  BUF_X1 U1280 ( .A(n2925), .Z(n11210) );
  BUF_X1 U1281 ( .A(n4297), .Z(n11084) );
  BUF_X1 U1282 ( .A(n4303), .Z(n11069) );
  BUF_X1 U1283 ( .A(n2797), .Z(n11348) );
  BUF_X1 U1284 ( .A(n2803), .Z(n11333) );
  BUF_X1 U1285 ( .A(n4334), .Z(n11003) );
  BUF_X1 U1286 ( .A(n2866), .Z(n11267) );
  BUF_X1 U1287 ( .A(n4328), .Z(n11018) );
  BUF_X1 U1288 ( .A(n4353), .Z(n10970) );
  BUF_X1 U1289 ( .A(n4356), .Z(n10961) );
  BUF_X1 U1290 ( .A(n4359), .Z(n10952) );
  BUF_X1 U1291 ( .A(n4365), .Z(n10937) );
  BUF_X1 U1292 ( .A(n2860), .Z(n11282) );
  BUF_X1 U1293 ( .A(n2917), .Z(n11234) );
  BUF_X1 U1294 ( .A(n2920), .Z(n11225) );
  BUF_X1 U1295 ( .A(n2923), .Z(n11216) );
  BUF_X1 U1296 ( .A(n2929), .Z(n11201) );
  BUF_X1 U1297 ( .A(n4339), .Z(n10988) );
  BUF_X1 U1298 ( .A(n2871), .Z(n11252) );
  BUF_X1 U1299 ( .A(n4295), .Z(n11090) );
  BUF_X1 U1300 ( .A(n4301), .Z(n11075) );
  BUF_X1 U1301 ( .A(n2795), .Z(n11354) );
  BUF_X1 U1302 ( .A(n2801), .Z(n11339) );
  BUF_X1 U1303 ( .A(n4296), .Z(n11087) );
  BUF_X1 U1304 ( .A(n4302), .Z(n11072) );
  BUF_X1 U1305 ( .A(n2796), .Z(n11351) );
  BUF_X1 U1306 ( .A(n2802), .Z(n11336) );
  BUF_X1 U1307 ( .A(n4332), .Z(n11009) );
  BUF_X1 U1308 ( .A(n2864), .Z(n11273) );
  BUF_X1 U1309 ( .A(n4323), .Z(n11033) );
  BUF_X1 U1310 ( .A(n4326), .Z(n11024) );
  BUF_X1 U1311 ( .A(n4351), .Z(n10976) );
  BUF_X1 U1312 ( .A(n4354), .Z(n10967) );
  BUF_X1 U1313 ( .A(n4363), .Z(n10943) );
  BUF_X1 U1314 ( .A(n2855), .Z(n11297) );
  BUF_X1 U1315 ( .A(n2858), .Z(n11288) );
  BUF_X1 U1316 ( .A(n2915), .Z(n11240) );
  BUF_X1 U1317 ( .A(n2918), .Z(n11231) );
  BUF_X1 U1318 ( .A(n2927), .Z(n11207) );
  BUF_X1 U1319 ( .A(n4333), .Z(n11006) );
  BUF_X1 U1320 ( .A(n2865), .Z(n11270) );
  BUF_X1 U1321 ( .A(n4352), .Z(n10973) );
  BUF_X1 U1322 ( .A(n4355), .Z(n10964) );
  BUF_X1 U1323 ( .A(n4358), .Z(n10955) );
  BUF_X1 U1324 ( .A(n2916), .Z(n11237) );
  BUF_X1 U1325 ( .A(n2919), .Z(n11228) );
  BUF_X1 U1326 ( .A(n2922), .Z(n11219) );
  BUF_X1 U1327 ( .A(n4337), .Z(n10994) );
  BUF_X1 U1328 ( .A(n4340), .Z(n10985) );
  BUF_X1 U1329 ( .A(n2869), .Z(n11258) );
  BUF_X1 U1330 ( .A(n2872), .Z(n11249) );
  BUF_X1 U1331 ( .A(n2490), .Z(n12419) );
  BUF_X1 U1332 ( .A(n2490), .Z(n12420) );
  BUF_X1 U1333 ( .A(n2490), .Z(n12421) );
  BUF_X1 U1334 ( .A(n2490), .Z(n12422) );
  BUF_X1 U1335 ( .A(n2490), .Z(n12423) );
  BUF_X1 U1336 ( .A(n2490), .Z(n12424) );
  BUF_X1 U1337 ( .A(n2490), .Z(n12425) );
  BUF_X1 U1338 ( .A(n12726), .Z(n12728) );
  BUF_X1 U1339 ( .A(n12730), .Z(n12725) );
  BUF_X1 U1340 ( .A(n12724), .Z(n12727) );
  BUF_X1 U1341 ( .A(n12722), .Z(n12726) );
  BUF_X1 U1342 ( .A(n12730), .Z(n12722) );
  BUF_X1 U1343 ( .A(n12730), .Z(n12721) );
  BUF_X1 U1344 ( .A(n12730), .Z(n12723) );
  BUF_X1 U1345 ( .A(n12721), .Z(n12724) );
  BUF_X1 U1346 ( .A(n12728), .Z(n12715) );
  BUF_X1 U1347 ( .A(n12727), .Z(n12716) );
  BUF_X1 U1348 ( .A(n12729), .Z(n12717) );
  BUF_X1 U1349 ( .A(n12714), .Z(n12718) );
  BUF_X1 U1350 ( .A(n12715), .Z(n12719) );
  BUF_X1 U1351 ( .A(n12716), .Z(n12720) );
  BUF_X1 U1352 ( .A(n12729), .Z(n12713) );
  BUF_X1 U1353 ( .A(n12725), .Z(n12714) );
  BUF_X1 U1354 ( .A(n12723), .Z(n12729) );
  NOR2_X1 U1355 ( .A1(n12771), .A2(N8436), .ZN(n5678) );
  NOR2_X1 U1356 ( .A1(n12775), .A2(N8580), .ZN(n4245) );
  NOR2_X1 U1357 ( .A1(n12770), .A2(n12771), .ZN(n5689) );
  NOR2_X1 U1358 ( .A1(n12774), .A2(n12775), .ZN(n4256) );
  AND2_X1 U1359 ( .A1(n2571), .A2(n12733), .ZN(n2574) );
  AND3_X1 U1360 ( .A1(n2615), .A2(n12733), .A3(N2172), .ZN(n2617) );
  AND3_X1 U1361 ( .A1(n12733), .A2(n12732), .A3(n2615), .ZN(n2715) );
  BUF_X1 U1362 ( .A(n4305), .Z(n11061) );
  BUF_X1 U1363 ( .A(n4308), .Z(n11052) );
  BUF_X1 U1364 ( .A(n4336), .Z(n10995) );
  BUF_X1 U1365 ( .A(n4367), .Z(n10929) );
  BUF_X1 U1366 ( .A(n4370), .Z(n10920) );
  BUF_X1 U1367 ( .A(n4398), .Z(n10863) );
  BUF_X1 U1368 ( .A(n4401), .Z(n10854) );
  BUF_X1 U1369 ( .A(n2805), .Z(n11325) );
  BUF_X1 U1370 ( .A(n2808), .Z(n11316) );
  BUF_X1 U1371 ( .A(n2868), .Z(n11259) );
  BUF_X1 U1372 ( .A(n2931), .Z(n11193) );
  BUF_X1 U1373 ( .A(n2934), .Z(n11184) );
  BUF_X1 U1374 ( .A(n2965), .Z(n11127) );
  BUF_X1 U1375 ( .A(n2968), .Z(n11118) );
  BUF_X1 U1376 ( .A(n4305), .Z(n11062) );
  BUF_X1 U1377 ( .A(n4308), .Z(n11053) );
  BUF_X1 U1378 ( .A(n4336), .Z(n10996) );
  BUF_X1 U1379 ( .A(n4367), .Z(n10930) );
  BUF_X1 U1380 ( .A(n4370), .Z(n10921) );
  BUF_X1 U1381 ( .A(n4398), .Z(n10864) );
  BUF_X1 U1382 ( .A(n4401), .Z(n10855) );
  BUF_X1 U1383 ( .A(n2805), .Z(n11326) );
  BUF_X1 U1384 ( .A(n2808), .Z(n11317) );
  BUF_X1 U1385 ( .A(n2868), .Z(n11260) );
  BUF_X1 U1386 ( .A(n2931), .Z(n11194) );
  BUF_X1 U1387 ( .A(n2934), .Z(n11185) );
  BUF_X1 U1388 ( .A(n2965), .Z(n11128) );
  BUF_X1 U1389 ( .A(n2968), .Z(n11119) );
  BUF_X1 U1390 ( .A(n4306), .Z(n11058) );
  BUF_X1 U1391 ( .A(n4309), .Z(n11049) );
  BUF_X1 U1392 ( .A(n4368), .Z(n10926) );
  BUF_X1 U1393 ( .A(n4371), .Z(n10917) );
  BUF_X1 U1394 ( .A(n4399), .Z(n10860) );
  BUF_X1 U1395 ( .A(n4402), .Z(n10851) );
  BUF_X1 U1396 ( .A(n2806), .Z(n11322) );
  BUF_X1 U1397 ( .A(n2809), .Z(n11313) );
  BUF_X1 U1398 ( .A(n2932), .Z(n11190) );
  BUF_X1 U1399 ( .A(n2938), .Z(n11181) );
  BUF_X1 U1400 ( .A(n2966), .Z(n11124) );
  BUF_X1 U1401 ( .A(n2969), .Z(n11115) );
  BUF_X1 U1402 ( .A(n4306), .Z(n11059) );
  BUF_X1 U1403 ( .A(n4309), .Z(n11050) );
  BUF_X1 U1404 ( .A(n4368), .Z(n10927) );
  BUF_X1 U1405 ( .A(n4371), .Z(n10918) );
  BUF_X1 U1406 ( .A(n4399), .Z(n10861) );
  BUF_X1 U1407 ( .A(n4402), .Z(n10852) );
  BUF_X1 U1408 ( .A(n2806), .Z(n11323) );
  BUF_X1 U1409 ( .A(n2809), .Z(n11314) );
  BUF_X1 U1410 ( .A(n2932), .Z(n11191) );
  BUF_X1 U1411 ( .A(n2938), .Z(n11182) );
  BUF_X1 U1412 ( .A(n2966), .Z(n11125) );
  BUF_X1 U1413 ( .A(n2969), .Z(n11116) );
  NAND2_X1 U1414 ( .A1(n5652), .A2(n5655), .ZN(n4297) );
  NAND2_X1 U1415 ( .A1(n5652), .A2(n5657), .ZN(n4295) );
  NAND2_X1 U1416 ( .A1(n5652), .A2(n5656), .ZN(n4296) );
  NAND2_X1 U1417 ( .A1(n5652), .A2(n5659), .ZN(n4303) );
  NAND2_X1 U1418 ( .A1(n5652), .A2(n5661), .ZN(n4301) );
  NAND2_X1 U1419 ( .A1(n5652), .A2(n5660), .ZN(n4302) );
  NAND2_X1 U1420 ( .A1(n4219), .A2(n4222), .ZN(n2797) );
  NAND2_X1 U1421 ( .A1(n4219), .A2(n4224), .ZN(n2795) );
  NAND2_X1 U1422 ( .A1(n4219), .A2(n4223), .ZN(n2796) );
  NAND2_X1 U1423 ( .A1(n4219), .A2(n4226), .ZN(n2803) );
  NAND2_X1 U1424 ( .A1(n4219), .A2(n4228), .ZN(n2801) );
  NAND2_X1 U1425 ( .A1(n4219), .A2(n4227), .ZN(n2802) );
  BUF_X1 U1426 ( .A(n4287), .Z(n11112) );
  BUF_X1 U1427 ( .A(n4349), .Z(n10980) );
  BUF_X1 U1428 ( .A(n4380), .Z(n10914) );
  BUF_X1 U1429 ( .A(n2787), .Z(n11376) );
  BUF_X1 U1430 ( .A(n2881), .Z(n11244) );
  BUF_X1 U1431 ( .A(n2947), .Z(n11178) );
  BUF_X1 U1432 ( .A(n4287), .Z(n11113) );
  BUF_X1 U1433 ( .A(n4349), .Z(n10981) );
  BUF_X1 U1434 ( .A(n4380), .Z(n10915) );
  BUF_X1 U1435 ( .A(n2787), .Z(n11377) );
  BUF_X1 U1436 ( .A(n2881), .Z(n11245) );
  BUF_X1 U1437 ( .A(n2947), .Z(n11179) );
  BUF_X1 U1438 ( .A(n4288), .Z(n11109) );
  BUF_X1 U1439 ( .A(n4319), .Z(n11043) );
  BUF_X1 U1440 ( .A(n4381), .Z(n10911) );
  BUF_X1 U1441 ( .A(n2788), .Z(n11373) );
  BUF_X1 U1442 ( .A(n2851), .Z(n11307) );
  BUF_X1 U1443 ( .A(n2948), .Z(n11175) );
  BUF_X1 U1444 ( .A(n4288), .Z(n11110) );
  BUF_X1 U1445 ( .A(n4319), .Z(n11044) );
  BUF_X1 U1446 ( .A(n4381), .Z(n10912) );
  BUF_X1 U1447 ( .A(n2788), .Z(n11374) );
  BUF_X1 U1448 ( .A(n2851), .Z(n11308) );
  BUF_X1 U1449 ( .A(n2948), .Z(n11176) );
  BUF_X1 U1450 ( .A(n4350), .Z(n10977) );
  BUF_X1 U1451 ( .A(n2914), .Z(n11241) );
  BUF_X1 U1452 ( .A(n4350), .Z(n10978) );
  BUF_X1 U1453 ( .A(n2914), .Z(n11242) );
  AND2_X1 U1454 ( .A1(n2730), .A2(n2717), .ZN(n2491) );
  BUF_X1 U1455 ( .A(n4329), .Z(n11013) );
  BUF_X1 U1456 ( .A(n4391), .Z(n10881) );
  BUF_X1 U1457 ( .A(n2861), .Z(n11277) );
  BUF_X1 U1458 ( .A(n2958), .Z(n11145) );
  BUF_X1 U1459 ( .A(n4329), .Z(n11014) );
  BUF_X1 U1460 ( .A(n4391), .Z(n10882) );
  BUF_X1 U1461 ( .A(n2861), .Z(n11278) );
  BUF_X1 U1462 ( .A(n2958), .Z(n11146) );
  BUF_X1 U1463 ( .A(n4304), .Z(n11064) );
  BUF_X1 U1464 ( .A(n4366), .Z(n10932) );
  BUF_X1 U1465 ( .A(n4369), .Z(n10923) );
  BUF_X1 U1466 ( .A(n4397), .Z(n10866) );
  BUF_X1 U1467 ( .A(n4400), .Z(n10857) );
  BUF_X1 U1468 ( .A(n2804), .Z(n11328) );
  BUF_X1 U1469 ( .A(n2930), .Z(n11196) );
  BUF_X1 U1470 ( .A(n2933), .Z(n11187) );
  BUF_X1 U1471 ( .A(n2964), .Z(n11130) );
  BUF_X1 U1472 ( .A(n2967), .Z(n11121) );
  BUF_X1 U1473 ( .A(n4304), .Z(n11065) );
  BUF_X1 U1474 ( .A(n4366), .Z(n10933) );
  BUF_X1 U1475 ( .A(n4369), .Z(n10924) );
  BUF_X1 U1476 ( .A(n4397), .Z(n10867) );
  BUF_X1 U1477 ( .A(n4400), .Z(n10858) );
  BUF_X1 U1478 ( .A(n2804), .Z(n11329) );
  BUF_X1 U1479 ( .A(n2930), .Z(n11197) );
  BUF_X1 U1480 ( .A(n2933), .Z(n11188) );
  BUF_X1 U1481 ( .A(n2964), .Z(n11131) );
  BUF_X1 U1482 ( .A(n2967), .Z(n11122) );
  BUF_X1 U1483 ( .A(n4299), .Z(n11076) );
  BUF_X1 U1484 ( .A(n4330), .Z(n11010) );
  BUF_X1 U1485 ( .A(n4392), .Z(n10878) );
  BUF_X1 U1486 ( .A(n2799), .Z(n11340) );
  BUF_X1 U1487 ( .A(n2862), .Z(n11274) );
  BUF_X1 U1488 ( .A(n2959), .Z(n11142) );
  BUF_X1 U1489 ( .A(n4299), .Z(n11077) );
  BUF_X1 U1490 ( .A(n4330), .Z(n11011) );
  BUF_X1 U1491 ( .A(n4392), .Z(n10879) );
  BUF_X1 U1492 ( .A(n2799), .Z(n11341) );
  BUF_X1 U1493 ( .A(n2862), .Z(n11275) );
  BUF_X1 U1494 ( .A(n2959), .Z(n11143) );
  BUF_X1 U1495 ( .A(n4390), .Z(n10884) );
  BUF_X1 U1496 ( .A(n4396), .Z(n10869) );
  BUF_X1 U1497 ( .A(n2957), .Z(n11148) );
  BUF_X1 U1498 ( .A(n2963), .Z(n11133) );
  BUF_X1 U1499 ( .A(n4390), .Z(n10885) );
  BUF_X1 U1500 ( .A(n4396), .Z(n10870) );
  BUF_X1 U1501 ( .A(n2957), .Z(n11149) );
  BUF_X1 U1502 ( .A(n2963), .Z(n11134) );
  BUF_X1 U1503 ( .A(n4291), .Z(n11100) );
  BUF_X1 U1504 ( .A(n4322), .Z(n11034) );
  BUF_X1 U1505 ( .A(n2791), .Z(n11364) );
  BUF_X1 U1506 ( .A(n2854), .Z(n11298) );
  BUF_X1 U1507 ( .A(n4291), .Z(n11101) );
  BUF_X1 U1508 ( .A(n4322), .Z(n11035) );
  BUF_X1 U1509 ( .A(n2791), .Z(n11365) );
  BUF_X1 U1510 ( .A(n2854), .Z(n11299) );
  BUF_X1 U1511 ( .A(n4294), .Z(n11091) );
  BUF_X1 U1512 ( .A(n4325), .Z(n11025) );
  BUF_X1 U1513 ( .A(n4384), .Z(n10902) );
  BUF_X1 U1514 ( .A(n4387), .Z(n10893) );
  BUF_X1 U1515 ( .A(n2794), .Z(n11355) );
  BUF_X1 U1516 ( .A(n2857), .Z(n11289) );
  BUF_X1 U1517 ( .A(n2951), .Z(n11166) );
  BUF_X1 U1518 ( .A(n2954), .Z(n11157) );
  BUF_X1 U1519 ( .A(n4294), .Z(n11092) );
  BUF_X1 U1520 ( .A(n4325), .Z(n11026) );
  BUF_X1 U1521 ( .A(n4384), .Z(n10903) );
  BUF_X1 U1522 ( .A(n4387), .Z(n10894) );
  BUF_X1 U1523 ( .A(n2794), .Z(n11356) );
  BUF_X1 U1524 ( .A(n2857), .Z(n11290) );
  BUF_X1 U1525 ( .A(n2951), .Z(n11167) );
  BUF_X1 U1526 ( .A(n2954), .Z(n11158) );
  BUF_X1 U1527 ( .A(n4385), .Z(n10899) );
  BUF_X1 U1528 ( .A(n4388), .Z(n10890) );
  BUF_X1 U1529 ( .A(n2952), .Z(n11163) );
  BUF_X1 U1530 ( .A(n2955), .Z(n11154) );
  BUF_X1 U1531 ( .A(n4385), .Z(n10900) );
  BUF_X1 U1532 ( .A(n4388), .Z(n10891) );
  BUF_X1 U1533 ( .A(n2952), .Z(n11164) );
  BUF_X1 U1534 ( .A(n2955), .Z(n11155) );
  BUF_X1 U1535 ( .A(n4386), .Z(n10896) );
  BUF_X1 U1536 ( .A(n4395), .Z(n10872) );
  BUF_X1 U1537 ( .A(n2953), .Z(n11160) );
  BUF_X1 U1538 ( .A(n2962), .Z(n11136) );
  BUF_X1 U1539 ( .A(n4386), .Z(n10897) );
  BUF_X1 U1540 ( .A(n4395), .Z(n10873) );
  BUF_X1 U1541 ( .A(n2953), .Z(n11161) );
  BUF_X1 U1542 ( .A(n2962), .Z(n11137) );
  BUF_X1 U1543 ( .A(n4389), .Z(n10887) );
  BUF_X1 U1544 ( .A(n2956), .Z(n11151) );
  BUF_X1 U1545 ( .A(n4389), .Z(n10888) );
  BUF_X1 U1546 ( .A(n2956), .Z(n11152) );
  BUF_X1 U1547 ( .A(n4289), .Z(n11106) );
  BUF_X1 U1548 ( .A(n4357), .Z(n10956) );
  BUF_X1 U1549 ( .A(n4394), .Z(n10875) );
  BUF_X1 U1550 ( .A(n2789), .Z(n11370) );
  BUF_X1 U1551 ( .A(n2921), .Z(n11220) );
  BUF_X1 U1552 ( .A(n2961), .Z(n11139) );
  BUF_X1 U1553 ( .A(n4289), .Z(n11107) );
  BUF_X1 U1554 ( .A(n4357), .Z(n10957) );
  BUF_X1 U1555 ( .A(n4394), .Z(n10876) );
  BUF_X1 U1556 ( .A(n2789), .Z(n11371) );
  BUF_X1 U1557 ( .A(n2921), .Z(n11221) );
  BUF_X1 U1558 ( .A(n2961), .Z(n11140) );
  BUF_X1 U1559 ( .A(n4292), .Z(n11097) );
  BUF_X1 U1560 ( .A(n4320), .Z(n11040) );
  BUF_X1 U1561 ( .A(n4382), .Z(n10908) );
  BUF_X1 U1562 ( .A(n2792), .Z(n11361) );
  BUF_X1 U1563 ( .A(n2852), .Z(n11304) );
  BUF_X1 U1564 ( .A(n2949), .Z(n11172) );
  BUF_X1 U1565 ( .A(n4292), .Z(n11098) );
  BUF_X1 U1566 ( .A(n4320), .Z(n11041) );
  BUF_X1 U1567 ( .A(n4382), .Z(n10909) );
  BUF_X1 U1568 ( .A(n2792), .Z(n11362) );
  BUF_X1 U1569 ( .A(n2852), .Z(n11305) );
  BUF_X1 U1570 ( .A(n2949), .Z(n11173) );
  BUF_X1 U1571 ( .A(n4321), .Z(n11037) );
  BUF_X1 U1572 ( .A(n4364), .Z(n10938) );
  BUF_X1 U1573 ( .A(n2853), .Z(n11301) );
  BUF_X1 U1574 ( .A(n2928), .Z(n11202) );
  BUF_X1 U1575 ( .A(n4321), .Z(n11038) );
  BUF_X1 U1576 ( .A(n4364), .Z(n10939) );
  BUF_X1 U1577 ( .A(n2853), .Z(n11302) );
  BUF_X1 U1578 ( .A(n2928), .Z(n11203) );
  BUF_X1 U1579 ( .A(n4290), .Z(n11103) );
  BUF_X1 U1580 ( .A(n4293), .Z(n11094) );
  BUF_X1 U1581 ( .A(n4324), .Z(n11028) );
  BUF_X1 U1582 ( .A(n4327), .Z(n11019) );
  BUF_X1 U1583 ( .A(n4383), .Z(n10905) );
  BUF_X1 U1584 ( .A(n2790), .Z(n11367) );
  BUF_X1 U1585 ( .A(n2793), .Z(n11358) );
  BUF_X1 U1586 ( .A(n2856), .Z(n11292) );
  BUF_X1 U1587 ( .A(n2859), .Z(n11283) );
  BUF_X1 U1588 ( .A(n2950), .Z(n11169) );
  BUF_X1 U1589 ( .A(n4290), .Z(n11104) );
  BUF_X1 U1590 ( .A(n4293), .Z(n11095) );
  BUF_X1 U1591 ( .A(n4324), .Z(n11029) );
  BUF_X1 U1592 ( .A(n4327), .Z(n11020) );
  BUF_X1 U1593 ( .A(n4383), .Z(n10906) );
  BUF_X1 U1594 ( .A(n2790), .Z(n11368) );
  BUF_X1 U1595 ( .A(n2793), .Z(n11359) );
  BUF_X1 U1596 ( .A(n2856), .Z(n11293) );
  BUF_X1 U1597 ( .A(n2859), .Z(n11284) );
  BUF_X1 U1598 ( .A(n2950), .Z(n11170) );
  BUF_X1 U1599 ( .A(n4287), .Z(n11114) );
  BUF_X1 U1600 ( .A(n4349), .Z(n10982) );
  BUF_X1 U1601 ( .A(n2787), .Z(n11378) );
  BUF_X1 U1602 ( .A(n2881), .Z(n11246) );
  BUF_X1 U1603 ( .A(n4380), .Z(n10916) );
  BUF_X1 U1604 ( .A(n2947), .Z(n11180) );
  BUF_X1 U1605 ( .A(n4288), .Z(n11111) );
  BUF_X1 U1606 ( .A(n4319), .Z(n11045) );
  BUF_X1 U1607 ( .A(n2788), .Z(n11375) );
  BUF_X1 U1608 ( .A(n2851), .Z(n11309) );
  BUF_X1 U1609 ( .A(n4381), .Z(n10913) );
  BUF_X1 U1610 ( .A(n2948), .Z(n11177) );
  BUF_X1 U1611 ( .A(n4350), .Z(n10979) );
  BUF_X1 U1612 ( .A(n2914), .Z(n11243) );
  BUF_X1 U1613 ( .A(n4391), .Z(n10883) );
  BUF_X1 U1614 ( .A(n2958), .Z(n11147) );
  BUF_X1 U1615 ( .A(n4329), .Z(n11015) );
  BUF_X1 U1616 ( .A(n2861), .Z(n11279) );
  BUF_X1 U1617 ( .A(n4304), .Z(n11066) );
  BUF_X1 U1618 ( .A(n4366), .Z(n10934) );
  BUF_X1 U1619 ( .A(n4369), .Z(n10925) );
  BUF_X1 U1620 ( .A(n4397), .Z(n10868) );
  BUF_X1 U1621 ( .A(n4400), .Z(n10859) );
  BUF_X1 U1622 ( .A(n2804), .Z(n11330) );
  BUF_X1 U1623 ( .A(n2930), .Z(n11198) );
  BUF_X1 U1624 ( .A(n2933), .Z(n11189) );
  BUF_X1 U1625 ( .A(n2964), .Z(n11132) );
  BUF_X1 U1626 ( .A(n2967), .Z(n11123) );
  BUF_X1 U1627 ( .A(n4299), .Z(n11078) );
  BUF_X1 U1628 ( .A(n4330), .Z(n11012) );
  BUF_X1 U1629 ( .A(n4392), .Z(n10880) );
  BUF_X1 U1630 ( .A(n2799), .Z(n11342) );
  BUF_X1 U1631 ( .A(n2862), .Z(n11276) );
  BUF_X1 U1632 ( .A(n2959), .Z(n11144) );
  BUF_X1 U1633 ( .A(n4390), .Z(n10886) );
  BUF_X1 U1634 ( .A(n4396), .Z(n10871) );
  BUF_X1 U1635 ( .A(n2957), .Z(n11150) );
  BUF_X1 U1636 ( .A(n2963), .Z(n11135) );
  BUF_X1 U1637 ( .A(n4291), .Z(n11102) );
  BUF_X1 U1638 ( .A(n4322), .Z(n11036) );
  BUF_X1 U1639 ( .A(n2791), .Z(n11366) );
  BUF_X1 U1640 ( .A(n2854), .Z(n11300) );
  BUF_X1 U1641 ( .A(n4294), .Z(n11093) );
  BUF_X1 U1642 ( .A(n4325), .Z(n11027) );
  BUF_X1 U1643 ( .A(n4384), .Z(n10904) );
  BUF_X1 U1644 ( .A(n4387), .Z(n10895) );
  BUF_X1 U1645 ( .A(n2794), .Z(n11357) );
  BUF_X1 U1646 ( .A(n2857), .Z(n11291) );
  BUF_X1 U1647 ( .A(n2951), .Z(n11168) );
  BUF_X1 U1648 ( .A(n2954), .Z(n11159) );
  BUF_X1 U1649 ( .A(n4305), .Z(n11063) );
  BUF_X1 U1650 ( .A(n4308), .Z(n11054) );
  BUF_X1 U1651 ( .A(n4336), .Z(n10997) );
  BUF_X1 U1652 ( .A(n4367), .Z(n10931) );
  BUF_X1 U1653 ( .A(n4370), .Z(n10922) );
  BUF_X1 U1654 ( .A(n4398), .Z(n10865) );
  BUF_X1 U1655 ( .A(n4401), .Z(n10856) );
  BUF_X1 U1656 ( .A(n2805), .Z(n11327) );
  BUF_X1 U1657 ( .A(n2808), .Z(n11318) );
  BUF_X1 U1658 ( .A(n2868), .Z(n11261) );
  BUF_X1 U1659 ( .A(n2931), .Z(n11195) );
  BUF_X1 U1660 ( .A(n2934), .Z(n11186) );
  BUF_X1 U1661 ( .A(n2965), .Z(n11129) );
  BUF_X1 U1662 ( .A(n2968), .Z(n11120) );
  BUF_X1 U1663 ( .A(n4385), .Z(n10901) );
  BUF_X1 U1664 ( .A(n4388), .Z(n10892) );
  BUF_X1 U1665 ( .A(n2952), .Z(n11165) );
  BUF_X1 U1666 ( .A(n2955), .Z(n11156) );
  BUF_X1 U1667 ( .A(n4386), .Z(n10898) );
  BUF_X1 U1668 ( .A(n4395), .Z(n10874) );
  BUF_X1 U1669 ( .A(n2953), .Z(n11162) );
  BUF_X1 U1670 ( .A(n2962), .Z(n11138) );
  BUF_X1 U1671 ( .A(n4389), .Z(n10889) );
  BUF_X1 U1672 ( .A(n2956), .Z(n11153) );
  BUF_X1 U1673 ( .A(n4357), .Z(n10958) );
  BUF_X1 U1674 ( .A(n4394), .Z(n10877) );
  BUF_X1 U1675 ( .A(n2921), .Z(n11222) );
  BUF_X1 U1676 ( .A(n2961), .Z(n11141) );
  BUF_X1 U1677 ( .A(n4289), .Z(n11108) );
  BUF_X1 U1678 ( .A(n2789), .Z(n11372) );
  BUF_X1 U1679 ( .A(n4292), .Z(n11099) );
  BUF_X1 U1680 ( .A(n4320), .Z(n11042) );
  BUF_X1 U1681 ( .A(n4382), .Z(n10910) );
  BUF_X1 U1682 ( .A(n2792), .Z(n11363) );
  BUF_X1 U1683 ( .A(n2852), .Z(n11306) );
  BUF_X1 U1684 ( .A(n2949), .Z(n11174) );
  BUF_X1 U1685 ( .A(n4364), .Z(n10940) );
  BUF_X1 U1686 ( .A(n2928), .Z(n11204) );
  BUF_X1 U1687 ( .A(n4321), .Z(n11039) );
  BUF_X1 U1688 ( .A(n2853), .Z(n11303) );
  BUF_X1 U1689 ( .A(n4290), .Z(n11105) );
  BUF_X1 U1690 ( .A(n4293), .Z(n11096) );
  BUF_X1 U1691 ( .A(n4324), .Z(n11030) );
  BUF_X1 U1692 ( .A(n4327), .Z(n11021) );
  BUF_X1 U1693 ( .A(n4383), .Z(n10907) );
  BUF_X1 U1694 ( .A(n2790), .Z(n11369) );
  BUF_X1 U1695 ( .A(n2793), .Z(n11360) );
  BUF_X1 U1696 ( .A(n2856), .Z(n11294) );
  BUF_X1 U1697 ( .A(n2859), .Z(n11285) );
  BUF_X1 U1698 ( .A(n2950), .Z(n11171) );
  AND2_X1 U1699 ( .A1(n2725), .A2(n2717), .ZN(n2582) );
  BUF_X1 U1700 ( .A(n4306), .Z(n11060) );
  BUF_X1 U1701 ( .A(n4309), .Z(n11051) );
  BUF_X1 U1702 ( .A(n4368), .Z(n10928) );
  BUF_X1 U1703 ( .A(n4371), .Z(n10919) );
  BUF_X1 U1704 ( .A(n4399), .Z(n10862) );
  BUF_X1 U1705 ( .A(n4402), .Z(n10853) );
  BUF_X1 U1706 ( .A(n2806), .Z(n11324) );
  BUF_X1 U1707 ( .A(n2809), .Z(n11315) );
  BUF_X1 U1708 ( .A(n2932), .Z(n11192) );
  BUF_X1 U1709 ( .A(n2938), .Z(n11183) );
  BUF_X1 U1710 ( .A(n2966), .Z(n11126) );
  BUF_X1 U1711 ( .A(n2969), .Z(n11117) );
  NAND2_X1 U1712 ( .A1(n5678), .A2(n5655), .ZN(n4334) );
  NAND2_X1 U1713 ( .A1(n5678), .A2(n5657), .ZN(n4332) );
  NAND2_X1 U1714 ( .A1(n5678), .A2(n5656), .ZN(n4333) );
  NAND2_X1 U1715 ( .A1(n4245), .A2(n4222), .ZN(n2866) );
  NAND2_X1 U1716 ( .A1(n4245), .A2(n4224), .ZN(n2864) );
  NAND2_X1 U1717 ( .A1(n4245), .A2(n4223), .ZN(n2865) );
  NAND2_X1 U1718 ( .A1(n2491), .A2(n2492), .ZN(n2490) );
  AND2_X1 U1719 ( .A1(n5652), .A2(n5653), .ZN(n5646) );
  AND2_X1 U1720 ( .A1(n4219), .A2(n4220), .ZN(n4213) );
  INV_X1 U1721 ( .A(N8436), .ZN(n12770) );
  INV_X1 U1722 ( .A(N8580), .ZN(n12774) );
  INV_X1 U1723 ( .A(N2172), .ZN(n12732) );
  AND2_X1 U1724 ( .A1(n5653), .A2(n5701), .ZN(n5690) );
  AND2_X1 U1725 ( .A1(n4220), .A2(n4268), .ZN(n4257) );
  AND2_X1 U1726 ( .A1(n5675), .A2(n5653), .ZN(n5674) );
  AND2_X1 U1727 ( .A1(n4242), .A2(n4220), .ZN(n4241) );
  NAND2_X1 U1728 ( .A1(n5689), .A2(n5655), .ZN(n4353) );
  NAND2_X1 U1729 ( .A1(n5689), .A2(n5656), .ZN(n4351) );
  NAND2_X1 U1730 ( .A1(n5689), .A2(n5657), .ZN(n4352) );
  NAND2_X1 U1731 ( .A1(n5689), .A2(n5663), .ZN(n4356) );
  NAND2_X1 U1732 ( .A1(n5689), .A2(n5661), .ZN(n4354) );
  NAND2_X1 U1733 ( .A1(n5689), .A2(n5659), .ZN(n4355) );
  NAND2_X1 U1734 ( .A1(n5689), .A2(n5665), .ZN(n4359) );
  NAND2_X1 U1735 ( .A1(n5689), .A2(n5660), .ZN(n4358) );
  NAND2_X1 U1736 ( .A1(n4256), .A2(n4222), .ZN(n2917) );
  NAND2_X1 U1737 ( .A1(n4256), .A2(n4223), .ZN(n2915) );
  NAND2_X1 U1738 ( .A1(n4256), .A2(n4224), .ZN(n2916) );
  NAND2_X1 U1739 ( .A1(n4256), .A2(n4230), .ZN(n2920) );
  NAND2_X1 U1740 ( .A1(n4256), .A2(n4228), .ZN(n2918) );
  NAND2_X1 U1741 ( .A1(n4256), .A2(n4226), .ZN(n2919) );
  NAND2_X1 U1742 ( .A1(n4256), .A2(n4232), .ZN(n2923) );
  NAND2_X1 U1743 ( .A1(n4256), .A2(n4227), .ZN(n2922) );
  NAND2_X1 U1744 ( .A1(n5675), .A2(n5655), .ZN(n4323) );
  NAND2_X1 U1745 ( .A1(n5675), .A2(n5657), .ZN(n4328) );
  NAND2_X1 U1746 ( .A1(n5675), .A2(n5663), .ZN(n4326) );
  NAND2_X1 U1747 ( .A1(n5675), .A2(n5656), .ZN(n4318) );
  NAND2_X1 U1748 ( .A1(n5675), .A2(n5661), .ZN(n4365) );
  NAND2_X1 U1749 ( .A1(n5675), .A2(n5665), .ZN(n4363) );
  NAND2_X1 U1750 ( .A1(n4242), .A2(n4222), .ZN(n2855) );
  NAND2_X1 U1751 ( .A1(n4242), .A2(n4224), .ZN(n2860) );
  NAND2_X1 U1752 ( .A1(n4242), .A2(n4230), .ZN(n2858) );
  NAND2_X1 U1753 ( .A1(n4242), .A2(n4223), .ZN(n2850) );
  NAND2_X1 U1754 ( .A1(n4242), .A2(n4228), .ZN(n2929) );
  NAND2_X1 U1755 ( .A1(n4242), .A2(n4232), .ZN(n2927) );
  AND2_X1 U1756 ( .A1(n5652), .A2(n5665), .ZN(n4307) );
  AND2_X1 U1757 ( .A1(n5652), .A2(n5663), .ZN(n4298) );
  AND2_X1 U1758 ( .A1(n4219), .A2(n4232), .ZN(n2807) );
  AND2_X1 U1759 ( .A1(n4219), .A2(n4230), .ZN(n2798) );
  AND3_X1 U1760 ( .A1(n5653), .A2(n12769), .A3(n5678), .ZN(n5664) );
  AND3_X1 U1761 ( .A1(n4220), .A2(n12773), .A3(n4245), .ZN(n4231) );
  AND2_X1 U1762 ( .A1(n5678), .A2(n5661), .ZN(n4335) );
  AND2_X1 U1763 ( .A1(n5678), .A2(n5663), .ZN(n4338) );
  AND2_X1 U1764 ( .A1(n4245), .A2(n4228), .ZN(n2867) );
  AND2_X1 U1765 ( .A1(n4245), .A2(n4230), .ZN(n2870) );
  AND2_X1 U1766 ( .A1(n5689), .A2(n5653), .ZN(n5687) );
  AND2_X1 U1767 ( .A1(n4256), .A2(n4220), .ZN(n4254) );
  AND2_X1 U1768 ( .A1(n5675), .A2(n5660), .ZN(n4360) );
  AND2_X1 U1769 ( .A1(n5675), .A2(n5659), .ZN(n4361) );
  AND2_X1 U1770 ( .A1(n4242), .A2(n4227), .ZN(n2924) );
  AND2_X1 U1771 ( .A1(n4242), .A2(n4226), .ZN(n2925) );
  AND2_X1 U1772 ( .A1(n5678), .A2(n5665), .ZN(n4337) );
  AND2_X1 U1773 ( .A1(n5678), .A2(n5660), .ZN(n4339) );
  AND2_X1 U1774 ( .A1(n5678), .A2(n5659), .ZN(n4340) );
  AND2_X1 U1775 ( .A1(n4245), .A2(n4232), .ZN(n2869) );
  AND2_X1 U1776 ( .A1(n4245), .A2(n4227), .ZN(n2871) );
  AND2_X1 U1777 ( .A1(n4245), .A2(n4226), .ZN(n2872) );
  INV_X1 U1778 ( .A(n12432), .ZN(n12730) );
  OAI22_X1 U1779 ( .A1(n10844), .A2(n12293), .B1(n12294), .B2(n14256), .ZN(
        n8779) );
  OAI22_X1 U1780 ( .A1(n10837), .A2(n12293), .B1(n12294), .B2(n14255), .ZN(
        n8778) );
  OAI22_X1 U1781 ( .A1(n10830), .A2(n12293), .B1(n12294), .B2(n14254), .ZN(
        n8777) );
  OAI22_X1 U1782 ( .A1(n10823), .A2(n12293), .B1(n12294), .B2(n14253), .ZN(
        n8776) );
  OAI22_X1 U1783 ( .A1(n10816), .A2(n12293), .B1(n12295), .B2(n14252), .ZN(
        n8775) );
  OAI22_X1 U1784 ( .A1(n10809), .A2(n12293), .B1(n12295), .B2(n14251), .ZN(
        n8774) );
  OAI22_X1 U1785 ( .A1(n10802), .A2(n12293), .B1(n12295), .B2(n14250), .ZN(
        n8773) );
  OAI22_X1 U1786 ( .A1(n10795), .A2(n12293), .B1(n12295), .B2(n14249), .ZN(
        n8772) );
  OAI22_X1 U1787 ( .A1(n10788), .A2(n12292), .B1(n12296), .B2(n14248), .ZN(
        n8771) );
  OAI22_X1 U1788 ( .A1(n10781), .A2(n12292), .B1(n12296), .B2(n14247), .ZN(
        n8770) );
  OAI22_X1 U1789 ( .A1(n10774), .A2(n12292), .B1(n12296), .B2(n14246), .ZN(
        n8769) );
  OAI22_X1 U1790 ( .A1(n10767), .A2(n12292), .B1(n12296), .B2(n14245), .ZN(
        n8768) );
  OAI22_X1 U1791 ( .A1(n10760), .A2(n12292), .B1(n12297), .B2(n14244), .ZN(
        n8767) );
  OAI22_X1 U1792 ( .A1(n10753), .A2(n12292), .B1(n12297), .B2(n14243), .ZN(
        n8766) );
  OAI22_X1 U1793 ( .A1(n10746), .A2(n12292), .B1(n12297), .B2(n14242), .ZN(
        n8765) );
  OAI22_X1 U1794 ( .A1(n10739), .A2(n12292), .B1(n12297), .B2(n14241), .ZN(
        n8764) );
  OAI22_X1 U1795 ( .A1(n10732), .A2(n12292), .B1(n12298), .B2(n14240), .ZN(
        n8763) );
  OAI22_X1 U1796 ( .A1(n10725), .A2(n12292), .B1(n12298), .B2(n14239), .ZN(
        n8762) );
  OAI22_X1 U1797 ( .A1(n10718), .A2(n12292), .B1(n12298), .B2(n14238), .ZN(
        n8761) );
  OAI22_X1 U1798 ( .A1(n10711), .A2(n12292), .B1(n12298), .B2(n14237), .ZN(
        n8760) );
  OAI22_X1 U1799 ( .A1(n10704), .A2(n12291), .B1(n12299), .B2(n14236), .ZN(
        n8759) );
  OAI22_X1 U1800 ( .A1(n10697), .A2(n12291), .B1(n12299), .B2(n14235), .ZN(
        n8758) );
  OAI22_X1 U1801 ( .A1(n10690), .A2(n12291), .B1(n12299), .B2(n14234), .ZN(
        n8757) );
  OAI22_X1 U1802 ( .A1(n10683), .A2(n12291), .B1(n12299), .B2(n14233), .ZN(
        n8756) );
  OAI22_X1 U1803 ( .A1(n10676), .A2(n12291), .B1(n12300), .B2(n14232), .ZN(
        n8755) );
  OAI22_X1 U1804 ( .A1(n10669), .A2(n12291), .B1(n12300), .B2(n14231), .ZN(
        n8754) );
  OAI22_X1 U1805 ( .A1(n10662), .A2(n12291), .B1(n12300), .B2(n14230), .ZN(
        n8753) );
  OAI22_X1 U1806 ( .A1(n10655), .A2(n12291), .B1(n12300), .B2(n14229), .ZN(
        n8752) );
  OAI22_X1 U1807 ( .A1(n10648), .A2(n12291), .B1(n12301), .B2(n14228), .ZN(
        n8751) );
  OAI22_X1 U1808 ( .A1(n10641), .A2(n12291), .B1(n12301), .B2(n14227), .ZN(
        n8750) );
  OAI22_X1 U1809 ( .A1(n10634), .A2(n12291), .B1(n12301), .B2(n14226), .ZN(
        n8749) );
  OAI22_X1 U1810 ( .A1(n10627), .A2(n12291), .B1(n12301), .B2(n14225), .ZN(
        n8748) );
  OAI22_X1 U1811 ( .A1(n10845), .A2(n12269), .B1(n12274), .B2(n14224), .ZN(
        n8715) );
  OAI22_X1 U1812 ( .A1(n10838), .A2(n12269), .B1(n12270), .B2(n14223), .ZN(
        n8714) );
  OAI22_X1 U1813 ( .A1(n10831), .A2(n12269), .B1(n12270), .B2(n14222), .ZN(
        n8713) );
  OAI22_X1 U1814 ( .A1(n10824), .A2(n12269), .B1(n12270), .B2(n14221), .ZN(
        n8712) );
  OAI22_X1 U1815 ( .A1(n10817), .A2(n12269), .B1(n12271), .B2(n14220), .ZN(
        n8711) );
  OAI22_X1 U1816 ( .A1(n10810), .A2(n12269), .B1(n12271), .B2(n14219), .ZN(
        n8710) );
  OAI22_X1 U1817 ( .A1(n10803), .A2(n12269), .B1(n12271), .B2(n14218), .ZN(
        n8709) );
  OAI22_X1 U1818 ( .A1(n10796), .A2(n12269), .B1(n12271), .B2(n14217), .ZN(
        n8708) );
  OAI22_X1 U1819 ( .A1(n10789), .A2(n12268), .B1(n12272), .B2(n14216), .ZN(
        n8707) );
  OAI22_X1 U1820 ( .A1(n10782), .A2(n12268), .B1(n12272), .B2(n14215), .ZN(
        n8706) );
  OAI22_X1 U1821 ( .A1(n10775), .A2(n12268), .B1(n12272), .B2(n14214), .ZN(
        n8705) );
  OAI22_X1 U1822 ( .A1(n10768), .A2(n12268), .B1(n12272), .B2(n14213), .ZN(
        n8704) );
  OAI22_X1 U1823 ( .A1(n10761), .A2(n12268), .B1(n12273), .B2(n14212), .ZN(
        n8703) );
  OAI22_X1 U1824 ( .A1(n10754), .A2(n12268), .B1(n12273), .B2(n14211), .ZN(
        n8702) );
  OAI22_X1 U1825 ( .A1(n10747), .A2(n12268), .B1(n12273), .B2(n14210), .ZN(
        n8701) );
  OAI22_X1 U1826 ( .A1(n10740), .A2(n12268), .B1(n12273), .B2(n14209), .ZN(
        n8700) );
  OAI22_X1 U1827 ( .A1(n10733), .A2(n12268), .B1(n12274), .B2(n14208), .ZN(
        n8699) );
  OAI22_X1 U1828 ( .A1(n10726), .A2(n12268), .B1(n12274), .B2(n14207), .ZN(
        n8698) );
  OAI22_X1 U1829 ( .A1(n10719), .A2(n12268), .B1(n12274), .B2(n14206), .ZN(
        n8697) );
  OAI22_X1 U1830 ( .A1(n10712), .A2(n12268), .B1(n12275), .B2(n14205), .ZN(
        n8696) );
  OAI22_X1 U1831 ( .A1(n10705), .A2(n12267), .B1(n12275), .B2(n14204), .ZN(
        n8695) );
  OAI22_X1 U1832 ( .A1(n10698), .A2(n12267), .B1(n12275), .B2(n14203), .ZN(
        n8694) );
  OAI22_X1 U1833 ( .A1(n10691), .A2(n12267), .B1(n12275), .B2(n14202), .ZN(
        n8693) );
  OAI22_X1 U1834 ( .A1(n10684), .A2(n12267), .B1(n12276), .B2(n14201), .ZN(
        n8692) );
  OAI22_X1 U1835 ( .A1(n10677), .A2(n12267), .B1(n12276), .B2(n14200), .ZN(
        n8691) );
  OAI22_X1 U1836 ( .A1(n10670), .A2(n12267), .B1(n12276), .B2(n14199), .ZN(
        n8690) );
  OAI22_X1 U1837 ( .A1(n10663), .A2(n12267), .B1(n12276), .B2(n14198), .ZN(
        n8689) );
  OAI22_X1 U1838 ( .A1(n10656), .A2(n12267), .B1(n12277), .B2(n14197), .ZN(
        n8688) );
  OAI22_X1 U1839 ( .A1(n10649), .A2(n12267), .B1(n12277), .B2(n14196), .ZN(
        n8687) );
  OAI22_X1 U1840 ( .A1(n10642), .A2(n12267), .B1(n12277), .B2(n14195), .ZN(
        n8686) );
  OAI22_X1 U1841 ( .A1(n10635), .A2(n12267), .B1(n12277), .B2(n14194), .ZN(
        n8685) );
  OAI22_X1 U1842 ( .A1(n10845), .A2(n12257), .B1(n12258), .B2(n14193), .ZN(
        n8683) );
  OAI22_X1 U1843 ( .A1(n10838), .A2(n12257), .B1(n12258), .B2(n14192), .ZN(
        n8682) );
  OAI22_X1 U1844 ( .A1(n10831), .A2(n12257), .B1(n12258), .B2(n14191), .ZN(
        n8681) );
  OAI22_X1 U1845 ( .A1(n10824), .A2(n12257), .B1(n12258), .B2(n14190), .ZN(
        n8680) );
  OAI22_X1 U1846 ( .A1(n10817), .A2(n12257), .B1(n12259), .B2(n14189), .ZN(
        n8679) );
  OAI22_X1 U1847 ( .A1(n10810), .A2(n12257), .B1(n12259), .B2(n14188), .ZN(
        n8678) );
  OAI22_X1 U1848 ( .A1(n10803), .A2(n12257), .B1(n12259), .B2(n14187), .ZN(
        n8677) );
  OAI22_X1 U1849 ( .A1(n10796), .A2(n12257), .B1(n12259), .B2(n14186), .ZN(
        n8676) );
  OAI22_X1 U1850 ( .A1(n10789), .A2(n12256), .B1(n12260), .B2(n14185), .ZN(
        n8675) );
  OAI22_X1 U1851 ( .A1(n10782), .A2(n12256), .B1(n12260), .B2(n14184), .ZN(
        n8674) );
  OAI22_X1 U1852 ( .A1(n10775), .A2(n12256), .B1(n12260), .B2(n14183), .ZN(
        n8673) );
  OAI22_X1 U1853 ( .A1(n10768), .A2(n12256), .B1(n12260), .B2(n14182), .ZN(
        n8672) );
  OAI22_X1 U1854 ( .A1(n10761), .A2(n12256), .B1(n12261), .B2(n14181), .ZN(
        n8671) );
  OAI22_X1 U1855 ( .A1(n10754), .A2(n12256), .B1(n12261), .B2(n14180), .ZN(
        n8670) );
  OAI22_X1 U1856 ( .A1(n10747), .A2(n12256), .B1(n12261), .B2(n14179), .ZN(
        n8669) );
  OAI22_X1 U1857 ( .A1(n10740), .A2(n12256), .B1(n12261), .B2(n14178), .ZN(
        n8668) );
  OAI22_X1 U1858 ( .A1(n10733), .A2(n12256), .B1(n12262), .B2(n14177), .ZN(
        n8667) );
  OAI22_X1 U1859 ( .A1(n10726), .A2(n12256), .B1(n12262), .B2(n14176), .ZN(
        n8666) );
  OAI22_X1 U1860 ( .A1(n10719), .A2(n12256), .B1(n12262), .B2(n14175), .ZN(
        n8665) );
  OAI22_X1 U1861 ( .A1(n10712), .A2(n12256), .B1(n12262), .B2(n14174), .ZN(
        n8664) );
  OAI22_X1 U1862 ( .A1(n10705), .A2(n12255), .B1(n12263), .B2(n14173), .ZN(
        n8663) );
  OAI22_X1 U1863 ( .A1(n10698), .A2(n12255), .B1(n12263), .B2(n14172), .ZN(
        n8662) );
  OAI22_X1 U1864 ( .A1(n10691), .A2(n12255), .B1(n12263), .B2(n14171), .ZN(
        n8661) );
  OAI22_X1 U1865 ( .A1(n10684), .A2(n12255), .B1(n12263), .B2(n14170), .ZN(
        n8660) );
  OAI22_X1 U1866 ( .A1(n10677), .A2(n12255), .B1(n12264), .B2(n14169), .ZN(
        n8659) );
  OAI22_X1 U1867 ( .A1(n10670), .A2(n12255), .B1(n12264), .B2(n14168), .ZN(
        n8658) );
  OAI22_X1 U1868 ( .A1(n10663), .A2(n12255), .B1(n12264), .B2(n14167), .ZN(
        n8657) );
  OAI22_X1 U1869 ( .A1(n10656), .A2(n12255), .B1(n12264), .B2(n14166), .ZN(
        n8656) );
  OAI22_X1 U1870 ( .A1(n10649), .A2(n12255), .B1(n12265), .B2(n14165), .ZN(
        n8655) );
  OAI22_X1 U1871 ( .A1(n10642), .A2(n12255), .B1(n12265), .B2(n14164), .ZN(
        n8654) );
  OAI22_X1 U1872 ( .A1(n10635), .A2(n12255), .B1(n12265), .B2(n14163), .ZN(
        n8653) );
  OAI22_X1 U1873 ( .A1(n10628), .A2(n12255), .B1(n12265), .B2(n14162), .ZN(
        n8652) );
  OAI22_X1 U1874 ( .A1(n10845), .A2(n12245), .B1(n12246), .B2(n14161), .ZN(
        n8651) );
  OAI22_X1 U1875 ( .A1(n10838), .A2(n12245), .B1(n12246), .B2(n14160), .ZN(
        n8650) );
  OAI22_X1 U1876 ( .A1(n10831), .A2(n12245), .B1(n12246), .B2(n14159), .ZN(
        n8649) );
  OAI22_X1 U1877 ( .A1(n10824), .A2(n12245), .B1(n12246), .B2(n14158), .ZN(
        n8648) );
  OAI22_X1 U1878 ( .A1(n10817), .A2(n12245), .B1(n12247), .B2(n14157), .ZN(
        n8647) );
  OAI22_X1 U1879 ( .A1(n10810), .A2(n12245), .B1(n12247), .B2(n14156), .ZN(
        n8646) );
  OAI22_X1 U1880 ( .A1(n10803), .A2(n12245), .B1(n12247), .B2(n14155), .ZN(
        n8645) );
  OAI22_X1 U1881 ( .A1(n10796), .A2(n12245), .B1(n12247), .B2(n14154), .ZN(
        n8644) );
  OAI22_X1 U1882 ( .A1(n10789), .A2(n12244), .B1(n12248), .B2(n14153), .ZN(
        n8643) );
  OAI22_X1 U1883 ( .A1(n10782), .A2(n12244), .B1(n12248), .B2(n14152), .ZN(
        n8642) );
  OAI22_X1 U1884 ( .A1(n10775), .A2(n12244), .B1(n12248), .B2(n14151), .ZN(
        n8641) );
  OAI22_X1 U1885 ( .A1(n10768), .A2(n12244), .B1(n12248), .B2(n14150), .ZN(
        n8640) );
  OAI22_X1 U1886 ( .A1(n10761), .A2(n12244), .B1(n12249), .B2(n14149), .ZN(
        n8639) );
  OAI22_X1 U1887 ( .A1(n10754), .A2(n12244), .B1(n12249), .B2(n14148), .ZN(
        n8638) );
  OAI22_X1 U1888 ( .A1(n10747), .A2(n12244), .B1(n12249), .B2(n14147), .ZN(
        n8637) );
  OAI22_X1 U1889 ( .A1(n10740), .A2(n12244), .B1(n12249), .B2(n14146), .ZN(
        n8636) );
  OAI22_X1 U1890 ( .A1(n10733), .A2(n12244), .B1(n12250), .B2(n14145), .ZN(
        n8635) );
  OAI22_X1 U1891 ( .A1(n10726), .A2(n12244), .B1(n12250), .B2(n14144), .ZN(
        n8634) );
  OAI22_X1 U1892 ( .A1(n10719), .A2(n12244), .B1(n12250), .B2(n14143), .ZN(
        n8633) );
  OAI22_X1 U1893 ( .A1(n10712), .A2(n12244), .B1(n12250), .B2(n14142), .ZN(
        n8632) );
  OAI22_X1 U1894 ( .A1(n10705), .A2(n12243), .B1(n12251), .B2(n14141), .ZN(
        n8631) );
  OAI22_X1 U1895 ( .A1(n10698), .A2(n12243), .B1(n12251), .B2(n14140), .ZN(
        n8630) );
  OAI22_X1 U1896 ( .A1(n10691), .A2(n12243), .B1(n12251), .B2(n14139), .ZN(
        n8629) );
  OAI22_X1 U1897 ( .A1(n10684), .A2(n12243), .B1(n12251), .B2(n14138), .ZN(
        n8628) );
  OAI22_X1 U1898 ( .A1(n10677), .A2(n12243), .B1(n12252), .B2(n14137), .ZN(
        n8627) );
  OAI22_X1 U1899 ( .A1(n10670), .A2(n12243), .B1(n12252), .B2(n14136), .ZN(
        n8626) );
  OAI22_X1 U1900 ( .A1(n10663), .A2(n12243), .B1(n12252), .B2(n14135), .ZN(
        n8625) );
  OAI22_X1 U1901 ( .A1(n10656), .A2(n12243), .B1(n12252), .B2(n14134), .ZN(
        n8624) );
  OAI22_X1 U1902 ( .A1(n10649), .A2(n12243), .B1(n12253), .B2(n14133), .ZN(
        n8623) );
  OAI22_X1 U1903 ( .A1(n10642), .A2(n12243), .B1(n12253), .B2(n14132), .ZN(
        n8622) );
  OAI22_X1 U1904 ( .A1(n10635), .A2(n12243), .B1(n12253), .B2(n14131), .ZN(
        n8621) );
  OAI22_X1 U1905 ( .A1(n10628), .A2(n12243), .B1(n12253), .B2(n14130), .ZN(
        n8620) );
  OAI22_X1 U1906 ( .A1(n10845), .A2(n12233), .B1(n12238), .B2(n14129), .ZN(
        n8619) );
  OAI22_X1 U1907 ( .A1(n10838), .A2(n12233), .B1(n12234), .B2(n14128), .ZN(
        n8618) );
  OAI22_X1 U1908 ( .A1(n10831), .A2(n12233), .B1(n12234), .B2(n14127), .ZN(
        n8617) );
  OAI22_X1 U1909 ( .A1(n10824), .A2(n12233), .B1(n12234), .B2(n14126), .ZN(
        n8616) );
  OAI22_X1 U1910 ( .A1(n10817), .A2(n12233), .B1(n12235), .B2(n14125), .ZN(
        n8615) );
  OAI22_X1 U1911 ( .A1(n10810), .A2(n12233), .B1(n12235), .B2(n14124), .ZN(
        n8614) );
  OAI22_X1 U1912 ( .A1(n10803), .A2(n12233), .B1(n12235), .B2(n14123), .ZN(
        n8613) );
  OAI22_X1 U1913 ( .A1(n10796), .A2(n12233), .B1(n12235), .B2(n14122), .ZN(
        n8612) );
  OAI22_X1 U1914 ( .A1(n10789), .A2(n12232), .B1(n12236), .B2(n14121), .ZN(
        n8611) );
  OAI22_X1 U1915 ( .A1(n10782), .A2(n12232), .B1(n12236), .B2(n14120), .ZN(
        n8610) );
  OAI22_X1 U1916 ( .A1(n10775), .A2(n12232), .B1(n12236), .B2(n14119), .ZN(
        n8609) );
  OAI22_X1 U1917 ( .A1(n10768), .A2(n12232), .B1(n12236), .B2(n14118), .ZN(
        n8608) );
  OAI22_X1 U1918 ( .A1(n10761), .A2(n12232), .B1(n12237), .B2(n14117), .ZN(
        n8607) );
  OAI22_X1 U1919 ( .A1(n10754), .A2(n12232), .B1(n12237), .B2(n14116), .ZN(
        n8606) );
  OAI22_X1 U1920 ( .A1(n10747), .A2(n12232), .B1(n12237), .B2(n14115), .ZN(
        n8605) );
  OAI22_X1 U1921 ( .A1(n10740), .A2(n12232), .B1(n12237), .B2(n14114), .ZN(
        n8604) );
  OAI22_X1 U1922 ( .A1(n10733), .A2(n12232), .B1(n12238), .B2(n14113), .ZN(
        n8603) );
  OAI22_X1 U1923 ( .A1(n10726), .A2(n12232), .B1(n12238), .B2(n14112), .ZN(
        n8602) );
  OAI22_X1 U1924 ( .A1(n10719), .A2(n12232), .B1(n12238), .B2(n14111), .ZN(
        n8601) );
  OAI22_X1 U1925 ( .A1(n10712), .A2(n12232), .B1(n12239), .B2(n14110), .ZN(
        n8600) );
  OAI22_X1 U1926 ( .A1(n10705), .A2(n12231), .B1(n12239), .B2(n14109), .ZN(
        n8599) );
  OAI22_X1 U1927 ( .A1(n10698), .A2(n12231), .B1(n12239), .B2(n14108), .ZN(
        n8598) );
  OAI22_X1 U1928 ( .A1(n10691), .A2(n12231), .B1(n12239), .B2(n14107), .ZN(
        n8597) );
  OAI22_X1 U1929 ( .A1(n10684), .A2(n12231), .B1(n12240), .B2(n14106), .ZN(
        n8596) );
  OAI22_X1 U1930 ( .A1(n10677), .A2(n12231), .B1(n12240), .B2(n14105), .ZN(
        n8595) );
  OAI22_X1 U1931 ( .A1(n10670), .A2(n12231), .B1(n12240), .B2(n14104), .ZN(
        n8594) );
  OAI22_X1 U1932 ( .A1(n10663), .A2(n12231), .B1(n12240), .B2(n14103), .ZN(
        n8593) );
  OAI22_X1 U1933 ( .A1(n10656), .A2(n12231), .B1(n12241), .B2(n14102), .ZN(
        n8592) );
  OAI22_X1 U1934 ( .A1(n10649), .A2(n12231), .B1(n12241), .B2(n14101), .ZN(
        n8591) );
  OAI22_X1 U1935 ( .A1(n10642), .A2(n12231), .B1(n12241), .B2(n14100), .ZN(
        n8590) );
  OAI22_X1 U1936 ( .A1(n10635), .A2(n12231), .B1(n12241), .B2(n14099), .ZN(
        n8589) );
  OAI22_X1 U1937 ( .A1(n10845), .A2(n12221), .B1(n12222), .B2(n14098), .ZN(
        n8587) );
  OAI22_X1 U1938 ( .A1(n10838), .A2(n12221), .B1(n12222), .B2(n14097), .ZN(
        n8586) );
  OAI22_X1 U1939 ( .A1(n10831), .A2(n12221), .B1(n12222), .B2(n14096), .ZN(
        n8585) );
  OAI22_X1 U1940 ( .A1(n10824), .A2(n12221), .B1(n12222), .B2(n14095), .ZN(
        n8584) );
  OAI22_X1 U1941 ( .A1(n10817), .A2(n12221), .B1(n12223), .B2(n14094), .ZN(
        n8583) );
  OAI22_X1 U1942 ( .A1(n10810), .A2(n12221), .B1(n12223), .B2(n14093), .ZN(
        n8582) );
  OAI22_X1 U1943 ( .A1(n10803), .A2(n12221), .B1(n12223), .B2(n14092), .ZN(
        n8581) );
  OAI22_X1 U1944 ( .A1(n10796), .A2(n12221), .B1(n12223), .B2(n14091), .ZN(
        n8580) );
  OAI22_X1 U1945 ( .A1(n10789), .A2(n12220), .B1(n12224), .B2(n14090), .ZN(
        n8579) );
  OAI22_X1 U1946 ( .A1(n10782), .A2(n12220), .B1(n12224), .B2(n14089), .ZN(
        n8578) );
  OAI22_X1 U1947 ( .A1(n10775), .A2(n12220), .B1(n12224), .B2(n14088), .ZN(
        n8577) );
  OAI22_X1 U1948 ( .A1(n10768), .A2(n12220), .B1(n12224), .B2(n14087), .ZN(
        n8576) );
  OAI22_X1 U1949 ( .A1(n10761), .A2(n12220), .B1(n12225), .B2(n14086), .ZN(
        n8575) );
  OAI22_X1 U1950 ( .A1(n10754), .A2(n12220), .B1(n12225), .B2(n14085), .ZN(
        n8574) );
  OAI22_X1 U1951 ( .A1(n10747), .A2(n12220), .B1(n12225), .B2(n14084), .ZN(
        n8573) );
  OAI22_X1 U1952 ( .A1(n10740), .A2(n12220), .B1(n12225), .B2(n14083), .ZN(
        n8572) );
  OAI22_X1 U1953 ( .A1(n10733), .A2(n12220), .B1(n12226), .B2(n14082), .ZN(
        n8571) );
  OAI22_X1 U1954 ( .A1(n10726), .A2(n12220), .B1(n12226), .B2(n14081), .ZN(
        n8570) );
  OAI22_X1 U1955 ( .A1(n10719), .A2(n12220), .B1(n12226), .B2(n14080), .ZN(
        n8569) );
  OAI22_X1 U1956 ( .A1(n10712), .A2(n12220), .B1(n12226), .B2(n14079), .ZN(
        n8568) );
  OAI22_X1 U1957 ( .A1(n10705), .A2(n12219), .B1(n12227), .B2(n14078), .ZN(
        n8567) );
  OAI22_X1 U1958 ( .A1(n10698), .A2(n12219), .B1(n12227), .B2(n14077), .ZN(
        n8566) );
  OAI22_X1 U1959 ( .A1(n10691), .A2(n12219), .B1(n12227), .B2(n14076), .ZN(
        n8565) );
  OAI22_X1 U1960 ( .A1(n10684), .A2(n12219), .B1(n12227), .B2(n14075), .ZN(
        n8564) );
  OAI22_X1 U1961 ( .A1(n10677), .A2(n12219), .B1(n12228), .B2(n14074), .ZN(
        n8563) );
  OAI22_X1 U1962 ( .A1(n10670), .A2(n12219), .B1(n12228), .B2(n14073), .ZN(
        n8562) );
  OAI22_X1 U1963 ( .A1(n10663), .A2(n12219), .B1(n12228), .B2(n14072), .ZN(
        n8561) );
  OAI22_X1 U1964 ( .A1(n10656), .A2(n12219), .B1(n12228), .B2(n14071), .ZN(
        n8560) );
  OAI22_X1 U1965 ( .A1(n10649), .A2(n12219), .B1(n12229), .B2(n14070), .ZN(
        n8559) );
  OAI22_X1 U1966 ( .A1(n10642), .A2(n12219), .B1(n12229), .B2(n14069), .ZN(
        n8558) );
  OAI22_X1 U1967 ( .A1(n10635), .A2(n12219), .B1(n12229), .B2(n14068), .ZN(
        n8557) );
  OAI22_X1 U1968 ( .A1(n10628), .A2(n12219), .B1(n12229), .B2(n14067), .ZN(
        n8556) );
  OAI22_X1 U1969 ( .A1(n10845), .A2(n12209), .B1(n12210), .B2(n14066), .ZN(
        n8555) );
  OAI22_X1 U1970 ( .A1(n10838), .A2(n12209), .B1(n12210), .B2(n14065), .ZN(
        n8554) );
  OAI22_X1 U1971 ( .A1(n10831), .A2(n12209), .B1(n12210), .B2(n14064), .ZN(
        n8553) );
  OAI22_X1 U1972 ( .A1(n10824), .A2(n12209), .B1(n12210), .B2(n14063), .ZN(
        n8552) );
  OAI22_X1 U1973 ( .A1(n10817), .A2(n12209), .B1(n12211), .B2(n14062), .ZN(
        n8551) );
  OAI22_X1 U1974 ( .A1(n10810), .A2(n12209), .B1(n12211), .B2(n14061), .ZN(
        n8550) );
  OAI22_X1 U1975 ( .A1(n10803), .A2(n12209), .B1(n12211), .B2(n14060), .ZN(
        n8549) );
  OAI22_X1 U1976 ( .A1(n10796), .A2(n12209), .B1(n12211), .B2(n14059), .ZN(
        n8548) );
  OAI22_X1 U1977 ( .A1(n10789), .A2(n12208), .B1(n12212), .B2(n14058), .ZN(
        n8547) );
  OAI22_X1 U1978 ( .A1(n10782), .A2(n12208), .B1(n12212), .B2(n14057), .ZN(
        n8546) );
  OAI22_X1 U1979 ( .A1(n10775), .A2(n12208), .B1(n12212), .B2(n14056), .ZN(
        n8545) );
  OAI22_X1 U1980 ( .A1(n10768), .A2(n12208), .B1(n12212), .B2(n14055), .ZN(
        n8544) );
  OAI22_X1 U1981 ( .A1(n10761), .A2(n12208), .B1(n12213), .B2(n14054), .ZN(
        n8543) );
  OAI22_X1 U1982 ( .A1(n10754), .A2(n12208), .B1(n12213), .B2(n14053), .ZN(
        n8542) );
  OAI22_X1 U1983 ( .A1(n10747), .A2(n12208), .B1(n12213), .B2(n14052), .ZN(
        n8541) );
  OAI22_X1 U1984 ( .A1(n10740), .A2(n12208), .B1(n12213), .B2(n14051), .ZN(
        n8540) );
  OAI22_X1 U1985 ( .A1(n10733), .A2(n12208), .B1(n12214), .B2(n14050), .ZN(
        n8539) );
  OAI22_X1 U1986 ( .A1(n10726), .A2(n12208), .B1(n12214), .B2(n14049), .ZN(
        n8538) );
  OAI22_X1 U1987 ( .A1(n10719), .A2(n12208), .B1(n12214), .B2(n14048), .ZN(
        n8537) );
  OAI22_X1 U1988 ( .A1(n10712), .A2(n12208), .B1(n12214), .B2(n14047), .ZN(
        n8536) );
  OAI22_X1 U1989 ( .A1(n10705), .A2(n12207), .B1(n12215), .B2(n14046), .ZN(
        n8535) );
  OAI22_X1 U1990 ( .A1(n10698), .A2(n12207), .B1(n12215), .B2(n14045), .ZN(
        n8534) );
  OAI22_X1 U1991 ( .A1(n10691), .A2(n12207), .B1(n12215), .B2(n14044), .ZN(
        n8533) );
  OAI22_X1 U1992 ( .A1(n10684), .A2(n12207), .B1(n12215), .B2(n14043), .ZN(
        n8532) );
  OAI22_X1 U1993 ( .A1(n10677), .A2(n12207), .B1(n12216), .B2(n14042), .ZN(
        n8531) );
  OAI22_X1 U1994 ( .A1(n10670), .A2(n12207), .B1(n12216), .B2(n14041), .ZN(
        n8530) );
  OAI22_X1 U1995 ( .A1(n10663), .A2(n12207), .B1(n12216), .B2(n14040), .ZN(
        n8529) );
  OAI22_X1 U1996 ( .A1(n10656), .A2(n12207), .B1(n12216), .B2(n14039), .ZN(
        n8528) );
  OAI22_X1 U1997 ( .A1(n10649), .A2(n12207), .B1(n12217), .B2(n14038), .ZN(
        n8527) );
  OAI22_X1 U1998 ( .A1(n10642), .A2(n12207), .B1(n12217), .B2(n14037), .ZN(
        n8526) );
  OAI22_X1 U1999 ( .A1(n10635), .A2(n12207), .B1(n12217), .B2(n14036), .ZN(
        n8525) );
  OAI22_X1 U2000 ( .A1(n10628), .A2(n12207), .B1(n12217), .B2(n14035), .ZN(
        n8524) );
  OAI22_X1 U2001 ( .A1(n10845), .A2(n12197), .B1(n12202), .B2(n14034), .ZN(
        n8523) );
  OAI22_X1 U2002 ( .A1(n10838), .A2(n12197), .B1(n12198), .B2(n14033), .ZN(
        n8522) );
  OAI22_X1 U2003 ( .A1(n10831), .A2(n12197), .B1(n12198), .B2(n14032), .ZN(
        n8521) );
  OAI22_X1 U2004 ( .A1(n10824), .A2(n12197), .B1(n12198), .B2(n14031), .ZN(
        n8520) );
  OAI22_X1 U2005 ( .A1(n10817), .A2(n12197), .B1(n12199), .B2(n14030), .ZN(
        n8519) );
  OAI22_X1 U2006 ( .A1(n10810), .A2(n12197), .B1(n12199), .B2(n14029), .ZN(
        n8518) );
  OAI22_X1 U2007 ( .A1(n10803), .A2(n12197), .B1(n12199), .B2(n14028), .ZN(
        n8517) );
  OAI22_X1 U2008 ( .A1(n10796), .A2(n12197), .B1(n12199), .B2(n14027), .ZN(
        n8516) );
  OAI22_X1 U2009 ( .A1(n10789), .A2(n12196), .B1(n12200), .B2(n14026), .ZN(
        n8515) );
  OAI22_X1 U2010 ( .A1(n10782), .A2(n12196), .B1(n12200), .B2(n14025), .ZN(
        n8514) );
  OAI22_X1 U2011 ( .A1(n10775), .A2(n12196), .B1(n12200), .B2(n14024), .ZN(
        n8513) );
  OAI22_X1 U2012 ( .A1(n10768), .A2(n12196), .B1(n12200), .B2(n14023), .ZN(
        n8512) );
  OAI22_X1 U2013 ( .A1(n10761), .A2(n12196), .B1(n12201), .B2(n14022), .ZN(
        n8511) );
  OAI22_X1 U2014 ( .A1(n10754), .A2(n12196), .B1(n12201), .B2(n14021), .ZN(
        n8510) );
  OAI22_X1 U2015 ( .A1(n10747), .A2(n12196), .B1(n12201), .B2(n14020), .ZN(
        n8509) );
  OAI22_X1 U2016 ( .A1(n10740), .A2(n12196), .B1(n12201), .B2(n14019), .ZN(
        n8508) );
  OAI22_X1 U2017 ( .A1(n10733), .A2(n12196), .B1(n12202), .B2(n14018), .ZN(
        n8507) );
  OAI22_X1 U2018 ( .A1(n10726), .A2(n12196), .B1(n12202), .B2(n14017), .ZN(
        n8506) );
  OAI22_X1 U2019 ( .A1(n10719), .A2(n12196), .B1(n12202), .B2(n14016), .ZN(
        n8505) );
  OAI22_X1 U2020 ( .A1(n10712), .A2(n12196), .B1(n12203), .B2(n14015), .ZN(
        n8504) );
  OAI22_X1 U2021 ( .A1(n10705), .A2(n12195), .B1(n12203), .B2(n14014), .ZN(
        n8503) );
  OAI22_X1 U2022 ( .A1(n10698), .A2(n12195), .B1(n12203), .B2(n14013), .ZN(
        n8502) );
  OAI22_X1 U2023 ( .A1(n10691), .A2(n12195), .B1(n12203), .B2(n14012), .ZN(
        n8501) );
  OAI22_X1 U2024 ( .A1(n10684), .A2(n12195), .B1(n12204), .B2(n14011), .ZN(
        n8500) );
  OAI22_X1 U2025 ( .A1(n10677), .A2(n12195), .B1(n12204), .B2(n14010), .ZN(
        n8499) );
  OAI22_X1 U2026 ( .A1(n10670), .A2(n12195), .B1(n12204), .B2(n14009), .ZN(
        n8498) );
  OAI22_X1 U2027 ( .A1(n10663), .A2(n12195), .B1(n12204), .B2(n14008), .ZN(
        n8497) );
  OAI22_X1 U2028 ( .A1(n10656), .A2(n12195), .B1(n12205), .B2(n14007), .ZN(
        n8496) );
  OAI22_X1 U2029 ( .A1(n10649), .A2(n12195), .B1(n12205), .B2(n14006), .ZN(
        n8495) );
  OAI22_X1 U2030 ( .A1(n10642), .A2(n12195), .B1(n12205), .B2(n14005), .ZN(
        n8494) );
  OAI22_X1 U2031 ( .A1(n10635), .A2(n12195), .B1(n12205), .B2(n14004), .ZN(
        n8493) );
  OAI22_X1 U2032 ( .A1(n10845), .A2(n12185), .B1(n12186), .B2(n14003), .ZN(
        n8491) );
  OAI22_X1 U2033 ( .A1(n10838), .A2(n12185), .B1(n12186), .B2(n14002), .ZN(
        n8490) );
  OAI22_X1 U2034 ( .A1(n10831), .A2(n12185), .B1(n12186), .B2(n14001), .ZN(
        n8489) );
  OAI22_X1 U2035 ( .A1(n10824), .A2(n12185), .B1(n12186), .B2(n14000), .ZN(
        n8488) );
  OAI22_X1 U2036 ( .A1(n10817), .A2(n12185), .B1(n12187), .B2(n13999), .ZN(
        n8487) );
  OAI22_X1 U2037 ( .A1(n10810), .A2(n12185), .B1(n12187), .B2(n13998), .ZN(
        n8486) );
  OAI22_X1 U2038 ( .A1(n10803), .A2(n12185), .B1(n12187), .B2(n13997), .ZN(
        n8485) );
  OAI22_X1 U2039 ( .A1(n10796), .A2(n12185), .B1(n12187), .B2(n13996), .ZN(
        n8484) );
  OAI22_X1 U2040 ( .A1(n10789), .A2(n12184), .B1(n12188), .B2(n13995), .ZN(
        n8483) );
  OAI22_X1 U2041 ( .A1(n10782), .A2(n12184), .B1(n12188), .B2(n13994), .ZN(
        n8482) );
  OAI22_X1 U2042 ( .A1(n10775), .A2(n12184), .B1(n12188), .B2(n13993), .ZN(
        n8481) );
  OAI22_X1 U2043 ( .A1(n10768), .A2(n12184), .B1(n12188), .B2(n13992), .ZN(
        n8480) );
  OAI22_X1 U2044 ( .A1(n10761), .A2(n12184), .B1(n12189), .B2(n13991), .ZN(
        n8479) );
  OAI22_X1 U2045 ( .A1(n10754), .A2(n12184), .B1(n12189), .B2(n13990), .ZN(
        n8478) );
  OAI22_X1 U2046 ( .A1(n10747), .A2(n12184), .B1(n12189), .B2(n13989), .ZN(
        n8477) );
  OAI22_X1 U2047 ( .A1(n10740), .A2(n12184), .B1(n12189), .B2(n13988), .ZN(
        n8476) );
  OAI22_X1 U2048 ( .A1(n10733), .A2(n12184), .B1(n12190), .B2(n13987), .ZN(
        n8475) );
  OAI22_X1 U2049 ( .A1(n10726), .A2(n12184), .B1(n12190), .B2(n13986), .ZN(
        n8474) );
  OAI22_X1 U2050 ( .A1(n10719), .A2(n12184), .B1(n12190), .B2(n13985), .ZN(
        n8473) );
  OAI22_X1 U2051 ( .A1(n10712), .A2(n12184), .B1(n12190), .B2(n13984), .ZN(
        n8472) );
  OAI22_X1 U2052 ( .A1(n10705), .A2(n12183), .B1(n12191), .B2(n13983), .ZN(
        n8471) );
  OAI22_X1 U2053 ( .A1(n10698), .A2(n12183), .B1(n12191), .B2(n13982), .ZN(
        n8470) );
  OAI22_X1 U2054 ( .A1(n10691), .A2(n12183), .B1(n12191), .B2(n13981), .ZN(
        n8469) );
  OAI22_X1 U2055 ( .A1(n10684), .A2(n12183), .B1(n12191), .B2(n13980), .ZN(
        n8468) );
  OAI22_X1 U2056 ( .A1(n10677), .A2(n12183), .B1(n12192), .B2(n13979), .ZN(
        n8467) );
  OAI22_X1 U2057 ( .A1(n10670), .A2(n12183), .B1(n12192), .B2(n13978), .ZN(
        n8466) );
  OAI22_X1 U2058 ( .A1(n10663), .A2(n12183), .B1(n12192), .B2(n13977), .ZN(
        n8465) );
  OAI22_X1 U2059 ( .A1(n10656), .A2(n12183), .B1(n12192), .B2(n13976), .ZN(
        n8464) );
  OAI22_X1 U2060 ( .A1(n10649), .A2(n12183), .B1(n12193), .B2(n13975), .ZN(
        n8463) );
  OAI22_X1 U2061 ( .A1(n10642), .A2(n12183), .B1(n12193), .B2(n13974), .ZN(
        n8462) );
  OAI22_X1 U2062 ( .A1(n10635), .A2(n12183), .B1(n12193), .B2(n13973), .ZN(
        n8461) );
  OAI22_X1 U2063 ( .A1(n10628), .A2(n12183), .B1(n12193), .B2(n13972), .ZN(
        n8460) );
  OAI22_X1 U2064 ( .A1(n10845), .A2(n12173), .B1(n12174), .B2(n13971), .ZN(
        n8459) );
  OAI22_X1 U2065 ( .A1(n10838), .A2(n12173), .B1(n12174), .B2(n13970), .ZN(
        n8458) );
  OAI22_X1 U2066 ( .A1(n10831), .A2(n12173), .B1(n12174), .B2(n13969), .ZN(
        n8457) );
  OAI22_X1 U2067 ( .A1(n10824), .A2(n12173), .B1(n12174), .B2(n13968), .ZN(
        n8456) );
  OAI22_X1 U2068 ( .A1(n10817), .A2(n12173), .B1(n12175), .B2(n13967), .ZN(
        n8455) );
  OAI22_X1 U2069 ( .A1(n10810), .A2(n12173), .B1(n12175), .B2(n13966), .ZN(
        n8454) );
  OAI22_X1 U2070 ( .A1(n10803), .A2(n12173), .B1(n12175), .B2(n13965), .ZN(
        n8453) );
  OAI22_X1 U2071 ( .A1(n10796), .A2(n12173), .B1(n12175), .B2(n13964), .ZN(
        n8452) );
  OAI22_X1 U2072 ( .A1(n10789), .A2(n12172), .B1(n12176), .B2(n13963), .ZN(
        n8451) );
  OAI22_X1 U2073 ( .A1(n10782), .A2(n12172), .B1(n12176), .B2(n13962), .ZN(
        n8450) );
  OAI22_X1 U2074 ( .A1(n10775), .A2(n12172), .B1(n12176), .B2(n13961), .ZN(
        n8449) );
  OAI22_X1 U2075 ( .A1(n10768), .A2(n12172), .B1(n12176), .B2(n13960), .ZN(
        n8448) );
  OAI22_X1 U2076 ( .A1(n10761), .A2(n12172), .B1(n12177), .B2(n13959), .ZN(
        n8447) );
  OAI22_X1 U2077 ( .A1(n10754), .A2(n12172), .B1(n12177), .B2(n13958), .ZN(
        n8446) );
  OAI22_X1 U2078 ( .A1(n10747), .A2(n12172), .B1(n12177), .B2(n13957), .ZN(
        n8445) );
  OAI22_X1 U2079 ( .A1(n10740), .A2(n12172), .B1(n12177), .B2(n13956), .ZN(
        n8444) );
  OAI22_X1 U2080 ( .A1(n10733), .A2(n12172), .B1(n12178), .B2(n13955), .ZN(
        n8443) );
  OAI22_X1 U2081 ( .A1(n10726), .A2(n12172), .B1(n12178), .B2(n13954), .ZN(
        n8442) );
  OAI22_X1 U2082 ( .A1(n10719), .A2(n12172), .B1(n12178), .B2(n13953), .ZN(
        n8441) );
  OAI22_X1 U2083 ( .A1(n10712), .A2(n12172), .B1(n12178), .B2(n13952), .ZN(
        n8440) );
  OAI22_X1 U2084 ( .A1(n10705), .A2(n12171), .B1(n12179), .B2(n13951), .ZN(
        n8439) );
  OAI22_X1 U2085 ( .A1(n10698), .A2(n12171), .B1(n12179), .B2(n13950), .ZN(
        n8438) );
  OAI22_X1 U2086 ( .A1(n10691), .A2(n12171), .B1(n12179), .B2(n13949), .ZN(
        n8437) );
  OAI22_X1 U2087 ( .A1(n10684), .A2(n12171), .B1(n12179), .B2(n13948), .ZN(
        n8436) );
  OAI22_X1 U2088 ( .A1(n10677), .A2(n12171), .B1(n12180), .B2(n13947), .ZN(
        n8435) );
  OAI22_X1 U2089 ( .A1(n10670), .A2(n12171), .B1(n12180), .B2(n13946), .ZN(
        n8434) );
  OAI22_X1 U2090 ( .A1(n10663), .A2(n12171), .B1(n12180), .B2(n13945), .ZN(
        n8433) );
  OAI22_X1 U2091 ( .A1(n10656), .A2(n12171), .B1(n12180), .B2(n13944), .ZN(
        n8432) );
  OAI22_X1 U2092 ( .A1(n10649), .A2(n12171), .B1(n12181), .B2(n13943), .ZN(
        n8431) );
  OAI22_X1 U2093 ( .A1(n10642), .A2(n12171), .B1(n12181), .B2(n13942), .ZN(
        n8430) );
  OAI22_X1 U2094 ( .A1(n10635), .A2(n12171), .B1(n12181), .B2(n13941), .ZN(
        n8429) );
  OAI22_X1 U2095 ( .A1(n10628), .A2(n12171), .B1(n12181), .B2(n13940), .ZN(
        n8428) );
  OAI22_X1 U2096 ( .A1(n10845), .A2(n12161), .B1(n12162), .B2(n13939), .ZN(
        n8427) );
  OAI22_X1 U2097 ( .A1(n10838), .A2(n12161), .B1(n12162), .B2(n13938), .ZN(
        n8426) );
  OAI22_X1 U2098 ( .A1(n10831), .A2(n12161), .B1(n12162), .B2(n13937), .ZN(
        n8425) );
  OAI22_X1 U2099 ( .A1(n10824), .A2(n12161), .B1(n12162), .B2(n13936), .ZN(
        n8424) );
  OAI22_X1 U2100 ( .A1(n10817), .A2(n12161), .B1(n12163), .B2(n13935), .ZN(
        n8423) );
  OAI22_X1 U2101 ( .A1(n10810), .A2(n12161), .B1(n12163), .B2(n13934), .ZN(
        n8422) );
  OAI22_X1 U2102 ( .A1(n10803), .A2(n12161), .B1(n12163), .B2(n13933), .ZN(
        n8421) );
  OAI22_X1 U2103 ( .A1(n10796), .A2(n12161), .B1(n12163), .B2(n13932), .ZN(
        n8420) );
  OAI22_X1 U2104 ( .A1(n10789), .A2(n12160), .B1(n12164), .B2(n13931), .ZN(
        n8419) );
  OAI22_X1 U2105 ( .A1(n10782), .A2(n12160), .B1(n12164), .B2(n13930), .ZN(
        n8418) );
  OAI22_X1 U2106 ( .A1(n10775), .A2(n12160), .B1(n12164), .B2(n13929), .ZN(
        n8417) );
  OAI22_X1 U2107 ( .A1(n10768), .A2(n12160), .B1(n12164), .B2(n13928), .ZN(
        n8416) );
  OAI22_X1 U2108 ( .A1(n10761), .A2(n12160), .B1(n12165), .B2(n13927), .ZN(
        n8415) );
  OAI22_X1 U2109 ( .A1(n10754), .A2(n12160), .B1(n12165), .B2(n13926), .ZN(
        n8414) );
  OAI22_X1 U2110 ( .A1(n10747), .A2(n12160), .B1(n12165), .B2(n13925), .ZN(
        n8413) );
  OAI22_X1 U2111 ( .A1(n10740), .A2(n12160), .B1(n12165), .B2(n13924), .ZN(
        n8412) );
  OAI22_X1 U2112 ( .A1(n10733), .A2(n12160), .B1(n12166), .B2(n13923), .ZN(
        n8411) );
  OAI22_X1 U2113 ( .A1(n10726), .A2(n12160), .B1(n12166), .B2(n13922), .ZN(
        n8410) );
  OAI22_X1 U2114 ( .A1(n10719), .A2(n12160), .B1(n12166), .B2(n13921), .ZN(
        n8409) );
  OAI22_X1 U2115 ( .A1(n10712), .A2(n12160), .B1(n12166), .B2(n13920), .ZN(
        n8408) );
  OAI22_X1 U2116 ( .A1(n10705), .A2(n12159), .B1(n12167), .B2(n13919), .ZN(
        n8407) );
  OAI22_X1 U2117 ( .A1(n10698), .A2(n12159), .B1(n12167), .B2(n13918), .ZN(
        n8406) );
  OAI22_X1 U2118 ( .A1(n10691), .A2(n12159), .B1(n12167), .B2(n13917), .ZN(
        n8405) );
  OAI22_X1 U2119 ( .A1(n10684), .A2(n12159), .B1(n12167), .B2(n13916), .ZN(
        n8404) );
  OAI22_X1 U2120 ( .A1(n10677), .A2(n12159), .B1(n12168), .B2(n13915), .ZN(
        n8403) );
  OAI22_X1 U2121 ( .A1(n10670), .A2(n12159), .B1(n12168), .B2(n13914), .ZN(
        n8402) );
  OAI22_X1 U2122 ( .A1(n10663), .A2(n12159), .B1(n12168), .B2(n13913), .ZN(
        n8401) );
  OAI22_X1 U2123 ( .A1(n10656), .A2(n12159), .B1(n12168), .B2(n13912), .ZN(
        n8400) );
  OAI22_X1 U2124 ( .A1(n10649), .A2(n12159), .B1(n12169), .B2(n13911), .ZN(
        n8399) );
  OAI22_X1 U2125 ( .A1(n10642), .A2(n12159), .B1(n12169), .B2(n13910), .ZN(
        n8398) );
  OAI22_X1 U2126 ( .A1(n10635), .A2(n12159), .B1(n12169), .B2(n13909), .ZN(
        n8397) );
  OAI22_X1 U2127 ( .A1(n10628), .A2(n12159), .B1(n12169), .B2(n13908), .ZN(
        n8396) );
  OAI22_X1 U2128 ( .A1(n10845), .A2(n12137), .B1(n12138), .B2(n13907), .ZN(
        n8363) );
  OAI22_X1 U2129 ( .A1(n10838), .A2(n12137), .B1(n12138), .B2(n13906), .ZN(
        n8362) );
  OAI22_X1 U2130 ( .A1(n10831), .A2(n12137), .B1(n12138), .B2(n13905), .ZN(
        n8361) );
  OAI22_X1 U2131 ( .A1(n10824), .A2(n12137), .B1(n12138), .B2(n13904), .ZN(
        n8360) );
  OAI22_X1 U2132 ( .A1(n10817), .A2(n12137), .B1(n12139), .B2(n13903), .ZN(
        n8359) );
  OAI22_X1 U2133 ( .A1(n10810), .A2(n12137), .B1(n12139), .B2(n13902), .ZN(
        n8358) );
  OAI22_X1 U2134 ( .A1(n10803), .A2(n12137), .B1(n12139), .B2(n13901), .ZN(
        n8357) );
  OAI22_X1 U2135 ( .A1(n10796), .A2(n12137), .B1(n12139), .B2(n13900), .ZN(
        n8356) );
  OAI22_X1 U2136 ( .A1(n10789), .A2(n12136), .B1(n12140), .B2(n13899), .ZN(
        n8355) );
  OAI22_X1 U2137 ( .A1(n10782), .A2(n12136), .B1(n12140), .B2(n13898), .ZN(
        n8354) );
  OAI22_X1 U2138 ( .A1(n10775), .A2(n12136), .B1(n12140), .B2(n13897), .ZN(
        n8353) );
  OAI22_X1 U2139 ( .A1(n10768), .A2(n12136), .B1(n12140), .B2(n13896), .ZN(
        n8352) );
  OAI22_X1 U2140 ( .A1(n10761), .A2(n12136), .B1(n12141), .B2(n13895), .ZN(
        n8351) );
  OAI22_X1 U2141 ( .A1(n10754), .A2(n12136), .B1(n12141), .B2(n13894), .ZN(
        n8350) );
  OAI22_X1 U2142 ( .A1(n10747), .A2(n12136), .B1(n12141), .B2(n13893), .ZN(
        n8349) );
  OAI22_X1 U2143 ( .A1(n10740), .A2(n12136), .B1(n12141), .B2(n13892), .ZN(
        n8348) );
  OAI22_X1 U2144 ( .A1(n10733), .A2(n12136), .B1(n12142), .B2(n13891), .ZN(
        n8347) );
  OAI22_X1 U2145 ( .A1(n10726), .A2(n12136), .B1(n12142), .B2(n13890), .ZN(
        n8346) );
  OAI22_X1 U2146 ( .A1(n10719), .A2(n12136), .B1(n12142), .B2(n13889), .ZN(
        n8345) );
  OAI22_X1 U2147 ( .A1(n10712), .A2(n12136), .B1(n12142), .B2(n13888), .ZN(
        n8344) );
  OAI22_X1 U2148 ( .A1(n10705), .A2(n12135), .B1(n12143), .B2(n13887), .ZN(
        n8343) );
  OAI22_X1 U2149 ( .A1(n10698), .A2(n12135), .B1(n12143), .B2(n13886), .ZN(
        n8342) );
  OAI22_X1 U2150 ( .A1(n10691), .A2(n12135), .B1(n12143), .B2(n13885), .ZN(
        n8341) );
  OAI22_X1 U2151 ( .A1(n10684), .A2(n12135), .B1(n12143), .B2(n13884), .ZN(
        n8340) );
  OAI22_X1 U2152 ( .A1(n10677), .A2(n12135), .B1(n12144), .B2(n13883), .ZN(
        n8339) );
  OAI22_X1 U2153 ( .A1(n10670), .A2(n12135), .B1(n12144), .B2(n13882), .ZN(
        n8338) );
  OAI22_X1 U2154 ( .A1(n10663), .A2(n12135), .B1(n12144), .B2(n13881), .ZN(
        n8337) );
  OAI22_X1 U2155 ( .A1(n10656), .A2(n12135), .B1(n12144), .B2(n13880), .ZN(
        n8336) );
  OAI22_X1 U2156 ( .A1(n10649), .A2(n12135), .B1(n12145), .B2(n13879), .ZN(
        n8335) );
  OAI22_X1 U2157 ( .A1(n10642), .A2(n12135), .B1(n12145), .B2(n13878), .ZN(
        n8334) );
  OAI22_X1 U2158 ( .A1(n10635), .A2(n12135), .B1(n12145), .B2(n13877), .ZN(
        n8333) );
  OAI22_X1 U2159 ( .A1(n10628), .A2(n12135), .B1(n12145), .B2(n13876), .ZN(
        n8332) );
  OAI22_X1 U2160 ( .A1(n10846), .A2(n12113), .B1(n12114), .B2(n13875), .ZN(
        n8299) );
  OAI22_X1 U2161 ( .A1(n10839), .A2(n12113), .B1(n12114), .B2(n13874), .ZN(
        n8298) );
  OAI22_X1 U2162 ( .A1(n10832), .A2(n12113), .B1(n12114), .B2(n13873), .ZN(
        n8297) );
  OAI22_X1 U2163 ( .A1(n10825), .A2(n12113), .B1(n12114), .B2(n13872), .ZN(
        n8296) );
  OAI22_X1 U2164 ( .A1(n10818), .A2(n12113), .B1(n12115), .B2(n13871), .ZN(
        n8295) );
  OAI22_X1 U2165 ( .A1(n10811), .A2(n12113), .B1(n12115), .B2(n13870), .ZN(
        n8294) );
  OAI22_X1 U2166 ( .A1(n10804), .A2(n12113), .B1(n12115), .B2(n13869), .ZN(
        n8293) );
  OAI22_X1 U2167 ( .A1(n10797), .A2(n12113), .B1(n12115), .B2(n13868), .ZN(
        n8292) );
  OAI22_X1 U2168 ( .A1(n10790), .A2(n12112), .B1(n12116), .B2(n13867), .ZN(
        n8291) );
  OAI22_X1 U2169 ( .A1(n10783), .A2(n12112), .B1(n12116), .B2(n13866), .ZN(
        n8290) );
  OAI22_X1 U2170 ( .A1(n10776), .A2(n12112), .B1(n12116), .B2(n13865), .ZN(
        n8289) );
  OAI22_X1 U2171 ( .A1(n10769), .A2(n12112), .B1(n12116), .B2(n13864), .ZN(
        n8288) );
  OAI22_X1 U2172 ( .A1(n10762), .A2(n12112), .B1(n12117), .B2(n13863), .ZN(
        n8287) );
  OAI22_X1 U2173 ( .A1(n10755), .A2(n12112), .B1(n12117), .B2(n13862), .ZN(
        n8286) );
  OAI22_X1 U2174 ( .A1(n10748), .A2(n12112), .B1(n12117), .B2(n13861), .ZN(
        n8285) );
  OAI22_X1 U2175 ( .A1(n10741), .A2(n12112), .B1(n12117), .B2(n13860), .ZN(
        n8284) );
  OAI22_X1 U2176 ( .A1(n10734), .A2(n12112), .B1(n12118), .B2(n13859), .ZN(
        n8283) );
  OAI22_X1 U2177 ( .A1(n10727), .A2(n12112), .B1(n12118), .B2(n13858), .ZN(
        n8282) );
  OAI22_X1 U2178 ( .A1(n10720), .A2(n12112), .B1(n12118), .B2(n13857), .ZN(
        n8281) );
  OAI22_X1 U2179 ( .A1(n10713), .A2(n12112), .B1(n12118), .B2(n13856), .ZN(
        n8280) );
  OAI22_X1 U2180 ( .A1(n10706), .A2(n12111), .B1(n12119), .B2(n13855), .ZN(
        n8279) );
  OAI22_X1 U2181 ( .A1(n10699), .A2(n12111), .B1(n12119), .B2(n13854), .ZN(
        n8278) );
  OAI22_X1 U2182 ( .A1(n10692), .A2(n12111), .B1(n12119), .B2(n13853), .ZN(
        n8277) );
  OAI22_X1 U2183 ( .A1(n10685), .A2(n12111), .B1(n12119), .B2(n13852), .ZN(
        n8276) );
  OAI22_X1 U2184 ( .A1(n10678), .A2(n12111), .B1(n12120), .B2(n13851), .ZN(
        n8275) );
  OAI22_X1 U2185 ( .A1(n10671), .A2(n12111), .B1(n12120), .B2(n13850), .ZN(
        n8274) );
  OAI22_X1 U2186 ( .A1(n10664), .A2(n12111), .B1(n12120), .B2(n13849), .ZN(
        n8273) );
  OAI22_X1 U2187 ( .A1(n10657), .A2(n12111), .B1(n12120), .B2(n13848), .ZN(
        n8272) );
  OAI22_X1 U2188 ( .A1(n10650), .A2(n12111), .B1(n12121), .B2(n13847), .ZN(
        n8271) );
  OAI22_X1 U2189 ( .A1(n10643), .A2(n12111), .B1(n12121), .B2(n13846), .ZN(
        n8270) );
  OAI22_X1 U2190 ( .A1(n10636), .A2(n12111), .B1(n12121), .B2(n13845), .ZN(
        n8269) );
  OAI22_X1 U2191 ( .A1(n10629), .A2(n12111), .B1(n12121), .B2(n13844), .ZN(
        n8268) );
  OAI22_X1 U2192 ( .A1(n10847), .A2(n11957), .B1(n11958), .B2(n13651), .ZN(
        n7883) );
  OAI22_X1 U2193 ( .A1(n10840), .A2(n11957), .B1(n11958), .B2(n13650), .ZN(
        n7882) );
  OAI22_X1 U2194 ( .A1(n10833), .A2(n11957), .B1(n11958), .B2(n13649), .ZN(
        n7881) );
  OAI22_X1 U2195 ( .A1(n10826), .A2(n11957), .B1(n11958), .B2(n13648), .ZN(
        n7880) );
  OAI22_X1 U2196 ( .A1(n10819), .A2(n11957), .B1(n11959), .B2(n13647), .ZN(
        n7879) );
  OAI22_X1 U2197 ( .A1(n10812), .A2(n11957), .B1(n11959), .B2(n13646), .ZN(
        n7878) );
  OAI22_X1 U2198 ( .A1(n10805), .A2(n11957), .B1(n11959), .B2(n13645), .ZN(
        n7877) );
  OAI22_X1 U2199 ( .A1(n10798), .A2(n11957), .B1(n11959), .B2(n13644), .ZN(
        n7876) );
  OAI22_X1 U2200 ( .A1(n10791), .A2(n11956), .B1(n11960), .B2(n13643), .ZN(
        n7875) );
  OAI22_X1 U2201 ( .A1(n10784), .A2(n11956), .B1(n11960), .B2(n13642), .ZN(
        n7874) );
  OAI22_X1 U2202 ( .A1(n10777), .A2(n11956), .B1(n11960), .B2(n13641), .ZN(
        n7873) );
  OAI22_X1 U2203 ( .A1(n10770), .A2(n11956), .B1(n11960), .B2(n13640), .ZN(
        n7872) );
  OAI22_X1 U2204 ( .A1(n10763), .A2(n11956), .B1(n11961), .B2(n13639), .ZN(
        n7871) );
  OAI22_X1 U2205 ( .A1(n10756), .A2(n11956), .B1(n11961), .B2(n13638), .ZN(
        n7870) );
  OAI22_X1 U2206 ( .A1(n10749), .A2(n11956), .B1(n11961), .B2(n13637), .ZN(
        n7869) );
  OAI22_X1 U2207 ( .A1(n10742), .A2(n11956), .B1(n11961), .B2(n13636), .ZN(
        n7868) );
  OAI22_X1 U2208 ( .A1(n10735), .A2(n11956), .B1(n11962), .B2(n13635), .ZN(
        n7867) );
  OAI22_X1 U2209 ( .A1(n10728), .A2(n11956), .B1(n11962), .B2(n13634), .ZN(
        n7866) );
  OAI22_X1 U2210 ( .A1(n10721), .A2(n11956), .B1(n11962), .B2(n13633), .ZN(
        n7865) );
  OAI22_X1 U2211 ( .A1(n10714), .A2(n11956), .B1(n11962), .B2(n13632), .ZN(
        n7864) );
  OAI22_X1 U2212 ( .A1(n10707), .A2(n11955), .B1(n11963), .B2(n13631), .ZN(
        n7863) );
  OAI22_X1 U2213 ( .A1(n10700), .A2(n11955), .B1(n11963), .B2(n13630), .ZN(
        n7862) );
  OAI22_X1 U2214 ( .A1(n10693), .A2(n11955), .B1(n11963), .B2(n13629), .ZN(
        n7861) );
  OAI22_X1 U2215 ( .A1(n10686), .A2(n11955), .B1(n11963), .B2(n13628), .ZN(
        n7860) );
  OAI22_X1 U2216 ( .A1(n10679), .A2(n11955), .B1(n11964), .B2(n13627), .ZN(
        n7859) );
  OAI22_X1 U2217 ( .A1(n10672), .A2(n11955), .B1(n11964), .B2(n13626), .ZN(
        n7858) );
  OAI22_X1 U2218 ( .A1(n10665), .A2(n11955), .B1(n11964), .B2(n13625), .ZN(
        n7857) );
  OAI22_X1 U2219 ( .A1(n10658), .A2(n11955), .B1(n11964), .B2(n13624), .ZN(
        n7856) );
  OAI22_X1 U2220 ( .A1(n10651), .A2(n11955), .B1(n11965), .B2(n13623), .ZN(
        n7855) );
  OAI22_X1 U2221 ( .A1(n10644), .A2(n11955), .B1(n11965), .B2(n13622), .ZN(
        n7854) );
  OAI22_X1 U2222 ( .A1(n10637), .A2(n11955), .B1(n11965), .B2(n13621), .ZN(
        n7853) );
  OAI22_X1 U2223 ( .A1(n10630), .A2(n11955), .B1(n11965), .B2(n13620), .ZN(
        n7852) );
  OAI22_X1 U2224 ( .A1(n10847), .A2(n11945), .B1(n11946), .B2(n13619), .ZN(
        n7851) );
  OAI22_X1 U2225 ( .A1(n10840), .A2(n11945), .B1(n11946), .B2(n13618), .ZN(
        n7850) );
  OAI22_X1 U2226 ( .A1(n10833), .A2(n11945), .B1(n11946), .B2(n13617), .ZN(
        n7849) );
  OAI22_X1 U2227 ( .A1(n10826), .A2(n11945), .B1(n11946), .B2(n13616), .ZN(
        n7848) );
  OAI22_X1 U2228 ( .A1(n10819), .A2(n11945), .B1(n11947), .B2(n13615), .ZN(
        n7847) );
  OAI22_X1 U2229 ( .A1(n10812), .A2(n11945), .B1(n11947), .B2(n13614), .ZN(
        n7846) );
  OAI22_X1 U2230 ( .A1(n10805), .A2(n11945), .B1(n11947), .B2(n13613), .ZN(
        n7845) );
  OAI22_X1 U2231 ( .A1(n10798), .A2(n11945), .B1(n11947), .B2(n13612), .ZN(
        n7844) );
  OAI22_X1 U2232 ( .A1(n10791), .A2(n11944), .B1(n11948), .B2(n13611), .ZN(
        n7843) );
  OAI22_X1 U2233 ( .A1(n10784), .A2(n11944), .B1(n11948), .B2(n13610), .ZN(
        n7842) );
  OAI22_X1 U2234 ( .A1(n10777), .A2(n11944), .B1(n11948), .B2(n13609), .ZN(
        n7841) );
  OAI22_X1 U2235 ( .A1(n10770), .A2(n11944), .B1(n11948), .B2(n13608), .ZN(
        n7840) );
  OAI22_X1 U2236 ( .A1(n10763), .A2(n11944), .B1(n11949), .B2(n13607), .ZN(
        n7839) );
  OAI22_X1 U2237 ( .A1(n10756), .A2(n11944), .B1(n11949), .B2(n13606), .ZN(
        n7838) );
  OAI22_X1 U2238 ( .A1(n10749), .A2(n11944), .B1(n11949), .B2(n13605), .ZN(
        n7837) );
  OAI22_X1 U2239 ( .A1(n10742), .A2(n11944), .B1(n11949), .B2(n13604), .ZN(
        n7836) );
  OAI22_X1 U2240 ( .A1(n10735), .A2(n11944), .B1(n11950), .B2(n13603), .ZN(
        n7835) );
  OAI22_X1 U2241 ( .A1(n10728), .A2(n11944), .B1(n11950), .B2(n13602), .ZN(
        n7834) );
  OAI22_X1 U2242 ( .A1(n10721), .A2(n11944), .B1(n11950), .B2(n13601), .ZN(
        n7833) );
  OAI22_X1 U2243 ( .A1(n10714), .A2(n11944), .B1(n11950), .B2(n13600), .ZN(
        n7832) );
  OAI22_X1 U2244 ( .A1(n10707), .A2(n11943), .B1(n11951), .B2(n13599), .ZN(
        n7831) );
  OAI22_X1 U2245 ( .A1(n10700), .A2(n11943), .B1(n11951), .B2(n13598), .ZN(
        n7830) );
  OAI22_X1 U2246 ( .A1(n10693), .A2(n11943), .B1(n11951), .B2(n13597), .ZN(
        n7829) );
  OAI22_X1 U2247 ( .A1(n10686), .A2(n11943), .B1(n11951), .B2(n13596), .ZN(
        n7828) );
  OAI22_X1 U2248 ( .A1(n10679), .A2(n11943), .B1(n11952), .B2(n13595), .ZN(
        n7827) );
  OAI22_X1 U2249 ( .A1(n10672), .A2(n11943), .B1(n11952), .B2(n13594), .ZN(
        n7826) );
  OAI22_X1 U2250 ( .A1(n10665), .A2(n11943), .B1(n11952), .B2(n13593), .ZN(
        n7825) );
  OAI22_X1 U2251 ( .A1(n10658), .A2(n11943), .B1(n11952), .B2(n13592), .ZN(
        n7824) );
  OAI22_X1 U2252 ( .A1(n10651), .A2(n11943), .B1(n11953), .B2(n13591), .ZN(
        n7823) );
  OAI22_X1 U2253 ( .A1(n10644), .A2(n11943), .B1(n11953), .B2(n13590), .ZN(
        n7822) );
  OAI22_X1 U2254 ( .A1(n10637), .A2(n11943), .B1(n11953), .B2(n13589), .ZN(
        n7821) );
  OAI22_X1 U2255 ( .A1(n10630), .A2(n11943), .B1(n11953), .B2(n13588), .ZN(
        n7820) );
  OAI22_X1 U2256 ( .A1(n10847), .A2(n11933), .B1(n11934), .B2(n13587), .ZN(
        n7819) );
  OAI22_X1 U2257 ( .A1(n10840), .A2(n11933), .B1(n11934), .B2(n13586), .ZN(
        n7818) );
  OAI22_X1 U2258 ( .A1(n10833), .A2(n11933), .B1(n11934), .B2(n13585), .ZN(
        n7817) );
  OAI22_X1 U2259 ( .A1(n10826), .A2(n11933), .B1(n11934), .B2(n13584), .ZN(
        n7816) );
  OAI22_X1 U2260 ( .A1(n10819), .A2(n11933), .B1(n11935), .B2(n13583), .ZN(
        n7815) );
  OAI22_X1 U2261 ( .A1(n10812), .A2(n11933), .B1(n11935), .B2(n13582), .ZN(
        n7814) );
  OAI22_X1 U2262 ( .A1(n10805), .A2(n11933), .B1(n11935), .B2(n13581), .ZN(
        n7813) );
  OAI22_X1 U2263 ( .A1(n10798), .A2(n11933), .B1(n11935), .B2(n13580), .ZN(
        n7812) );
  OAI22_X1 U2264 ( .A1(n10791), .A2(n11932), .B1(n11936), .B2(n13579), .ZN(
        n7811) );
  OAI22_X1 U2265 ( .A1(n10784), .A2(n11932), .B1(n11936), .B2(n13578), .ZN(
        n7810) );
  OAI22_X1 U2266 ( .A1(n10777), .A2(n11932), .B1(n11936), .B2(n13577), .ZN(
        n7809) );
  OAI22_X1 U2267 ( .A1(n10770), .A2(n11932), .B1(n11936), .B2(n13576), .ZN(
        n7808) );
  OAI22_X1 U2268 ( .A1(n10763), .A2(n11932), .B1(n11937), .B2(n13575), .ZN(
        n7807) );
  OAI22_X1 U2269 ( .A1(n10756), .A2(n11932), .B1(n11937), .B2(n13574), .ZN(
        n7806) );
  OAI22_X1 U2270 ( .A1(n10749), .A2(n11932), .B1(n11937), .B2(n13573), .ZN(
        n7805) );
  OAI22_X1 U2271 ( .A1(n10742), .A2(n11932), .B1(n11937), .B2(n13572), .ZN(
        n7804) );
  OAI22_X1 U2272 ( .A1(n10735), .A2(n11932), .B1(n11938), .B2(n13571), .ZN(
        n7803) );
  OAI22_X1 U2273 ( .A1(n10728), .A2(n11932), .B1(n11938), .B2(n13570), .ZN(
        n7802) );
  OAI22_X1 U2274 ( .A1(n10721), .A2(n11932), .B1(n11938), .B2(n13569), .ZN(
        n7801) );
  OAI22_X1 U2275 ( .A1(n10714), .A2(n11932), .B1(n11938), .B2(n13568), .ZN(
        n7800) );
  OAI22_X1 U2276 ( .A1(n10707), .A2(n11931), .B1(n11939), .B2(n13567), .ZN(
        n7799) );
  OAI22_X1 U2277 ( .A1(n10700), .A2(n11931), .B1(n11939), .B2(n13566), .ZN(
        n7798) );
  OAI22_X1 U2278 ( .A1(n10693), .A2(n11931), .B1(n11939), .B2(n13565), .ZN(
        n7797) );
  OAI22_X1 U2279 ( .A1(n10686), .A2(n11931), .B1(n11939), .B2(n13564), .ZN(
        n7796) );
  OAI22_X1 U2280 ( .A1(n10679), .A2(n11931), .B1(n11940), .B2(n13563), .ZN(
        n7795) );
  OAI22_X1 U2281 ( .A1(n10672), .A2(n11931), .B1(n11940), .B2(n13562), .ZN(
        n7794) );
  OAI22_X1 U2282 ( .A1(n10665), .A2(n11931), .B1(n11940), .B2(n13561), .ZN(
        n7793) );
  OAI22_X1 U2283 ( .A1(n10658), .A2(n11931), .B1(n11940), .B2(n13560), .ZN(
        n7792) );
  OAI22_X1 U2284 ( .A1(n10651), .A2(n11931), .B1(n11941), .B2(n13559), .ZN(
        n7791) );
  OAI22_X1 U2285 ( .A1(n10644), .A2(n11931), .B1(n11941), .B2(n13558), .ZN(
        n7790) );
  OAI22_X1 U2286 ( .A1(n10637), .A2(n11931), .B1(n11941), .B2(n13557), .ZN(
        n7789) );
  OAI22_X1 U2287 ( .A1(n10630), .A2(n11931), .B1(n11941), .B2(n13556), .ZN(
        n7788) );
  OAI22_X1 U2288 ( .A1(n10847), .A2(n11897), .B1(n11898), .B2(n13491), .ZN(
        n7723) );
  OAI22_X1 U2289 ( .A1(n10840), .A2(n11897), .B1(n11898), .B2(n13490), .ZN(
        n7722) );
  OAI22_X1 U2290 ( .A1(n10833), .A2(n11897), .B1(n11898), .B2(n13489), .ZN(
        n7721) );
  OAI22_X1 U2291 ( .A1(n10826), .A2(n11897), .B1(n11898), .B2(n13488), .ZN(
        n7720) );
  OAI22_X1 U2292 ( .A1(n10819), .A2(n11897), .B1(n11899), .B2(n13487), .ZN(
        n7719) );
  OAI22_X1 U2293 ( .A1(n10812), .A2(n11897), .B1(n11899), .B2(n13486), .ZN(
        n7718) );
  OAI22_X1 U2294 ( .A1(n10805), .A2(n11897), .B1(n11899), .B2(n13485), .ZN(
        n7717) );
  OAI22_X1 U2295 ( .A1(n10798), .A2(n11897), .B1(n11899), .B2(n13484), .ZN(
        n7716) );
  OAI22_X1 U2296 ( .A1(n10791), .A2(n11896), .B1(n11900), .B2(n13483), .ZN(
        n7715) );
  OAI22_X1 U2297 ( .A1(n10784), .A2(n11896), .B1(n11900), .B2(n13482), .ZN(
        n7714) );
  OAI22_X1 U2298 ( .A1(n10777), .A2(n11896), .B1(n11900), .B2(n13481), .ZN(
        n7713) );
  OAI22_X1 U2299 ( .A1(n10770), .A2(n11896), .B1(n11900), .B2(n13480), .ZN(
        n7712) );
  OAI22_X1 U2300 ( .A1(n10763), .A2(n11896), .B1(n11901), .B2(n13479), .ZN(
        n7711) );
  OAI22_X1 U2301 ( .A1(n10756), .A2(n11896), .B1(n11901), .B2(n13478), .ZN(
        n7710) );
  OAI22_X1 U2302 ( .A1(n10749), .A2(n11896), .B1(n11901), .B2(n13477), .ZN(
        n7709) );
  OAI22_X1 U2303 ( .A1(n10742), .A2(n11896), .B1(n11901), .B2(n13476), .ZN(
        n7708) );
  OAI22_X1 U2304 ( .A1(n10735), .A2(n11896), .B1(n11902), .B2(n13475), .ZN(
        n7707) );
  OAI22_X1 U2305 ( .A1(n10728), .A2(n11896), .B1(n11902), .B2(n13474), .ZN(
        n7706) );
  OAI22_X1 U2306 ( .A1(n10721), .A2(n11896), .B1(n11902), .B2(n13473), .ZN(
        n7705) );
  OAI22_X1 U2307 ( .A1(n10714), .A2(n11896), .B1(n11902), .B2(n13472), .ZN(
        n7704) );
  OAI22_X1 U2308 ( .A1(n10707), .A2(n11895), .B1(n11903), .B2(n13471), .ZN(
        n7703) );
  OAI22_X1 U2309 ( .A1(n10700), .A2(n11895), .B1(n11903), .B2(n13470), .ZN(
        n7702) );
  OAI22_X1 U2310 ( .A1(n10693), .A2(n11895), .B1(n11903), .B2(n13469), .ZN(
        n7701) );
  OAI22_X1 U2311 ( .A1(n10686), .A2(n11895), .B1(n11903), .B2(n13468), .ZN(
        n7700) );
  OAI22_X1 U2312 ( .A1(n10679), .A2(n11895), .B1(n11904), .B2(n13467), .ZN(
        n7699) );
  OAI22_X1 U2313 ( .A1(n10672), .A2(n11895), .B1(n11904), .B2(n13466), .ZN(
        n7698) );
  OAI22_X1 U2314 ( .A1(n10665), .A2(n11895), .B1(n11904), .B2(n13465), .ZN(
        n7697) );
  OAI22_X1 U2315 ( .A1(n10658), .A2(n11895), .B1(n11904), .B2(n13464), .ZN(
        n7696) );
  OAI22_X1 U2316 ( .A1(n10651), .A2(n11895), .B1(n11905), .B2(n13463), .ZN(
        n7695) );
  OAI22_X1 U2317 ( .A1(n10644), .A2(n11895), .B1(n11905), .B2(n13462), .ZN(
        n7694) );
  OAI22_X1 U2318 ( .A1(n10637), .A2(n11895), .B1(n11905), .B2(n13461), .ZN(
        n7693) );
  OAI22_X1 U2319 ( .A1(n10630), .A2(n11895), .B1(n11905), .B2(n13460), .ZN(
        n7692) );
  OAI22_X1 U2320 ( .A1(n10847), .A2(n11873), .B1(n11874), .B2(n13459), .ZN(
        n7659) );
  OAI22_X1 U2321 ( .A1(n10840), .A2(n11873), .B1(n11874), .B2(n13458), .ZN(
        n7658) );
  OAI22_X1 U2322 ( .A1(n10833), .A2(n11873), .B1(n11874), .B2(n13457), .ZN(
        n7657) );
  OAI22_X1 U2323 ( .A1(n10826), .A2(n11873), .B1(n11874), .B2(n13456), .ZN(
        n7656) );
  OAI22_X1 U2324 ( .A1(n10819), .A2(n11873), .B1(n11875), .B2(n13455), .ZN(
        n7655) );
  OAI22_X1 U2325 ( .A1(n10812), .A2(n11873), .B1(n11875), .B2(n13454), .ZN(
        n7654) );
  OAI22_X1 U2326 ( .A1(n10805), .A2(n11873), .B1(n11875), .B2(n13453), .ZN(
        n7653) );
  OAI22_X1 U2327 ( .A1(n10798), .A2(n11873), .B1(n11875), .B2(n13452), .ZN(
        n7652) );
  OAI22_X1 U2328 ( .A1(n10791), .A2(n11872), .B1(n11876), .B2(n13451), .ZN(
        n7651) );
  OAI22_X1 U2329 ( .A1(n10784), .A2(n11872), .B1(n11876), .B2(n13450), .ZN(
        n7650) );
  OAI22_X1 U2330 ( .A1(n10777), .A2(n11872), .B1(n11876), .B2(n13449), .ZN(
        n7649) );
  OAI22_X1 U2331 ( .A1(n10770), .A2(n11872), .B1(n11876), .B2(n13448), .ZN(
        n7648) );
  OAI22_X1 U2332 ( .A1(n10763), .A2(n11872), .B1(n11877), .B2(n13447), .ZN(
        n7647) );
  OAI22_X1 U2333 ( .A1(n10756), .A2(n11872), .B1(n11877), .B2(n13446), .ZN(
        n7646) );
  OAI22_X1 U2334 ( .A1(n10749), .A2(n11872), .B1(n11877), .B2(n13445), .ZN(
        n7645) );
  OAI22_X1 U2335 ( .A1(n10742), .A2(n11872), .B1(n11877), .B2(n13444), .ZN(
        n7644) );
  OAI22_X1 U2336 ( .A1(n10735), .A2(n11872), .B1(n11878), .B2(n13443), .ZN(
        n7643) );
  OAI22_X1 U2337 ( .A1(n10728), .A2(n11872), .B1(n11878), .B2(n13442), .ZN(
        n7642) );
  OAI22_X1 U2338 ( .A1(n10721), .A2(n11872), .B1(n11878), .B2(n13441), .ZN(
        n7641) );
  OAI22_X1 U2339 ( .A1(n10714), .A2(n11872), .B1(n11878), .B2(n13440), .ZN(
        n7640) );
  OAI22_X1 U2340 ( .A1(n10707), .A2(n11871), .B1(n11879), .B2(n13439), .ZN(
        n7639) );
  OAI22_X1 U2341 ( .A1(n10700), .A2(n11871), .B1(n11879), .B2(n13438), .ZN(
        n7638) );
  OAI22_X1 U2342 ( .A1(n10693), .A2(n11871), .B1(n11879), .B2(n13437), .ZN(
        n7637) );
  OAI22_X1 U2343 ( .A1(n10686), .A2(n11871), .B1(n11879), .B2(n13436), .ZN(
        n7636) );
  OAI22_X1 U2344 ( .A1(n10679), .A2(n11871), .B1(n11880), .B2(n13435), .ZN(
        n7635) );
  OAI22_X1 U2345 ( .A1(n10672), .A2(n11871), .B1(n11880), .B2(n13434), .ZN(
        n7634) );
  OAI22_X1 U2346 ( .A1(n10665), .A2(n11871), .B1(n11880), .B2(n13433), .ZN(
        n7633) );
  OAI22_X1 U2347 ( .A1(n10658), .A2(n11871), .B1(n11880), .B2(n13432), .ZN(
        n7632) );
  OAI22_X1 U2348 ( .A1(n10651), .A2(n11871), .B1(n11881), .B2(n13431), .ZN(
        n7631) );
  OAI22_X1 U2349 ( .A1(n10644), .A2(n11871), .B1(n11881), .B2(n13430), .ZN(
        n7630) );
  OAI22_X1 U2350 ( .A1(n10637), .A2(n11871), .B1(n11881), .B2(n13429), .ZN(
        n7629) );
  OAI22_X1 U2351 ( .A1(n10630), .A2(n11871), .B1(n11881), .B2(n13428), .ZN(
        n7628) );
  OAI22_X1 U2352 ( .A1(n10847), .A2(n11849), .B1(n11850), .B2(n13427), .ZN(
        n7595) );
  OAI22_X1 U2353 ( .A1(n10840), .A2(n11849), .B1(n11850), .B2(n13426), .ZN(
        n7594) );
  OAI22_X1 U2354 ( .A1(n10833), .A2(n11849), .B1(n11850), .B2(n13425), .ZN(
        n7593) );
  OAI22_X1 U2355 ( .A1(n10826), .A2(n11849), .B1(n11850), .B2(n13424), .ZN(
        n7592) );
  OAI22_X1 U2356 ( .A1(n10819), .A2(n11849), .B1(n11851), .B2(n13423), .ZN(
        n7591) );
  OAI22_X1 U2357 ( .A1(n10812), .A2(n11849), .B1(n11851), .B2(n13422), .ZN(
        n7590) );
  OAI22_X1 U2358 ( .A1(n10805), .A2(n11849), .B1(n11851), .B2(n13421), .ZN(
        n7589) );
  OAI22_X1 U2359 ( .A1(n10798), .A2(n11849), .B1(n11851), .B2(n13420), .ZN(
        n7588) );
  OAI22_X1 U2360 ( .A1(n10791), .A2(n11848), .B1(n11852), .B2(n13419), .ZN(
        n7587) );
  OAI22_X1 U2361 ( .A1(n10784), .A2(n11848), .B1(n11852), .B2(n13418), .ZN(
        n7586) );
  OAI22_X1 U2362 ( .A1(n10777), .A2(n11848), .B1(n11852), .B2(n13417), .ZN(
        n7585) );
  OAI22_X1 U2363 ( .A1(n10770), .A2(n11848), .B1(n11852), .B2(n13416), .ZN(
        n7584) );
  OAI22_X1 U2364 ( .A1(n10763), .A2(n11848), .B1(n11853), .B2(n13415), .ZN(
        n7583) );
  OAI22_X1 U2365 ( .A1(n10756), .A2(n11848), .B1(n11853), .B2(n13414), .ZN(
        n7582) );
  OAI22_X1 U2366 ( .A1(n10749), .A2(n11848), .B1(n11853), .B2(n13413), .ZN(
        n7581) );
  OAI22_X1 U2367 ( .A1(n10742), .A2(n11848), .B1(n11853), .B2(n13412), .ZN(
        n7580) );
  OAI22_X1 U2368 ( .A1(n10735), .A2(n11848), .B1(n11854), .B2(n13411), .ZN(
        n7579) );
  OAI22_X1 U2369 ( .A1(n10728), .A2(n11848), .B1(n11854), .B2(n13410), .ZN(
        n7578) );
  OAI22_X1 U2370 ( .A1(n10721), .A2(n11848), .B1(n11854), .B2(n13409), .ZN(
        n7577) );
  OAI22_X1 U2371 ( .A1(n10714), .A2(n11848), .B1(n11854), .B2(n13408), .ZN(
        n7576) );
  OAI22_X1 U2372 ( .A1(n10707), .A2(n11847), .B1(n11855), .B2(n13407), .ZN(
        n7575) );
  OAI22_X1 U2373 ( .A1(n10700), .A2(n11847), .B1(n11855), .B2(n13406), .ZN(
        n7574) );
  OAI22_X1 U2374 ( .A1(n10693), .A2(n11847), .B1(n11855), .B2(n13405), .ZN(
        n7573) );
  OAI22_X1 U2375 ( .A1(n10686), .A2(n11847), .B1(n11855), .B2(n13404), .ZN(
        n7572) );
  OAI22_X1 U2376 ( .A1(n10679), .A2(n11847), .B1(n11856), .B2(n13403), .ZN(
        n7571) );
  OAI22_X1 U2377 ( .A1(n10672), .A2(n11847), .B1(n11856), .B2(n13402), .ZN(
        n7570) );
  OAI22_X1 U2378 ( .A1(n10665), .A2(n11847), .B1(n11856), .B2(n13401), .ZN(
        n7569) );
  OAI22_X1 U2379 ( .A1(n10658), .A2(n11847), .B1(n11856), .B2(n13400), .ZN(
        n7568) );
  OAI22_X1 U2380 ( .A1(n10651), .A2(n11847), .B1(n11857), .B2(n13399), .ZN(
        n7567) );
  OAI22_X1 U2381 ( .A1(n10644), .A2(n11847), .B1(n11857), .B2(n13398), .ZN(
        n7566) );
  OAI22_X1 U2382 ( .A1(n10637), .A2(n11847), .B1(n11857), .B2(n13397), .ZN(
        n7565) );
  OAI22_X1 U2383 ( .A1(n10630), .A2(n11847), .B1(n11857), .B2(n13396), .ZN(
        n7564) );
  OAI22_X1 U2384 ( .A1(n10848), .A2(n11693), .B1(n11694), .B2(n13203), .ZN(
        n7179) );
  OAI22_X1 U2385 ( .A1(n10841), .A2(n11693), .B1(n11694), .B2(n13202), .ZN(
        n7178) );
  OAI22_X1 U2386 ( .A1(n10834), .A2(n11693), .B1(n11694), .B2(n13201), .ZN(
        n7177) );
  OAI22_X1 U2387 ( .A1(n10827), .A2(n11693), .B1(n11694), .B2(n13200), .ZN(
        n7176) );
  OAI22_X1 U2388 ( .A1(n10820), .A2(n11693), .B1(n11695), .B2(n13199), .ZN(
        n7175) );
  OAI22_X1 U2389 ( .A1(n10813), .A2(n11693), .B1(n11695), .B2(n13198), .ZN(
        n7174) );
  OAI22_X1 U2390 ( .A1(n10806), .A2(n11693), .B1(n11695), .B2(n13197), .ZN(
        n7173) );
  OAI22_X1 U2391 ( .A1(n10799), .A2(n11693), .B1(n11695), .B2(n13196), .ZN(
        n7172) );
  OAI22_X1 U2392 ( .A1(n10792), .A2(n11692), .B1(n11696), .B2(n13195), .ZN(
        n7171) );
  OAI22_X1 U2393 ( .A1(n10785), .A2(n11692), .B1(n11696), .B2(n13194), .ZN(
        n7170) );
  OAI22_X1 U2394 ( .A1(n10778), .A2(n11692), .B1(n11696), .B2(n13193), .ZN(
        n7169) );
  OAI22_X1 U2395 ( .A1(n10771), .A2(n11692), .B1(n11696), .B2(n13192), .ZN(
        n7168) );
  OAI22_X1 U2396 ( .A1(n10764), .A2(n11692), .B1(n11697), .B2(n13191), .ZN(
        n7167) );
  OAI22_X1 U2397 ( .A1(n10757), .A2(n11692), .B1(n11697), .B2(n13190), .ZN(
        n7166) );
  OAI22_X1 U2398 ( .A1(n10750), .A2(n11692), .B1(n11697), .B2(n13189), .ZN(
        n7165) );
  OAI22_X1 U2399 ( .A1(n10743), .A2(n11692), .B1(n11697), .B2(n13188), .ZN(
        n7164) );
  OAI22_X1 U2400 ( .A1(n10736), .A2(n11692), .B1(n11698), .B2(n13187), .ZN(
        n7163) );
  OAI22_X1 U2401 ( .A1(n10729), .A2(n11692), .B1(n11698), .B2(n13186), .ZN(
        n7162) );
  OAI22_X1 U2402 ( .A1(n10722), .A2(n11692), .B1(n11698), .B2(n13185), .ZN(
        n7161) );
  OAI22_X1 U2403 ( .A1(n10715), .A2(n11692), .B1(n11698), .B2(n13184), .ZN(
        n7160) );
  OAI22_X1 U2404 ( .A1(n10708), .A2(n11691), .B1(n11699), .B2(n13183), .ZN(
        n7159) );
  OAI22_X1 U2405 ( .A1(n10701), .A2(n11691), .B1(n11699), .B2(n13182), .ZN(
        n7158) );
  OAI22_X1 U2406 ( .A1(n10694), .A2(n11691), .B1(n11699), .B2(n13181), .ZN(
        n7157) );
  OAI22_X1 U2407 ( .A1(n10687), .A2(n11691), .B1(n11699), .B2(n13180), .ZN(
        n7156) );
  OAI22_X1 U2408 ( .A1(n10680), .A2(n11691), .B1(n11700), .B2(n13179), .ZN(
        n7155) );
  OAI22_X1 U2409 ( .A1(n10673), .A2(n11691), .B1(n11700), .B2(n13178), .ZN(
        n7154) );
  OAI22_X1 U2410 ( .A1(n10666), .A2(n11691), .B1(n11700), .B2(n13177), .ZN(
        n7153) );
  OAI22_X1 U2411 ( .A1(n10659), .A2(n11691), .B1(n11700), .B2(n13176), .ZN(
        n7152) );
  OAI22_X1 U2412 ( .A1(n10652), .A2(n11691), .B1(n11701), .B2(n13175), .ZN(
        n7151) );
  OAI22_X1 U2413 ( .A1(n10645), .A2(n11691), .B1(n11701), .B2(n13174), .ZN(
        n7150) );
  OAI22_X1 U2414 ( .A1(n10638), .A2(n11691), .B1(n11701), .B2(n13173), .ZN(
        n7149) );
  OAI22_X1 U2415 ( .A1(n10631), .A2(n11691), .B1(n11701), .B2(n13172), .ZN(
        n7148) );
  OAI22_X1 U2416 ( .A1(n10848), .A2(n11681), .B1(n11682), .B2(n13171), .ZN(
        n7147) );
  OAI22_X1 U2417 ( .A1(n10841), .A2(n11681), .B1(n11682), .B2(n13170), .ZN(
        n7146) );
  OAI22_X1 U2418 ( .A1(n10834), .A2(n11681), .B1(n11682), .B2(n13169), .ZN(
        n7145) );
  OAI22_X1 U2419 ( .A1(n10827), .A2(n11681), .B1(n11682), .B2(n13168), .ZN(
        n7144) );
  OAI22_X1 U2420 ( .A1(n10820), .A2(n11681), .B1(n11683), .B2(n13167), .ZN(
        n7143) );
  OAI22_X1 U2421 ( .A1(n10813), .A2(n11681), .B1(n11683), .B2(n13166), .ZN(
        n7142) );
  OAI22_X1 U2422 ( .A1(n10806), .A2(n11681), .B1(n11683), .B2(n13165), .ZN(
        n7141) );
  OAI22_X1 U2423 ( .A1(n10799), .A2(n11681), .B1(n11683), .B2(n13164), .ZN(
        n7140) );
  OAI22_X1 U2424 ( .A1(n10792), .A2(n11680), .B1(n11684), .B2(n13163), .ZN(
        n7139) );
  OAI22_X1 U2425 ( .A1(n10785), .A2(n11680), .B1(n11684), .B2(n13162), .ZN(
        n7138) );
  OAI22_X1 U2426 ( .A1(n10778), .A2(n11680), .B1(n11684), .B2(n13161), .ZN(
        n7137) );
  OAI22_X1 U2427 ( .A1(n10771), .A2(n11680), .B1(n11684), .B2(n13160), .ZN(
        n7136) );
  OAI22_X1 U2428 ( .A1(n10764), .A2(n11680), .B1(n11685), .B2(n13159), .ZN(
        n7135) );
  OAI22_X1 U2429 ( .A1(n10757), .A2(n11680), .B1(n11685), .B2(n13158), .ZN(
        n7134) );
  OAI22_X1 U2430 ( .A1(n10750), .A2(n11680), .B1(n11685), .B2(n13157), .ZN(
        n7133) );
  OAI22_X1 U2431 ( .A1(n10743), .A2(n11680), .B1(n11685), .B2(n13156), .ZN(
        n7132) );
  OAI22_X1 U2432 ( .A1(n10736), .A2(n11680), .B1(n11686), .B2(n13155), .ZN(
        n7131) );
  OAI22_X1 U2433 ( .A1(n10729), .A2(n11680), .B1(n11686), .B2(n13154), .ZN(
        n7130) );
  OAI22_X1 U2434 ( .A1(n10722), .A2(n11680), .B1(n11686), .B2(n13153), .ZN(
        n7129) );
  OAI22_X1 U2435 ( .A1(n10715), .A2(n11680), .B1(n11686), .B2(n13152), .ZN(
        n7128) );
  OAI22_X1 U2436 ( .A1(n10708), .A2(n11679), .B1(n11687), .B2(n13151), .ZN(
        n7127) );
  OAI22_X1 U2437 ( .A1(n10701), .A2(n11679), .B1(n11687), .B2(n13150), .ZN(
        n7126) );
  OAI22_X1 U2438 ( .A1(n10694), .A2(n11679), .B1(n11687), .B2(n13149), .ZN(
        n7125) );
  OAI22_X1 U2439 ( .A1(n10687), .A2(n11679), .B1(n11687), .B2(n13148), .ZN(
        n7124) );
  OAI22_X1 U2440 ( .A1(n10680), .A2(n11679), .B1(n11688), .B2(n13147), .ZN(
        n7123) );
  OAI22_X1 U2441 ( .A1(n10673), .A2(n11679), .B1(n11688), .B2(n13146), .ZN(
        n7122) );
  OAI22_X1 U2442 ( .A1(n10666), .A2(n11679), .B1(n11688), .B2(n13145), .ZN(
        n7121) );
  OAI22_X1 U2443 ( .A1(n10659), .A2(n11679), .B1(n11688), .B2(n13144), .ZN(
        n7120) );
  OAI22_X1 U2444 ( .A1(n10652), .A2(n11679), .B1(n11689), .B2(n13143), .ZN(
        n7119) );
  OAI22_X1 U2445 ( .A1(n10645), .A2(n11679), .B1(n11689), .B2(n13142), .ZN(
        n7118) );
  OAI22_X1 U2446 ( .A1(n10638), .A2(n11679), .B1(n11689), .B2(n13141), .ZN(
        n7117) );
  OAI22_X1 U2447 ( .A1(n10631), .A2(n11679), .B1(n11689), .B2(n13140), .ZN(
        n7116) );
  OAI22_X1 U2448 ( .A1(n10848), .A2(n11669), .B1(n11670), .B2(n13139), .ZN(
        n7115) );
  OAI22_X1 U2449 ( .A1(n10841), .A2(n11669), .B1(n11670), .B2(n13138), .ZN(
        n7114) );
  OAI22_X1 U2450 ( .A1(n10834), .A2(n11669), .B1(n11670), .B2(n13137), .ZN(
        n7113) );
  OAI22_X1 U2451 ( .A1(n10827), .A2(n11669), .B1(n11670), .B2(n13136), .ZN(
        n7112) );
  OAI22_X1 U2452 ( .A1(n10820), .A2(n11669), .B1(n11671), .B2(n13135), .ZN(
        n7111) );
  OAI22_X1 U2453 ( .A1(n10813), .A2(n11669), .B1(n11671), .B2(n13134), .ZN(
        n7110) );
  OAI22_X1 U2454 ( .A1(n10806), .A2(n11669), .B1(n11671), .B2(n13133), .ZN(
        n7109) );
  OAI22_X1 U2455 ( .A1(n10799), .A2(n11669), .B1(n11671), .B2(n13132), .ZN(
        n7108) );
  OAI22_X1 U2456 ( .A1(n10792), .A2(n11668), .B1(n11672), .B2(n13131), .ZN(
        n7107) );
  OAI22_X1 U2457 ( .A1(n10785), .A2(n11668), .B1(n11672), .B2(n13130), .ZN(
        n7106) );
  OAI22_X1 U2458 ( .A1(n10778), .A2(n11668), .B1(n11672), .B2(n13129), .ZN(
        n7105) );
  OAI22_X1 U2459 ( .A1(n10771), .A2(n11668), .B1(n11672), .B2(n13128), .ZN(
        n7104) );
  OAI22_X1 U2460 ( .A1(n10764), .A2(n11668), .B1(n11673), .B2(n13127), .ZN(
        n7103) );
  OAI22_X1 U2461 ( .A1(n10757), .A2(n11668), .B1(n11673), .B2(n13126), .ZN(
        n7102) );
  OAI22_X1 U2462 ( .A1(n10750), .A2(n11668), .B1(n11673), .B2(n13125), .ZN(
        n7101) );
  OAI22_X1 U2463 ( .A1(n10743), .A2(n11668), .B1(n11673), .B2(n13124), .ZN(
        n7100) );
  OAI22_X1 U2464 ( .A1(n10736), .A2(n11668), .B1(n11674), .B2(n13123), .ZN(
        n7099) );
  OAI22_X1 U2465 ( .A1(n10729), .A2(n11668), .B1(n11674), .B2(n13122), .ZN(
        n7098) );
  OAI22_X1 U2466 ( .A1(n10722), .A2(n11668), .B1(n11674), .B2(n13121), .ZN(
        n7097) );
  OAI22_X1 U2467 ( .A1(n10715), .A2(n11668), .B1(n11674), .B2(n13120), .ZN(
        n7096) );
  OAI22_X1 U2468 ( .A1(n10708), .A2(n11667), .B1(n11675), .B2(n13119), .ZN(
        n7095) );
  OAI22_X1 U2469 ( .A1(n10701), .A2(n11667), .B1(n11675), .B2(n13118), .ZN(
        n7094) );
  OAI22_X1 U2470 ( .A1(n10694), .A2(n11667), .B1(n11675), .B2(n13117), .ZN(
        n7093) );
  OAI22_X1 U2471 ( .A1(n10687), .A2(n11667), .B1(n11675), .B2(n13116), .ZN(
        n7092) );
  OAI22_X1 U2472 ( .A1(n10680), .A2(n11667), .B1(n11676), .B2(n13115), .ZN(
        n7091) );
  OAI22_X1 U2473 ( .A1(n10673), .A2(n11667), .B1(n11676), .B2(n13114), .ZN(
        n7090) );
  OAI22_X1 U2474 ( .A1(n10666), .A2(n11667), .B1(n11676), .B2(n13113), .ZN(
        n7089) );
  OAI22_X1 U2475 ( .A1(n10659), .A2(n11667), .B1(n11676), .B2(n13112), .ZN(
        n7088) );
  OAI22_X1 U2476 ( .A1(n10652), .A2(n11667), .B1(n11677), .B2(n13111), .ZN(
        n7087) );
  OAI22_X1 U2477 ( .A1(n10645), .A2(n11667), .B1(n11677), .B2(n13110), .ZN(
        n7086) );
  OAI22_X1 U2478 ( .A1(n10638), .A2(n11667), .B1(n11677), .B2(n13109), .ZN(
        n7085) );
  OAI22_X1 U2479 ( .A1(n10631), .A2(n11667), .B1(n11677), .B2(n13108), .ZN(
        n7084) );
  OAI22_X1 U2480 ( .A1(n10640), .A2(n11475), .B1(n11485), .B2(n12787), .ZN(
        n6573) );
  OAI22_X1 U2481 ( .A1(n10633), .A2(n11475), .B1(n11485), .B2(n12786), .ZN(
        n6572) );
  OAI22_X1 U2482 ( .A1(n10647), .A2(n11439), .B1(n11449), .B2(n12785), .ZN(
        n6478) );
  OAI22_X1 U2483 ( .A1(n10640), .A2(n11439), .B1(n11449), .B2(n12784), .ZN(
        n6477) );
  OAI22_X1 U2484 ( .A1(n10633), .A2(n11439), .B1(n11449), .B2(n12783), .ZN(
        n6476) );
  OAI22_X1 U2485 ( .A1(n10647), .A2(n11403), .B1(n11413), .B2(n12782), .ZN(
        n6382) );
  OAI22_X1 U2486 ( .A1(n10640), .A2(n11403), .B1(n11413), .B2(n12781), .ZN(
        n6381) );
  OAI22_X1 U2487 ( .A1(n10633), .A2(n11403), .B1(n11413), .B2(n12780), .ZN(
        n6380) );
  INV_X1 U2488 ( .A(n2478), .ZN(n14517) );
  INV_X1 U2489 ( .A(n2481), .ZN(n12777) );
  NAND2_X1 U2490 ( .A1(n10625), .A2(n10626), .ZN(n2487) );
  INV_X1 U2491 ( .A(n2477), .ZN(n12778) );
  AOI21_X1 U2492 ( .B1(n10625), .B2(n2478), .A(n2479), .ZN(n2477) );
  AOI21_X1 U2493 ( .B1(n2480), .B2(n2481), .A(n10625), .ZN(n2479) );
  AOI222_X1 U2494 ( .A1(n11064), .A2(n12979), .B1(n11061), .B2(n12915), .C1(
        n11058), .C2(n13043), .ZN(n5639) );
  AOI222_X1 U2495 ( .A1(n10866), .A2(n14448), .B1(n10863), .B2(n14384), .C1(
        n10860), .C2(n14512), .ZN(n5694) );
  AOI222_X1 U2496 ( .A1(n11328), .A2(n12979), .B1(n11325), .B2(n12915), .C1(
        n11322), .C2(n13043), .ZN(n4206) );
  AOI222_X1 U2497 ( .A1(n11130), .A2(n14448), .B1(n11127), .B2(n14384), .C1(
        n11124), .C2(n14512), .ZN(n4261) );
  AOI222_X1 U2498 ( .A1(n11064), .A2(n12978), .B1(n11061), .B2(n12914), .C1(
        n11058), .C2(n13042), .ZN(n5598) );
  AOI222_X1 U2499 ( .A1(n10866), .A2(n14447), .B1(n10863), .B2(n14383), .C1(
        n10860), .C2(n14511), .ZN(n5625) );
  AOI222_X1 U2500 ( .A1(n11328), .A2(n12978), .B1(n11325), .B2(n12914), .C1(
        n11322), .C2(n13042), .ZN(n4165) );
  AOI222_X1 U2501 ( .A1(n11130), .A2(n14447), .B1(n11127), .B2(n14383), .C1(
        n11124), .C2(n14511), .ZN(n4192) );
  AOI222_X1 U2502 ( .A1(n11064), .A2(n12977), .B1(n11061), .B2(n12913), .C1(
        n11058), .C2(n13041), .ZN(n5557) );
  AOI222_X1 U2503 ( .A1(n10866), .A2(n14446), .B1(n10863), .B2(n14382), .C1(
        n10860), .C2(n14510), .ZN(n5584) );
  AOI222_X1 U2504 ( .A1(n11328), .A2(n12977), .B1(n11325), .B2(n12913), .C1(
        n11322), .C2(n13041), .ZN(n4124) );
  AOI222_X1 U2505 ( .A1(n11130), .A2(n14446), .B1(n11127), .B2(n14382), .C1(
        n11124), .C2(n14510), .ZN(n4151) );
  AOI222_X1 U2506 ( .A1(n11064), .A2(n12976), .B1(n11061), .B2(n12912), .C1(
        n11058), .C2(n13040), .ZN(n5516) );
  AOI222_X1 U2507 ( .A1(n10866), .A2(n14445), .B1(n10863), .B2(n14381), .C1(
        n10860), .C2(n14509), .ZN(n5543) );
  AOI222_X1 U2508 ( .A1(n11328), .A2(n12976), .B1(n11325), .B2(n12912), .C1(
        n11322), .C2(n13040), .ZN(n4083) );
  AOI222_X1 U2509 ( .A1(n11130), .A2(n14445), .B1(n11127), .B2(n14381), .C1(
        n11124), .C2(n14509), .ZN(n4110) );
  AOI222_X1 U2510 ( .A1(n11064), .A2(n12975), .B1(n11061), .B2(n12911), .C1(
        n11058), .C2(n13039), .ZN(n5475) );
  AOI222_X1 U2511 ( .A1(n10866), .A2(n14444), .B1(n10863), .B2(n14380), .C1(
        n10860), .C2(n14508), .ZN(n5502) );
  AOI222_X1 U2512 ( .A1(n11328), .A2(n12975), .B1(n11325), .B2(n12911), .C1(
        n11322), .C2(n13039), .ZN(n4042) );
  AOI222_X1 U2513 ( .A1(n11130), .A2(n14444), .B1(n11127), .B2(n14380), .C1(
        n11124), .C2(n14508), .ZN(n4069) );
  AOI222_X1 U2514 ( .A1(n11064), .A2(n12974), .B1(n11061), .B2(n12910), .C1(
        n11058), .C2(n13038), .ZN(n5434) );
  AOI222_X1 U2515 ( .A1(n10866), .A2(n14443), .B1(n10863), .B2(n14379), .C1(
        n10860), .C2(n14507), .ZN(n5461) );
  AOI222_X1 U2516 ( .A1(n11328), .A2(n12974), .B1(n11325), .B2(n12910), .C1(
        n11322), .C2(n13038), .ZN(n4001) );
  AOI222_X1 U2517 ( .A1(n11130), .A2(n14443), .B1(n11127), .B2(n14379), .C1(
        n11124), .C2(n14507), .ZN(n4028) );
  AOI222_X1 U2518 ( .A1(n11064), .A2(n12973), .B1(n11061), .B2(n12909), .C1(
        n11058), .C2(n13037), .ZN(n5393) );
  AOI222_X1 U2519 ( .A1(n10866), .A2(n14442), .B1(n10863), .B2(n14378), .C1(
        n10860), .C2(n14506), .ZN(n5420) );
  AOI222_X1 U2520 ( .A1(n11328), .A2(n12973), .B1(n11325), .B2(n12909), .C1(
        n11322), .C2(n13037), .ZN(n3960) );
  AOI222_X1 U2521 ( .A1(n11130), .A2(n14442), .B1(n11127), .B2(n14378), .C1(
        n11124), .C2(n14506), .ZN(n3987) );
  AOI222_X1 U2522 ( .A1(n11064), .A2(n12972), .B1(n11061), .B2(n12908), .C1(
        n11058), .C2(n13036), .ZN(n5352) );
  AOI222_X1 U2523 ( .A1(n10866), .A2(n14441), .B1(n10863), .B2(n14377), .C1(
        n10860), .C2(n14505), .ZN(n5379) );
  AOI222_X1 U2524 ( .A1(n11328), .A2(n12972), .B1(n11325), .B2(n12908), .C1(
        n11322), .C2(n13036), .ZN(n3919) );
  AOI222_X1 U2525 ( .A1(n11130), .A2(n14441), .B1(n11127), .B2(n14377), .C1(
        n11124), .C2(n14505), .ZN(n3946) );
  AOI222_X1 U2526 ( .A1(n11064), .A2(n12971), .B1(n11061), .B2(n12907), .C1(
        n11058), .C2(n13035), .ZN(n5311) );
  AOI222_X1 U2527 ( .A1(n10866), .A2(n14440), .B1(n10863), .B2(n14376), .C1(
        n10860), .C2(n14504), .ZN(n5338) );
  AOI222_X1 U2528 ( .A1(n11328), .A2(n12971), .B1(n11325), .B2(n12907), .C1(
        n11322), .C2(n13035), .ZN(n3878) );
  AOI222_X1 U2529 ( .A1(n11130), .A2(n14440), .B1(n11127), .B2(n14376), .C1(
        n11124), .C2(n14504), .ZN(n3905) );
  AOI222_X1 U2530 ( .A1(n11064), .A2(n12970), .B1(n11061), .B2(n12906), .C1(
        n11058), .C2(n13034), .ZN(n5270) );
  AOI222_X1 U2531 ( .A1(n10866), .A2(n14439), .B1(n10863), .B2(n14375), .C1(
        n10860), .C2(n14503), .ZN(n5297) );
  AOI222_X1 U2532 ( .A1(n11328), .A2(n12970), .B1(n11325), .B2(n12906), .C1(
        n11322), .C2(n13034), .ZN(n3837) );
  AOI222_X1 U2533 ( .A1(n11130), .A2(n14439), .B1(n11127), .B2(n14375), .C1(
        n11124), .C2(n14503), .ZN(n3864) );
  AOI222_X1 U2534 ( .A1(n11064), .A2(n12969), .B1(n11061), .B2(n12905), .C1(
        n11058), .C2(n13033), .ZN(n5229) );
  AOI222_X1 U2535 ( .A1(n10866), .A2(n14438), .B1(n10863), .B2(n14374), .C1(
        n10860), .C2(n14502), .ZN(n5256) );
  AOI222_X1 U2536 ( .A1(n11328), .A2(n12969), .B1(n11325), .B2(n12905), .C1(
        n11322), .C2(n13033), .ZN(n3796) );
  AOI222_X1 U2537 ( .A1(n11130), .A2(n14438), .B1(n11127), .B2(n14374), .C1(
        n11124), .C2(n14502), .ZN(n3823) );
  AOI222_X1 U2538 ( .A1(n11064), .A2(n12968), .B1(n11061), .B2(n12904), .C1(
        n11058), .C2(n13032), .ZN(n5188) );
  AOI222_X1 U2539 ( .A1(n10866), .A2(n14437), .B1(n10863), .B2(n14373), .C1(
        n10860), .C2(n14501), .ZN(n5215) );
  AOI222_X1 U2540 ( .A1(n11328), .A2(n12968), .B1(n11325), .B2(n12904), .C1(
        n11322), .C2(n13032), .ZN(n3755) );
  AOI222_X1 U2541 ( .A1(n11130), .A2(n14437), .B1(n11127), .B2(n14373), .C1(
        n11124), .C2(n14501), .ZN(n3782) );
  AOI222_X1 U2542 ( .A1(n11065), .A2(n12967), .B1(n11062), .B2(n12903), .C1(
        n11059), .C2(n13031), .ZN(n5147) );
  AOI222_X1 U2543 ( .A1(n10867), .A2(n14436), .B1(n10864), .B2(n14372), .C1(
        n10861), .C2(n14500), .ZN(n5174) );
  AOI222_X1 U2544 ( .A1(n11329), .A2(n12967), .B1(n11326), .B2(n12903), .C1(
        n11323), .C2(n13031), .ZN(n3714) );
  AOI222_X1 U2545 ( .A1(n11131), .A2(n14436), .B1(n11128), .B2(n14372), .C1(
        n11125), .C2(n14500), .ZN(n3741) );
  AOI222_X1 U2546 ( .A1(n11065), .A2(n12966), .B1(n11062), .B2(n12902), .C1(
        n11059), .C2(n13030), .ZN(n5106) );
  AOI222_X1 U2547 ( .A1(n10867), .A2(n14435), .B1(n10864), .B2(n14371), .C1(
        n10861), .C2(n14499), .ZN(n5133) );
  AOI222_X1 U2548 ( .A1(n11329), .A2(n12966), .B1(n11326), .B2(n12902), .C1(
        n11323), .C2(n13030), .ZN(n3673) );
  AOI222_X1 U2549 ( .A1(n11131), .A2(n14435), .B1(n11128), .B2(n14371), .C1(
        n11125), .C2(n14499), .ZN(n3700) );
  AOI222_X1 U2550 ( .A1(n11065), .A2(n12965), .B1(n11062), .B2(n12901), .C1(
        n11059), .C2(n13029), .ZN(n5065) );
  AOI222_X1 U2551 ( .A1(n10867), .A2(n14434), .B1(n10864), .B2(n14370), .C1(
        n10861), .C2(n14498), .ZN(n5092) );
  AOI222_X1 U2552 ( .A1(n11329), .A2(n12965), .B1(n11326), .B2(n12901), .C1(
        n11323), .C2(n13029), .ZN(n3632) );
  AOI222_X1 U2553 ( .A1(n11131), .A2(n14434), .B1(n11128), .B2(n14370), .C1(
        n11125), .C2(n14498), .ZN(n3659) );
  AOI222_X1 U2554 ( .A1(n11065), .A2(n12964), .B1(n11062), .B2(n12900), .C1(
        n11059), .C2(n13028), .ZN(n5024) );
  AOI222_X1 U2555 ( .A1(n10867), .A2(n14433), .B1(n10864), .B2(n14369), .C1(
        n10861), .C2(n14497), .ZN(n5051) );
  AOI222_X1 U2556 ( .A1(n11329), .A2(n12964), .B1(n11326), .B2(n12900), .C1(
        n11323), .C2(n13028), .ZN(n3591) );
  AOI222_X1 U2557 ( .A1(n11131), .A2(n14433), .B1(n11128), .B2(n14369), .C1(
        n11125), .C2(n14497), .ZN(n3618) );
  AOI222_X1 U2558 ( .A1(n11065), .A2(n12963), .B1(n11062), .B2(n12899), .C1(
        n11059), .C2(n13027), .ZN(n4983) );
  AOI222_X1 U2559 ( .A1(n10867), .A2(n14432), .B1(n10864), .B2(n14368), .C1(
        n10861), .C2(n14496), .ZN(n5010) );
  AOI222_X1 U2560 ( .A1(n11329), .A2(n12963), .B1(n11326), .B2(n12899), .C1(
        n11323), .C2(n13027), .ZN(n3550) );
  AOI222_X1 U2561 ( .A1(n11131), .A2(n14432), .B1(n11128), .B2(n14368), .C1(
        n11125), .C2(n14496), .ZN(n3577) );
  AOI222_X1 U2562 ( .A1(n11065), .A2(n12962), .B1(n11062), .B2(n12898), .C1(
        n11059), .C2(n13026), .ZN(n4942) );
  AOI222_X1 U2563 ( .A1(n10867), .A2(n14431), .B1(n10864), .B2(n14367), .C1(
        n10861), .C2(n14495), .ZN(n4969) );
  AOI222_X1 U2564 ( .A1(n11329), .A2(n12962), .B1(n11326), .B2(n12898), .C1(
        n11323), .C2(n13026), .ZN(n3509) );
  AOI222_X1 U2565 ( .A1(n11131), .A2(n14431), .B1(n11128), .B2(n14367), .C1(
        n11125), .C2(n14495), .ZN(n3536) );
  AOI222_X1 U2566 ( .A1(n11065), .A2(n12961), .B1(n11062), .B2(n12897), .C1(
        n11059), .C2(n13025), .ZN(n4901) );
  AOI222_X1 U2567 ( .A1(n10867), .A2(n14430), .B1(n10864), .B2(n14366), .C1(
        n10861), .C2(n14494), .ZN(n4928) );
  AOI222_X1 U2568 ( .A1(n11329), .A2(n12961), .B1(n11326), .B2(n12897), .C1(
        n11323), .C2(n13025), .ZN(n3468) );
  AOI222_X1 U2569 ( .A1(n11131), .A2(n14430), .B1(n11128), .B2(n14366), .C1(
        n11125), .C2(n14494), .ZN(n3495) );
  AOI222_X1 U2570 ( .A1(n11065), .A2(n12960), .B1(n11062), .B2(n12896), .C1(
        n11059), .C2(n13024), .ZN(n4860) );
  AOI222_X1 U2571 ( .A1(n10867), .A2(n14429), .B1(n10864), .B2(n14365), .C1(
        n10861), .C2(n14493), .ZN(n4887) );
  AOI222_X1 U2572 ( .A1(n11329), .A2(n12960), .B1(n11326), .B2(n12896), .C1(
        n11323), .C2(n13024), .ZN(n3427) );
  AOI222_X1 U2573 ( .A1(n11131), .A2(n14429), .B1(n11128), .B2(n14365), .C1(
        n11125), .C2(n14493), .ZN(n3454) );
  AOI222_X1 U2574 ( .A1(n11065), .A2(n12959), .B1(n11062), .B2(n12895), .C1(
        n11059), .C2(n13023), .ZN(n4819) );
  AOI222_X1 U2575 ( .A1(n10867), .A2(n14428), .B1(n10864), .B2(n14364), .C1(
        n10861), .C2(n14492), .ZN(n4846) );
  AOI222_X1 U2576 ( .A1(n11329), .A2(n12959), .B1(n11326), .B2(n12895), .C1(
        n11323), .C2(n13023), .ZN(n3386) );
  AOI222_X1 U2577 ( .A1(n11131), .A2(n14428), .B1(n11128), .B2(n14364), .C1(
        n11125), .C2(n14492), .ZN(n3413) );
  AOI222_X1 U2578 ( .A1(n11065), .A2(n12958), .B1(n11062), .B2(n12894), .C1(
        n11059), .C2(n13022), .ZN(n4778) );
  AOI222_X1 U2579 ( .A1(n10867), .A2(n14427), .B1(n10864), .B2(n14363), .C1(
        n10861), .C2(n14491), .ZN(n4805) );
  AOI222_X1 U2580 ( .A1(n11329), .A2(n12958), .B1(n11326), .B2(n12894), .C1(
        n11323), .C2(n13022), .ZN(n3345) );
  AOI222_X1 U2581 ( .A1(n11131), .A2(n14427), .B1(n11128), .B2(n14363), .C1(
        n11125), .C2(n14491), .ZN(n3372) );
  AOI222_X1 U2582 ( .A1(n11065), .A2(n12957), .B1(n11062), .B2(n12893), .C1(
        n11059), .C2(n13021), .ZN(n4737) );
  AOI222_X1 U2583 ( .A1(n10867), .A2(n14426), .B1(n10864), .B2(n14362), .C1(
        n10861), .C2(n14490), .ZN(n4764) );
  AOI222_X1 U2584 ( .A1(n11329), .A2(n12957), .B1(n11326), .B2(n12893), .C1(
        n11323), .C2(n13021), .ZN(n3304) );
  AOI222_X1 U2585 ( .A1(n11131), .A2(n14426), .B1(n11128), .B2(n14362), .C1(
        n11125), .C2(n14490), .ZN(n3331) );
  AOI222_X1 U2586 ( .A1(n11065), .A2(n12956), .B1(n11062), .B2(n12892), .C1(
        n11059), .C2(n13020), .ZN(n4696) );
  AOI222_X1 U2587 ( .A1(n10867), .A2(n14425), .B1(n10864), .B2(n14361), .C1(
        n10861), .C2(n14489), .ZN(n4723) );
  AOI222_X1 U2588 ( .A1(n11329), .A2(n12956), .B1(n11326), .B2(n12892), .C1(
        n11323), .C2(n13020), .ZN(n3263) );
  AOI222_X1 U2589 ( .A1(n11131), .A2(n14425), .B1(n11128), .B2(n14361), .C1(
        n11125), .C2(n14489), .ZN(n3290) );
  AOI222_X1 U2590 ( .A1(n11066), .A2(n12955), .B1(n11063), .B2(n12891), .C1(
        n11060), .C2(n13019), .ZN(n4655) );
  AOI222_X1 U2591 ( .A1(n10868), .A2(n14424), .B1(n10865), .B2(n14360), .C1(
        n10862), .C2(n14488), .ZN(n4682) );
  AOI222_X1 U2592 ( .A1(n11330), .A2(n12955), .B1(n11327), .B2(n12891), .C1(
        n11324), .C2(n13019), .ZN(n3222) );
  AOI222_X1 U2593 ( .A1(n11132), .A2(n14424), .B1(n11129), .B2(n14360), .C1(
        n11126), .C2(n14488), .ZN(n3249) );
  AOI222_X1 U2594 ( .A1(n11066), .A2(n12954), .B1(n11063), .B2(n12890), .C1(
        n11060), .C2(n13018), .ZN(n4614) );
  AOI222_X1 U2595 ( .A1(n10868), .A2(n14423), .B1(n10865), .B2(n14359), .C1(
        n10862), .C2(n14487), .ZN(n4641) );
  AOI222_X1 U2596 ( .A1(n11330), .A2(n12954), .B1(n11327), .B2(n12890), .C1(
        n11324), .C2(n13018), .ZN(n3181) );
  AOI222_X1 U2597 ( .A1(n11132), .A2(n14423), .B1(n11129), .B2(n14359), .C1(
        n11126), .C2(n14487), .ZN(n3208) );
  AOI222_X1 U2598 ( .A1(n11066), .A2(n12953), .B1(n11063), .B2(n12889), .C1(
        n11060), .C2(n13017), .ZN(n4573) );
  AOI222_X1 U2599 ( .A1(n10868), .A2(n14422), .B1(n10865), .B2(n14358), .C1(
        n10862), .C2(n14486), .ZN(n4600) );
  AOI222_X1 U2600 ( .A1(n11330), .A2(n12953), .B1(n11327), .B2(n12889), .C1(
        n11324), .C2(n13017), .ZN(n3140) );
  AOI222_X1 U2601 ( .A1(n11132), .A2(n14422), .B1(n11129), .B2(n14358), .C1(
        n11126), .C2(n14486), .ZN(n3167) );
  AOI222_X1 U2602 ( .A1(n11066), .A2(n12952), .B1(n11063), .B2(n12888), .C1(
        n11060), .C2(n13016), .ZN(n4532) );
  AOI222_X1 U2603 ( .A1(n10868), .A2(n14421), .B1(n10865), .B2(n14357), .C1(
        n10862), .C2(n14485), .ZN(n4559) );
  AOI222_X1 U2604 ( .A1(n11330), .A2(n12952), .B1(n11327), .B2(n12888), .C1(
        n11324), .C2(n13016), .ZN(n3099) );
  AOI222_X1 U2605 ( .A1(n11132), .A2(n14421), .B1(n11129), .B2(n14357), .C1(
        n11126), .C2(n14485), .ZN(n3126) );
  AOI222_X1 U2606 ( .A1(n11066), .A2(n12951), .B1(n11063), .B2(n12887), .C1(
        n11060), .C2(n13015), .ZN(n4491) );
  AOI222_X1 U2607 ( .A1(n10868), .A2(n14420), .B1(n10865), .B2(n14356), .C1(
        n10862), .C2(n14484), .ZN(n4518) );
  AOI222_X1 U2608 ( .A1(n11330), .A2(n12951), .B1(n11327), .B2(n12887), .C1(
        n11324), .C2(n13015), .ZN(n3058) );
  AOI222_X1 U2609 ( .A1(n11132), .A2(n14420), .B1(n11129), .B2(n14356), .C1(
        n11126), .C2(n14484), .ZN(n3085) );
  AOI222_X1 U2610 ( .A1(n11066), .A2(n12950), .B1(n11063), .B2(n12886), .C1(
        n11060), .C2(n13014), .ZN(n4450) );
  AOI222_X1 U2611 ( .A1(n10868), .A2(n14419), .B1(n10865), .B2(n14355), .C1(
        n10862), .C2(n14483), .ZN(n4477) );
  AOI222_X1 U2612 ( .A1(n11330), .A2(n12950), .B1(n11327), .B2(n12886), .C1(
        n11324), .C2(n13014), .ZN(n3017) );
  AOI222_X1 U2613 ( .A1(n11132), .A2(n14419), .B1(n11129), .B2(n14355), .C1(
        n11126), .C2(n14483), .ZN(n3044) );
  AOI222_X1 U2614 ( .A1(n11066), .A2(n12949), .B1(n11063), .B2(n12885), .C1(
        n11060), .C2(n13013), .ZN(n4409) );
  AOI222_X1 U2615 ( .A1(n10868), .A2(n14418), .B1(n10865), .B2(n14354), .C1(
        n10862), .C2(n14482), .ZN(n4436) );
  AOI222_X1 U2616 ( .A1(n11330), .A2(n12949), .B1(n11327), .B2(n12885), .C1(
        n11324), .C2(n13013), .ZN(n2976) );
  AOI222_X1 U2617 ( .A1(n11132), .A2(n14418), .B1(n11129), .B2(n14354), .C1(
        n11126), .C2(n14482), .ZN(n3003) );
  AOI222_X1 U2618 ( .A1(n11066), .A2(n12948), .B1(n11063), .B2(n12884), .C1(
        n11060), .C2(n13012), .ZN(n4280) );
  AOI222_X1 U2619 ( .A1(n10868), .A2(n14417), .B1(n10865), .B2(n14353), .C1(
        n10862), .C2(n14481), .ZN(n4373) );
  AOI222_X1 U2620 ( .A1(n11330), .A2(n12948), .B1(n11327), .B2(n12884), .C1(
        n11324), .C2(n13012), .ZN(n2748) );
  AOI222_X1 U2621 ( .A1(n11132), .A2(n14417), .B1(n11129), .B2(n14353), .C1(
        n11126), .C2(n14481), .ZN(n2940) );
  OAI222_X1 U2622 ( .A1(n14042), .A2(n10910), .B1(n14074), .B2(n10907), .C1(
        n14010), .C2(n10904), .ZN(n4687) );
  OAI222_X1 U2623 ( .A1(n14042), .A2(n11174), .B1(n14074), .B2(n11171), .C1(
        n14010), .C2(n11168), .ZN(n3254) );
  OAI222_X1 U2624 ( .A1(n14041), .A2(n10910), .B1(n14073), .B2(n10907), .C1(
        n14009), .C2(n10904), .ZN(n4646) );
  OAI222_X1 U2625 ( .A1(n14041), .A2(n11174), .B1(n14073), .B2(n11171), .C1(
        n14009), .C2(n11168), .ZN(n3213) );
  OAI222_X1 U2626 ( .A1(n14040), .A2(n10910), .B1(n14072), .B2(n10907), .C1(
        n14008), .C2(n10904), .ZN(n4605) );
  OAI222_X1 U2627 ( .A1(n14040), .A2(n11174), .B1(n14072), .B2(n11171), .C1(
        n14008), .C2(n11168), .ZN(n3172) );
  OAI222_X1 U2628 ( .A1(n14039), .A2(n10910), .B1(n14071), .B2(n10907), .C1(
        n14007), .C2(n10904), .ZN(n4564) );
  OAI222_X1 U2629 ( .A1(n14039), .A2(n11174), .B1(n14071), .B2(n11171), .C1(
        n14007), .C2(n11168), .ZN(n3131) );
  OAI222_X1 U2630 ( .A1(n14038), .A2(n10910), .B1(n14070), .B2(n10907), .C1(
        n14006), .C2(n10904), .ZN(n4523) );
  OAI222_X1 U2631 ( .A1(n14038), .A2(n11174), .B1(n14070), .B2(n11171), .C1(
        n14006), .C2(n11168), .ZN(n3090) );
  OAI222_X1 U2632 ( .A1(n14037), .A2(n10910), .B1(n14069), .B2(n10907), .C1(
        n14005), .C2(n10904), .ZN(n4482) );
  OAI222_X1 U2633 ( .A1(n14037), .A2(n11174), .B1(n14069), .B2(n11171), .C1(
        n14005), .C2(n11168), .ZN(n3049) );
  OAI222_X1 U2634 ( .A1(n14036), .A2(n10910), .B1(n14068), .B2(n10907), .C1(
        n14004), .C2(n10904), .ZN(n4441) );
  OAI222_X1 U2635 ( .A1(n14036), .A2(n11174), .B1(n14068), .B2(n11171), .C1(
        n14004), .C2(n11168), .ZN(n3008) );
  OAI222_X1 U2636 ( .A1(n14066), .A2(n10908), .B1(n14098), .B2(n10905), .C1(
        n14034), .C2(n10902), .ZN(n5699) );
  OAI222_X1 U2637 ( .A1(n14066), .A2(n11172), .B1(n14098), .B2(n11169), .C1(
        n14034), .C2(n11166), .ZN(n4266) );
  OAI222_X1 U2638 ( .A1(n14065), .A2(n10908), .B1(n14097), .B2(n10905), .C1(
        n14033), .C2(n10902), .ZN(n5630) );
  OAI222_X1 U2639 ( .A1(n14065), .A2(n11172), .B1(n14097), .B2(n11169), .C1(
        n14033), .C2(n11166), .ZN(n4197) );
  OAI222_X1 U2640 ( .A1(n14064), .A2(n10908), .B1(n14096), .B2(n10905), .C1(
        n14032), .C2(n10902), .ZN(n5589) );
  OAI222_X1 U2641 ( .A1(n14064), .A2(n11172), .B1(n14096), .B2(n11169), .C1(
        n14032), .C2(n11166), .ZN(n4156) );
  OAI222_X1 U2642 ( .A1(n14063), .A2(n10908), .B1(n14095), .B2(n10905), .C1(
        n14031), .C2(n10902), .ZN(n5548) );
  OAI222_X1 U2643 ( .A1(n14063), .A2(n11172), .B1(n14095), .B2(n11169), .C1(
        n14031), .C2(n11166), .ZN(n4115) );
  OAI222_X1 U2644 ( .A1(n14062), .A2(n10908), .B1(n14094), .B2(n10905), .C1(
        n14030), .C2(n10902), .ZN(n5507) );
  OAI222_X1 U2645 ( .A1(n14062), .A2(n11172), .B1(n14094), .B2(n11169), .C1(
        n14030), .C2(n11166), .ZN(n4074) );
  OAI222_X1 U2646 ( .A1(n14061), .A2(n10908), .B1(n14093), .B2(n10905), .C1(
        n14029), .C2(n10902), .ZN(n5466) );
  OAI222_X1 U2647 ( .A1(n14061), .A2(n11172), .B1(n14093), .B2(n11169), .C1(
        n14029), .C2(n11166), .ZN(n4033) );
  OAI222_X1 U2648 ( .A1(n14060), .A2(n10908), .B1(n14092), .B2(n10905), .C1(
        n14028), .C2(n10902), .ZN(n5425) );
  OAI222_X1 U2649 ( .A1(n14060), .A2(n11172), .B1(n14092), .B2(n11169), .C1(
        n14028), .C2(n11166), .ZN(n3992) );
  OAI222_X1 U2650 ( .A1(n14059), .A2(n10908), .B1(n14091), .B2(n10905), .C1(
        n14027), .C2(n10902), .ZN(n5384) );
  OAI222_X1 U2651 ( .A1(n14059), .A2(n11172), .B1(n14091), .B2(n11169), .C1(
        n14027), .C2(n11166), .ZN(n3951) );
  OAI222_X1 U2652 ( .A1(n14058), .A2(n10908), .B1(n14090), .B2(n10905), .C1(
        n14026), .C2(n10902), .ZN(n5343) );
  OAI222_X1 U2653 ( .A1(n14058), .A2(n11172), .B1(n14090), .B2(n11169), .C1(
        n14026), .C2(n11166), .ZN(n3910) );
  OAI222_X1 U2654 ( .A1(n14057), .A2(n10908), .B1(n14089), .B2(n10905), .C1(
        n14025), .C2(n10902), .ZN(n5302) );
  OAI222_X1 U2655 ( .A1(n14057), .A2(n11172), .B1(n14089), .B2(n11169), .C1(
        n14025), .C2(n11166), .ZN(n3869) );
  OAI222_X1 U2656 ( .A1(n14056), .A2(n10908), .B1(n14088), .B2(n10905), .C1(
        n14024), .C2(n10902), .ZN(n5261) );
  OAI222_X1 U2657 ( .A1(n14056), .A2(n11172), .B1(n14088), .B2(n11169), .C1(
        n14024), .C2(n11166), .ZN(n3828) );
  OAI222_X1 U2658 ( .A1(n14055), .A2(n10908), .B1(n14087), .B2(n10905), .C1(
        n14023), .C2(n10902), .ZN(n5220) );
  OAI222_X1 U2659 ( .A1(n14055), .A2(n11172), .B1(n14087), .B2(n11169), .C1(
        n14023), .C2(n11166), .ZN(n3787) );
  OAI222_X1 U2660 ( .A1(n14054), .A2(n10909), .B1(n14086), .B2(n10906), .C1(
        n14022), .C2(n10903), .ZN(n5179) );
  OAI222_X1 U2661 ( .A1(n14054), .A2(n11173), .B1(n14086), .B2(n11170), .C1(
        n14022), .C2(n11167), .ZN(n3746) );
  OAI222_X1 U2662 ( .A1(n14053), .A2(n10909), .B1(n14085), .B2(n10906), .C1(
        n14021), .C2(n10903), .ZN(n5138) );
  OAI222_X1 U2663 ( .A1(n14053), .A2(n11173), .B1(n14085), .B2(n11170), .C1(
        n14021), .C2(n11167), .ZN(n3705) );
  OAI222_X1 U2664 ( .A1(n14052), .A2(n10909), .B1(n14084), .B2(n10906), .C1(
        n14020), .C2(n10903), .ZN(n5097) );
  OAI222_X1 U2665 ( .A1(n14052), .A2(n11173), .B1(n14084), .B2(n11170), .C1(
        n14020), .C2(n11167), .ZN(n3664) );
  OAI222_X1 U2666 ( .A1(n14051), .A2(n10909), .B1(n14083), .B2(n10906), .C1(
        n14019), .C2(n10903), .ZN(n5056) );
  OAI222_X1 U2667 ( .A1(n14051), .A2(n11173), .B1(n14083), .B2(n11170), .C1(
        n14019), .C2(n11167), .ZN(n3623) );
  OAI222_X1 U2668 ( .A1(n14050), .A2(n10909), .B1(n14082), .B2(n10906), .C1(
        n14018), .C2(n10903), .ZN(n5015) );
  OAI222_X1 U2669 ( .A1(n14050), .A2(n11173), .B1(n14082), .B2(n11170), .C1(
        n14018), .C2(n11167), .ZN(n3582) );
  OAI222_X1 U2670 ( .A1(n14049), .A2(n10909), .B1(n14081), .B2(n10906), .C1(
        n14017), .C2(n10903), .ZN(n4974) );
  OAI222_X1 U2671 ( .A1(n14049), .A2(n11173), .B1(n14081), .B2(n11170), .C1(
        n14017), .C2(n11167), .ZN(n3541) );
  OAI222_X1 U2672 ( .A1(n14048), .A2(n10909), .B1(n14080), .B2(n10906), .C1(
        n14016), .C2(n10903), .ZN(n4933) );
  OAI222_X1 U2673 ( .A1(n14048), .A2(n11173), .B1(n14080), .B2(n11170), .C1(
        n14016), .C2(n11167), .ZN(n3500) );
  OAI222_X1 U2674 ( .A1(n14047), .A2(n10909), .B1(n14079), .B2(n10906), .C1(
        n14015), .C2(n10903), .ZN(n4892) );
  OAI222_X1 U2675 ( .A1(n14047), .A2(n11173), .B1(n14079), .B2(n11170), .C1(
        n14015), .C2(n11167), .ZN(n3459) );
  OAI222_X1 U2676 ( .A1(n14046), .A2(n10909), .B1(n14078), .B2(n10906), .C1(
        n14014), .C2(n10903), .ZN(n4851) );
  OAI222_X1 U2677 ( .A1(n14046), .A2(n11173), .B1(n14078), .B2(n11170), .C1(
        n14014), .C2(n11167), .ZN(n3418) );
  OAI222_X1 U2678 ( .A1(n14045), .A2(n10909), .B1(n14077), .B2(n10906), .C1(
        n14013), .C2(n10903), .ZN(n4810) );
  OAI222_X1 U2679 ( .A1(n14045), .A2(n11173), .B1(n14077), .B2(n11170), .C1(
        n14013), .C2(n11167), .ZN(n3377) );
  OAI222_X1 U2680 ( .A1(n14044), .A2(n10909), .B1(n14076), .B2(n10906), .C1(
        n14012), .C2(n10903), .ZN(n4769) );
  OAI222_X1 U2681 ( .A1(n14044), .A2(n11173), .B1(n14076), .B2(n11170), .C1(
        n14012), .C2(n11167), .ZN(n3336) );
  OAI222_X1 U2682 ( .A1(n14043), .A2(n10909), .B1(n14075), .B2(n10906), .C1(
        n14011), .C2(n10903), .ZN(n4728) );
  OAI222_X1 U2683 ( .A1(n14043), .A2(n11173), .B1(n14075), .B2(n11170), .C1(
        n14011), .C2(n11167), .ZN(n3295) );
  OAI222_X1 U2684 ( .A1(n13147), .A2(n11009), .B1(n13179), .B2(n11006), .C1(
        n13115), .C2(n11003), .ZN(n4671) );
  OAI222_X1 U2685 ( .A1(n13147), .A2(n11273), .B1(n13179), .B2(n11270), .C1(
        n13115), .C2(n11267), .ZN(n3238) );
  OAI222_X1 U2686 ( .A1(n13146), .A2(n11009), .B1(n13178), .B2(n11006), .C1(
        n13114), .C2(n11003), .ZN(n4630) );
  OAI222_X1 U2687 ( .A1(n13146), .A2(n11273), .B1(n13178), .B2(n11270), .C1(
        n13114), .C2(n11267), .ZN(n3197) );
  OAI222_X1 U2688 ( .A1(n13145), .A2(n11009), .B1(n13177), .B2(n11006), .C1(
        n13113), .C2(n11003), .ZN(n4589) );
  OAI222_X1 U2689 ( .A1(n13145), .A2(n11273), .B1(n13177), .B2(n11270), .C1(
        n13113), .C2(n11267), .ZN(n3156) );
  OAI222_X1 U2690 ( .A1(n13144), .A2(n11009), .B1(n13176), .B2(n11006), .C1(
        n13112), .C2(n11003), .ZN(n4548) );
  OAI222_X1 U2691 ( .A1(n13144), .A2(n11273), .B1(n13176), .B2(n11270), .C1(
        n13112), .C2(n11267), .ZN(n3115) );
  OAI222_X1 U2692 ( .A1(n13143), .A2(n11009), .B1(n13175), .B2(n11006), .C1(
        n13111), .C2(n11003), .ZN(n4507) );
  OAI222_X1 U2693 ( .A1(n13143), .A2(n11273), .B1(n13175), .B2(n11270), .C1(
        n13111), .C2(n11267), .ZN(n3074) );
  OAI222_X1 U2694 ( .A1(n13142), .A2(n11009), .B1(n13174), .B2(n11006), .C1(
        n13110), .C2(n11003), .ZN(n4466) );
  OAI222_X1 U2695 ( .A1(n13142), .A2(n11273), .B1(n13174), .B2(n11270), .C1(
        n13110), .C2(n11267), .ZN(n3033) );
  OAI222_X1 U2696 ( .A1(n13141), .A2(n11009), .B1(n13173), .B2(n11006), .C1(
        n13109), .C2(n11003), .ZN(n4425) );
  OAI222_X1 U2697 ( .A1(n13141), .A2(n11273), .B1(n13173), .B2(n11270), .C1(
        n13109), .C2(n11267), .ZN(n2992) );
  OAI222_X1 U2698 ( .A1(n13140), .A2(n11009), .B1(n13172), .B2(n11006), .C1(
        n13108), .C2(n11003), .ZN(n4331) );
  OAI222_X1 U2699 ( .A1(n13140), .A2(n11273), .B1(n13172), .B2(n11270), .C1(
        n13108), .C2(n11267), .ZN(n2863) );
  OAI222_X1 U2700 ( .A1(n13171), .A2(n11007), .B1(n13203), .B2(n11004), .C1(
        n13139), .C2(n11001), .ZN(n5677) );
  OAI222_X1 U2701 ( .A1(n13171), .A2(n11271), .B1(n13203), .B2(n11268), .C1(
        n13139), .C2(n11265), .ZN(n4244) );
  OAI222_X1 U2702 ( .A1(n13170), .A2(n11007), .B1(n13202), .B2(n11004), .C1(
        n13138), .C2(n11001), .ZN(n5614) );
  OAI222_X1 U2703 ( .A1(n13170), .A2(n11271), .B1(n13202), .B2(n11268), .C1(
        n13138), .C2(n11265), .ZN(n4181) );
  OAI222_X1 U2704 ( .A1(n13169), .A2(n11007), .B1(n13201), .B2(n11004), .C1(
        n13137), .C2(n11001), .ZN(n5573) );
  OAI222_X1 U2705 ( .A1(n13169), .A2(n11271), .B1(n13201), .B2(n11268), .C1(
        n13137), .C2(n11265), .ZN(n4140) );
  OAI222_X1 U2706 ( .A1(n13168), .A2(n11007), .B1(n13200), .B2(n11004), .C1(
        n13136), .C2(n11001), .ZN(n5532) );
  OAI222_X1 U2707 ( .A1(n13168), .A2(n11271), .B1(n13200), .B2(n11268), .C1(
        n13136), .C2(n11265), .ZN(n4099) );
  OAI222_X1 U2708 ( .A1(n13167), .A2(n11007), .B1(n13199), .B2(n11004), .C1(
        n13135), .C2(n11001), .ZN(n5491) );
  OAI222_X1 U2709 ( .A1(n13167), .A2(n11271), .B1(n13199), .B2(n11268), .C1(
        n13135), .C2(n11265), .ZN(n4058) );
  OAI222_X1 U2710 ( .A1(n13166), .A2(n11007), .B1(n13198), .B2(n11004), .C1(
        n13134), .C2(n11001), .ZN(n5450) );
  OAI222_X1 U2711 ( .A1(n13166), .A2(n11271), .B1(n13198), .B2(n11268), .C1(
        n13134), .C2(n11265), .ZN(n4017) );
  OAI222_X1 U2712 ( .A1(n13165), .A2(n11007), .B1(n13197), .B2(n11004), .C1(
        n13133), .C2(n11001), .ZN(n5409) );
  OAI222_X1 U2713 ( .A1(n13165), .A2(n11271), .B1(n13197), .B2(n11268), .C1(
        n13133), .C2(n11265), .ZN(n3976) );
  OAI222_X1 U2714 ( .A1(n13164), .A2(n11007), .B1(n13196), .B2(n11004), .C1(
        n13132), .C2(n11001), .ZN(n5368) );
  OAI222_X1 U2715 ( .A1(n13164), .A2(n11271), .B1(n13196), .B2(n11268), .C1(
        n13132), .C2(n11265), .ZN(n3935) );
  OAI222_X1 U2716 ( .A1(n13163), .A2(n11007), .B1(n13195), .B2(n11004), .C1(
        n13131), .C2(n11001), .ZN(n5327) );
  OAI222_X1 U2717 ( .A1(n13163), .A2(n11271), .B1(n13195), .B2(n11268), .C1(
        n13131), .C2(n11265), .ZN(n3894) );
  OAI222_X1 U2718 ( .A1(n13162), .A2(n11007), .B1(n13194), .B2(n11004), .C1(
        n13130), .C2(n11001), .ZN(n5286) );
  OAI222_X1 U2719 ( .A1(n13162), .A2(n11271), .B1(n13194), .B2(n11268), .C1(
        n13130), .C2(n11265), .ZN(n3853) );
  OAI222_X1 U2720 ( .A1(n13161), .A2(n11007), .B1(n13193), .B2(n11004), .C1(
        n13129), .C2(n11001), .ZN(n5245) );
  OAI222_X1 U2721 ( .A1(n13161), .A2(n11271), .B1(n13193), .B2(n11268), .C1(
        n13129), .C2(n11265), .ZN(n3812) );
  OAI222_X1 U2722 ( .A1(n13160), .A2(n11007), .B1(n13192), .B2(n11004), .C1(
        n13128), .C2(n11001), .ZN(n5204) );
  OAI222_X1 U2723 ( .A1(n13160), .A2(n11271), .B1(n13192), .B2(n11268), .C1(
        n13128), .C2(n11265), .ZN(n3771) );
  OAI222_X1 U2724 ( .A1(n13159), .A2(n11008), .B1(n13191), .B2(n11005), .C1(
        n13127), .C2(n11002), .ZN(n5163) );
  OAI222_X1 U2725 ( .A1(n13159), .A2(n11272), .B1(n13191), .B2(n11269), .C1(
        n13127), .C2(n11266), .ZN(n3730) );
  OAI222_X1 U2726 ( .A1(n13158), .A2(n11008), .B1(n13190), .B2(n11005), .C1(
        n13126), .C2(n11002), .ZN(n5122) );
  OAI222_X1 U2727 ( .A1(n13158), .A2(n11272), .B1(n13190), .B2(n11269), .C1(
        n13126), .C2(n11266), .ZN(n3689) );
  OAI222_X1 U2728 ( .A1(n13157), .A2(n11008), .B1(n13189), .B2(n11005), .C1(
        n13125), .C2(n11002), .ZN(n5081) );
  OAI222_X1 U2729 ( .A1(n13157), .A2(n11272), .B1(n13189), .B2(n11269), .C1(
        n13125), .C2(n11266), .ZN(n3648) );
  OAI222_X1 U2730 ( .A1(n13156), .A2(n11008), .B1(n13188), .B2(n11005), .C1(
        n13124), .C2(n11002), .ZN(n5040) );
  OAI222_X1 U2731 ( .A1(n13156), .A2(n11272), .B1(n13188), .B2(n11269), .C1(
        n13124), .C2(n11266), .ZN(n3607) );
  OAI222_X1 U2732 ( .A1(n13155), .A2(n11008), .B1(n13187), .B2(n11005), .C1(
        n13123), .C2(n11002), .ZN(n4999) );
  OAI222_X1 U2733 ( .A1(n13155), .A2(n11272), .B1(n13187), .B2(n11269), .C1(
        n13123), .C2(n11266), .ZN(n3566) );
  OAI222_X1 U2734 ( .A1(n13154), .A2(n11008), .B1(n13186), .B2(n11005), .C1(
        n13122), .C2(n11002), .ZN(n4958) );
  OAI222_X1 U2735 ( .A1(n13154), .A2(n11272), .B1(n13186), .B2(n11269), .C1(
        n13122), .C2(n11266), .ZN(n3525) );
  OAI222_X1 U2736 ( .A1(n13153), .A2(n11008), .B1(n13185), .B2(n11005), .C1(
        n13121), .C2(n11002), .ZN(n4917) );
  OAI222_X1 U2737 ( .A1(n13153), .A2(n11272), .B1(n13185), .B2(n11269), .C1(
        n13121), .C2(n11266), .ZN(n3484) );
  OAI222_X1 U2738 ( .A1(n13152), .A2(n11008), .B1(n13184), .B2(n11005), .C1(
        n13120), .C2(n11002), .ZN(n4876) );
  OAI222_X1 U2739 ( .A1(n13152), .A2(n11272), .B1(n13184), .B2(n11269), .C1(
        n13120), .C2(n11266), .ZN(n3443) );
  OAI222_X1 U2740 ( .A1(n13151), .A2(n11008), .B1(n13183), .B2(n11005), .C1(
        n13119), .C2(n11002), .ZN(n4835) );
  OAI222_X1 U2741 ( .A1(n13151), .A2(n11272), .B1(n13183), .B2(n11269), .C1(
        n13119), .C2(n11266), .ZN(n3402) );
  OAI222_X1 U2742 ( .A1(n13150), .A2(n11008), .B1(n13182), .B2(n11005), .C1(
        n13118), .C2(n11002), .ZN(n4794) );
  OAI222_X1 U2743 ( .A1(n13150), .A2(n11272), .B1(n13182), .B2(n11269), .C1(
        n13118), .C2(n11266), .ZN(n3361) );
  OAI222_X1 U2744 ( .A1(n13149), .A2(n11008), .B1(n13181), .B2(n11005), .C1(
        n13117), .C2(n11002), .ZN(n4753) );
  OAI222_X1 U2745 ( .A1(n13149), .A2(n11272), .B1(n13181), .B2(n11269), .C1(
        n13117), .C2(n11266), .ZN(n3320) );
  OAI222_X1 U2746 ( .A1(n13148), .A2(n11008), .B1(n13180), .B2(n11005), .C1(
        n13116), .C2(n11002), .ZN(n4712) );
  OAI222_X1 U2747 ( .A1(n13148), .A2(n11272), .B1(n13180), .B2(n11269), .C1(
        n13116), .C2(n11266), .ZN(n3279) );
  OAI222_X1 U2748 ( .A1(n13467), .A2(n11024), .B1(n13403), .B2(n11021), .C1(
        n13435), .C2(n11018), .ZN(n4667) );
  OAI222_X1 U2749 ( .A1(n13467), .A2(n11288), .B1(n13403), .B2(n11285), .C1(
        n13435), .C2(n11282), .ZN(n3234) );
  OAI222_X1 U2750 ( .A1(n13466), .A2(n11024), .B1(n13402), .B2(n11021), .C1(
        n13434), .C2(n11018), .ZN(n4626) );
  OAI222_X1 U2751 ( .A1(n13466), .A2(n11288), .B1(n13402), .B2(n11285), .C1(
        n13434), .C2(n11282), .ZN(n3193) );
  OAI222_X1 U2752 ( .A1(n13465), .A2(n11024), .B1(n13401), .B2(n11021), .C1(
        n13433), .C2(n11018), .ZN(n4585) );
  OAI222_X1 U2753 ( .A1(n13465), .A2(n11288), .B1(n13401), .B2(n11285), .C1(
        n13433), .C2(n11282), .ZN(n3152) );
  OAI222_X1 U2754 ( .A1(n13464), .A2(n11024), .B1(n13400), .B2(n11021), .C1(
        n13432), .C2(n11018), .ZN(n4544) );
  OAI222_X1 U2755 ( .A1(n13464), .A2(n11288), .B1(n13400), .B2(n11285), .C1(
        n13432), .C2(n11282), .ZN(n3111) );
  OAI222_X1 U2756 ( .A1(n13463), .A2(n11024), .B1(n13399), .B2(n11021), .C1(
        n13431), .C2(n11018), .ZN(n4503) );
  OAI222_X1 U2757 ( .A1(n13463), .A2(n11288), .B1(n13399), .B2(n11285), .C1(
        n13431), .C2(n11282), .ZN(n3070) );
  OAI222_X1 U2758 ( .A1(n13462), .A2(n11024), .B1(n13398), .B2(n11021), .C1(
        n13430), .C2(n11018), .ZN(n4462) );
  OAI222_X1 U2759 ( .A1(n13462), .A2(n11288), .B1(n13398), .B2(n11285), .C1(
        n13430), .C2(n11282), .ZN(n3029) );
  OAI222_X1 U2760 ( .A1(n13461), .A2(n11024), .B1(n13397), .B2(n11021), .C1(
        n13429), .C2(n11018), .ZN(n4421) );
  OAI222_X1 U2761 ( .A1(n13461), .A2(n11288), .B1(n13397), .B2(n11285), .C1(
        n13429), .C2(n11282), .ZN(n2988) );
  OAI222_X1 U2762 ( .A1(n13460), .A2(n11024), .B1(n13396), .B2(n11021), .C1(
        n13428), .C2(n11018), .ZN(n4314) );
  OAI222_X1 U2763 ( .A1(n13460), .A2(n11288), .B1(n13396), .B2(n11285), .C1(
        n13428), .C2(n11282), .ZN(n2814) );
  OAI222_X1 U2764 ( .A1(n13491), .A2(n11022), .B1(n13427), .B2(n11019), .C1(
        n13459), .C2(n11016), .ZN(n5670) );
  OAI222_X1 U2765 ( .A1(n13491), .A2(n11286), .B1(n13427), .B2(n11283), .C1(
        n13459), .C2(n11280), .ZN(n4237) );
  OAI222_X1 U2766 ( .A1(n13490), .A2(n11022), .B1(n13426), .B2(n11019), .C1(
        n13458), .C2(n11016), .ZN(n5610) );
  OAI222_X1 U2767 ( .A1(n13490), .A2(n11286), .B1(n13426), .B2(n11283), .C1(
        n13458), .C2(n11280), .ZN(n4177) );
  OAI222_X1 U2768 ( .A1(n13489), .A2(n11022), .B1(n13425), .B2(n11019), .C1(
        n13457), .C2(n11016), .ZN(n5569) );
  OAI222_X1 U2769 ( .A1(n13489), .A2(n11286), .B1(n13425), .B2(n11283), .C1(
        n13457), .C2(n11280), .ZN(n4136) );
  OAI222_X1 U2770 ( .A1(n13488), .A2(n11022), .B1(n13424), .B2(n11019), .C1(
        n13456), .C2(n11016), .ZN(n5528) );
  OAI222_X1 U2771 ( .A1(n13488), .A2(n11286), .B1(n13424), .B2(n11283), .C1(
        n13456), .C2(n11280), .ZN(n4095) );
  OAI222_X1 U2772 ( .A1(n13487), .A2(n11022), .B1(n13423), .B2(n11019), .C1(
        n13455), .C2(n11016), .ZN(n5487) );
  OAI222_X1 U2773 ( .A1(n13487), .A2(n11286), .B1(n13423), .B2(n11283), .C1(
        n13455), .C2(n11280), .ZN(n4054) );
  OAI222_X1 U2774 ( .A1(n13486), .A2(n11022), .B1(n13422), .B2(n11019), .C1(
        n13454), .C2(n11016), .ZN(n5446) );
  OAI222_X1 U2775 ( .A1(n13486), .A2(n11286), .B1(n13422), .B2(n11283), .C1(
        n13454), .C2(n11280), .ZN(n4013) );
  OAI222_X1 U2776 ( .A1(n13485), .A2(n11022), .B1(n13421), .B2(n11019), .C1(
        n13453), .C2(n11016), .ZN(n5405) );
  OAI222_X1 U2777 ( .A1(n13485), .A2(n11286), .B1(n13421), .B2(n11283), .C1(
        n13453), .C2(n11280), .ZN(n3972) );
  OAI222_X1 U2778 ( .A1(n13484), .A2(n11022), .B1(n13420), .B2(n11019), .C1(
        n13452), .C2(n11016), .ZN(n5364) );
  OAI222_X1 U2779 ( .A1(n13484), .A2(n11286), .B1(n13420), .B2(n11283), .C1(
        n13452), .C2(n11280), .ZN(n3931) );
  OAI222_X1 U2780 ( .A1(n13483), .A2(n11022), .B1(n13419), .B2(n11019), .C1(
        n13451), .C2(n11016), .ZN(n5323) );
  OAI222_X1 U2781 ( .A1(n13483), .A2(n11286), .B1(n13419), .B2(n11283), .C1(
        n13451), .C2(n11280), .ZN(n3890) );
  OAI222_X1 U2782 ( .A1(n13482), .A2(n11022), .B1(n13418), .B2(n11019), .C1(
        n13450), .C2(n11016), .ZN(n5282) );
  OAI222_X1 U2783 ( .A1(n13482), .A2(n11286), .B1(n13418), .B2(n11283), .C1(
        n13450), .C2(n11280), .ZN(n3849) );
  OAI222_X1 U2784 ( .A1(n13481), .A2(n11022), .B1(n13417), .B2(n11019), .C1(
        n13449), .C2(n11016), .ZN(n5241) );
  OAI222_X1 U2785 ( .A1(n13481), .A2(n11286), .B1(n13417), .B2(n11283), .C1(
        n13449), .C2(n11280), .ZN(n3808) );
  OAI222_X1 U2786 ( .A1(n13480), .A2(n11022), .B1(n13416), .B2(n11019), .C1(
        n13448), .C2(n11016), .ZN(n5200) );
  OAI222_X1 U2787 ( .A1(n13480), .A2(n11286), .B1(n13416), .B2(n11283), .C1(
        n13448), .C2(n11280), .ZN(n3767) );
  OAI222_X1 U2788 ( .A1(n13479), .A2(n11023), .B1(n13415), .B2(n11020), .C1(
        n13447), .C2(n11017), .ZN(n5159) );
  OAI222_X1 U2789 ( .A1(n13479), .A2(n11287), .B1(n13415), .B2(n11284), .C1(
        n13447), .C2(n11281), .ZN(n3726) );
  OAI222_X1 U2790 ( .A1(n13478), .A2(n11023), .B1(n13414), .B2(n11020), .C1(
        n13446), .C2(n11017), .ZN(n5118) );
  OAI222_X1 U2791 ( .A1(n13478), .A2(n11287), .B1(n13414), .B2(n11284), .C1(
        n13446), .C2(n11281), .ZN(n3685) );
  OAI222_X1 U2792 ( .A1(n13477), .A2(n11023), .B1(n13413), .B2(n11020), .C1(
        n13445), .C2(n11017), .ZN(n5077) );
  OAI222_X1 U2793 ( .A1(n13477), .A2(n11287), .B1(n13413), .B2(n11284), .C1(
        n13445), .C2(n11281), .ZN(n3644) );
  OAI222_X1 U2794 ( .A1(n13476), .A2(n11023), .B1(n13412), .B2(n11020), .C1(
        n13444), .C2(n11017), .ZN(n5036) );
  OAI222_X1 U2795 ( .A1(n13476), .A2(n11287), .B1(n13412), .B2(n11284), .C1(
        n13444), .C2(n11281), .ZN(n3603) );
  OAI222_X1 U2796 ( .A1(n13475), .A2(n11023), .B1(n13411), .B2(n11020), .C1(
        n13443), .C2(n11017), .ZN(n4995) );
  OAI222_X1 U2797 ( .A1(n13475), .A2(n11287), .B1(n13411), .B2(n11284), .C1(
        n13443), .C2(n11281), .ZN(n3562) );
  OAI222_X1 U2798 ( .A1(n13474), .A2(n11023), .B1(n13410), .B2(n11020), .C1(
        n13442), .C2(n11017), .ZN(n4954) );
  OAI222_X1 U2799 ( .A1(n13474), .A2(n11287), .B1(n13410), .B2(n11284), .C1(
        n13442), .C2(n11281), .ZN(n3521) );
  OAI222_X1 U2800 ( .A1(n13473), .A2(n11023), .B1(n13409), .B2(n11020), .C1(
        n13441), .C2(n11017), .ZN(n4913) );
  OAI222_X1 U2801 ( .A1(n13473), .A2(n11287), .B1(n13409), .B2(n11284), .C1(
        n13441), .C2(n11281), .ZN(n3480) );
  OAI222_X1 U2802 ( .A1(n13472), .A2(n11023), .B1(n13408), .B2(n11020), .C1(
        n13440), .C2(n11017), .ZN(n4872) );
  OAI222_X1 U2803 ( .A1(n13472), .A2(n11287), .B1(n13408), .B2(n11284), .C1(
        n13440), .C2(n11281), .ZN(n3439) );
  OAI222_X1 U2804 ( .A1(n13471), .A2(n11023), .B1(n13407), .B2(n11020), .C1(
        n13439), .C2(n11017), .ZN(n4831) );
  OAI222_X1 U2805 ( .A1(n13471), .A2(n11287), .B1(n13407), .B2(n11284), .C1(
        n13439), .C2(n11281), .ZN(n3398) );
  OAI222_X1 U2806 ( .A1(n13470), .A2(n11023), .B1(n13406), .B2(n11020), .C1(
        n13438), .C2(n11017), .ZN(n4790) );
  OAI222_X1 U2807 ( .A1(n13470), .A2(n11287), .B1(n13406), .B2(n11284), .C1(
        n13438), .C2(n11281), .ZN(n3357) );
  OAI222_X1 U2808 ( .A1(n13469), .A2(n11023), .B1(n13405), .B2(n11020), .C1(
        n13437), .C2(n11017), .ZN(n4749) );
  OAI222_X1 U2809 ( .A1(n13469), .A2(n11287), .B1(n13405), .B2(n11284), .C1(
        n13437), .C2(n11281), .ZN(n3316) );
  OAI222_X1 U2810 ( .A1(n13468), .A2(n11023), .B1(n13404), .B2(n11020), .C1(
        n13436), .C2(n11017), .ZN(n4708) );
  OAI222_X1 U2811 ( .A1(n13468), .A2(n11287), .B1(n13404), .B2(n11284), .C1(
        n13436), .C2(n11281), .ZN(n3275) );
  AOI222_X1 U2812 ( .A1(n10857), .A2(n14320), .B1(n10854), .B2(n14352), .C1(
        n10851), .C2(n14416), .ZN(n5693) );
  AOI222_X1 U2813 ( .A1(n11121), .A2(n14320), .B1(n11118), .B2(n14352), .C1(
        n11115), .C2(n14416), .ZN(n4260) );
  AOI222_X1 U2814 ( .A1(n10857), .A2(n14319), .B1(n10854), .B2(n14351), .C1(
        n10851), .C2(n14415), .ZN(n5624) );
  AOI222_X1 U2815 ( .A1(n11121), .A2(n14319), .B1(n11118), .B2(n14351), .C1(
        n11115), .C2(n14415), .ZN(n4191) );
  AOI222_X1 U2816 ( .A1(n10857), .A2(n14318), .B1(n10854), .B2(n14350), .C1(
        n10851), .C2(n14414), .ZN(n5583) );
  AOI222_X1 U2817 ( .A1(n11121), .A2(n14318), .B1(n11118), .B2(n14350), .C1(
        n11115), .C2(n14414), .ZN(n4150) );
  AOI222_X1 U2818 ( .A1(n10857), .A2(n14317), .B1(n10854), .B2(n14349), .C1(
        n10851), .C2(n14413), .ZN(n5542) );
  AOI222_X1 U2819 ( .A1(n11121), .A2(n14317), .B1(n11118), .B2(n14349), .C1(
        n11115), .C2(n14413), .ZN(n4109) );
  AOI222_X1 U2820 ( .A1(n10857), .A2(n14316), .B1(n10854), .B2(n14348), .C1(
        n10851), .C2(n14412), .ZN(n5501) );
  AOI222_X1 U2821 ( .A1(n11121), .A2(n14316), .B1(n11118), .B2(n14348), .C1(
        n11115), .C2(n14412), .ZN(n4068) );
  AOI222_X1 U2822 ( .A1(n10857), .A2(n14315), .B1(n10854), .B2(n14347), .C1(
        n10851), .C2(n14411), .ZN(n5460) );
  AOI222_X1 U2823 ( .A1(n11121), .A2(n14315), .B1(n11118), .B2(n14347), .C1(
        n11115), .C2(n14411), .ZN(n4027) );
  AOI222_X1 U2824 ( .A1(n10857), .A2(n14314), .B1(n10854), .B2(n14346), .C1(
        n10851), .C2(n14410), .ZN(n5419) );
  AOI222_X1 U2825 ( .A1(n11121), .A2(n14314), .B1(n11118), .B2(n14346), .C1(
        n11115), .C2(n14410), .ZN(n3986) );
  AOI222_X1 U2826 ( .A1(n10857), .A2(n14313), .B1(n10854), .B2(n14345), .C1(
        n10851), .C2(n14409), .ZN(n5378) );
  AOI222_X1 U2827 ( .A1(n11121), .A2(n14313), .B1(n11118), .B2(n14345), .C1(
        n11115), .C2(n14409), .ZN(n3945) );
  AOI222_X1 U2828 ( .A1(n10857), .A2(n14312), .B1(n10854), .B2(n14344), .C1(
        n10851), .C2(n14408), .ZN(n5337) );
  AOI222_X1 U2829 ( .A1(n11121), .A2(n14312), .B1(n11118), .B2(n14344), .C1(
        n11115), .C2(n14408), .ZN(n3904) );
  AOI222_X1 U2830 ( .A1(n10857), .A2(n14311), .B1(n10854), .B2(n14343), .C1(
        n10851), .C2(n14407), .ZN(n5296) );
  AOI222_X1 U2831 ( .A1(n11121), .A2(n14311), .B1(n11118), .B2(n14343), .C1(
        n11115), .C2(n14407), .ZN(n3863) );
  AOI222_X1 U2832 ( .A1(n10857), .A2(n14310), .B1(n10854), .B2(n14342), .C1(
        n10851), .C2(n14406), .ZN(n5255) );
  AOI222_X1 U2833 ( .A1(n11121), .A2(n14310), .B1(n11118), .B2(n14342), .C1(
        n11115), .C2(n14406), .ZN(n3822) );
  AOI222_X1 U2834 ( .A1(n10857), .A2(n14309), .B1(n10854), .B2(n14341), .C1(
        n10851), .C2(n14405), .ZN(n5214) );
  AOI222_X1 U2835 ( .A1(n11121), .A2(n14309), .B1(n11118), .B2(n14341), .C1(
        n11115), .C2(n14405), .ZN(n3781) );
  AOI222_X1 U2836 ( .A1(n10858), .A2(n14308), .B1(n10855), .B2(n14340), .C1(
        n10852), .C2(n14404), .ZN(n5173) );
  AOI222_X1 U2837 ( .A1(n11122), .A2(n14308), .B1(n11119), .B2(n14340), .C1(
        n11116), .C2(n14404), .ZN(n3740) );
  AOI222_X1 U2838 ( .A1(n10858), .A2(n14307), .B1(n10855), .B2(n14339), .C1(
        n10852), .C2(n14403), .ZN(n5132) );
  AOI222_X1 U2839 ( .A1(n11122), .A2(n14307), .B1(n11119), .B2(n14339), .C1(
        n11116), .C2(n14403), .ZN(n3699) );
  AOI222_X1 U2840 ( .A1(n10858), .A2(n14306), .B1(n10855), .B2(n14338), .C1(
        n10852), .C2(n14402), .ZN(n5091) );
  AOI222_X1 U2841 ( .A1(n11122), .A2(n14306), .B1(n11119), .B2(n14338), .C1(
        n11116), .C2(n14402), .ZN(n3658) );
  AOI222_X1 U2842 ( .A1(n10858), .A2(n14305), .B1(n10855), .B2(n14337), .C1(
        n10852), .C2(n14401), .ZN(n5050) );
  AOI222_X1 U2843 ( .A1(n11122), .A2(n14305), .B1(n11119), .B2(n14337), .C1(
        n11116), .C2(n14401), .ZN(n3617) );
  AOI222_X1 U2844 ( .A1(n10858), .A2(n14304), .B1(n10855), .B2(n14336), .C1(
        n10852), .C2(n14400), .ZN(n5009) );
  AOI222_X1 U2845 ( .A1(n11122), .A2(n14304), .B1(n11119), .B2(n14336), .C1(
        n11116), .C2(n14400), .ZN(n3576) );
  AOI222_X1 U2846 ( .A1(n10858), .A2(n14303), .B1(n10855), .B2(n14335), .C1(
        n10852), .C2(n14399), .ZN(n4968) );
  AOI222_X1 U2847 ( .A1(n11122), .A2(n14303), .B1(n11119), .B2(n14335), .C1(
        n11116), .C2(n14399), .ZN(n3535) );
  AOI222_X1 U2848 ( .A1(n10858), .A2(n14302), .B1(n10855), .B2(n14334), .C1(
        n10852), .C2(n14398), .ZN(n4927) );
  AOI222_X1 U2849 ( .A1(n11122), .A2(n14302), .B1(n11119), .B2(n14334), .C1(
        n11116), .C2(n14398), .ZN(n3494) );
  AOI222_X1 U2850 ( .A1(n10858), .A2(n14301), .B1(n10855), .B2(n14333), .C1(
        n10852), .C2(n14397), .ZN(n4886) );
  AOI222_X1 U2851 ( .A1(n11122), .A2(n14301), .B1(n11119), .B2(n14333), .C1(
        n11116), .C2(n14397), .ZN(n3453) );
  AOI222_X1 U2852 ( .A1(n10858), .A2(n14300), .B1(n10855), .B2(n14332), .C1(
        n10852), .C2(n14396), .ZN(n4845) );
  AOI222_X1 U2853 ( .A1(n11122), .A2(n14300), .B1(n11119), .B2(n14332), .C1(
        n11116), .C2(n14396), .ZN(n3412) );
  AOI222_X1 U2854 ( .A1(n10858), .A2(n14299), .B1(n10855), .B2(n14331), .C1(
        n10852), .C2(n14395), .ZN(n4804) );
  AOI222_X1 U2855 ( .A1(n11122), .A2(n14299), .B1(n11119), .B2(n14331), .C1(
        n11116), .C2(n14395), .ZN(n3371) );
  AOI222_X1 U2856 ( .A1(n10858), .A2(n14298), .B1(n10855), .B2(n14330), .C1(
        n10852), .C2(n14394), .ZN(n4763) );
  AOI222_X1 U2857 ( .A1(n11122), .A2(n14298), .B1(n11119), .B2(n14330), .C1(
        n11116), .C2(n14394), .ZN(n3330) );
  AOI222_X1 U2858 ( .A1(n10858), .A2(n14297), .B1(n10855), .B2(n14329), .C1(
        n10852), .C2(n14393), .ZN(n4722) );
  AOI222_X1 U2859 ( .A1(n11122), .A2(n14297), .B1(n11119), .B2(n14329), .C1(
        n11116), .C2(n14393), .ZN(n3289) );
  AOI222_X1 U2860 ( .A1(n10859), .A2(n14296), .B1(n10856), .B2(n14328), .C1(
        n10853), .C2(n14392), .ZN(n4681) );
  AOI222_X1 U2861 ( .A1(n11123), .A2(n14296), .B1(n11120), .B2(n14328), .C1(
        n11117), .C2(n14392), .ZN(n3248) );
  AOI222_X1 U2862 ( .A1(n10859), .A2(n14295), .B1(n10856), .B2(n14327), .C1(
        n10853), .C2(n14391), .ZN(n4640) );
  AOI222_X1 U2863 ( .A1(n11123), .A2(n14295), .B1(n11120), .B2(n14327), .C1(
        n11117), .C2(n14391), .ZN(n3207) );
  AOI222_X1 U2864 ( .A1(n10859), .A2(n14294), .B1(n10856), .B2(n14326), .C1(
        n10853), .C2(n14390), .ZN(n4599) );
  AOI222_X1 U2865 ( .A1(n11123), .A2(n14294), .B1(n11120), .B2(n14326), .C1(
        n11117), .C2(n14390), .ZN(n3166) );
  AOI222_X1 U2866 ( .A1(n10859), .A2(n14293), .B1(n10856), .B2(n14325), .C1(
        n10853), .C2(n14389), .ZN(n4558) );
  AOI222_X1 U2867 ( .A1(n11123), .A2(n14293), .B1(n11120), .B2(n14325), .C1(
        n11117), .C2(n14389), .ZN(n3125) );
  AOI222_X1 U2868 ( .A1(n10859), .A2(n14292), .B1(n10856), .B2(n14324), .C1(
        n10853), .C2(n14388), .ZN(n4517) );
  AOI222_X1 U2869 ( .A1(n11123), .A2(n14292), .B1(n11120), .B2(n14324), .C1(
        n11117), .C2(n14388), .ZN(n3084) );
  AOI222_X1 U2870 ( .A1(n10859), .A2(n14291), .B1(n10856), .B2(n14323), .C1(
        n10853), .C2(n14387), .ZN(n4476) );
  AOI222_X1 U2871 ( .A1(n11123), .A2(n14291), .B1(n11120), .B2(n14323), .C1(
        n11117), .C2(n14387), .ZN(n3043) );
  AOI222_X1 U2872 ( .A1(n10859), .A2(n14290), .B1(n10856), .B2(n14322), .C1(
        n10853), .C2(n14386), .ZN(n4435) );
  AOI222_X1 U2873 ( .A1(n11123), .A2(n14290), .B1(n11120), .B2(n14322), .C1(
        n11117), .C2(n14386), .ZN(n3002) );
  AOI222_X1 U2874 ( .A1(n10859), .A2(n14289), .B1(n10856), .B2(n14321), .C1(
        n10853), .C2(n14385), .ZN(n4372) );
  AOI222_X1 U2875 ( .A1(n11123), .A2(n14289), .B1(n11120), .B2(n14321), .C1(
        n11117), .C2(n14385), .ZN(n2939) );
  NOR3_X1 U2876 ( .A1(n14514), .A2(n12769), .A3(n12771), .ZN(n5706) );
  NOR3_X1 U2877 ( .A1(n14516), .A2(n12773), .A3(n12775), .ZN(n4273) );
  NOR2_X1 U2878 ( .A1(n2597), .A2(N2173), .ZN(n2615) );
  BUF_X1 U2879 ( .A(n12768), .Z(n10844) );
  BUF_X1 U2880 ( .A(n12767), .Z(n10837) );
  BUF_X1 U2881 ( .A(n12766), .Z(n10830) );
  BUF_X1 U2882 ( .A(n12765), .Z(n10823) );
  BUF_X1 U2883 ( .A(n12764), .Z(n10816) );
  BUF_X1 U2884 ( .A(n12763), .Z(n10809) );
  BUF_X1 U2885 ( .A(n12762), .Z(n10802) );
  BUF_X1 U2886 ( .A(n12761), .Z(n10795) );
  BUF_X1 U2887 ( .A(n12760), .Z(n10788) );
  BUF_X1 U2888 ( .A(n12759), .Z(n10781) );
  BUF_X1 U2889 ( .A(n12758), .Z(n10774) );
  BUF_X1 U2890 ( .A(n12757), .Z(n10767) );
  BUF_X1 U2891 ( .A(n12756), .Z(n10760) );
  BUF_X1 U2892 ( .A(n12755), .Z(n10753) );
  BUF_X1 U2893 ( .A(n12754), .Z(n10746) );
  BUF_X1 U2894 ( .A(n12753), .Z(n10739) );
  BUF_X1 U2895 ( .A(n12752), .Z(n10732) );
  BUF_X1 U2896 ( .A(n12751), .Z(n10725) );
  BUF_X1 U2897 ( .A(n12750), .Z(n10718) );
  BUF_X1 U2898 ( .A(n12749), .Z(n10711) );
  BUF_X1 U2899 ( .A(n12748), .Z(n10704) );
  BUF_X1 U2900 ( .A(n12747), .Z(n10697) );
  BUF_X1 U2901 ( .A(n12746), .Z(n10690) );
  BUF_X1 U2902 ( .A(n12745), .Z(n10683) );
  BUF_X1 U2903 ( .A(n12744), .Z(n10676) );
  BUF_X1 U2904 ( .A(n12743), .Z(n10669) );
  BUF_X1 U2905 ( .A(n12742), .Z(n10662) );
  BUF_X1 U2906 ( .A(n12741), .Z(n10655) );
  BUF_X1 U2907 ( .A(n12740), .Z(n10648) );
  BUF_X1 U2908 ( .A(n12739), .Z(n10641) );
  BUF_X1 U2909 ( .A(n12738), .Z(n10634) );
  BUF_X1 U2910 ( .A(n12737), .Z(n10627) );
  BUF_X1 U2911 ( .A(n12768), .Z(n10845) );
  BUF_X1 U2912 ( .A(n12767), .Z(n10838) );
  BUF_X1 U2913 ( .A(n12766), .Z(n10831) );
  BUF_X1 U2914 ( .A(n12765), .Z(n10824) );
  BUF_X1 U2915 ( .A(n12764), .Z(n10817) );
  BUF_X1 U2916 ( .A(n12763), .Z(n10810) );
  BUF_X1 U2917 ( .A(n12762), .Z(n10803) );
  BUF_X1 U2918 ( .A(n12761), .Z(n10796) );
  BUF_X1 U2919 ( .A(n12760), .Z(n10789) );
  BUF_X1 U2920 ( .A(n12759), .Z(n10782) );
  BUF_X1 U2921 ( .A(n12758), .Z(n10775) );
  BUF_X1 U2922 ( .A(n12757), .Z(n10768) );
  BUF_X1 U2923 ( .A(n12756), .Z(n10761) );
  BUF_X1 U2924 ( .A(n12755), .Z(n10754) );
  BUF_X1 U2925 ( .A(n12754), .Z(n10747) );
  BUF_X1 U2926 ( .A(n12753), .Z(n10740) );
  BUF_X1 U2927 ( .A(n12752), .Z(n10733) );
  BUF_X1 U2928 ( .A(n12751), .Z(n10726) );
  BUF_X1 U2929 ( .A(n12750), .Z(n10719) );
  BUF_X1 U2930 ( .A(n12749), .Z(n10712) );
  BUF_X1 U2931 ( .A(n12748), .Z(n10705) );
  BUF_X1 U2932 ( .A(n12747), .Z(n10698) );
  BUF_X1 U2933 ( .A(n12746), .Z(n10691) );
  BUF_X1 U2934 ( .A(n12745), .Z(n10684) );
  BUF_X1 U2935 ( .A(n12744), .Z(n10677) );
  BUF_X1 U2936 ( .A(n12743), .Z(n10670) );
  BUF_X1 U2937 ( .A(n12742), .Z(n10663) );
  BUF_X1 U2938 ( .A(n12741), .Z(n10656) );
  BUF_X1 U2939 ( .A(n12740), .Z(n10649) );
  BUF_X1 U2940 ( .A(n12739), .Z(n10642) );
  BUF_X1 U2941 ( .A(n12738), .Z(n10635) );
  BUF_X1 U2942 ( .A(n12737), .Z(n10628) );
  BUF_X1 U2943 ( .A(n12768), .Z(n10846) );
  BUF_X1 U2944 ( .A(n12767), .Z(n10839) );
  BUF_X1 U2945 ( .A(n12766), .Z(n10832) );
  BUF_X1 U2946 ( .A(n12765), .Z(n10825) );
  BUF_X1 U2947 ( .A(n12764), .Z(n10818) );
  BUF_X1 U2948 ( .A(n12763), .Z(n10811) );
  BUF_X1 U2949 ( .A(n12762), .Z(n10804) );
  BUF_X1 U2950 ( .A(n12761), .Z(n10797) );
  BUF_X1 U2951 ( .A(n12760), .Z(n10790) );
  BUF_X1 U2952 ( .A(n12759), .Z(n10783) );
  BUF_X1 U2953 ( .A(n12758), .Z(n10776) );
  BUF_X1 U2954 ( .A(n12757), .Z(n10769) );
  BUF_X1 U2955 ( .A(n12756), .Z(n10762) );
  BUF_X1 U2956 ( .A(n12755), .Z(n10755) );
  BUF_X1 U2957 ( .A(n12754), .Z(n10748) );
  BUF_X1 U2958 ( .A(n12753), .Z(n10741) );
  BUF_X1 U2959 ( .A(n12752), .Z(n10734) );
  BUF_X1 U2960 ( .A(n12751), .Z(n10727) );
  BUF_X1 U2961 ( .A(n12750), .Z(n10720) );
  BUF_X1 U2962 ( .A(n12749), .Z(n10713) );
  BUF_X1 U2963 ( .A(n12748), .Z(n10706) );
  BUF_X1 U2964 ( .A(n12747), .Z(n10699) );
  BUF_X1 U2965 ( .A(n12746), .Z(n10692) );
  BUF_X1 U2966 ( .A(n12745), .Z(n10685) );
  BUF_X1 U2967 ( .A(n12744), .Z(n10678) );
  BUF_X1 U2968 ( .A(n12743), .Z(n10671) );
  BUF_X1 U2969 ( .A(n12742), .Z(n10664) );
  BUF_X1 U2970 ( .A(n12741), .Z(n10657) );
  BUF_X1 U2971 ( .A(n12740), .Z(n10650) );
  BUF_X1 U2972 ( .A(n12739), .Z(n10643) );
  BUF_X1 U2973 ( .A(n12738), .Z(n10636) );
  BUF_X1 U2974 ( .A(n12737), .Z(n10629) );
  BUF_X1 U2975 ( .A(n12768), .Z(n10847) );
  BUF_X1 U2976 ( .A(n12767), .Z(n10840) );
  BUF_X1 U2977 ( .A(n12766), .Z(n10833) );
  BUF_X1 U2978 ( .A(n12765), .Z(n10826) );
  BUF_X1 U2979 ( .A(n12764), .Z(n10819) );
  BUF_X1 U2980 ( .A(n12763), .Z(n10812) );
  BUF_X1 U2981 ( .A(n12762), .Z(n10805) );
  BUF_X1 U2982 ( .A(n12761), .Z(n10798) );
  BUF_X1 U2983 ( .A(n12760), .Z(n10791) );
  BUF_X1 U2984 ( .A(n12759), .Z(n10784) );
  BUF_X1 U2985 ( .A(n12758), .Z(n10777) );
  BUF_X1 U2986 ( .A(n12757), .Z(n10770) );
  BUF_X1 U2987 ( .A(n12756), .Z(n10763) );
  BUF_X1 U2988 ( .A(n12755), .Z(n10756) );
  BUF_X1 U2989 ( .A(n12754), .Z(n10749) );
  BUF_X1 U2990 ( .A(n12753), .Z(n10742) );
  BUF_X1 U2991 ( .A(n12752), .Z(n10735) );
  BUF_X1 U2992 ( .A(n12751), .Z(n10728) );
  BUF_X1 U2993 ( .A(n12750), .Z(n10721) );
  BUF_X1 U2994 ( .A(n12749), .Z(n10714) );
  BUF_X1 U2995 ( .A(n12748), .Z(n10707) );
  BUF_X1 U2996 ( .A(n12747), .Z(n10700) );
  BUF_X1 U2997 ( .A(n12746), .Z(n10693) );
  BUF_X1 U2998 ( .A(n12745), .Z(n10686) );
  BUF_X1 U2999 ( .A(n12744), .Z(n10679) );
  BUF_X1 U3000 ( .A(n12743), .Z(n10672) );
  BUF_X1 U3001 ( .A(n12742), .Z(n10665) );
  BUF_X1 U3002 ( .A(n12741), .Z(n10658) );
  BUF_X1 U3003 ( .A(n12740), .Z(n10651) );
  BUF_X1 U3004 ( .A(n12739), .Z(n10644) );
  BUF_X1 U3005 ( .A(n12738), .Z(n10637) );
  BUF_X1 U3006 ( .A(n12737), .Z(n10630) );
  BUF_X1 U3007 ( .A(n12768), .Z(n10848) );
  BUF_X1 U3008 ( .A(n12767), .Z(n10841) );
  BUF_X1 U3009 ( .A(n12766), .Z(n10834) );
  BUF_X1 U3010 ( .A(n12765), .Z(n10827) );
  BUF_X1 U3011 ( .A(n12764), .Z(n10820) );
  BUF_X1 U3012 ( .A(n12763), .Z(n10813) );
  BUF_X1 U3013 ( .A(n12762), .Z(n10806) );
  BUF_X1 U3014 ( .A(n12761), .Z(n10799) );
  BUF_X1 U3015 ( .A(n12760), .Z(n10792) );
  BUF_X1 U3016 ( .A(n12759), .Z(n10785) );
  BUF_X1 U3017 ( .A(n12758), .Z(n10778) );
  BUF_X1 U3018 ( .A(n12757), .Z(n10771) );
  BUF_X1 U3019 ( .A(n12756), .Z(n10764) );
  BUF_X1 U3020 ( .A(n12755), .Z(n10757) );
  BUF_X1 U3021 ( .A(n12754), .Z(n10750) );
  BUF_X1 U3022 ( .A(n12753), .Z(n10743) );
  BUF_X1 U3023 ( .A(n12752), .Z(n10736) );
  BUF_X1 U3024 ( .A(n12751), .Z(n10729) );
  BUF_X1 U3025 ( .A(n12750), .Z(n10722) );
  BUF_X1 U3026 ( .A(n12749), .Z(n10715) );
  BUF_X1 U3027 ( .A(n12748), .Z(n10708) );
  BUF_X1 U3028 ( .A(n12747), .Z(n10701) );
  BUF_X1 U3029 ( .A(n12746), .Z(n10694) );
  BUF_X1 U3030 ( .A(n12745), .Z(n10687) );
  BUF_X1 U3031 ( .A(n12744), .Z(n10680) );
  BUF_X1 U3032 ( .A(n12743), .Z(n10673) );
  BUF_X1 U3033 ( .A(n12742), .Z(n10666) );
  BUF_X1 U3034 ( .A(n12741), .Z(n10659) );
  BUF_X1 U3035 ( .A(n12740), .Z(n10652) );
  BUF_X1 U3036 ( .A(n12739), .Z(n10645) );
  BUF_X1 U3037 ( .A(n12738), .Z(n10638) );
  BUF_X1 U3038 ( .A(n12737), .Z(n10631) );
  BUF_X1 U3039 ( .A(n12768), .Z(n10849) );
  BUF_X1 U3040 ( .A(n12767), .Z(n10842) );
  BUF_X1 U3041 ( .A(n12766), .Z(n10835) );
  BUF_X1 U3042 ( .A(n12765), .Z(n10828) );
  BUF_X1 U3043 ( .A(n12764), .Z(n10821) );
  BUF_X1 U3044 ( .A(n12763), .Z(n10814) );
  BUF_X1 U3045 ( .A(n12762), .Z(n10807) );
  BUF_X1 U3046 ( .A(n12761), .Z(n10800) );
  BUF_X1 U3047 ( .A(n12760), .Z(n10793) );
  BUF_X1 U3048 ( .A(n12759), .Z(n10786) );
  BUF_X1 U3049 ( .A(n12758), .Z(n10779) );
  BUF_X1 U3050 ( .A(n12757), .Z(n10772) );
  BUF_X1 U3051 ( .A(n12756), .Z(n10765) );
  BUF_X1 U3052 ( .A(n12755), .Z(n10758) );
  BUF_X1 U3053 ( .A(n12754), .Z(n10751) );
  BUF_X1 U3054 ( .A(n12753), .Z(n10744) );
  BUF_X1 U3055 ( .A(n12752), .Z(n10737) );
  BUF_X1 U3056 ( .A(n12751), .Z(n10730) );
  BUF_X1 U3057 ( .A(n12750), .Z(n10723) );
  BUF_X1 U3058 ( .A(n12749), .Z(n10716) );
  BUF_X1 U3059 ( .A(n12748), .Z(n10709) );
  BUF_X1 U3060 ( .A(n12747), .Z(n10702) );
  BUF_X1 U3061 ( .A(n12746), .Z(n10695) );
  BUF_X1 U3062 ( .A(n12745), .Z(n10688) );
  BUF_X1 U3063 ( .A(n12744), .Z(n10681) );
  BUF_X1 U3064 ( .A(n12743), .Z(n10674) );
  BUF_X1 U3065 ( .A(n12742), .Z(n10667) );
  BUF_X1 U3066 ( .A(n12741), .Z(n10660) );
  BUF_X1 U3067 ( .A(n12740), .Z(n10653) );
  BUF_X1 U3068 ( .A(n12739), .Z(n10646) );
  BUF_X1 U3069 ( .A(n12738), .Z(n10639) );
  BUF_X1 U3070 ( .A(n12737), .Z(n10632) );
  AND2_X1 U3071 ( .A1(N2171), .A2(n2571), .ZN(n2492) );
  NOR3_X1 U3072 ( .A1(n2597), .A2(N2172), .A3(n12731), .ZN(n2571) );
  INV_X1 U3073 ( .A(N2173), .ZN(n12731) );
  NOR2_X1 U3074 ( .A1(n14514), .A2(N8434), .ZN(n5653) );
  NOR2_X1 U3075 ( .A1(n14516), .A2(N8578), .ZN(n4220) );
  BUF_X1 U3076 ( .A(n12768), .Z(n10850) );
  BUF_X1 U3077 ( .A(n12767), .Z(n10843) );
  BUF_X1 U3078 ( .A(n12766), .Z(n10836) );
  BUF_X1 U3079 ( .A(n12765), .Z(n10829) );
  BUF_X1 U3080 ( .A(n12764), .Z(n10822) );
  BUF_X1 U3081 ( .A(n12763), .Z(n10815) );
  BUF_X1 U3082 ( .A(n12762), .Z(n10808) );
  BUF_X1 U3083 ( .A(n12761), .Z(n10801) );
  BUF_X1 U3084 ( .A(n12760), .Z(n10794) );
  BUF_X1 U3085 ( .A(n12759), .Z(n10787) );
  BUF_X1 U3086 ( .A(n12758), .Z(n10780) );
  BUF_X1 U3087 ( .A(n12757), .Z(n10773) );
  BUF_X1 U3088 ( .A(n12756), .Z(n10766) );
  BUF_X1 U3089 ( .A(n12755), .Z(n10759) );
  BUF_X1 U3090 ( .A(n12754), .Z(n10752) );
  BUF_X1 U3091 ( .A(n12753), .Z(n10745) );
  BUF_X1 U3092 ( .A(n12752), .Z(n10738) );
  BUF_X1 U3093 ( .A(n12751), .Z(n10731) );
  BUF_X1 U3094 ( .A(n12750), .Z(n10724) );
  BUF_X1 U3095 ( .A(n12749), .Z(n10717) );
  BUF_X1 U3096 ( .A(n12748), .Z(n10710) );
  BUF_X1 U3097 ( .A(n12747), .Z(n10703) );
  BUF_X1 U3098 ( .A(n12746), .Z(n10696) );
  BUF_X1 U3099 ( .A(n12745), .Z(n10689) );
  BUF_X1 U3100 ( .A(n12744), .Z(n10682) );
  BUF_X1 U3101 ( .A(n12743), .Z(n10675) );
  BUF_X1 U3102 ( .A(n12742), .Z(n10668) );
  BUF_X1 U3103 ( .A(n12741), .Z(n10661) );
  BUF_X1 U3104 ( .A(n12740), .Z(n10654) );
  BUF_X1 U3105 ( .A(n12739), .Z(n10647) );
  BUF_X1 U3106 ( .A(n12738), .Z(n10640) );
  BUF_X1 U3107 ( .A(n12737), .Z(n10633) );
  AND2_X1 U3108 ( .A1(n2719), .A2(n2730), .ZN(n2494) );
  AND2_X1 U3109 ( .A1(n2721), .A2(n2730), .ZN(n2496) );
  AND2_X1 U3110 ( .A1(n2723), .A2(n2730), .ZN(n2498) );
  AND2_X1 U3111 ( .A1(n2735), .A2(n2717), .ZN(n2500) );
  AND2_X1 U3112 ( .A1(n2735), .A2(n2719), .ZN(n2566) );
  AND2_X1 U3113 ( .A1(n2735), .A2(n2721), .ZN(n2568) );
  AND2_X1 U3114 ( .A1(n2735), .A2(n2723), .ZN(n2570) );
  NAND2_X1 U3115 ( .A1(N8437), .A2(n5659), .ZN(n4389) );
  NAND2_X1 U3116 ( .A1(N8581), .A2(n4226), .ZN(n2956) );
  INV_X1 U3117 ( .A(N8437), .ZN(n12769) );
  INV_X1 U3118 ( .A(N8581), .ZN(n12773) );
  NOR2_X1 U3119 ( .A1(n12734), .A2(N2170), .ZN(n2730) );
  NOR2_X1 U3120 ( .A1(n12735), .A2(n12736), .ZN(n2717) );
  NOR2_X1 U3121 ( .A1(n14514), .A2(n12772), .ZN(n5702) );
  NOR2_X1 U3122 ( .A1(n14516), .A2(n12776), .ZN(n4269) );
  AND2_X1 U3123 ( .A1(n5647), .A2(n5703), .ZN(n5655) );
  AND2_X1 U3124 ( .A1(n5647), .A2(n5702), .ZN(n5657) );
  AND2_X1 U3125 ( .A1(n4214), .A2(n4270), .ZN(n4222) );
  AND2_X1 U3126 ( .A1(n4214), .A2(n4269), .ZN(n4224) );
  AND2_X1 U3127 ( .A1(n5649), .A2(n5703), .ZN(n5656) );
  AND2_X1 U3128 ( .A1(n4216), .A2(n4270), .ZN(n4223) );
  INV_X1 U3129 ( .A(N8435), .ZN(n12771) );
  INV_X1 U3130 ( .A(N8579), .ZN(n12775) );
  AND2_X1 U3131 ( .A1(n2716), .A2(n2717), .ZN(n2573) );
  AND2_X1 U3132 ( .A1(n2716), .A2(n2719), .ZN(n2576) );
  AND2_X1 U3133 ( .A1(n2716), .A2(n2721), .ZN(n2578) );
  AND2_X1 U3134 ( .A1(n2716), .A2(n2723), .ZN(n2580) );
  AND2_X1 U3135 ( .A1(n2725), .A2(n2719), .ZN(n2584) );
  AND2_X1 U3136 ( .A1(n2725), .A2(n2721), .ZN(n2586) );
  AND2_X1 U3137 ( .A1(n2725), .A2(n2723), .ZN(n2588) );
  AND2_X1 U3138 ( .A1(n5651), .A2(n5703), .ZN(n5661) );
  AND2_X1 U3139 ( .A1(n4218), .A2(n4270), .ZN(n4228) );
  NAND2_X1 U3140 ( .A1(n5655), .A2(N8437), .ZN(n4385) );
  NAND2_X1 U3141 ( .A1(n5657), .A2(N8437), .ZN(n4386) );
  NAND2_X1 U3142 ( .A1(n5656), .A2(N8437), .ZN(n4390) );
  NAND2_X1 U3143 ( .A1(n5663), .A2(N8437), .ZN(n4388) );
  NAND2_X1 U3144 ( .A1(n5661), .A2(N8437), .ZN(n4396) );
  NAND2_X1 U3145 ( .A1(n5665), .A2(N8437), .ZN(n4395) );
  NAND2_X1 U3146 ( .A1(n4222), .A2(N8581), .ZN(n2952) );
  NAND2_X1 U3147 ( .A1(n4224), .A2(N8581), .ZN(n2953) );
  NAND2_X1 U3148 ( .A1(n4223), .A2(N8581), .ZN(n2957) );
  NAND2_X1 U3149 ( .A1(n4230), .A2(N8581), .ZN(n2955) );
  NAND2_X1 U3150 ( .A1(n4228), .A2(N8581), .ZN(n2963) );
  NAND2_X1 U3151 ( .A1(n4232), .A2(N8581), .ZN(n2962) );
  NAND4_X1 U3152 ( .A1(n5638), .A2(n5639), .A3(n5640), .A4(n5641), .ZN(n5637)
         );
  AOI221_X1 U3153 ( .B1(n11079), .B2(n12819), .C1(n11076), .C2(n13011), .A(
        n5658), .ZN(n5640) );
  NOR4_X1 U3154 ( .A1(n5642), .A2(n5643), .A3(n5644), .A4(n5645), .ZN(n5641)
         );
  AOI222_X1 U3155 ( .A1(n11055), .A2(n12851), .B1(n11052), .B2(n12883), .C1(
        n11049), .C2(n12947), .ZN(n5638) );
  NAND4_X1 U3156 ( .A1(n4205), .A2(n4206), .A3(n4207), .A4(n4208), .ZN(n4204)
         );
  AOI221_X1 U3157 ( .B1(n11343), .B2(n12819), .C1(n11340), .C2(n13011), .A(
        n4225), .ZN(n4207) );
  NOR4_X1 U3158 ( .A1(n4209), .A2(n4210), .A3(n4211), .A4(n4212), .ZN(n4208)
         );
  AOI222_X1 U3159 ( .A1(n11319), .A2(n12851), .B1(n11316), .B2(n12883), .C1(
        n11313), .C2(n12947), .ZN(n4205) );
  NAND4_X1 U3160 ( .A1(n5597), .A2(n5598), .A3(n5599), .A4(n5600), .ZN(n5596)
         );
  AOI221_X1 U3161 ( .B1(n11079), .B2(n12818), .C1(n11076), .C2(n13010), .A(
        n5605), .ZN(n5599) );
  NOR4_X1 U3162 ( .A1(n5601), .A2(n5602), .A3(n5603), .A4(n5604), .ZN(n5600)
         );
  AOI222_X1 U3163 ( .A1(n11055), .A2(n12850), .B1(n11052), .B2(n12882), .C1(
        n11049), .C2(n12946), .ZN(n5597) );
  NAND4_X1 U3164 ( .A1(n4164), .A2(n4165), .A3(n4166), .A4(n4167), .ZN(n4163)
         );
  AOI221_X1 U3165 ( .B1(n11343), .B2(n12818), .C1(n11340), .C2(n13010), .A(
        n4172), .ZN(n4166) );
  NOR4_X1 U3166 ( .A1(n4168), .A2(n4169), .A3(n4170), .A4(n4171), .ZN(n4167)
         );
  AOI222_X1 U3167 ( .A1(n11319), .A2(n12850), .B1(n11316), .B2(n12882), .C1(
        n11313), .C2(n12946), .ZN(n4164) );
  NAND4_X1 U3168 ( .A1(n5556), .A2(n5557), .A3(n5558), .A4(n5559), .ZN(n5555)
         );
  AOI221_X1 U3169 ( .B1(n11079), .B2(n12817), .C1(n11076), .C2(n13009), .A(
        n5564), .ZN(n5558) );
  NOR4_X1 U3170 ( .A1(n5560), .A2(n5561), .A3(n5562), .A4(n5563), .ZN(n5559)
         );
  AOI222_X1 U3171 ( .A1(n11055), .A2(n12849), .B1(n11052), .B2(n12881), .C1(
        n11049), .C2(n12945), .ZN(n5556) );
  NAND4_X1 U3172 ( .A1(n4123), .A2(n4124), .A3(n4125), .A4(n4126), .ZN(n4122)
         );
  AOI221_X1 U3173 ( .B1(n11343), .B2(n12817), .C1(n11340), .C2(n13009), .A(
        n4131), .ZN(n4125) );
  NOR4_X1 U3174 ( .A1(n4127), .A2(n4128), .A3(n4129), .A4(n4130), .ZN(n4126)
         );
  AOI222_X1 U3175 ( .A1(n11319), .A2(n12849), .B1(n11316), .B2(n12881), .C1(
        n11313), .C2(n12945), .ZN(n4123) );
  NAND4_X1 U3176 ( .A1(n5515), .A2(n5516), .A3(n5517), .A4(n5518), .ZN(n5514)
         );
  AOI221_X1 U3177 ( .B1(n11079), .B2(n12816), .C1(n11076), .C2(n13008), .A(
        n5523), .ZN(n5517) );
  NOR4_X1 U3178 ( .A1(n5519), .A2(n5520), .A3(n5521), .A4(n5522), .ZN(n5518)
         );
  AOI222_X1 U3179 ( .A1(n11055), .A2(n12848), .B1(n11052), .B2(n12880), .C1(
        n11049), .C2(n12944), .ZN(n5515) );
  NAND4_X1 U3180 ( .A1(n4082), .A2(n4083), .A3(n4084), .A4(n4085), .ZN(n4081)
         );
  AOI221_X1 U3181 ( .B1(n11343), .B2(n12816), .C1(n11340), .C2(n13008), .A(
        n4090), .ZN(n4084) );
  NOR4_X1 U3182 ( .A1(n4086), .A2(n4087), .A3(n4088), .A4(n4089), .ZN(n4085)
         );
  AOI222_X1 U3183 ( .A1(n11319), .A2(n12848), .B1(n11316), .B2(n12880), .C1(
        n11313), .C2(n12944), .ZN(n4082) );
  NAND4_X1 U3184 ( .A1(n5474), .A2(n5475), .A3(n5476), .A4(n5477), .ZN(n5473)
         );
  AOI221_X1 U3185 ( .B1(n11079), .B2(n12815), .C1(n11076), .C2(n13007), .A(
        n5482), .ZN(n5476) );
  NOR4_X1 U3186 ( .A1(n5478), .A2(n5479), .A3(n5480), .A4(n5481), .ZN(n5477)
         );
  AOI222_X1 U3187 ( .A1(n11055), .A2(n12847), .B1(n11052), .B2(n12879), .C1(
        n11049), .C2(n12943), .ZN(n5474) );
  NAND4_X1 U3188 ( .A1(n4041), .A2(n4042), .A3(n4043), .A4(n4044), .ZN(n4040)
         );
  AOI221_X1 U3189 ( .B1(n11343), .B2(n12815), .C1(n11340), .C2(n13007), .A(
        n4049), .ZN(n4043) );
  NOR4_X1 U3190 ( .A1(n4045), .A2(n4046), .A3(n4047), .A4(n4048), .ZN(n4044)
         );
  AOI222_X1 U3191 ( .A1(n11319), .A2(n12847), .B1(n11316), .B2(n12879), .C1(
        n11313), .C2(n12943), .ZN(n4041) );
  NAND4_X1 U3192 ( .A1(n5433), .A2(n5434), .A3(n5435), .A4(n5436), .ZN(n5432)
         );
  AOI221_X1 U3193 ( .B1(n11079), .B2(n12814), .C1(n11076), .C2(n13006), .A(
        n5441), .ZN(n5435) );
  NOR4_X1 U3194 ( .A1(n5437), .A2(n5438), .A3(n5439), .A4(n5440), .ZN(n5436)
         );
  AOI222_X1 U3195 ( .A1(n11055), .A2(n12846), .B1(n11052), .B2(n12878), .C1(
        n11049), .C2(n12942), .ZN(n5433) );
  NAND4_X1 U3196 ( .A1(n4000), .A2(n4001), .A3(n4002), .A4(n4003), .ZN(n3999)
         );
  AOI221_X1 U3197 ( .B1(n11343), .B2(n12814), .C1(n11340), .C2(n13006), .A(
        n4008), .ZN(n4002) );
  NOR4_X1 U3198 ( .A1(n4004), .A2(n4005), .A3(n4006), .A4(n4007), .ZN(n4003)
         );
  AOI222_X1 U3199 ( .A1(n11319), .A2(n12846), .B1(n11316), .B2(n12878), .C1(
        n11313), .C2(n12942), .ZN(n4000) );
  NAND4_X1 U3200 ( .A1(n5392), .A2(n5393), .A3(n5394), .A4(n5395), .ZN(n5391)
         );
  AOI221_X1 U3201 ( .B1(n11079), .B2(n12813), .C1(n11076), .C2(n13005), .A(
        n5400), .ZN(n5394) );
  NOR4_X1 U3202 ( .A1(n5396), .A2(n5397), .A3(n5398), .A4(n5399), .ZN(n5395)
         );
  AOI222_X1 U3203 ( .A1(n11055), .A2(n12845), .B1(n11052), .B2(n12877), .C1(
        n11049), .C2(n12941), .ZN(n5392) );
  NAND4_X1 U3204 ( .A1(n3959), .A2(n3960), .A3(n3961), .A4(n3962), .ZN(n3958)
         );
  AOI221_X1 U3205 ( .B1(n11343), .B2(n12813), .C1(n11340), .C2(n13005), .A(
        n3967), .ZN(n3961) );
  NOR4_X1 U3206 ( .A1(n3963), .A2(n3964), .A3(n3965), .A4(n3966), .ZN(n3962)
         );
  AOI222_X1 U3207 ( .A1(n11319), .A2(n12845), .B1(n11316), .B2(n12877), .C1(
        n11313), .C2(n12941), .ZN(n3959) );
  NAND4_X1 U3208 ( .A1(n5351), .A2(n5352), .A3(n5353), .A4(n5354), .ZN(n5350)
         );
  AOI221_X1 U3209 ( .B1(n11079), .B2(n12812), .C1(n11076), .C2(n13004), .A(
        n5359), .ZN(n5353) );
  NOR4_X1 U3210 ( .A1(n5355), .A2(n5356), .A3(n5357), .A4(n5358), .ZN(n5354)
         );
  AOI222_X1 U3211 ( .A1(n11055), .A2(n12844), .B1(n11052), .B2(n12876), .C1(
        n11049), .C2(n12940), .ZN(n5351) );
  NAND4_X1 U3212 ( .A1(n3918), .A2(n3919), .A3(n3920), .A4(n3921), .ZN(n3917)
         );
  AOI221_X1 U3213 ( .B1(n11343), .B2(n12812), .C1(n11340), .C2(n13004), .A(
        n3926), .ZN(n3920) );
  NOR4_X1 U3214 ( .A1(n3922), .A2(n3923), .A3(n3924), .A4(n3925), .ZN(n3921)
         );
  AOI222_X1 U3215 ( .A1(n11319), .A2(n12844), .B1(n11316), .B2(n12876), .C1(
        n11313), .C2(n12940), .ZN(n3918) );
  NAND4_X1 U3216 ( .A1(n5310), .A2(n5311), .A3(n5312), .A4(n5313), .ZN(n5309)
         );
  AOI221_X1 U3217 ( .B1(n11079), .B2(n12811), .C1(n11076), .C2(n13003), .A(
        n5318), .ZN(n5312) );
  NOR4_X1 U3218 ( .A1(n5314), .A2(n5315), .A3(n5316), .A4(n5317), .ZN(n5313)
         );
  AOI222_X1 U3219 ( .A1(n11055), .A2(n12843), .B1(n11052), .B2(n12875), .C1(
        n11049), .C2(n12939), .ZN(n5310) );
  NAND4_X1 U3220 ( .A1(n3877), .A2(n3878), .A3(n3879), .A4(n3880), .ZN(n3876)
         );
  AOI221_X1 U3221 ( .B1(n11343), .B2(n12811), .C1(n11340), .C2(n13003), .A(
        n3885), .ZN(n3879) );
  NOR4_X1 U3222 ( .A1(n3881), .A2(n3882), .A3(n3883), .A4(n3884), .ZN(n3880)
         );
  AOI222_X1 U3223 ( .A1(n11319), .A2(n12843), .B1(n11316), .B2(n12875), .C1(
        n11313), .C2(n12939), .ZN(n3877) );
  NAND4_X1 U3224 ( .A1(n5269), .A2(n5270), .A3(n5271), .A4(n5272), .ZN(n5268)
         );
  AOI221_X1 U3225 ( .B1(n11079), .B2(n12810), .C1(n11076), .C2(n13002), .A(
        n5277), .ZN(n5271) );
  NOR4_X1 U3226 ( .A1(n5273), .A2(n5274), .A3(n5275), .A4(n5276), .ZN(n5272)
         );
  AOI222_X1 U3227 ( .A1(n11055), .A2(n12842), .B1(n11052), .B2(n12874), .C1(
        n11049), .C2(n12938), .ZN(n5269) );
  NAND4_X1 U3228 ( .A1(n3836), .A2(n3837), .A3(n3838), .A4(n3839), .ZN(n3835)
         );
  AOI221_X1 U3229 ( .B1(n11343), .B2(n12810), .C1(n11340), .C2(n13002), .A(
        n3844), .ZN(n3838) );
  NOR4_X1 U3230 ( .A1(n3840), .A2(n3841), .A3(n3842), .A4(n3843), .ZN(n3839)
         );
  AOI222_X1 U3231 ( .A1(n11319), .A2(n12842), .B1(n11316), .B2(n12874), .C1(
        n11313), .C2(n12938), .ZN(n3836) );
  NAND4_X1 U3232 ( .A1(n5228), .A2(n5229), .A3(n5230), .A4(n5231), .ZN(n5227)
         );
  AOI221_X1 U3233 ( .B1(n11079), .B2(n12809), .C1(n11076), .C2(n13001), .A(
        n5236), .ZN(n5230) );
  NOR4_X1 U3234 ( .A1(n5232), .A2(n5233), .A3(n5234), .A4(n5235), .ZN(n5231)
         );
  AOI222_X1 U3235 ( .A1(n11055), .A2(n12841), .B1(n11052), .B2(n12873), .C1(
        n11049), .C2(n12937), .ZN(n5228) );
  NAND4_X1 U3236 ( .A1(n3795), .A2(n3796), .A3(n3797), .A4(n3798), .ZN(n3794)
         );
  AOI221_X1 U3237 ( .B1(n11343), .B2(n12809), .C1(n11340), .C2(n13001), .A(
        n3803), .ZN(n3797) );
  NOR4_X1 U3238 ( .A1(n3799), .A2(n3800), .A3(n3801), .A4(n3802), .ZN(n3798)
         );
  AOI222_X1 U3239 ( .A1(n11319), .A2(n12841), .B1(n11316), .B2(n12873), .C1(
        n11313), .C2(n12937), .ZN(n3795) );
  NAND4_X1 U3240 ( .A1(n5187), .A2(n5188), .A3(n5189), .A4(n5190), .ZN(n5186)
         );
  AOI221_X1 U3241 ( .B1(n11079), .B2(n12808), .C1(n11076), .C2(n13000), .A(
        n5195), .ZN(n5189) );
  NOR4_X1 U3242 ( .A1(n5191), .A2(n5192), .A3(n5193), .A4(n5194), .ZN(n5190)
         );
  AOI222_X1 U3243 ( .A1(n11055), .A2(n12840), .B1(n11052), .B2(n12872), .C1(
        n11049), .C2(n12936), .ZN(n5187) );
  NAND4_X1 U3244 ( .A1(n3754), .A2(n3755), .A3(n3756), .A4(n3757), .ZN(n3753)
         );
  AOI221_X1 U3245 ( .B1(n11343), .B2(n12808), .C1(n11340), .C2(n13000), .A(
        n3762), .ZN(n3756) );
  NOR4_X1 U3246 ( .A1(n3758), .A2(n3759), .A3(n3760), .A4(n3761), .ZN(n3757)
         );
  AOI222_X1 U3247 ( .A1(n11319), .A2(n12840), .B1(n11316), .B2(n12872), .C1(
        n11313), .C2(n12936), .ZN(n3754) );
  NAND4_X1 U3248 ( .A1(n5146), .A2(n5147), .A3(n5148), .A4(n5149), .ZN(n5145)
         );
  AOI221_X1 U3249 ( .B1(n11080), .B2(n12807), .C1(n11077), .C2(n12999), .A(
        n5154), .ZN(n5148) );
  NOR4_X1 U3250 ( .A1(n5150), .A2(n5151), .A3(n5152), .A4(n5153), .ZN(n5149)
         );
  AOI222_X1 U3251 ( .A1(n11056), .A2(n12839), .B1(n11053), .B2(n12871), .C1(
        n11050), .C2(n12935), .ZN(n5146) );
  NAND4_X1 U3252 ( .A1(n3713), .A2(n3714), .A3(n3715), .A4(n3716), .ZN(n3712)
         );
  AOI221_X1 U3253 ( .B1(n11344), .B2(n12807), .C1(n11341), .C2(n12999), .A(
        n3721), .ZN(n3715) );
  NOR4_X1 U3254 ( .A1(n3717), .A2(n3718), .A3(n3719), .A4(n3720), .ZN(n3716)
         );
  AOI222_X1 U3255 ( .A1(n11320), .A2(n12839), .B1(n11317), .B2(n12871), .C1(
        n11314), .C2(n12935), .ZN(n3713) );
  NAND4_X1 U3256 ( .A1(n5105), .A2(n5106), .A3(n5107), .A4(n5108), .ZN(n5104)
         );
  AOI221_X1 U3257 ( .B1(n11080), .B2(n12806), .C1(n11077), .C2(n12998), .A(
        n5113), .ZN(n5107) );
  NOR4_X1 U3258 ( .A1(n5109), .A2(n5110), .A3(n5111), .A4(n5112), .ZN(n5108)
         );
  AOI222_X1 U3259 ( .A1(n11056), .A2(n12838), .B1(n11053), .B2(n12870), .C1(
        n11050), .C2(n12934), .ZN(n5105) );
  NAND4_X1 U3260 ( .A1(n3672), .A2(n3673), .A3(n3674), .A4(n3675), .ZN(n3671)
         );
  AOI221_X1 U3261 ( .B1(n11344), .B2(n12806), .C1(n11341), .C2(n12998), .A(
        n3680), .ZN(n3674) );
  NOR4_X1 U3262 ( .A1(n3676), .A2(n3677), .A3(n3678), .A4(n3679), .ZN(n3675)
         );
  AOI222_X1 U3263 ( .A1(n11320), .A2(n12838), .B1(n11317), .B2(n12870), .C1(
        n11314), .C2(n12934), .ZN(n3672) );
  NAND4_X1 U3264 ( .A1(n5064), .A2(n5065), .A3(n5066), .A4(n5067), .ZN(n5063)
         );
  AOI221_X1 U3265 ( .B1(n11080), .B2(n12805), .C1(n11077), .C2(n12997), .A(
        n5072), .ZN(n5066) );
  NOR4_X1 U3266 ( .A1(n5068), .A2(n5069), .A3(n5070), .A4(n5071), .ZN(n5067)
         );
  AOI222_X1 U3267 ( .A1(n11056), .A2(n12837), .B1(n11053), .B2(n12869), .C1(
        n11050), .C2(n12933), .ZN(n5064) );
  NAND4_X1 U3268 ( .A1(n3631), .A2(n3632), .A3(n3633), .A4(n3634), .ZN(n3630)
         );
  AOI221_X1 U3269 ( .B1(n11344), .B2(n12805), .C1(n11341), .C2(n12997), .A(
        n3639), .ZN(n3633) );
  NOR4_X1 U3270 ( .A1(n3635), .A2(n3636), .A3(n3637), .A4(n3638), .ZN(n3634)
         );
  AOI222_X1 U3271 ( .A1(n11320), .A2(n12837), .B1(n11317), .B2(n12869), .C1(
        n11314), .C2(n12933), .ZN(n3631) );
  NAND4_X1 U3272 ( .A1(n5023), .A2(n5024), .A3(n5025), .A4(n5026), .ZN(n5022)
         );
  AOI221_X1 U3273 ( .B1(n11080), .B2(n12804), .C1(n11077), .C2(n12996), .A(
        n5031), .ZN(n5025) );
  NOR4_X1 U3274 ( .A1(n5027), .A2(n5028), .A3(n5029), .A4(n5030), .ZN(n5026)
         );
  AOI222_X1 U3275 ( .A1(n11056), .A2(n12836), .B1(n11053), .B2(n12868), .C1(
        n11050), .C2(n12932), .ZN(n5023) );
  NAND4_X1 U3276 ( .A1(n3590), .A2(n3591), .A3(n3592), .A4(n3593), .ZN(n3589)
         );
  AOI221_X1 U3277 ( .B1(n11344), .B2(n12804), .C1(n11341), .C2(n12996), .A(
        n3598), .ZN(n3592) );
  NOR4_X1 U3278 ( .A1(n3594), .A2(n3595), .A3(n3596), .A4(n3597), .ZN(n3593)
         );
  AOI222_X1 U3279 ( .A1(n11320), .A2(n12836), .B1(n11317), .B2(n12868), .C1(
        n11314), .C2(n12932), .ZN(n3590) );
  NAND4_X1 U3280 ( .A1(n4982), .A2(n4983), .A3(n4984), .A4(n4985), .ZN(n4981)
         );
  AOI221_X1 U3281 ( .B1(n11080), .B2(n12803), .C1(n11077), .C2(n12995), .A(
        n4990), .ZN(n4984) );
  NOR4_X1 U3282 ( .A1(n4986), .A2(n4987), .A3(n4988), .A4(n4989), .ZN(n4985)
         );
  AOI222_X1 U3283 ( .A1(n11056), .A2(n12835), .B1(n11053), .B2(n12867), .C1(
        n11050), .C2(n12931), .ZN(n4982) );
  NAND4_X1 U3284 ( .A1(n3549), .A2(n3550), .A3(n3551), .A4(n3552), .ZN(n3548)
         );
  AOI221_X1 U3285 ( .B1(n11344), .B2(n12803), .C1(n11341), .C2(n12995), .A(
        n3557), .ZN(n3551) );
  NOR4_X1 U3286 ( .A1(n3553), .A2(n3554), .A3(n3555), .A4(n3556), .ZN(n3552)
         );
  AOI222_X1 U3287 ( .A1(n11320), .A2(n12835), .B1(n11317), .B2(n12867), .C1(
        n11314), .C2(n12931), .ZN(n3549) );
  NAND4_X1 U3288 ( .A1(n4941), .A2(n4942), .A3(n4943), .A4(n4944), .ZN(n4940)
         );
  AOI221_X1 U3289 ( .B1(n11080), .B2(n12802), .C1(n11077), .C2(n12994), .A(
        n4949), .ZN(n4943) );
  NOR4_X1 U3290 ( .A1(n4945), .A2(n4946), .A3(n4947), .A4(n4948), .ZN(n4944)
         );
  AOI222_X1 U3291 ( .A1(n11056), .A2(n12834), .B1(n11053), .B2(n12866), .C1(
        n11050), .C2(n12930), .ZN(n4941) );
  NAND4_X1 U3292 ( .A1(n3508), .A2(n3509), .A3(n3510), .A4(n3511), .ZN(n3507)
         );
  AOI221_X1 U3293 ( .B1(n11344), .B2(n12802), .C1(n11341), .C2(n12994), .A(
        n3516), .ZN(n3510) );
  NOR4_X1 U3294 ( .A1(n3512), .A2(n3513), .A3(n3514), .A4(n3515), .ZN(n3511)
         );
  AOI222_X1 U3295 ( .A1(n11320), .A2(n12834), .B1(n11317), .B2(n12866), .C1(
        n11314), .C2(n12930), .ZN(n3508) );
  NAND4_X1 U3296 ( .A1(n4900), .A2(n4901), .A3(n4902), .A4(n4903), .ZN(n4899)
         );
  AOI221_X1 U3297 ( .B1(n11080), .B2(n12801), .C1(n11077), .C2(n12993), .A(
        n4908), .ZN(n4902) );
  NOR4_X1 U3298 ( .A1(n4904), .A2(n4905), .A3(n4906), .A4(n4907), .ZN(n4903)
         );
  AOI222_X1 U3299 ( .A1(n11056), .A2(n12833), .B1(n11053), .B2(n12865), .C1(
        n11050), .C2(n12929), .ZN(n4900) );
  NAND4_X1 U3300 ( .A1(n3467), .A2(n3468), .A3(n3469), .A4(n3470), .ZN(n3466)
         );
  AOI221_X1 U3301 ( .B1(n11344), .B2(n12801), .C1(n11341), .C2(n12993), .A(
        n3475), .ZN(n3469) );
  NOR4_X1 U3302 ( .A1(n3471), .A2(n3472), .A3(n3473), .A4(n3474), .ZN(n3470)
         );
  AOI222_X1 U3303 ( .A1(n11320), .A2(n12833), .B1(n11317), .B2(n12865), .C1(
        n11314), .C2(n12929), .ZN(n3467) );
  NAND4_X1 U3304 ( .A1(n4859), .A2(n4860), .A3(n4861), .A4(n4862), .ZN(n4858)
         );
  AOI221_X1 U3305 ( .B1(n11080), .B2(n12800), .C1(n11077), .C2(n12992), .A(
        n4867), .ZN(n4861) );
  NOR4_X1 U3306 ( .A1(n4863), .A2(n4864), .A3(n4865), .A4(n4866), .ZN(n4862)
         );
  AOI222_X1 U3307 ( .A1(n11056), .A2(n12832), .B1(n11053), .B2(n12864), .C1(
        n11050), .C2(n12928), .ZN(n4859) );
  NAND4_X1 U3308 ( .A1(n3426), .A2(n3427), .A3(n3428), .A4(n3429), .ZN(n3425)
         );
  AOI221_X1 U3309 ( .B1(n11344), .B2(n12800), .C1(n11341), .C2(n12992), .A(
        n3434), .ZN(n3428) );
  NOR4_X1 U3310 ( .A1(n3430), .A2(n3431), .A3(n3432), .A4(n3433), .ZN(n3429)
         );
  AOI222_X1 U3311 ( .A1(n11320), .A2(n12832), .B1(n11317), .B2(n12864), .C1(
        n11314), .C2(n12928), .ZN(n3426) );
  NAND4_X1 U3312 ( .A1(n4818), .A2(n4819), .A3(n4820), .A4(n4821), .ZN(n4817)
         );
  AOI221_X1 U3313 ( .B1(n11080), .B2(n12799), .C1(n11077), .C2(n12991), .A(
        n4826), .ZN(n4820) );
  NOR4_X1 U3314 ( .A1(n4822), .A2(n4823), .A3(n4824), .A4(n4825), .ZN(n4821)
         );
  AOI222_X1 U3315 ( .A1(n11056), .A2(n12831), .B1(n11053), .B2(n12863), .C1(
        n11050), .C2(n12927), .ZN(n4818) );
  NAND4_X1 U3316 ( .A1(n3385), .A2(n3386), .A3(n3387), .A4(n3388), .ZN(n3384)
         );
  AOI221_X1 U3317 ( .B1(n11344), .B2(n12799), .C1(n11341), .C2(n12991), .A(
        n3393), .ZN(n3387) );
  NOR4_X1 U3318 ( .A1(n3389), .A2(n3390), .A3(n3391), .A4(n3392), .ZN(n3388)
         );
  AOI222_X1 U3319 ( .A1(n11320), .A2(n12831), .B1(n11317), .B2(n12863), .C1(
        n11314), .C2(n12927), .ZN(n3385) );
  NAND4_X1 U3320 ( .A1(n4777), .A2(n4778), .A3(n4779), .A4(n4780), .ZN(n4776)
         );
  AOI221_X1 U3321 ( .B1(n11080), .B2(n12798), .C1(n11077), .C2(n12990), .A(
        n4785), .ZN(n4779) );
  NOR4_X1 U3322 ( .A1(n4781), .A2(n4782), .A3(n4783), .A4(n4784), .ZN(n4780)
         );
  AOI222_X1 U3323 ( .A1(n11056), .A2(n12830), .B1(n11053), .B2(n12862), .C1(
        n11050), .C2(n12926), .ZN(n4777) );
  NAND4_X1 U3324 ( .A1(n3344), .A2(n3345), .A3(n3346), .A4(n3347), .ZN(n3343)
         );
  AOI221_X1 U3325 ( .B1(n11344), .B2(n12798), .C1(n11341), .C2(n12990), .A(
        n3352), .ZN(n3346) );
  NOR4_X1 U3326 ( .A1(n3348), .A2(n3349), .A3(n3350), .A4(n3351), .ZN(n3347)
         );
  AOI222_X1 U3327 ( .A1(n11320), .A2(n12830), .B1(n11317), .B2(n12862), .C1(
        n11314), .C2(n12926), .ZN(n3344) );
  NAND4_X1 U3328 ( .A1(n4736), .A2(n4737), .A3(n4738), .A4(n4739), .ZN(n4735)
         );
  AOI221_X1 U3329 ( .B1(n11080), .B2(n12797), .C1(n11077), .C2(n12989), .A(
        n4744), .ZN(n4738) );
  NOR4_X1 U3330 ( .A1(n4740), .A2(n4741), .A3(n4742), .A4(n4743), .ZN(n4739)
         );
  AOI222_X1 U3331 ( .A1(n11056), .A2(n12829), .B1(n11053), .B2(n12861), .C1(
        n11050), .C2(n12925), .ZN(n4736) );
  NAND4_X1 U3332 ( .A1(n3303), .A2(n3304), .A3(n3305), .A4(n3306), .ZN(n3302)
         );
  AOI221_X1 U3333 ( .B1(n11344), .B2(n12797), .C1(n11341), .C2(n12989), .A(
        n3311), .ZN(n3305) );
  NOR4_X1 U3334 ( .A1(n3307), .A2(n3308), .A3(n3309), .A4(n3310), .ZN(n3306)
         );
  AOI222_X1 U3335 ( .A1(n11320), .A2(n12829), .B1(n11317), .B2(n12861), .C1(
        n11314), .C2(n12925), .ZN(n3303) );
  NAND4_X1 U3336 ( .A1(n4695), .A2(n4696), .A3(n4697), .A4(n4698), .ZN(n4694)
         );
  AOI221_X1 U3337 ( .B1(n11080), .B2(n12796), .C1(n11077), .C2(n12988), .A(
        n4703), .ZN(n4697) );
  NOR4_X1 U3338 ( .A1(n4699), .A2(n4700), .A3(n4701), .A4(n4702), .ZN(n4698)
         );
  AOI222_X1 U3339 ( .A1(n11056), .A2(n12828), .B1(n11053), .B2(n12860), .C1(
        n11050), .C2(n12924), .ZN(n4695) );
  NAND4_X1 U3340 ( .A1(n3262), .A2(n3263), .A3(n3264), .A4(n3265), .ZN(n3261)
         );
  AOI221_X1 U3341 ( .B1(n11344), .B2(n12796), .C1(n11341), .C2(n12988), .A(
        n3270), .ZN(n3264) );
  NOR4_X1 U3342 ( .A1(n3266), .A2(n3267), .A3(n3268), .A4(n3269), .ZN(n3265)
         );
  AOI222_X1 U3343 ( .A1(n11320), .A2(n12828), .B1(n11317), .B2(n12860), .C1(
        n11314), .C2(n12924), .ZN(n3262) );
  NAND4_X1 U3344 ( .A1(n4654), .A2(n4655), .A3(n4656), .A4(n4657), .ZN(n4653)
         );
  AOI221_X1 U3345 ( .B1(n11081), .B2(n12795), .C1(n11078), .C2(n12987), .A(
        n4662), .ZN(n4656) );
  NOR4_X1 U3346 ( .A1(n4658), .A2(n4659), .A3(n4660), .A4(n4661), .ZN(n4657)
         );
  AOI222_X1 U3347 ( .A1(n11057), .A2(n12827), .B1(n11054), .B2(n12859), .C1(
        n11051), .C2(n12923), .ZN(n4654) );
  NAND4_X1 U3348 ( .A1(n3221), .A2(n3222), .A3(n3223), .A4(n3224), .ZN(n3220)
         );
  AOI221_X1 U3349 ( .B1(n11345), .B2(n12795), .C1(n11342), .C2(n12987), .A(
        n3229), .ZN(n3223) );
  NOR4_X1 U3350 ( .A1(n3225), .A2(n3226), .A3(n3227), .A4(n3228), .ZN(n3224)
         );
  AOI222_X1 U3351 ( .A1(n11321), .A2(n12827), .B1(n11318), .B2(n12859), .C1(
        n11315), .C2(n12923), .ZN(n3221) );
  NAND4_X1 U3352 ( .A1(n4613), .A2(n4614), .A3(n4615), .A4(n4616), .ZN(n4612)
         );
  AOI221_X1 U3353 ( .B1(n11081), .B2(n12794), .C1(n11078), .C2(n12986), .A(
        n4621), .ZN(n4615) );
  NOR4_X1 U3354 ( .A1(n4617), .A2(n4618), .A3(n4619), .A4(n4620), .ZN(n4616)
         );
  AOI222_X1 U3355 ( .A1(n11057), .A2(n12826), .B1(n11054), .B2(n12858), .C1(
        n11051), .C2(n12922), .ZN(n4613) );
  NAND4_X1 U3356 ( .A1(n3180), .A2(n3181), .A3(n3182), .A4(n3183), .ZN(n3179)
         );
  AOI221_X1 U3357 ( .B1(n11345), .B2(n12794), .C1(n11342), .C2(n12986), .A(
        n3188), .ZN(n3182) );
  NOR4_X1 U3358 ( .A1(n3184), .A2(n3185), .A3(n3186), .A4(n3187), .ZN(n3183)
         );
  AOI222_X1 U3359 ( .A1(n11321), .A2(n12826), .B1(n11318), .B2(n12858), .C1(
        n11315), .C2(n12922), .ZN(n3180) );
  NAND4_X1 U3360 ( .A1(n4572), .A2(n4573), .A3(n4574), .A4(n4575), .ZN(n4571)
         );
  AOI221_X1 U3361 ( .B1(n11081), .B2(n12793), .C1(n11078), .C2(n12985), .A(
        n4580), .ZN(n4574) );
  NOR4_X1 U3362 ( .A1(n4576), .A2(n4577), .A3(n4578), .A4(n4579), .ZN(n4575)
         );
  AOI222_X1 U3363 ( .A1(n11057), .A2(n12825), .B1(n11054), .B2(n12857), .C1(
        n11051), .C2(n12921), .ZN(n4572) );
  NAND4_X1 U3364 ( .A1(n3139), .A2(n3140), .A3(n3141), .A4(n3142), .ZN(n3138)
         );
  AOI221_X1 U3365 ( .B1(n11345), .B2(n12793), .C1(n11342), .C2(n12985), .A(
        n3147), .ZN(n3141) );
  NOR4_X1 U3366 ( .A1(n3143), .A2(n3144), .A3(n3145), .A4(n3146), .ZN(n3142)
         );
  AOI222_X1 U3367 ( .A1(n11321), .A2(n12825), .B1(n11318), .B2(n12857), .C1(
        n11315), .C2(n12921), .ZN(n3139) );
  NAND4_X1 U3368 ( .A1(n4531), .A2(n4532), .A3(n4533), .A4(n4534), .ZN(n4530)
         );
  AOI221_X1 U3369 ( .B1(n11081), .B2(n12792), .C1(n11078), .C2(n12984), .A(
        n4539), .ZN(n4533) );
  NOR4_X1 U3370 ( .A1(n4535), .A2(n4536), .A3(n4537), .A4(n4538), .ZN(n4534)
         );
  AOI222_X1 U3371 ( .A1(n11057), .A2(n12824), .B1(n11054), .B2(n12856), .C1(
        n11051), .C2(n12920), .ZN(n4531) );
  NAND4_X1 U3372 ( .A1(n3098), .A2(n3099), .A3(n3100), .A4(n3101), .ZN(n3097)
         );
  AOI221_X1 U3373 ( .B1(n11345), .B2(n12792), .C1(n11342), .C2(n12984), .A(
        n3106), .ZN(n3100) );
  NOR4_X1 U3374 ( .A1(n3102), .A2(n3103), .A3(n3104), .A4(n3105), .ZN(n3101)
         );
  AOI222_X1 U3375 ( .A1(n11321), .A2(n12824), .B1(n11318), .B2(n12856), .C1(
        n11315), .C2(n12920), .ZN(n3098) );
  NAND4_X1 U3376 ( .A1(n4490), .A2(n4491), .A3(n4492), .A4(n4493), .ZN(n4489)
         );
  AOI221_X1 U3377 ( .B1(n11081), .B2(n12791), .C1(n11078), .C2(n12983), .A(
        n4498), .ZN(n4492) );
  NOR4_X1 U3378 ( .A1(n4494), .A2(n4495), .A3(n4496), .A4(n4497), .ZN(n4493)
         );
  AOI222_X1 U3379 ( .A1(n11057), .A2(n12823), .B1(n11054), .B2(n12855), .C1(
        n11051), .C2(n12919), .ZN(n4490) );
  NAND4_X1 U3380 ( .A1(n3057), .A2(n3058), .A3(n3059), .A4(n3060), .ZN(n3056)
         );
  AOI221_X1 U3381 ( .B1(n11345), .B2(n12791), .C1(n11342), .C2(n12983), .A(
        n3065), .ZN(n3059) );
  NOR4_X1 U3382 ( .A1(n3061), .A2(n3062), .A3(n3063), .A4(n3064), .ZN(n3060)
         );
  AOI222_X1 U3383 ( .A1(n11321), .A2(n12823), .B1(n11318), .B2(n12855), .C1(
        n11315), .C2(n12919), .ZN(n3057) );
  NAND4_X1 U3384 ( .A1(n4449), .A2(n4450), .A3(n4451), .A4(n4452), .ZN(n4448)
         );
  AOI221_X1 U3385 ( .B1(n11081), .B2(n12790), .C1(n11078), .C2(n12982), .A(
        n4457), .ZN(n4451) );
  NOR4_X1 U3386 ( .A1(n4453), .A2(n4454), .A3(n4455), .A4(n4456), .ZN(n4452)
         );
  AOI222_X1 U3387 ( .A1(n11057), .A2(n12822), .B1(n11054), .B2(n12854), .C1(
        n11051), .C2(n12918), .ZN(n4449) );
  NAND4_X1 U3388 ( .A1(n3016), .A2(n3017), .A3(n3018), .A4(n3019), .ZN(n3015)
         );
  AOI221_X1 U3389 ( .B1(n11345), .B2(n12790), .C1(n11342), .C2(n12982), .A(
        n3024), .ZN(n3018) );
  NOR4_X1 U3390 ( .A1(n3020), .A2(n3021), .A3(n3022), .A4(n3023), .ZN(n3019)
         );
  AOI222_X1 U3391 ( .A1(n11321), .A2(n12822), .B1(n11318), .B2(n12854), .C1(
        n11315), .C2(n12918), .ZN(n3016) );
  NAND4_X1 U3392 ( .A1(n4408), .A2(n4409), .A3(n4410), .A4(n4411), .ZN(n4407)
         );
  AOI221_X1 U3393 ( .B1(n11081), .B2(n12789), .C1(n11078), .C2(n12981), .A(
        n4416), .ZN(n4410) );
  NOR4_X1 U3394 ( .A1(n4412), .A2(n4413), .A3(n4414), .A4(n4415), .ZN(n4411)
         );
  AOI222_X1 U3395 ( .A1(n11057), .A2(n12821), .B1(n11054), .B2(n12853), .C1(
        n11051), .C2(n12917), .ZN(n4408) );
  NAND4_X1 U3396 ( .A1(n2975), .A2(n2976), .A3(n2977), .A4(n2978), .ZN(n2974)
         );
  AOI221_X1 U3397 ( .B1(n11345), .B2(n12789), .C1(n11342), .C2(n12981), .A(
        n2983), .ZN(n2977) );
  NOR4_X1 U3398 ( .A1(n2979), .A2(n2980), .A3(n2981), .A4(n2982), .ZN(n2978)
         );
  AOI222_X1 U3399 ( .A1(n11321), .A2(n12821), .B1(n11318), .B2(n12853), .C1(
        n11315), .C2(n12917), .ZN(n2975) );
  NAND4_X1 U3400 ( .A1(n4279), .A2(n4280), .A3(n4281), .A4(n4282), .ZN(n4278)
         );
  AOI221_X1 U3401 ( .B1(n11081), .B2(n12788), .C1(n11078), .C2(n12980), .A(
        n4300), .ZN(n4281) );
  NOR4_X1 U3402 ( .A1(n4283), .A2(n4284), .A3(n4285), .A4(n4286), .ZN(n4282)
         );
  AOI222_X1 U3403 ( .A1(n11057), .A2(n12820), .B1(n11054), .B2(n12852), .C1(
        n11051), .C2(n12916), .ZN(n4279) );
  NAND4_X1 U3404 ( .A1(n2747), .A2(n2748), .A3(n2749), .A4(n2750), .ZN(n2746)
         );
  AOI221_X1 U3405 ( .B1(n11345), .B2(n12788), .C1(n11342), .C2(n12980), .A(
        n2800), .ZN(n2749) );
  NOR4_X1 U3406 ( .A1(n2751), .A2(n2752), .A3(n2753), .A4(n2786), .ZN(n2750)
         );
  AOI222_X1 U3407 ( .A1(n11321), .A2(n12820), .B1(n11318), .B2(n12852), .C1(
        n11315), .C2(n12916), .ZN(n2747) );
  AND2_X1 U3408 ( .A1(n5650), .A2(n5703), .ZN(n5659) );
  AND2_X1 U3409 ( .A1(n4217), .A2(n4270), .ZN(n4226) );
  AND2_X1 U3410 ( .A1(n5649), .A2(n5702), .ZN(n5663) );
  AND2_X1 U3411 ( .A1(n4216), .A2(n4269), .ZN(n4230) );
  AND2_X1 U3412 ( .A1(n5651), .A2(n5702), .ZN(n5665) );
  AND2_X1 U3413 ( .A1(n4218), .A2(n4269), .ZN(n4232) );
  AND2_X1 U3414 ( .A1(n5652), .A2(n5654), .ZN(n5648) );
  AND2_X1 U3415 ( .A1(n4219), .A2(n4221), .ZN(n4215) );
  AND2_X1 U3416 ( .A1(n5702), .A2(n5650), .ZN(n5660) );
  AND2_X1 U3417 ( .A1(n4269), .A2(n4217), .ZN(n4227) );
  NAND2_X1 U3418 ( .A1(n5705), .A2(n5647), .ZN(n4394) );
  NAND2_X1 U3419 ( .A1(n4272), .A2(n4214), .ZN(n2961) );
  AND2_X1 U3420 ( .A1(n5654), .A2(n5701), .ZN(n5688) );
  AND2_X1 U3421 ( .A1(n4221), .A2(n4268), .ZN(n4255) );
  NOR2_X1 U3422 ( .A1(n12769), .A2(N8435), .ZN(n5701) );
  NOR2_X1 U3423 ( .A1(n12773), .A2(N8579), .ZN(n4268) );
  AND2_X1 U3424 ( .A1(n5675), .A2(n5654), .ZN(n5676) );
  AND2_X1 U3425 ( .A1(n4242), .A2(n4221), .ZN(n4243) );
  INV_X1 U3426 ( .A(N2171), .ZN(n12733) );
  NAND2_X1 U3427 ( .A1(n5648), .A2(n5647), .ZN(n4287) );
  NAND2_X1 U3428 ( .A1(n5646), .A2(n5647), .ZN(n4288) );
  NAND2_X1 U3429 ( .A1(n5674), .A2(n5647), .ZN(n4319) );
  NAND2_X1 U3430 ( .A1(n5690), .A2(n5647), .ZN(n4357) );
  NAND2_X1 U3431 ( .A1(n5688), .A2(n5647), .ZN(n4349) );
  NAND2_X1 U3432 ( .A1(n5692), .A2(n5647), .ZN(n4364) );
  NAND2_X1 U3433 ( .A1(n4215), .A2(n4214), .ZN(n2787) );
  NAND2_X1 U3434 ( .A1(n4213), .A2(n4214), .ZN(n2788) );
  NAND2_X1 U3435 ( .A1(n4241), .A2(n4214), .ZN(n2851) );
  NAND2_X1 U3436 ( .A1(n4257), .A2(n4214), .ZN(n2921) );
  NAND2_X1 U3437 ( .A1(n4255), .A2(n4214), .ZN(n2881) );
  NAND2_X1 U3438 ( .A1(n4259), .A2(n4214), .ZN(n2928) );
  BUF_X1 U3439 ( .A(N8735), .Z(n12427) );
  BUF_X1 U3440 ( .A(N8702), .Z(n12430) );
  BUF_X1 U3441 ( .A(N8702), .Z(n12429) );
  BUF_X1 U3442 ( .A(N8735), .Z(n12426) );
  NAND2_X1 U3443 ( .A1(n5648), .A2(n5649), .ZN(n4291) );
  NAND2_X1 U3444 ( .A1(n5646), .A2(n5649), .ZN(n4289) );
  NAND2_X1 U3445 ( .A1(n5676), .A2(n5649), .ZN(n4322) );
  NAND2_X1 U3446 ( .A1(n5674), .A2(n5649), .ZN(n4321) );
  NAND2_X1 U3447 ( .A1(n5688), .A2(n5649), .ZN(n4380) );
  NAND2_X1 U3448 ( .A1(n5690), .A2(n5649), .ZN(n4381) );
  NAND2_X1 U3449 ( .A1(n4215), .A2(n4216), .ZN(n2791) );
  NAND2_X1 U3450 ( .A1(n4213), .A2(n4216), .ZN(n2789) );
  NAND2_X1 U3451 ( .A1(n4243), .A2(n4216), .ZN(n2854) );
  NAND2_X1 U3452 ( .A1(n4241), .A2(n4216), .ZN(n2853) );
  NAND2_X1 U3453 ( .A1(n4255), .A2(n4216), .ZN(n2947) );
  NAND2_X1 U3454 ( .A1(n4257), .A2(n4216), .ZN(n2948) );
  INV_X1 U3455 ( .A(N8434), .ZN(n12772) );
  INV_X1 U3456 ( .A(N8578), .ZN(n12776) );
  BUF_X1 U3457 ( .A(N8702), .Z(n12431) );
  BUF_X1 U3458 ( .A(N8735), .Z(n12428) );
  NAND2_X1 U3459 ( .A1(n5648), .A2(n5651), .ZN(n4292) );
  NAND2_X1 U3460 ( .A1(n5646), .A2(n5651), .ZN(n4293) );
  NAND2_X1 U3461 ( .A1(n5676), .A2(n5651), .ZN(n4324) );
  NAND2_X1 U3462 ( .A1(n5674), .A2(n5651), .ZN(n4327) );
  NAND2_X1 U3463 ( .A1(n5687), .A2(n5651), .ZN(n4350) );
  NAND2_X1 U3464 ( .A1(n5688), .A2(n5651), .ZN(n4383) );
  NAND2_X1 U3465 ( .A1(n4215), .A2(n4218), .ZN(n2792) );
  NAND2_X1 U3466 ( .A1(n4213), .A2(n4218), .ZN(n2793) );
  NAND2_X1 U3467 ( .A1(n4243), .A2(n4218), .ZN(n2856) );
  NAND2_X1 U3468 ( .A1(n4241), .A2(n4218), .ZN(n2859) );
  NAND2_X1 U3469 ( .A1(n4254), .A2(n4218), .ZN(n2914) );
  NAND2_X1 U3470 ( .A1(n4255), .A2(n4218), .ZN(n2950) );
  NAND2_X1 U3471 ( .A1(n5648), .A2(n5650), .ZN(n4290) );
  NAND2_X1 U3472 ( .A1(n5646), .A2(n5650), .ZN(n4294) );
  NAND2_X1 U3473 ( .A1(n5676), .A2(n5650), .ZN(n4320) );
  NAND2_X1 U3474 ( .A1(n5674), .A2(n5650), .ZN(n4325) );
  NAND2_X1 U3475 ( .A1(n5688), .A2(n5650), .ZN(n4384) );
  NAND2_X1 U3476 ( .A1(n5690), .A2(n5650), .ZN(n4382) );
  NAND2_X1 U3477 ( .A1(n4215), .A2(n4217), .ZN(n2790) );
  NAND2_X1 U3478 ( .A1(n4213), .A2(n4217), .ZN(n2794) );
  NAND2_X1 U3479 ( .A1(n4243), .A2(n4217), .ZN(n2852) );
  NAND2_X1 U3480 ( .A1(n4241), .A2(n4217), .ZN(n2857) );
  NAND2_X1 U3481 ( .A1(n4255), .A2(n4217), .ZN(n2951) );
  NAND2_X1 U3482 ( .A1(n4257), .A2(n4217), .ZN(n2949) );
  AND2_X1 U3483 ( .A1(n5660), .A2(N8437), .ZN(n4391) );
  AND2_X1 U3484 ( .A1(n4227), .A2(N8581), .ZN(n2958) );
  NAND2_X1 U3485 ( .A1(n5651), .A2(n5690), .ZN(n4387) );
  NAND2_X1 U3486 ( .A1(n4218), .A2(n4257), .ZN(n2954) );
  AND3_X1 U3487 ( .A1(n5654), .A2(n12769), .A3(n5678), .ZN(n5662) );
  AND3_X1 U3488 ( .A1(n4221), .A2(n12773), .A3(n4245), .ZN(n4229) );
  AND2_X1 U3489 ( .A1(n5689), .A2(n5654), .ZN(n5692) );
  AND2_X1 U3490 ( .A1(n4256), .A2(n4221), .ZN(n4259) );
  AND2_X1 U3491 ( .A1(n5705), .A2(n5651), .ZN(n4392) );
  AND2_X1 U3492 ( .A1(n4272), .A2(n4218), .ZN(n2959) );
  AND2_X1 U3493 ( .A1(n5687), .A2(n5647), .ZN(n4369) );
  AND2_X1 U3494 ( .A1(n5706), .A2(n5647), .ZN(n4400) );
  AND2_X1 U3495 ( .A1(n4254), .A2(n4214), .ZN(n2933) );
  AND2_X1 U3496 ( .A1(n4273), .A2(n4214), .ZN(n2967) );
  AND2_X1 U3497 ( .A1(n5664), .A2(n5649), .ZN(n4304) );
  AND2_X1 U3498 ( .A1(n4231), .A2(n4216), .ZN(n2804) );
  AND2_X1 U3499 ( .A1(n5706), .A2(n5650), .ZN(n4397) );
  AND2_X1 U3500 ( .A1(n4273), .A2(n4217), .ZN(n2964) );
  AND2_X1 U3501 ( .A1(n5664), .A2(n5651), .ZN(n4329) );
  AND2_X1 U3502 ( .A1(n5662), .A2(n5651), .ZN(n4330) );
  AND2_X1 U3503 ( .A1(n4231), .A2(n4218), .ZN(n2861) );
  AND2_X1 U3504 ( .A1(n4229), .A2(n4218), .ZN(n2862) );
  AND2_X1 U3505 ( .A1(n5662), .A2(n5650), .ZN(n4299) );
  AND2_X1 U3506 ( .A1(n5692), .A2(n5650), .ZN(n4366) );
  AND2_X1 U3507 ( .A1(n4229), .A2(n4217), .ZN(n2799) );
  AND2_X1 U3508 ( .A1(n4259), .A2(n4217), .ZN(n2930) );
  AND2_X1 U3509 ( .A1(N2170), .A2(n12734), .ZN(n2725) );
  BUF_X1 U3510 ( .A(RESET), .Z(n12432) );
  INV_X1 U3511 ( .A(n2740), .ZN(\r480/A[3] ) );
  INV_X1 U3512 ( .A(n2739), .ZN(\r486/A[3] ) );
  INV_X1 U3513 ( .A(n2741), .ZN(\r472/B[3] ) );
  AND2_X1 U3514 ( .A1(n5705), .A2(n5649), .ZN(n4401) );
  AND2_X1 U3515 ( .A1(n5705), .A2(n5650), .ZN(n4402) );
  AND2_X1 U3516 ( .A1(n4272), .A2(n4216), .ZN(n2968) );
  AND2_X1 U3517 ( .A1(n4272), .A2(n4217), .ZN(n2969) );
  AND2_X1 U3518 ( .A1(n5664), .A2(n5647), .ZN(n4305) );
  AND2_X1 U3519 ( .A1(n5662), .A2(n5647), .ZN(n4308) );
  AND2_X1 U3520 ( .A1(n5676), .A2(n5647), .ZN(n4336) );
  AND2_X1 U3521 ( .A1(n4231), .A2(n4214), .ZN(n2805) );
  AND2_X1 U3522 ( .A1(n4229), .A2(n4214), .ZN(n2808) );
  AND2_X1 U3523 ( .A1(n4243), .A2(n4214), .ZN(n2868) );
  AND2_X1 U3524 ( .A1(n5706), .A2(n5649), .ZN(n4398) );
  AND2_X1 U3525 ( .A1(n5706), .A2(n5651), .ZN(n4399) );
  AND2_X1 U3526 ( .A1(n4273), .A2(n4216), .ZN(n2965) );
  AND2_X1 U3527 ( .A1(n4273), .A2(n4218), .ZN(n2966) );
  AND2_X1 U3528 ( .A1(n5662), .A2(n5649), .ZN(n4309) );
  AND2_X1 U3529 ( .A1(n5687), .A2(n5649), .ZN(n4370) );
  AND2_X1 U3530 ( .A1(n5692), .A2(n5649), .ZN(n4371) );
  AND2_X1 U3531 ( .A1(n4229), .A2(n4216), .ZN(n2809) );
  AND2_X1 U3532 ( .A1(n4254), .A2(n4216), .ZN(n2934) );
  AND2_X1 U3533 ( .A1(n4259), .A2(n4216), .ZN(n2938) );
  AND2_X1 U3534 ( .A1(n5692), .A2(n5651), .ZN(n4367) );
  AND2_X1 U3535 ( .A1(n4259), .A2(n4218), .ZN(n2931) );
  AND2_X1 U3536 ( .A1(n5664), .A2(n5650), .ZN(n4306) );
  AND2_X1 U3537 ( .A1(n5687), .A2(n5650), .ZN(n4368) );
  AND2_X1 U3538 ( .A1(n4231), .A2(n4217), .ZN(n2806) );
  AND2_X1 U3539 ( .A1(n4254), .A2(n4217), .ZN(n2932) );
  NOR2_X1 U3540 ( .A1(n5633), .A2(n12663), .ZN(N8703) );
  NOR4_X1 U3541 ( .A1(n5634), .A2(n5635), .A3(n5636), .A4(n5637), .ZN(n5633)
         );
  NAND4_X1 U3542 ( .A1(n5693), .A2(n5694), .A3(n5695), .A4(n5696), .ZN(n5634)
         );
  NAND4_X1 U3543 ( .A1(n5679), .A2(n5680), .A3(n5681), .A4(n5682), .ZN(n5635)
         );
  NOR2_X1 U3544 ( .A1(n4200), .A2(n12671), .ZN(N8736) );
  NOR4_X1 U3545 ( .A1(n4201), .A2(n4202), .A3(n4203), .A4(n4204), .ZN(n4200)
         );
  NAND4_X1 U3546 ( .A1(n4260), .A2(n4261), .A3(n4262), .A4(n4263), .ZN(n4201)
         );
  NAND4_X1 U3547 ( .A1(n4246), .A2(n4247), .A3(n4248), .A4(n4249), .ZN(n4202)
         );
  NOR2_X1 U3548 ( .A1(n5592), .A2(n12663), .ZN(N8704) );
  NOR4_X1 U3549 ( .A1(n5593), .A2(n5594), .A3(n5595), .A4(n5596), .ZN(n5592)
         );
  NAND4_X1 U3550 ( .A1(n5624), .A2(n5625), .A3(n5626), .A4(n5627), .ZN(n5593)
         );
  NAND4_X1 U3551 ( .A1(n5615), .A2(n5616), .A3(n5617), .A4(n5618), .ZN(n5594)
         );
  NOR2_X1 U3552 ( .A1(n4159), .A2(n12671), .ZN(N8737) );
  NOR4_X1 U3553 ( .A1(n4160), .A2(n4161), .A3(n4162), .A4(n4163), .ZN(n4159)
         );
  NAND4_X1 U3554 ( .A1(n4191), .A2(n4192), .A3(n4193), .A4(n4194), .ZN(n4160)
         );
  NAND4_X1 U3555 ( .A1(n4182), .A2(n4183), .A3(n4184), .A4(n4185), .ZN(n4161)
         );
  NOR2_X1 U3556 ( .A1(n5551), .A2(n12663), .ZN(N8705) );
  NOR4_X1 U3557 ( .A1(n5552), .A2(n5553), .A3(n5554), .A4(n5555), .ZN(n5551)
         );
  NAND4_X1 U3558 ( .A1(n5583), .A2(n5584), .A3(n5585), .A4(n5586), .ZN(n5552)
         );
  NAND4_X1 U3559 ( .A1(n5574), .A2(n5575), .A3(n5576), .A4(n5577), .ZN(n5553)
         );
  NOR2_X1 U3560 ( .A1(n4118), .A2(n12671), .ZN(N8738) );
  NOR4_X1 U3561 ( .A1(n4119), .A2(n4120), .A3(n4121), .A4(n4122), .ZN(n4118)
         );
  NAND4_X1 U3562 ( .A1(n4150), .A2(n4151), .A3(n4152), .A4(n4153), .ZN(n4119)
         );
  NAND4_X1 U3563 ( .A1(n4141), .A2(n4142), .A3(n4143), .A4(n4144), .ZN(n4120)
         );
  NOR2_X1 U3564 ( .A1(n5510), .A2(n12663), .ZN(N8706) );
  NOR4_X1 U3565 ( .A1(n5511), .A2(n5512), .A3(n5513), .A4(n5514), .ZN(n5510)
         );
  NAND4_X1 U3566 ( .A1(n5542), .A2(n5543), .A3(n5544), .A4(n5545), .ZN(n5511)
         );
  NAND4_X1 U3567 ( .A1(n5533), .A2(n5534), .A3(n5535), .A4(n5536), .ZN(n5512)
         );
  NOR2_X1 U3568 ( .A1(n4077), .A2(n12672), .ZN(N8739) );
  NOR4_X1 U3569 ( .A1(n4078), .A2(n4079), .A3(n4080), .A4(n4081), .ZN(n4077)
         );
  NAND4_X1 U3570 ( .A1(n4109), .A2(n4110), .A3(n4111), .A4(n4112), .ZN(n4078)
         );
  NAND4_X1 U3571 ( .A1(n4100), .A2(n4101), .A3(n4102), .A4(n4103), .ZN(n4079)
         );
  NOR2_X1 U3572 ( .A1(n5469), .A2(n12664), .ZN(N8707) );
  NOR4_X1 U3573 ( .A1(n5470), .A2(n5471), .A3(n5472), .A4(n5473), .ZN(n5469)
         );
  NAND4_X1 U3574 ( .A1(n5501), .A2(n5502), .A3(n5503), .A4(n5504), .ZN(n5470)
         );
  NAND4_X1 U3575 ( .A1(n5492), .A2(n5493), .A3(n5494), .A4(n5495), .ZN(n5471)
         );
  NOR2_X1 U3576 ( .A1(n4036), .A2(n12672), .ZN(N8740) );
  NOR4_X1 U3577 ( .A1(n4037), .A2(n4038), .A3(n4039), .A4(n4040), .ZN(n4036)
         );
  NAND4_X1 U3578 ( .A1(n4068), .A2(n4069), .A3(n4070), .A4(n4071), .ZN(n4037)
         );
  NAND4_X1 U3579 ( .A1(n4059), .A2(n4060), .A3(n4061), .A4(n4062), .ZN(n4038)
         );
  NOR2_X1 U3580 ( .A1(n5428), .A2(n12664), .ZN(N8708) );
  NOR4_X1 U3581 ( .A1(n5429), .A2(n5430), .A3(n5431), .A4(n5432), .ZN(n5428)
         );
  NAND4_X1 U3582 ( .A1(n5460), .A2(n5461), .A3(n5462), .A4(n5463), .ZN(n5429)
         );
  NAND4_X1 U3583 ( .A1(n5451), .A2(n5452), .A3(n5453), .A4(n5454), .ZN(n5430)
         );
  NOR2_X1 U3584 ( .A1(n3995), .A2(n12672), .ZN(N8741) );
  NOR4_X1 U3585 ( .A1(n3996), .A2(n3997), .A3(n3998), .A4(n3999), .ZN(n3995)
         );
  NAND4_X1 U3586 ( .A1(n4027), .A2(n4028), .A3(n4029), .A4(n4030), .ZN(n3996)
         );
  NAND4_X1 U3587 ( .A1(n4018), .A2(n4019), .A3(n4020), .A4(n4021), .ZN(n3997)
         );
  NOR2_X1 U3588 ( .A1(n5387), .A2(n12664), .ZN(N8709) );
  NOR4_X1 U3589 ( .A1(n5388), .A2(n5389), .A3(n5390), .A4(n5391), .ZN(n5387)
         );
  NAND4_X1 U3590 ( .A1(n5419), .A2(n5420), .A3(n5421), .A4(n5422), .ZN(n5388)
         );
  NAND4_X1 U3591 ( .A1(n5410), .A2(n5411), .A3(n5412), .A4(n5413), .ZN(n5389)
         );
  NOR2_X1 U3592 ( .A1(n3954), .A2(n12672), .ZN(N8742) );
  NOR4_X1 U3593 ( .A1(n3955), .A2(n3956), .A3(n3957), .A4(n3958), .ZN(n3954)
         );
  NAND4_X1 U3594 ( .A1(n3986), .A2(n3987), .A3(n3988), .A4(n3989), .ZN(n3955)
         );
  NAND4_X1 U3595 ( .A1(n3977), .A2(n3978), .A3(n3979), .A4(n3980), .ZN(n3956)
         );
  NOR2_X1 U3596 ( .A1(n5346), .A2(n12664), .ZN(N8710) );
  NOR4_X1 U3597 ( .A1(n5347), .A2(n5348), .A3(n5349), .A4(n5350), .ZN(n5346)
         );
  NAND4_X1 U3598 ( .A1(n5378), .A2(n5379), .A3(n5380), .A4(n5381), .ZN(n5347)
         );
  NAND4_X1 U3599 ( .A1(n5369), .A2(n5370), .A3(n5371), .A4(n5372), .ZN(n5348)
         );
  NOR2_X1 U3600 ( .A1(n3913), .A2(n12673), .ZN(N8743) );
  NOR4_X1 U3601 ( .A1(n3914), .A2(n3915), .A3(n3916), .A4(n3917), .ZN(n3913)
         );
  NAND4_X1 U3602 ( .A1(n3945), .A2(n3946), .A3(n3947), .A4(n3948), .ZN(n3914)
         );
  NAND4_X1 U3603 ( .A1(n3936), .A2(n3937), .A3(n3938), .A4(n3939), .ZN(n3915)
         );
  NOR2_X1 U3604 ( .A1(n5305), .A2(n12665), .ZN(N8711) );
  NOR4_X1 U3605 ( .A1(n5306), .A2(n5307), .A3(n5308), .A4(n5309), .ZN(n5305)
         );
  NAND4_X1 U3606 ( .A1(n5337), .A2(n5338), .A3(n5339), .A4(n5340), .ZN(n5306)
         );
  NAND4_X1 U3607 ( .A1(n5328), .A2(n5329), .A3(n5330), .A4(n5331), .ZN(n5307)
         );
  NOR2_X1 U3608 ( .A1(n3872), .A2(n12673), .ZN(N8744) );
  NOR4_X1 U3609 ( .A1(n3873), .A2(n3874), .A3(n3875), .A4(n3876), .ZN(n3872)
         );
  NAND4_X1 U3610 ( .A1(n3904), .A2(n3905), .A3(n3906), .A4(n3907), .ZN(n3873)
         );
  NAND4_X1 U3611 ( .A1(n3895), .A2(n3896), .A3(n3897), .A4(n3898), .ZN(n3874)
         );
  NOR2_X1 U3612 ( .A1(n5264), .A2(n12665), .ZN(N8712) );
  NOR4_X1 U3613 ( .A1(n5265), .A2(n5266), .A3(n5267), .A4(n5268), .ZN(n5264)
         );
  NAND4_X1 U3614 ( .A1(n5296), .A2(n5297), .A3(n5298), .A4(n5299), .ZN(n5265)
         );
  NAND4_X1 U3615 ( .A1(n5287), .A2(n5288), .A3(n5289), .A4(n5290), .ZN(n5266)
         );
  NOR2_X1 U3616 ( .A1(n3831), .A2(n12673), .ZN(N8745) );
  NOR4_X1 U3617 ( .A1(n3832), .A2(n3833), .A3(n3834), .A4(n3835), .ZN(n3831)
         );
  NAND4_X1 U3618 ( .A1(n3863), .A2(n3864), .A3(n3865), .A4(n3866), .ZN(n3832)
         );
  NAND4_X1 U3619 ( .A1(n3854), .A2(n3855), .A3(n3856), .A4(n3857), .ZN(n3833)
         );
  NOR2_X1 U3620 ( .A1(n5223), .A2(n12665), .ZN(N8713) );
  NOR4_X1 U3621 ( .A1(n5224), .A2(n5225), .A3(n5226), .A4(n5227), .ZN(n5223)
         );
  NAND4_X1 U3622 ( .A1(n5255), .A2(n5256), .A3(n5257), .A4(n5258), .ZN(n5224)
         );
  NAND4_X1 U3623 ( .A1(n5246), .A2(n5247), .A3(n5248), .A4(n5249), .ZN(n5225)
         );
  NOR2_X1 U3624 ( .A1(n3790), .A2(n12673), .ZN(N8746) );
  NOR4_X1 U3625 ( .A1(n3791), .A2(n3792), .A3(n3793), .A4(n3794), .ZN(n3790)
         );
  NAND4_X1 U3626 ( .A1(n3822), .A2(n3823), .A3(n3824), .A4(n3825), .ZN(n3791)
         );
  NAND4_X1 U3627 ( .A1(n3813), .A2(n3814), .A3(n3815), .A4(n3816), .ZN(n3792)
         );
  NOR2_X1 U3628 ( .A1(n5182), .A2(n12665), .ZN(N8714) );
  NOR4_X1 U3629 ( .A1(n5183), .A2(n5184), .A3(n5185), .A4(n5186), .ZN(n5182)
         );
  NAND4_X1 U3630 ( .A1(n5214), .A2(n5215), .A3(n5216), .A4(n5217), .ZN(n5183)
         );
  NAND4_X1 U3631 ( .A1(n5205), .A2(n5206), .A3(n5207), .A4(n5208), .ZN(n5184)
         );
  NOR2_X1 U3632 ( .A1(n3749), .A2(n12674), .ZN(N8747) );
  NOR4_X1 U3633 ( .A1(n3750), .A2(n3751), .A3(n3752), .A4(n3753), .ZN(n3749)
         );
  NAND4_X1 U3634 ( .A1(n3781), .A2(n3782), .A3(n3783), .A4(n3784), .ZN(n3750)
         );
  NAND4_X1 U3635 ( .A1(n3772), .A2(n3773), .A3(n3774), .A4(n3775), .ZN(n3751)
         );
  NOR2_X1 U3636 ( .A1(n5141), .A2(n12666), .ZN(N8715) );
  NOR4_X1 U3637 ( .A1(n5142), .A2(n5143), .A3(n5144), .A4(n5145), .ZN(n5141)
         );
  NAND4_X1 U3638 ( .A1(n5173), .A2(n5174), .A3(n5175), .A4(n5176), .ZN(n5142)
         );
  NAND4_X1 U3639 ( .A1(n5164), .A2(n5165), .A3(n5166), .A4(n5167), .ZN(n5143)
         );
  NOR2_X1 U3640 ( .A1(n3708), .A2(n12674), .ZN(N8748) );
  NOR4_X1 U3641 ( .A1(n3709), .A2(n3710), .A3(n3711), .A4(n3712), .ZN(n3708)
         );
  NAND4_X1 U3642 ( .A1(n3740), .A2(n3741), .A3(n3742), .A4(n3743), .ZN(n3709)
         );
  NAND4_X1 U3643 ( .A1(n3731), .A2(n3732), .A3(n3733), .A4(n3734), .ZN(n3710)
         );
  NOR2_X1 U3644 ( .A1(n5100), .A2(n12666), .ZN(N8716) );
  NOR4_X1 U3645 ( .A1(n5101), .A2(n5102), .A3(n5103), .A4(n5104), .ZN(n5100)
         );
  NAND4_X1 U3646 ( .A1(n5132), .A2(n5133), .A3(n5134), .A4(n5135), .ZN(n5101)
         );
  NAND4_X1 U3647 ( .A1(n5123), .A2(n5124), .A3(n5125), .A4(n5126), .ZN(n5102)
         );
  NOR2_X1 U3648 ( .A1(n3667), .A2(n12674), .ZN(N8749) );
  NOR4_X1 U3649 ( .A1(n3668), .A2(n3669), .A3(n3670), .A4(n3671), .ZN(n3667)
         );
  NAND4_X1 U3650 ( .A1(n3699), .A2(n3700), .A3(n3701), .A4(n3702), .ZN(n3668)
         );
  NAND4_X1 U3651 ( .A1(n3690), .A2(n3691), .A3(n3692), .A4(n3693), .ZN(n3669)
         );
  NOR2_X1 U3652 ( .A1(n5059), .A2(n12666), .ZN(N8717) );
  NOR4_X1 U3653 ( .A1(n5060), .A2(n5061), .A3(n5062), .A4(n5063), .ZN(n5059)
         );
  NAND4_X1 U3654 ( .A1(n5091), .A2(n5092), .A3(n5093), .A4(n5094), .ZN(n5060)
         );
  NAND4_X1 U3655 ( .A1(n5082), .A2(n5083), .A3(n5084), .A4(n5085), .ZN(n5061)
         );
  NOR2_X1 U3656 ( .A1(n3626), .A2(n12674), .ZN(N8750) );
  NOR4_X1 U3657 ( .A1(n3627), .A2(n3628), .A3(n3629), .A4(n3630), .ZN(n3626)
         );
  NAND4_X1 U3658 ( .A1(n3658), .A2(n3659), .A3(n3660), .A4(n3661), .ZN(n3627)
         );
  NAND4_X1 U3659 ( .A1(n3649), .A2(n3650), .A3(n3651), .A4(n3652), .ZN(n3628)
         );
  NOR2_X1 U3660 ( .A1(n5018), .A2(n12666), .ZN(N8718) );
  NOR4_X1 U3661 ( .A1(n5019), .A2(n5020), .A3(n5021), .A4(n5022), .ZN(n5018)
         );
  NAND4_X1 U3662 ( .A1(n5050), .A2(n5051), .A3(n5052), .A4(n5053), .ZN(n5019)
         );
  NAND4_X1 U3663 ( .A1(n5041), .A2(n5042), .A3(n5043), .A4(n5044), .ZN(n5020)
         );
  NOR2_X1 U3664 ( .A1(n3585), .A2(n12675), .ZN(N8751) );
  NOR4_X1 U3665 ( .A1(n3586), .A2(n3587), .A3(n3588), .A4(n3589), .ZN(n3585)
         );
  NAND4_X1 U3666 ( .A1(n3617), .A2(n3618), .A3(n3619), .A4(n3620), .ZN(n3586)
         );
  NAND4_X1 U3667 ( .A1(n3608), .A2(n3609), .A3(n3610), .A4(n3611), .ZN(n3587)
         );
  NOR2_X1 U3668 ( .A1(n4977), .A2(n12667), .ZN(N8719) );
  NOR4_X1 U3669 ( .A1(n4978), .A2(n4979), .A3(n4980), .A4(n4981), .ZN(n4977)
         );
  NAND4_X1 U3670 ( .A1(n5009), .A2(n5010), .A3(n5011), .A4(n5012), .ZN(n4978)
         );
  NAND4_X1 U3671 ( .A1(n5000), .A2(n5001), .A3(n5002), .A4(n5003), .ZN(n4979)
         );
  NOR2_X1 U3672 ( .A1(n3544), .A2(n12675), .ZN(N8752) );
  NOR4_X1 U3673 ( .A1(n3545), .A2(n3546), .A3(n3547), .A4(n3548), .ZN(n3544)
         );
  NAND4_X1 U3674 ( .A1(n3576), .A2(n3577), .A3(n3578), .A4(n3579), .ZN(n3545)
         );
  NAND4_X1 U3675 ( .A1(n3567), .A2(n3568), .A3(n3569), .A4(n3570), .ZN(n3546)
         );
  NOR2_X1 U3676 ( .A1(n4936), .A2(n12667), .ZN(N8720) );
  NOR4_X1 U3677 ( .A1(n4937), .A2(n4938), .A3(n4939), .A4(n4940), .ZN(n4936)
         );
  NAND4_X1 U3678 ( .A1(n4968), .A2(n4969), .A3(n4970), .A4(n4971), .ZN(n4937)
         );
  NAND4_X1 U3679 ( .A1(n4959), .A2(n4960), .A3(n4961), .A4(n4962), .ZN(n4938)
         );
  NOR2_X1 U3680 ( .A1(n3503), .A2(n12675), .ZN(N8753) );
  NOR4_X1 U3681 ( .A1(n3504), .A2(n3505), .A3(n3506), .A4(n3507), .ZN(n3503)
         );
  NAND4_X1 U3682 ( .A1(n3535), .A2(n3536), .A3(n3537), .A4(n3538), .ZN(n3504)
         );
  NAND4_X1 U3683 ( .A1(n3526), .A2(n3527), .A3(n3528), .A4(n3529), .ZN(n3505)
         );
  NOR2_X1 U3684 ( .A1(n4895), .A2(n12667), .ZN(N8721) );
  NOR4_X1 U3685 ( .A1(n4896), .A2(n4897), .A3(n4898), .A4(n4899), .ZN(n4895)
         );
  NAND4_X1 U3686 ( .A1(n4927), .A2(n4928), .A3(n4929), .A4(n4930), .ZN(n4896)
         );
  NAND4_X1 U3687 ( .A1(n4918), .A2(n4919), .A3(n4920), .A4(n4921), .ZN(n4897)
         );
  NOR2_X1 U3688 ( .A1(n3462), .A2(n12675), .ZN(N8754) );
  NOR4_X1 U3689 ( .A1(n3463), .A2(n3464), .A3(n3465), .A4(n3466), .ZN(n3462)
         );
  NAND4_X1 U3690 ( .A1(n3494), .A2(n3495), .A3(n3496), .A4(n3497), .ZN(n3463)
         );
  NAND4_X1 U3691 ( .A1(n3485), .A2(n3486), .A3(n3487), .A4(n3488), .ZN(n3464)
         );
  NOR2_X1 U3692 ( .A1(n4854), .A2(n12667), .ZN(N8722) );
  NOR4_X1 U3693 ( .A1(n4855), .A2(n4856), .A3(n4857), .A4(n4858), .ZN(n4854)
         );
  NAND4_X1 U3694 ( .A1(n4886), .A2(n4887), .A3(n4888), .A4(n4889), .ZN(n4855)
         );
  NAND4_X1 U3695 ( .A1(n4877), .A2(n4878), .A3(n4879), .A4(n4880), .ZN(n4856)
         );
  NOR2_X1 U3696 ( .A1(n3421), .A2(n12676), .ZN(N8755) );
  NOR4_X1 U3697 ( .A1(n3422), .A2(n3423), .A3(n3424), .A4(n3425), .ZN(n3421)
         );
  NAND4_X1 U3698 ( .A1(n3453), .A2(n3454), .A3(n3455), .A4(n3456), .ZN(n3422)
         );
  NAND4_X1 U3699 ( .A1(n3444), .A2(n3445), .A3(n3446), .A4(n3447), .ZN(n3423)
         );
  NOR2_X1 U3700 ( .A1(n4813), .A2(n12668), .ZN(N8723) );
  NOR4_X1 U3701 ( .A1(n4814), .A2(n4815), .A3(n4816), .A4(n4817), .ZN(n4813)
         );
  NAND4_X1 U3702 ( .A1(n4845), .A2(n4846), .A3(n4847), .A4(n4848), .ZN(n4814)
         );
  NAND4_X1 U3703 ( .A1(n4836), .A2(n4837), .A3(n4838), .A4(n4839), .ZN(n4815)
         );
  NOR2_X1 U3704 ( .A1(n3380), .A2(n12676), .ZN(N8756) );
  NOR4_X1 U3705 ( .A1(n3381), .A2(n3382), .A3(n3383), .A4(n3384), .ZN(n3380)
         );
  NAND4_X1 U3706 ( .A1(n3412), .A2(n3413), .A3(n3414), .A4(n3415), .ZN(n3381)
         );
  NAND4_X1 U3707 ( .A1(n3403), .A2(n3404), .A3(n3405), .A4(n3406), .ZN(n3382)
         );
  NOR2_X1 U3708 ( .A1(n4772), .A2(n12668), .ZN(N8724) );
  NOR4_X1 U3709 ( .A1(n4773), .A2(n4774), .A3(n4775), .A4(n4776), .ZN(n4772)
         );
  NAND4_X1 U3710 ( .A1(n4804), .A2(n4805), .A3(n4806), .A4(n4807), .ZN(n4773)
         );
  NAND4_X1 U3711 ( .A1(n4795), .A2(n4796), .A3(n4797), .A4(n4798), .ZN(n4774)
         );
  NOR2_X1 U3712 ( .A1(n3339), .A2(n12676), .ZN(N8757) );
  NOR4_X1 U3713 ( .A1(n3340), .A2(n3341), .A3(n3342), .A4(n3343), .ZN(n3339)
         );
  NAND4_X1 U3714 ( .A1(n3371), .A2(n3372), .A3(n3373), .A4(n3374), .ZN(n3340)
         );
  NAND4_X1 U3715 ( .A1(n3362), .A2(n3363), .A3(n3364), .A4(n3365), .ZN(n3341)
         );
  NOR2_X1 U3716 ( .A1(n4731), .A2(n12668), .ZN(N8725) );
  NOR4_X1 U3717 ( .A1(n4732), .A2(n4733), .A3(n4734), .A4(n4735), .ZN(n4731)
         );
  NAND4_X1 U3718 ( .A1(n4763), .A2(n4764), .A3(n4765), .A4(n4766), .ZN(n4732)
         );
  NAND4_X1 U3719 ( .A1(n4754), .A2(n4755), .A3(n4756), .A4(n4757), .ZN(n4733)
         );
  NOR2_X1 U3720 ( .A1(n3298), .A2(n12676), .ZN(N8758) );
  NOR4_X1 U3721 ( .A1(n3299), .A2(n3300), .A3(n3301), .A4(n3302), .ZN(n3298)
         );
  NAND4_X1 U3722 ( .A1(n3330), .A2(n3331), .A3(n3332), .A4(n3333), .ZN(n3299)
         );
  NAND4_X1 U3723 ( .A1(n3321), .A2(n3322), .A3(n3323), .A4(n3324), .ZN(n3300)
         );
  NOR2_X1 U3724 ( .A1(n4690), .A2(n12668), .ZN(N8726) );
  NOR4_X1 U3725 ( .A1(n4691), .A2(n4692), .A3(n4693), .A4(n4694), .ZN(n4690)
         );
  NAND4_X1 U3726 ( .A1(n4722), .A2(n4723), .A3(n4724), .A4(n4725), .ZN(n4691)
         );
  NAND4_X1 U3727 ( .A1(n4713), .A2(n4714), .A3(n4715), .A4(n4716), .ZN(n4692)
         );
  NOR2_X1 U3728 ( .A1(n3257), .A2(n12677), .ZN(N8759) );
  NOR4_X1 U3729 ( .A1(n3258), .A2(n3259), .A3(n3260), .A4(n3261), .ZN(n3257)
         );
  NAND4_X1 U3730 ( .A1(n3289), .A2(n3290), .A3(n3291), .A4(n3292), .ZN(n3258)
         );
  NAND4_X1 U3731 ( .A1(n3280), .A2(n3281), .A3(n3282), .A4(n3283), .ZN(n3259)
         );
  NOR2_X1 U3732 ( .A1(n4649), .A2(n12669), .ZN(N8727) );
  NOR4_X1 U3733 ( .A1(n4650), .A2(n4651), .A3(n4652), .A4(n4653), .ZN(n4649)
         );
  NAND4_X1 U3734 ( .A1(n4681), .A2(n4682), .A3(n4683), .A4(n4684), .ZN(n4650)
         );
  NAND4_X1 U3735 ( .A1(n4672), .A2(n4673), .A3(n4674), .A4(n4675), .ZN(n4651)
         );
  NOR2_X1 U3736 ( .A1(n3216), .A2(n12677), .ZN(N8760) );
  NOR4_X1 U3737 ( .A1(n3217), .A2(n3218), .A3(n3219), .A4(n3220), .ZN(n3216)
         );
  NAND4_X1 U3738 ( .A1(n3248), .A2(n3249), .A3(n3250), .A4(n3251), .ZN(n3217)
         );
  NAND4_X1 U3739 ( .A1(n3239), .A2(n3240), .A3(n3241), .A4(n3242), .ZN(n3218)
         );
  NOR2_X1 U3740 ( .A1(n4608), .A2(n12669), .ZN(N8728) );
  NOR4_X1 U3741 ( .A1(n4609), .A2(n4610), .A3(n4611), .A4(n4612), .ZN(n4608)
         );
  NAND4_X1 U3742 ( .A1(n4640), .A2(n4641), .A3(n4642), .A4(n4643), .ZN(n4609)
         );
  NAND4_X1 U3743 ( .A1(n4631), .A2(n4632), .A3(n4633), .A4(n4634), .ZN(n4610)
         );
  NOR2_X1 U3744 ( .A1(n3175), .A2(n12677), .ZN(N8761) );
  NOR4_X1 U3745 ( .A1(n3176), .A2(n3177), .A3(n3178), .A4(n3179), .ZN(n3175)
         );
  NAND4_X1 U3746 ( .A1(n3207), .A2(n3208), .A3(n3209), .A4(n3210), .ZN(n3176)
         );
  NAND4_X1 U3747 ( .A1(n3198), .A2(n3199), .A3(n3200), .A4(n3201), .ZN(n3177)
         );
  NOR2_X1 U3748 ( .A1(n4567), .A2(n12669), .ZN(N8729) );
  NOR4_X1 U3749 ( .A1(n4568), .A2(n4569), .A3(n4570), .A4(n4571), .ZN(n4567)
         );
  NAND4_X1 U3750 ( .A1(n4599), .A2(n4600), .A3(n4601), .A4(n4602), .ZN(n4568)
         );
  NAND4_X1 U3751 ( .A1(n4590), .A2(n4591), .A3(n4592), .A4(n4593), .ZN(n4569)
         );
  NOR2_X1 U3752 ( .A1(n3134), .A2(n12677), .ZN(N8762) );
  NOR4_X1 U3753 ( .A1(n3135), .A2(n3136), .A3(n3137), .A4(n3138), .ZN(n3134)
         );
  NAND4_X1 U3754 ( .A1(n3166), .A2(n3167), .A3(n3168), .A4(n3169), .ZN(n3135)
         );
  NAND4_X1 U3755 ( .A1(n3157), .A2(n3158), .A3(n3159), .A4(n3160), .ZN(n3136)
         );
  NOR2_X1 U3756 ( .A1(n4526), .A2(n12669), .ZN(N8730) );
  NOR4_X1 U3757 ( .A1(n4527), .A2(n4528), .A3(n4529), .A4(n4530), .ZN(n4526)
         );
  NAND4_X1 U3758 ( .A1(n4558), .A2(n4559), .A3(n4560), .A4(n4561), .ZN(n4527)
         );
  NAND4_X1 U3759 ( .A1(n4549), .A2(n4550), .A3(n4551), .A4(n4552), .ZN(n4528)
         );
  NOR2_X1 U3760 ( .A1(n3093), .A2(n12678), .ZN(N8763) );
  NOR4_X1 U3761 ( .A1(n3094), .A2(n3095), .A3(n3096), .A4(n3097), .ZN(n3093)
         );
  NAND4_X1 U3762 ( .A1(n3125), .A2(n3126), .A3(n3127), .A4(n3128), .ZN(n3094)
         );
  NAND4_X1 U3763 ( .A1(n3116), .A2(n3117), .A3(n3118), .A4(n3119), .ZN(n3095)
         );
  NOR2_X1 U3764 ( .A1(n4485), .A2(n12670), .ZN(N8731) );
  NOR4_X1 U3765 ( .A1(n4486), .A2(n4487), .A3(n4488), .A4(n4489), .ZN(n4485)
         );
  NAND4_X1 U3766 ( .A1(n4517), .A2(n4518), .A3(n4519), .A4(n4520), .ZN(n4486)
         );
  NAND4_X1 U3767 ( .A1(n4508), .A2(n4509), .A3(n4510), .A4(n4511), .ZN(n4487)
         );
  NOR2_X1 U3768 ( .A1(n3052), .A2(n12678), .ZN(N8764) );
  NOR4_X1 U3769 ( .A1(n3053), .A2(n3054), .A3(n3055), .A4(n3056), .ZN(n3052)
         );
  NAND4_X1 U3770 ( .A1(n3084), .A2(n3085), .A3(n3086), .A4(n3087), .ZN(n3053)
         );
  NAND4_X1 U3771 ( .A1(n3075), .A2(n3076), .A3(n3077), .A4(n3078), .ZN(n3054)
         );
  NOR2_X1 U3772 ( .A1(n4444), .A2(n12670), .ZN(N8732) );
  NOR4_X1 U3773 ( .A1(n4445), .A2(n4446), .A3(n4447), .A4(n4448), .ZN(n4444)
         );
  NAND4_X1 U3774 ( .A1(n4476), .A2(n4477), .A3(n4478), .A4(n4479), .ZN(n4445)
         );
  NAND4_X1 U3775 ( .A1(n4467), .A2(n4468), .A3(n4469), .A4(n4470), .ZN(n4446)
         );
  NOR2_X1 U3776 ( .A1(n3011), .A2(n12678), .ZN(N8765) );
  NOR4_X1 U3777 ( .A1(n3012), .A2(n3013), .A3(n3014), .A4(n3015), .ZN(n3011)
         );
  NAND4_X1 U3778 ( .A1(n3043), .A2(n3044), .A3(n3045), .A4(n3046), .ZN(n3012)
         );
  NAND4_X1 U3779 ( .A1(n3034), .A2(n3035), .A3(n3036), .A4(n3037), .ZN(n3013)
         );
  NOR2_X1 U3780 ( .A1(n4403), .A2(n12670), .ZN(N8733) );
  NOR4_X1 U3781 ( .A1(n4404), .A2(n4405), .A3(n4406), .A4(n4407), .ZN(n4403)
         );
  NAND4_X1 U3782 ( .A1(n4435), .A2(n4436), .A3(n4437), .A4(n4438), .ZN(n4404)
         );
  NAND4_X1 U3783 ( .A1(n4426), .A2(n4427), .A3(n4428), .A4(n4429), .ZN(n4405)
         );
  NOR2_X1 U3784 ( .A1(n2970), .A2(n12678), .ZN(N8766) );
  NOR4_X1 U3785 ( .A1(n2971), .A2(n2972), .A3(n2973), .A4(n2974), .ZN(n2970)
         );
  NAND4_X1 U3786 ( .A1(n3002), .A2(n3003), .A3(n3004), .A4(n3005), .ZN(n2971)
         );
  NAND4_X1 U3787 ( .A1(n2993), .A2(n2994), .A3(n2995), .A4(n2996), .ZN(n2972)
         );
  NOR2_X1 U3788 ( .A1(n4274), .A2(n12670), .ZN(N8734) );
  NOR4_X1 U3789 ( .A1(n4275), .A2(n4276), .A3(n4277), .A4(n4278), .ZN(n4274)
         );
  NAND4_X1 U3790 ( .A1(n4372), .A2(n4373), .A3(n4374), .A4(n4375), .ZN(n4275)
         );
  NAND4_X1 U3791 ( .A1(n4341), .A2(n4342), .A3(n4343), .A4(n4344), .ZN(n4276)
         );
  NOR2_X1 U3792 ( .A1(n2742), .A2(n12671), .ZN(N8767) );
  NOR4_X1 U3793 ( .A1(n2743), .A2(n2744), .A3(n2745), .A4(n2746), .ZN(n2742)
         );
  NAND4_X1 U3794 ( .A1(n2939), .A2(n2940), .A3(n2941), .A4(n2942), .ZN(n2743)
         );
  NAND4_X1 U3795 ( .A1(n2873), .A2(n2874), .A3(n2875), .A4(n2876), .ZN(n2744)
         );
  OAI222_X1 U3796 ( .A1(n12779), .A2(n2481), .B1(n2482), .B2(n2480), .C1(n2936), .C2(n14517), .ZN(n9133) );
  INV_X1 U3797 ( .A(n2482), .ZN(n12779) );
  XNOR2_X1 U3798 ( .A(n10626), .B(n2937), .ZN(n2482) );
  OAI21_X1 U3799 ( .B1(RETRN), .B2(CALL), .A(ENABLE), .ZN(n2478) );
  OR3_X1 U3800 ( .A1(n10626), .A2(n2935), .A3(n10625), .ZN(n2489) );
  OAI221_X1 U3801 ( .B1(n2483), .B2(n2484), .C1(n2935), .C2(n2485), .A(n2486), 
        .ZN(n9132) );
  NAND2_X1 U3802 ( .A1(RETRN), .A2(n14517), .ZN(n2484) );
  NAND4_X1 U3803 ( .A1(n12777), .A2(n2935), .A3(n10626), .A4(n10625), .ZN(
        n2486) );
  AOI211_X1 U3804 ( .C1(n12777), .C2(n2487), .A(n2478), .B(n2488), .ZN(n2485)
         );
  OAI22_X1 U3805 ( .A1(n10844), .A2(n12317), .B1(n10511), .B2(n12318), .ZN(
        n8843) );
  OAI22_X1 U3806 ( .A1(n10837), .A2(n12317), .B1(n10479), .B2(n12318), .ZN(
        n8842) );
  OAI22_X1 U3807 ( .A1(n10830), .A2(n12317), .B1(n10447), .B2(n12318), .ZN(
        n8841) );
  OAI22_X1 U3808 ( .A1(n10823), .A2(n12317), .B1(n10415), .B2(n12318), .ZN(
        n8840) );
  OAI22_X1 U3809 ( .A1(n10816), .A2(n12317), .B1(n10380), .B2(n12319), .ZN(
        n8839) );
  OAI22_X1 U3810 ( .A1(n10809), .A2(n12317), .B1(n10348), .B2(n12319), .ZN(
        n8838) );
  OAI22_X1 U3811 ( .A1(n10802), .A2(n12317), .B1(n10316), .B2(n12319), .ZN(
        n8837) );
  OAI22_X1 U3812 ( .A1(n10795), .A2(n12317), .B1(n10281), .B2(n12319), .ZN(
        n8836) );
  OAI22_X1 U3813 ( .A1(n10788), .A2(n12316), .B1(n10249), .B2(n12320), .ZN(
        n8835) );
  OAI22_X1 U3814 ( .A1(n10781), .A2(n12316), .B1(n10217), .B2(n12320), .ZN(
        n8834) );
  OAI22_X1 U3815 ( .A1(n10774), .A2(n12316), .B1(n10183), .B2(n12320), .ZN(
        n8833) );
  OAI22_X1 U3816 ( .A1(n10767), .A2(n12316), .B1(n10151), .B2(n12320), .ZN(
        n8832) );
  OAI22_X1 U3817 ( .A1(n10760), .A2(n12316), .B1(n10119), .B2(n12321), .ZN(
        n8831) );
  OAI22_X1 U3818 ( .A1(n10753), .A2(n12316), .B1(n10087), .B2(n12321), .ZN(
        n8830) );
  OAI22_X1 U3819 ( .A1(n10746), .A2(n12316), .B1(n10055), .B2(n12321), .ZN(
        n8829) );
  OAI22_X1 U3820 ( .A1(n10739), .A2(n12316), .B1(n10023), .B2(n12321), .ZN(
        n8828) );
  OAI22_X1 U3821 ( .A1(n10732), .A2(n12316), .B1(n9661), .B2(n12322), .ZN(
        n8827) );
  OAI22_X1 U3822 ( .A1(n10725), .A2(n12316), .B1(n9629), .B2(n12322), .ZN(
        n8826) );
  OAI22_X1 U3823 ( .A1(n10718), .A2(n12316), .B1(n9597), .B2(n12322), .ZN(
        n8825) );
  OAI22_X1 U3824 ( .A1(n10711), .A2(n12316), .B1(n9263), .B2(n12322), .ZN(
        n8824) );
  OAI22_X1 U3825 ( .A1(n10704), .A2(n12315), .B1(n9199), .B2(n12323), .ZN(
        n8823) );
  OAI22_X1 U3826 ( .A1(n10697), .A2(n12315), .B1(n9167), .B2(n12323), .ZN(
        n8822) );
  OAI22_X1 U3827 ( .A1(n10690), .A2(n12315), .B1(n9135), .B2(n12323), .ZN(
        n8821) );
  OAI22_X1 U3828 ( .A1(n10683), .A2(n12315), .B1(n6000), .B2(n12323), .ZN(
        n8820) );
  OAI22_X1 U3829 ( .A1(n10676), .A2(n12315), .B1(n5936), .B2(n12324), .ZN(
        n8819) );
  OAI22_X1 U3830 ( .A1(n10669), .A2(n12315), .B1(n5904), .B2(n12324), .ZN(
        n8818) );
  OAI22_X1 U3831 ( .A1(n10662), .A2(n12315), .B1(n5872), .B2(n12324), .ZN(
        n8817) );
  OAI22_X1 U3832 ( .A1(n10655), .A2(n12315), .B1(n5840), .B2(n12324), .ZN(
        n8816) );
  OAI22_X1 U3833 ( .A1(n10648), .A2(n12315), .B1(n5808), .B2(n12325), .ZN(
        n8815) );
  OAI22_X1 U3834 ( .A1(n10641), .A2(n12315), .B1(n5776), .B2(n12325), .ZN(
        n8814) );
  OAI22_X1 U3835 ( .A1(n10634), .A2(n12315), .B1(n5744), .B2(n12325), .ZN(
        n8813) );
  OAI22_X1 U3836 ( .A1(n10627), .A2(n12315), .B1(n5712), .B2(n12325), .ZN(
        n8812) );
  OAI22_X1 U3837 ( .A1(n10628), .A2(n12267), .B1(n996), .B2(n12270), .ZN(n8684) );
  OAI22_X1 U3838 ( .A1(n10628), .A2(n12231), .B1(n997), .B2(n12234), .ZN(n8588) );
  OAI22_X1 U3839 ( .A1(n10628), .A2(n12195), .B1(n998), .B2(n12198), .ZN(n8492) );
  OAI22_X1 U3840 ( .A1(n10846), .A2(n12089), .B1(n10516), .B2(n12090), .ZN(
        n8235) );
  OAI22_X1 U3841 ( .A1(n10839), .A2(n12089), .B1(n10484), .B2(n12090), .ZN(
        n8234) );
  OAI22_X1 U3842 ( .A1(n10832), .A2(n12089), .B1(n10452), .B2(n12090), .ZN(
        n8233) );
  OAI22_X1 U3843 ( .A1(n10825), .A2(n12089), .B1(n10420), .B2(n12090), .ZN(
        n8232) );
  OAI22_X1 U3844 ( .A1(n10818), .A2(n12089), .B1(n10385), .B2(n12091), .ZN(
        n8231) );
  OAI22_X1 U3845 ( .A1(n10811), .A2(n12089), .B1(n10353), .B2(n12091), .ZN(
        n8230) );
  OAI22_X1 U3846 ( .A1(n10804), .A2(n12089), .B1(n10321), .B2(n12091), .ZN(
        n8229) );
  OAI22_X1 U3847 ( .A1(n10797), .A2(n12089), .B1(n10286), .B2(n12091), .ZN(
        n8228) );
  OAI22_X1 U3848 ( .A1(n10790), .A2(n12088), .B1(n10254), .B2(n12092), .ZN(
        n8227) );
  OAI22_X1 U3849 ( .A1(n10783), .A2(n12088), .B1(n10222), .B2(n12092), .ZN(
        n8226) );
  OAI22_X1 U3850 ( .A1(n10776), .A2(n12088), .B1(n10188), .B2(n12092), .ZN(
        n8225) );
  OAI22_X1 U3851 ( .A1(n10769), .A2(n12088), .B1(n10156), .B2(n12092), .ZN(
        n8224) );
  OAI22_X1 U3852 ( .A1(n10762), .A2(n12088), .B1(n10124), .B2(n12093), .ZN(
        n8223) );
  OAI22_X1 U3853 ( .A1(n10755), .A2(n12088), .B1(n10092), .B2(n12093), .ZN(
        n8222) );
  OAI22_X1 U3854 ( .A1(n10748), .A2(n12088), .B1(n10060), .B2(n12093), .ZN(
        n8221) );
  OAI22_X1 U3855 ( .A1(n10741), .A2(n12088), .B1(n10028), .B2(n12093), .ZN(
        n8220) );
  OAI22_X1 U3856 ( .A1(n10734), .A2(n12088), .B1(n9698), .B2(n12094), .ZN(
        n8219) );
  OAI22_X1 U3857 ( .A1(n10727), .A2(n12088), .B1(n9634), .B2(n12094), .ZN(
        n8218) );
  OAI22_X1 U3858 ( .A1(n10720), .A2(n12088), .B1(n9602), .B2(n12094), .ZN(
        n8217) );
  OAI22_X1 U3859 ( .A1(n10713), .A2(n12088), .B1(n9570), .B2(n12094), .ZN(
        n8216) );
  OAI22_X1 U3860 ( .A1(n10706), .A2(n12087), .B1(n9204), .B2(n12095), .ZN(
        n8215) );
  OAI22_X1 U3861 ( .A1(n10699), .A2(n12087), .B1(n9172), .B2(n12095), .ZN(
        n8214) );
  OAI22_X1 U3862 ( .A1(n10692), .A2(n12087), .B1(n9140), .B2(n12095), .ZN(
        n8213) );
  OAI22_X1 U3863 ( .A1(n10685), .A2(n12087), .B1(n6005), .B2(n12095), .ZN(
        n8212) );
  OAI22_X1 U3864 ( .A1(n10678), .A2(n12087), .B1(n5941), .B2(n12096), .ZN(
        n8211) );
  OAI22_X1 U3865 ( .A1(n10671), .A2(n12087), .B1(n5909), .B2(n12096), .ZN(
        n8210) );
  OAI22_X1 U3866 ( .A1(n10664), .A2(n12087), .B1(n5877), .B2(n12096), .ZN(
        n8209) );
  OAI22_X1 U3867 ( .A1(n10657), .A2(n12087), .B1(n5845), .B2(n12096), .ZN(
        n8208) );
  OAI22_X1 U3868 ( .A1(n10650), .A2(n12087), .B1(n5813), .B2(n12097), .ZN(
        n8207) );
  OAI22_X1 U3869 ( .A1(n10643), .A2(n12087), .B1(n5781), .B2(n12097), .ZN(
        n8206) );
  OAI22_X1 U3870 ( .A1(n10636), .A2(n12087), .B1(n5749), .B2(n12097), .ZN(
        n8205) );
  OAI22_X1 U3871 ( .A1(n10629), .A2(n12087), .B1(n5717), .B2(n12097), .ZN(
        n8204) );
  OAI22_X1 U3872 ( .A1(n10846), .A2(n12053), .B1(n10519), .B2(n12054), .ZN(
        n8139) );
  OAI22_X1 U3873 ( .A1(n10839), .A2(n12053), .B1(n10487), .B2(n12054), .ZN(
        n8138) );
  OAI22_X1 U3874 ( .A1(n10832), .A2(n12053), .B1(n10455), .B2(n12054), .ZN(
        n8137) );
  OAI22_X1 U3875 ( .A1(n10825), .A2(n12053), .B1(n10423), .B2(n12054), .ZN(
        n8136) );
  OAI22_X1 U3876 ( .A1(n10818), .A2(n12053), .B1(n10388), .B2(n12055), .ZN(
        n8135) );
  OAI22_X1 U3877 ( .A1(n10811), .A2(n12053), .B1(n10356), .B2(n12055), .ZN(
        n8134) );
  OAI22_X1 U3878 ( .A1(n10804), .A2(n12053), .B1(n10324), .B2(n12055), .ZN(
        n8133) );
  OAI22_X1 U3879 ( .A1(n10797), .A2(n12053), .B1(n10289), .B2(n12055), .ZN(
        n8132) );
  OAI22_X1 U3880 ( .A1(n10790), .A2(n12052), .B1(n10257), .B2(n12056), .ZN(
        n8131) );
  OAI22_X1 U3881 ( .A1(n10783), .A2(n12052), .B1(n10225), .B2(n12056), .ZN(
        n8130) );
  OAI22_X1 U3882 ( .A1(n10776), .A2(n12052), .B1(n10191), .B2(n12056), .ZN(
        n8129) );
  OAI22_X1 U3883 ( .A1(n10769), .A2(n12052), .B1(n10159), .B2(n12056), .ZN(
        n8128) );
  OAI22_X1 U3884 ( .A1(n10762), .A2(n12052), .B1(n10127), .B2(n12057), .ZN(
        n8127) );
  OAI22_X1 U3885 ( .A1(n10755), .A2(n12052), .B1(n10095), .B2(n12057), .ZN(
        n8126) );
  OAI22_X1 U3886 ( .A1(n10748), .A2(n12052), .B1(n10063), .B2(n12057), .ZN(
        n8125) );
  OAI22_X1 U3887 ( .A1(n10741), .A2(n12052), .B1(n10031), .B2(n12057), .ZN(
        n8124) );
  OAI22_X1 U3888 ( .A1(n10734), .A2(n12052), .B1(n9701), .B2(n12058), .ZN(
        n8123) );
  OAI22_X1 U3889 ( .A1(n10727), .A2(n12052), .B1(n9637), .B2(n12058), .ZN(
        n8122) );
  OAI22_X1 U3890 ( .A1(n10720), .A2(n12052), .B1(n9605), .B2(n12058), .ZN(
        n8121) );
  OAI22_X1 U3891 ( .A1(n10713), .A2(n12052), .B1(n9573), .B2(n12058), .ZN(
        n8120) );
  OAI22_X1 U3892 ( .A1(n10706), .A2(n12051), .B1(n9207), .B2(n12059), .ZN(
        n8119) );
  OAI22_X1 U3893 ( .A1(n10699), .A2(n12051), .B1(n9175), .B2(n12059), .ZN(
        n8118) );
  OAI22_X1 U3894 ( .A1(n10692), .A2(n12051), .B1(n9143), .B2(n12059), .ZN(
        n8117) );
  OAI22_X1 U3895 ( .A1(n10685), .A2(n12051), .B1(n6008), .B2(n12059), .ZN(
        n8116) );
  OAI22_X1 U3896 ( .A1(n10678), .A2(n12051), .B1(n5944), .B2(n12060), .ZN(
        n8115) );
  OAI22_X1 U3897 ( .A1(n10671), .A2(n12051), .B1(n5912), .B2(n12060), .ZN(
        n8114) );
  OAI22_X1 U3898 ( .A1(n10664), .A2(n12051), .B1(n5880), .B2(n12060), .ZN(
        n8113) );
  OAI22_X1 U3899 ( .A1(n10657), .A2(n12051), .B1(n5848), .B2(n12060), .ZN(
        n8112) );
  OAI22_X1 U3900 ( .A1(n10650), .A2(n12051), .B1(n5816), .B2(n12061), .ZN(
        n8111) );
  OAI22_X1 U3901 ( .A1(n10643), .A2(n12051), .B1(n5784), .B2(n12061), .ZN(
        n8110) );
  OAI22_X1 U3902 ( .A1(n10636), .A2(n12051), .B1(n5752), .B2(n12061), .ZN(
        n8109) );
  OAI22_X1 U3903 ( .A1(n10629), .A2(n12051), .B1(n5720), .B2(n12061), .ZN(
        n8108) );
  OAI22_X1 U3904 ( .A1(n10847), .A2(n11825), .B1(n10524), .B2(n11826), .ZN(
        n7531) );
  OAI22_X1 U3905 ( .A1(n10840), .A2(n11825), .B1(n10492), .B2(n11826), .ZN(
        n7530) );
  OAI22_X1 U3906 ( .A1(n10833), .A2(n11825), .B1(n10460), .B2(n11826), .ZN(
        n7529) );
  OAI22_X1 U3907 ( .A1(n10826), .A2(n11825), .B1(n10428), .B2(n11826), .ZN(
        n7528) );
  OAI22_X1 U3908 ( .A1(n10819), .A2(n11825), .B1(n10393), .B2(n11827), .ZN(
        n7527) );
  OAI22_X1 U3909 ( .A1(n10812), .A2(n11825), .B1(n10361), .B2(n11827), .ZN(
        n7526) );
  OAI22_X1 U3910 ( .A1(n10805), .A2(n11825), .B1(n10329), .B2(n11827), .ZN(
        n7525) );
  OAI22_X1 U3911 ( .A1(n10798), .A2(n11825), .B1(n10294), .B2(n11827), .ZN(
        n7524) );
  OAI22_X1 U3912 ( .A1(n10791), .A2(n11824), .B1(n10262), .B2(n11828), .ZN(
        n7523) );
  OAI22_X1 U3913 ( .A1(n10784), .A2(n11824), .B1(n10230), .B2(n11828), .ZN(
        n7522) );
  OAI22_X1 U3914 ( .A1(n10777), .A2(n11824), .B1(n10196), .B2(n11828), .ZN(
        n7521) );
  OAI22_X1 U3915 ( .A1(n10770), .A2(n11824), .B1(n10164), .B2(n11828), .ZN(
        n7520) );
  OAI22_X1 U3916 ( .A1(n10763), .A2(n11824), .B1(n10132), .B2(n11829), .ZN(
        n7519) );
  OAI22_X1 U3917 ( .A1(n10756), .A2(n11824), .B1(n10100), .B2(n11829), .ZN(
        n7518) );
  OAI22_X1 U3918 ( .A1(n10749), .A2(n11824), .B1(n10068), .B2(n11829), .ZN(
        n7517) );
  OAI22_X1 U3919 ( .A1(n10742), .A2(n11824), .B1(n10036), .B2(n11829), .ZN(
        n7516) );
  OAI22_X1 U3920 ( .A1(n10735), .A2(n11824), .B1(n10004), .B2(n11830), .ZN(
        n7515) );
  OAI22_X1 U3921 ( .A1(n10728), .A2(n11824), .B1(n9642), .B2(n11830), .ZN(
        n7514) );
  OAI22_X1 U3922 ( .A1(n10721), .A2(n11824), .B1(n9610), .B2(n11830), .ZN(
        n7513) );
  OAI22_X1 U3923 ( .A1(n10714), .A2(n11824), .B1(n9578), .B2(n11830), .ZN(
        n7512) );
  OAI22_X1 U3924 ( .A1(n10707), .A2(n11823), .B1(n9212), .B2(n11831), .ZN(
        n7511) );
  OAI22_X1 U3925 ( .A1(n10700), .A2(n11823), .B1(n9180), .B2(n11831), .ZN(
        n7510) );
  OAI22_X1 U3926 ( .A1(n10693), .A2(n11823), .B1(n9148), .B2(n11831), .ZN(
        n7509) );
  OAI22_X1 U3927 ( .A1(n10686), .A2(n11823), .B1(n6044), .B2(n11831), .ZN(
        n7508) );
  OAI22_X1 U3928 ( .A1(n10679), .A2(n11823), .B1(n5981), .B2(n11832), .ZN(
        n7507) );
  OAI22_X1 U3929 ( .A1(n10672), .A2(n11823), .B1(n5917), .B2(n11832), .ZN(
        n7506) );
  OAI22_X1 U3930 ( .A1(n10665), .A2(n11823), .B1(n5885), .B2(n11832), .ZN(
        n7505) );
  OAI22_X1 U3931 ( .A1(n10658), .A2(n11823), .B1(n5853), .B2(n11832), .ZN(
        n7504) );
  OAI22_X1 U3932 ( .A1(n10651), .A2(n11823), .B1(n5821), .B2(n11833), .ZN(
        n7503) );
  OAI22_X1 U3933 ( .A1(n10644), .A2(n11823), .B1(n5789), .B2(n11833), .ZN(
        n7502) );
  OAI22_X1 U3934 ( .A1(n10637), .A2(n11823), .B1(n5757), .B2(n11833), .ZN(
        n7501) );
  OAI22_X1 U3935 ( .A1(n10630), .A2(n11823), .B1(n5725), .B2(n11833), .ZN(
        n7500) );
  OAI22_X1 U3936 ( .A1(n10848), .A2(n11789), .B1(n10527), .B2(n11790), .ZN(
        n7435) );
  OAI22_X1 U3937 ( .A1(n10841), .A2(n11789), .B1(n10495), .B2(n11790), .ZN(
        n7434) );
  OAI22_X1 U3938 ( .A1(n10834), .A2(n11789), .B1(n10463), .B2(n11790), .ZN(
        n7433) );
  OAI22_X1 U3939 ( .A1(n10827), .A2(n11789), .B1(n10431), .B2(n11790), .ZN(
        n7432) );
  OAI22_X1 U3940 ( .A1(n10820), .A2(n11789), .B1(n10396), .B2(n11791), .ZN(
        n7431) );
  OAI22_X1 U3941 ( .A1(n10813), .A2(n11789), .B1(n10364), .B2(n11791), .ZN(
        n7430) );
  OAI22_X1 U3942 ( .A1(n10806), .A2(n11789), .B1(n10332), .B2(n11791), .ZN(
        n7429) );
  OAI22_X1 U3943 ( .A1(n10799), .A2(n11789), .B1(n10297), .B2(n11791), .ZN(
        n7428) );
  OAI22_X1 U3944 ( .A1(n10792), .A2(n11788), .B1(n10265), .B2(n11792), .ZN(
        n7427) );
  OAI22_X1 U3945 ( .A1(n10785), .A2(n11788), .B1(n10233), .B2(n11792), .ZN(
        n7426) );
  OAI22_X1 U3946 ( .A1(n10778), .A2(n11788), .B1(n10199), .B2(n11792), .ZN(
        n7425) );
  OAI22_X1 U3947 ( .A1(n10771), .A2(n11788), .B1(n10167), .B2(n11792), .ZN(
        n7424) );
  OAI22_X1 U3948 ( .A1(n10764), .A2(n11788), .B1(n10135), .B2(n11793), .ZN(
        n7423) );
  OAI22_X1 U3949 ( .A1(n10757), .A2(n11788), .B1(n10103), .B2(n11793), .ZN(
        n7422) );
  OAI22_X1 U3950 ( .A1(n10750), .A2(n11788), .B1(n10071), .B2(n11793), .ZN(
        n7421) );
  OAI22_X1 U3951 ( .A1(n10743), .A2(n11788), .B1(n10039), .B2(n11793), .ZN(
        n7420) );
  OAI22_X1 U3952 ( .A1(n10736), .A2(n11788), .B1(n10007), .B2(n11794), .ZN(
        n7419) );
  OAI22_X1 U3953 ( .A1(n10729), .A2(n11788), .B1(n9645), .B2(n11794), .ZN(
        n7418) );
  OAI22_X1 U3954 ( .A1(n10722), .A2(n11788), .B1(n9613), .B2(n11794), .ZN(
        n7417) );
  OAI22_X1 U3955 ( .A1(n10715), .A2(n11788), .B1(n9581), .B2(n11794), .ZN(
        n7416) );
  OAI22_X1 U3956 ( .A1(n10708), .A2(n11787), .B1(n9215), .B2(n11795), .ZN(
        n7415) );
  OAI22_X1 U3957 ( .A1(n10701), .A2(n11787), .B1(n9183), .B2(n11795), .ZN(
        n7414) );
  OAI22_X1 U3958 ( .A1(n10694), .A2(n11787), .B1(n9151), .B2(n11795), .ZN(
        n7413) );
  OAI22_X1 U3959 ( .A1(n10687), .A2(n11787), .B1(n6301), .B2(n11795), .ZN(
        n7412) );
  OAI22_X1 U3960 ( .A1(n10680), .A2(n11787), .B1(n5984), .B2(n11796), .ZN(
        n7411) );
  OAI22_X1 U3961 ( .A1(n10673), .A2(n11787), .B1(n5920), .B2(n11796), .ZN(
        n7410) );
  OAI22_X1 U3962 ( .A1(n10666), .A2(n11787), .B1(n5888), .B2(n11796), .ZN(
        n7409) );
  OAI22_X1 U3963 ( .A1(n10659), .A2(n11787), .B1(n5856), .B2(n11796), .ZN(
        n7408) );
  OAI22_X1 U3964 ( .A1(n10652), .A2(n11787), .B1(n5824), .B2(n11797), .ZN(
        n7407) );
  OAI22_X1 U3965 ( .A1(n10645), .A2(n11787), .B1(n5792), .B2(n11797), .ZN(
        n7406) );
  OAI22_X1 U3966 ( .A1(n10638), .A2(n11787), .B1(n5760), .B2(n11797), .ZN(
        n7405) );
  OAI22_X1 U3967 ( .A1(n10631), .A2(n11787), .B1(n5728), .B2(n11797), .ZN(
        n7404) );
  OAI22_X1 U3968 ( .A1(n10849), .A2(n11525), .B1(n10535), .B2(n11526), .ZN(
        n6731) );
  OAI22_X1 U3969 ( .A1(n10842), .A2(n11525), .B1(n10503), .B2(n11526), .ZN(
        n6730) );
  OAI22_X1 U3970 ( .A1(n10835), .A2(n11525), .B1(n10471), .B2(n11526), .ZN(
        n6729) );
  OAI22_X1 U3971 ( .A1(n10828), .A2(n11525), .B1(n10439), .B2(n11526), .ZN(
        n6728) );
  OAI22_X1 U3972 ( .A1(n10821), .A2(n11525), .B1(n10407), .B2(n11527), .ZN(
        n6727) );
  OAI22_X1 U3973 ( .A1(n10814), .A2(n11525), .B1(n10372), .B2(n11527), .ZN(
        n6726) );
  OAI22_X1 U3974 ( .A1(n10807), .A2(n11525), .B1(n10340), .B2(n11527), .ZN(
        n6725) );
  OAI22_X1 U3975 ( .A1(n10800), .A2(n11525), .B1(n10308), .B2(n11527), .ZN(
        n6724) );
  OAI22_X1 U3976 ( .A1(n10793), .A2(n11524), .B1(n10273), .B2(n11528), .ZN(
        n6723) );
  OAI22_X1 U3977 ( .A1(n10786), .A2(n11524), .B1(n10241), .B2(n11528), .ZN(
        n6722) );
  OAI22_X1 U3978 ( .A1(n10779), .A2(n11524), .B1(n10209), .B2(n11528), .ZN(
        n6721) );
  OAI22_X1 U3979 ( .A1(n10772), .A2(n11524), .B1(n10175), .B2(n11528), .ZN(
        n6720) );
  OAI22_X1 U3980 ( .A1(n10765), .A2(n11524), .B1(n10143), .B2(n11529), .ZN(
        n6719) );
  OAI22_X1 U3981 ( .A1(n10758), .A2(n11524), .B1(n10111), .B2(n11529), .ZN(
        n6718) );
  OAI22_X1 U3982 ( .A1(n10751), .A2(n11524), .B1(n10079), .B2(n11529), .ZN(
        n6717) );
  OAI22_X1 U3983 ( .A1(n10744), .A2(n11524), .B1(n10047), .B2(n11529), .ZN(
        n6716) );
  OAI22_X1 U3984 ( .A1(n10737), .A2(n11524), .B1(n10015), .B2(n11530), .ZN(
        n6715) );
  OAI22_X1 U3985 ( .A1(n10730), .A2(n11524), .B1(n9653), .B2(n11530), .ZN(
        n6714) );
  OAI22_X1 U3986 ( .A1(n10723), .A2(n11524), .B1(n9621), .B2(n11530), .ZN(
        n6713) );
  OAI22_X1 U3987 ( .A1(n10716), .A2(n11524), .B1(n9589), .B2(n11530), .ZN(
        n6712) );
  OAI22_X1 U3988 ( .A1(n10709), .A2(n11523), .B1(n9255), .B2(n11531), .ZN(
        n6711) );
  OAI22_X1 U3989 ( .A1(n10702), .A2(n11523), .B1(n9191), .B2(n11531), .ZN(
        n6710) );
  OAI22_X1 U3990 ( .A1(n10695), .A2(n11523), .B1(n9159), .B2(n11531), .ZN(
        n6709) );
  OAI22_X1 U3991 ( .A1(n10688), .A2(n11523), .B1(n6309), .B2(n11531), .ZN(
        n6708) );
  OAI22_X1 U3992 ( .A1(n10681), .A2(n11523), .B1(n5992), .B2(n11532), .ZN(
        n6707) );
  OAI22_X1 U3993 ( .A1(n10674), .A2(n11523), .B1(n5928), .B2(n11532), .ZN(
        n6706) );
  OAI22_X1 U3994 ( .A1(n10667), .A2(n11523), .B1(n5896), .B2(n11532), .ZN(
        n6705) );
  OAI22_X1 U3995 ( .A1(n10660), .A2(n11523), .B1(n5864), .B2(n11532), .ZN(
        n6704) );
  OAI22_X1 U3996 ( .A1(n10653), .A2(n11523), .B1(n5832), .B2(n11533), .ZN(
        n6703) );
  OAI22_X1 U3997 ( .A1(n10646), .A2(n11523), .B1(n5800), .B2(n11533), .ZN(
        n6702) );
  OAI22_X1 U3998 ( .A1(n10639), .A2(n11523), .B1(n5768), .B2(n11533), .ZN(
        n6701) );
  OAI22_X1 U3999 ( .A1(n10632), .A2(n11523), .B1(n5736), .B2(n11533), .ZN(
        n6700) );
  OAI22_X1 U4000 ( .A1(n10850), .A2(n11477), .B1(n1409), .B2(n11478), .ZN(
        n6603) );
  OAI22_X1 U4001 ( .A1(n10843), .A2(n11477), .B1(n1397), .B2(n11478), .ZN(
        n6602) );
  OAI22_X1 U4002 ( .A1(n10836), .A2(n11477), .B1(n1385), .B2(n11478), .ZN(
        n6601) );
  OAI22_X1 U4003 ( .A1(n10829), .A2(n11477), .B1(n1341), .B2(n11478), .ZN(
        n6600) );
  OAI22_X1 U4004 ( .A1(n10822), .A2(n11477), .B1(n1329), .B2(n11479), .ZN(
        n6599) );
  OAI22_X1 U4005 ( .A1(n10815), .A2(n11477), .B1(n1317), .B2(n11479), .ZN(
        n6598) );
  OAI22_X1 U4006 ( .A1(n10808), .A2(n11477), .B1(n1305), .B2(n11479), .ZN(
        n6597) );
  OAI22_X1 U4007 ( .A1(n10801), .A2(n11477), .B1(n1293), .B2(n11479), .ZN(
        n6596) );
  OAI22_X1 U4008 ( .A1(n10794), .A2(n11476), .B1(n1281), .B2(n11480), .ZN(
        n6595) );
  OAI22_X1 U4009 ( .A1(n10787), .A2(n11476), .B1(n1269), .B2(n11480), .ZN(
        n6594) );
  OAI22_X1 U4010 ( .A1(n10780), .A2(n11476), .B1(n1257), .B2(n11480), .ZN(
        n6593) );
  OAI22_X1 U4011 ( .A1(n10773), .A2(n11476), .B1(n1245), .B2(n11480), .ZN(
        n6592) );
  OAI22_X1 U4012 ( .A1(n10766), .A2(n11476), .B1(n1233), .B2(n11481), .ZN(
        n6591) );
  OAI22_X1 U4013 ( .A1(n10759), .A2(n11476), .B1(n1221), .B2(n11481), .ZN(
        n6590) );
  OAI22_X1 U4014 ( .A1(n10752), .A2(n11476), .B1(n1209), .B2(n11481), .ZN(
        n6589) );
  OAI22_X1 U4015 ( .A1(n10745), .A2(n11476), .B1(n1197), .B2(n11481), .ZN(
        n6588) );
  OAI22_X1 U4016 ( .A1(n10738), .A2(n11476), .B1(n1185), .B2(n11482), .ZN(
        n6587) );
  OAI22_X1 U4017 ( .A1(n10731), .A2(n11476), .B1(n1173), .B2(n11482), .ZN(
        n6586) );
  OAI22_X1 U4018 ( .A1(n10724), .A2(n11476), .B1(n1161), .B2(n11482), .ZN(
        n6585) );
  OAI22_X1 U4019 ( .A1(n10717), .A2(n11476), .B1(n1149), .B2(n11482), .ZN(
        n6584) );
  OAI22_X1 U4020 ( .A1(n10710), .A2(n11475), .B1(n1137), .B2(n11483), .ZN(
        n6583) );
  OAI22_X1 U4021 ( .A1(n10703), .A2(n11475), .B1(n1125), .B2(n11483), .ZN(
        n6582) );
  OAI22_X1 U4022 ( .A1(n10696), .A2(n11475), .B1(n1113), .B2(n11483), .ZN(
        n6581) );
  OAI22_X1 U4023 ( .A1(n10689), .A2(n11475), .B1(n1101), .B2(n11483), .ZN(
        n6580) );
  OAI22_X1 U4024 ( .A1(n10682), .A2(n11475), .B1(n1089), .B2(n11484), .ZN(
        n6579) );
  OAI22_X1 U4025 ( .A1(n10675), .A2(n11475), .B1(n1077), .B2(n11484), .ZN(
        n6578) );
  OAI22_X1 U4026 ( .A1(n10668), .A2(n11475), .B1(n1065), .B2(n11484), .ZN(
        n6577) );
  OAI22_X1 U4027 ( .A1(n10661), .A2(n11475), .B1(n1053), .B2(n11484), .ZN(
        n6576) );
  OAI22_X1 U4028 ( .A1(n10654), .A2(n11475), .B1(n1041), .B2(n11485), .ZN(
        n6575) );
  OAI22_X1 U4029 ( .A1(n10647), .A2(n11475), .B1(n1029), .B2(n11485), .ZN(
        n6574) );
  OAI22_X1 U4030 ( .A1(n10850), .A2(n11441), .B1(n1442), .B2(n11442), .ZN(
        n6507) );
  OAI22_X1 U4031 ( .A1(n10843), .A2(n11441), .B1(n1398), .B2(n11442), .ZN(
        n6506) );
  OAI22_X1 U4032 ( .A1(n10836), .A2(n11441), .B1(n1386), .B2(n11442), .ZN(
        n6505) );
  OAI22_X1 U4033 ( .A1(n10829), .A2(n11441), .B1(n1342), .B2(n11442), .ZN(
        n6504) );
  OAI22_X1 U4034 ( .A1(n10822), .A2(n11441), .B1(n1330), .B2(n11443), .ZN(
        n6503) );
  OAI22_X1 U4035 ( .A1(n10815), .A2(n11441), .B1(n1318), .B2(n11443), .ZN(
        n6502) );
  OAI22_X1 U4036 ( .A1(n10808), .A2(n11441), .B1(n1306), .B2(n11443), .ZN(
        n6501) );
  OAI22_X1 U4037 ( .A1(n10801), .A2(n11441), .B1(n1294), .B2(n11443), .ZN(
        n6500) );
  OAI22_X1 U4038 ( .A1(n10794), .A2(n11440), .B1(n1282), .B2(n11444), .ZN(
        n6499) );
  OAI22_X1 U4039 ( .A1(n10787), .A2(n11440), .B1(n1270), .B2(n11444), .ZN(
        n6498) );
  OAI22_X1 U4040 ( .A1(n10780), .A2(n11440), .B1(n1258), .B2(n11444), .ZN(
        n6497) );
  OAI22_X1 U4041 ( .A1(n10773), .A2(n11440), .B1(n1246), .B2(n11444), .ZN(
        n6496) );
  OAI22_X1 U4042 ( .A1(n10766), .A2(n11440), .B1(n1234), .B2(n11445), .ZN(
        n6495) );
  OAI22_X1 U4043 ( .A1(n10759), .A2(n11440), .B1(n1222), .B2(n11445), .ZN(
        n6494) );
  OAI22_X1 U4044 ( .A1(n10752), .A2(n11440), .B1(n1210), .B2(n11445), .ZN(
        n6493) );
  OAI22_X1 U4045 ( .A1(n10745), .A2(n11440), .B1(n1198), .B2(n11445), .ZN(
        n6492) );
  OAI22_X1 U4046 ( .A1(n10738), .A2(n11440), .B1(n1186), .B2(n11446), .ZN(
        n6491) );
  OAI22_X1 U4047 ( .A1(n10731), .A2(n11440), .B1(n1174), .B2(n11446), .ZN(
        n6490) );
  OAI22_X1 U4048 ( .A1(n10724), .A2(n11440), .B1(n1162), .B2(n11446), .ZN(
        n6489) );
  OAI22_X1 U4049 ( .A1(n10717), .A2(n11440), .B1(n1150), .B2(n11446), .ZN(
        n6488) );
  OAI22_X1 U4050 ( .A1(n10710), .A2(n11439), .B1(n1138), .B2(n11447), .ZN(
        n6487) );
  OAI22_X1 U4051 ( .A1(n10703), .A2(n11439), .B1(n1126), .B2(n11447), .ZN(
        n6486) );
  OAI22_X1 U4052 ( .A1(n10696), .A2(n11439), .B1(n1114), .B2(n11447), .ZN(
        n6485) );
  OAI22_X1 U4053 ( .A1(n10689), .A2(n11439), .B1(n1102), .B2(n11447), .ZN(
        n6484) );
  OAI22_X1 U4054 ( .A1(n10682), .A2(n11439), .B1(n1090), .B2(n11448), .ZN(
        n6483) );
  OAI22_X1 U4055 ( .A1(n10675), .A2(n11439), .B1(n1078), .B2(n11448), .ZN(
        n6482) );
  OAI22_X1 U4056 ( .A1(n10668), .A2(n11439), .B1(n1066), .B2(n11448), .ZN(
        n6481) );
  OAI22_X1 U4057 ( .A1(n10661), .A2(n11439), .B1(n1054), .B2(n11448), .ZN(
        n6480) );
  OAI22_X1 U4058 ( .A1(n10654), .A2(n11439), .B1(n1042), .B2(n11449), .ZN(
        n6479) );
  OAI22_X1 U4059 ( .A1(n10850), .A2(n11405), .B1(n1443), .B2(n11406), .ZN(
        n6411) );
  OAI22_X1 U4060 ( .A1(n10843), .A2(n11405), .B1(n1399), .B2(n11406), .ZN(
        n6410) );
  OAI22_X1 U4061 ( .A1(n10836), .A2(n11405), .B1(n1387), .B2(n11406), .ZN(
        n6409) );
  OAI22_X1 U4062 ( .A1(n10829), .A2(n11405), .B1(n1343), .B2(n11406), .ZN(
        n6408) );
  OAI22_X1 U4063 ( .A1(n10822), .A2(n11405), .B1(n1331), .B2(n11407), .ZN(
        n6407) );
  OAI22_X1 U4064 ( .A1(n10815), .A2(n11405), .B1(n1319), .B2(n11407), .ZN(
        n6406) );
  OAI22_X1 U4065 ( .A1(n10808), .A2(n11405), .B1(n1307), .B2(n11407), .ZN(
        n6405) );
  OAI22_X1 U4066 ( .A1(n10801), .A2(n11405), .B1(n1295), .B2(n11407), .ZN(
        n6404) );
  OAI22_X1 U4067 ( .A1(n10794), .A2(n11404), .B1(n1283), .B2(n11408), .ZN(
        n6403) );
  OAI22_X1 U4068 ( .A1(n10787), .A2(n11404), .B1(n1271), .B2(n11408), .ZN(
        n6402) );
  OAI22_X1 U4069 ( .A1(n10780), .A2(n11404), .B1(n1259), .B2(n11408), .ZN(
        n6401) );
  OAI22_X1 U4070 ( .A1(n10773), .A2(n11404), .B1(n1247), .B2(n11408), .ZN(
        n6400) );
  OAI22_X1 U4071 ( .A1(n10766), .A2(n11404), .B1(n1235), .B2(n11409), .ZN(
        n6399) );
  OAI22_X1 U4072 ( .A1(n10759), .A2(n11404), .B1(n1223), .B2(n11409), .ZN(
        n6398) );
  OAI22_X1 U4073 ( .A1(n10752), .A2(n11404), .B1(n1211), .B2(n11409), .ZN(
        n6397) );
  OAI22_X1 U4074 ( .A1(n10745), .A2(n11404), .B1(n1199), .B2(n11409), .ZN(
        n6396) );
  OAI22_X1 U4075 ( .A1(n10738), .A2(n11404), .B1(n1187), .B2(n11410), .ZN(
        n6395) );
  OAI22_X1 U4076 ( .A1(n10731), .A2(n11404), .B1(n1175), .B2(n11410), .ZN(
        n6394) );
  OAI22_X1 U4077 ( .A1(n10724), .A2(n11404), .B1(n1163), .B2(n11410), .ZN(
        n6393) );
  OAI22_X1 U4078 ( .A1(n10717), .A2(n11404), .B1(n1151), .B2(n11410), .ZN(
        n6392) );
  OAI22_X1 U4079 ( .A1(n10710), .A2(n11403), .B1(n1139), .B2(n11411), .ZN(
        n6391) );
  OAI22_X1 U4080 ( .A1(n10703), .A2(n11403), .B1(n1127), .B2(n11411), .ZN(
        n6390) );
  OAI22_X1 U4081 ( .A1(n10696), .A2(n11403), .B1(n1115), .B2(n11411), .ZN(
        n6389) );
  OAI22_X1 U4082 ( .A1(n10689), .A2(n11403), .B1(n1103), .B2(n11411), .ZN(
        n6388) );
  OAI22_X1 U4083 ( .A1(n10682), .A2(n11403), .B1(n1091), .B2(n11412), .ZN(
        n6387) );
  OAI22_X1 U4084 ( .A1(n10675), .A2(n11403), .B1(n1079), .B2(n11412), .ZN(
        n6386) );
  OAI22_X1 U4085 ( .A1(n10668), .A2(n11403), .B1(n1067), .B2(n11412), .ZN(
        n6385) );
  OAI22_X1 U4086 ( .A1(n10661), .A2(n11403), .B1(n1055), .B2(n11412), .ZN(
        n6384) );
  OAI22_X1 U4087 ( .A1(n10654), .A2(n11403), .B1(n1043), .B2(n11413), .ZN(
        n6383) );
  OAI22_X1 U4088 ( .A1(n10844), .A2(n12329), .B1(n10509), .B2(n12330), .ZN(
        n8875) );
  OAI22_X1 U4089 ( .A1(n10837), .A2(n12329), .B1(n10477), .B2(n12330), .ZN(
        n8874) );
  OAI22_X1 U4090 ( .A1(n10830), .A2(n12329), .B1(n10445), .B2(n12330), .ZN(
        n8873) );
  OAI22_X1 U4091 ( .A1(n10823), .A2(n12329), .B1(n10413), .B2(n12330), .ZN(
        n8872) );
  OAI22_X1 U4092 ( .A1(n10816), .A2(n12329), .B1(n10378), .B2(n12331), .ZN(
        n8871) );
  OAI22_X1 U4093 ( .A1(n10809), .A2(n12329), .B1(n10346), .B2(n12331), .ZN(
        n8870) );
  OAI22_X1 U4094 ( .A1(n10802), .A2(n12329), .B1(n10314), .B2(n12331), .ZN(
        n8869) );
  OAI22_X1 U4095 ( .A1(n10795), .A2(n12329), .B1(n10279), .B2(n12331), .ZN(
        n8868) );
  OAI22_X1 U4096 ( .A1(n10788), .A2(n12328), .B1(n10247), .B2(n12332), .ZN(
        n8867) );
  OAI22_X1 U4097 ( .A1(n10781), .A2(n12328), .B1(n10215), .B2(n12332), .ZN(
        n8866) );
  OAI22_X1 U4098 ( .A1(n10774), .A2(n12328), .B1(n10181), .B2(n12332), .ZN(
        n8865) );
  OAI22_X1 U4099 ( .A1(n10767), .A2(n12328), .B1(n10149), .B2(n12332), .ZN(
        n8864) );
  OAI22_X1 U4100 ( .A1(n10760), .A2(n12328), .B1(n10117), .B2(n12333), .ZN(
        n8863) );
  OAI22_X1 U4101 ( .A1(n10753), .A2(n12328), .B1(n10085), .B2(n12333), .ZN(
        n8862) );
  OAI22_X1 U4102 ( .A1(n10746), .A2(n12328), .B1(n10053), .B2(n12333), .ZN(
        n8861) );
  OAI22_X1 U4103 ( .A1(n10739), .A2(n12328), .B1(n10021), .B2(n12333), .ZN(
        n8860) );
  OAI22_X1 U4104 ( .A1(n10732), .A2(n12328), .B1(n9659), .B2(n12334), .ZN(
        n8859) );
  OAI22_X1 U4105 ( .A1(n10725), .A2(n12328), .B1(n9627), .B2(n12334), .ZN(
        n8858) );
  OAI22_X1 U4106 ( .A1(n10718), .A2(n12328), .B1(n9595), .B2(n12334), .ZN(
        n8857) );
  OAI22_X1 U4107 ( .A1(n10711), .A2(n12328), .B1(n9261), .B2(n12334), .ZN(
        n8856) );
  OAI22_X1 U4108 ( .A1(n10704), .A2(n12327), .B1(n9197), .B2(n12335), .ZN(
        n8855) );
  OAI22_X1 U4109 ( .A1(n10697), .A2(n12327), .B1(n9165), .B2(n12335), .ZN(
        n8854) );
  OAI22_X1 U4110 ( .A1(n10690), .A2(n12327), .B1(n6315), .B2(n12335), .ZN(
        n8853) );
  OAI22_X1 U4111 ( .A1(n10683), .A2(n12327), .B1(n5998), .B2(n12335), .ZN(
        n8852) );
  OAI22_X1 U4112 ( .A1(n10676), .A2(n12327), .B1(n5934), .B2(n12336), .ZN(
        n8851) );
  OAI22_X1 U4113 ( .A1(n10669), .A2(n12327), .B1(n5902), .B2(n12336), .ZN(
        n8850) );
  OAI22_X1 U4114 ( .A1(n10662), .A2(n12327), .B1(n5870), .B2(n12336), .ZN(
        n8849) );
  OAI22_X1 U4115 ( .A1(n10655), .A2(n12327), .B1(n5838), .B2(n12336), .ZN(
        n8848) );
  OAI22_X1 U4116 ( .A1(n10648), .A2(n12327), .B1(n5806), .B2(n12337), .ZN(
        n8847) );
  OAI22_X1 U4117 ( .A1(n10641), .A2(n12327), .B1(n5774), .B2(n12337), .ZN(
        n8846) );
  OAI22_X1 U4118 ( .A1(n10634), .A2(n12327), .B1(n5742), .B2(n12337), .ZN(
        n8845) );
  OAI22_X1 U4119 ( .A1(n10627), .A2(n12327), .B1(n5710), .B2(n12337), .ZN(
        n8844) );
  OAI22_X1 U4120 ( .A1(n10846), .A2(n12101), .B1(n10514), .B2(n12102), .ZN(
        n8267) );
  OAI22_X1 U4121 ( .A1(n10839), .A2(n12101), .B1(n10482), .B2(n12102), .ZN(
        n8266) );
  OAI22_X1 U4122 ( .A1(n10832), .A2(n12101), .B1(n10450), .B2(n12102), .ZN(
        n8265) );
  OAI22_X1 U4123 ( .A1(n10825), .A2(n12101), .B1(n10418), .B2(n12102), .ZN(
        n8264) );
  OAI22_X1 U4124 ( .A1(n10818), .A2(n12101), .B1(n10383), .B2(n12103), .ZN(
        n8263) );
  OAI22_X1 U4125 ( .A1(n10811), .A2(n12101), .B1(n10351), .B2(n12103), .ZN(
        n8262) );
  OAI22_X1 U4126 ( .A1(n10804), .A2(n12101), .B1(n10319), .B2(n12103), .ZN(
        n8261) );
  OAI22_X1 U4127 ( .A1(n10797), .A2(n12101), .B1(n10284), .B2(n12103), .ZN(
        n8260) );
  OAI22_X1 U4128 ( .A1(n10790), .A2(n12100), .B1(n10252), .B2(n12104), .ZN(
        n8259) );
  OAI22_X1 U4129 ( .A1(n10783), .A2(n12100), .B1(n10220), .B2(n12104), .ZN(
        n8258) );
  OAI22_X1 U4130 ( .A1(n10776), .A2(n12100), .B1(n10186), .B2(n12104), .ZN(
        n8257) );
  OAI22_X1 U4131 ( .A1(n10769), .A2(n12100), .B1(n10154), .B2(n12104), .ZN(
        n8256) );
  OAI22_X1 U4132 ( .A1(n10762), .A2(n12100), .B1(n10122), .B2(n12105), .ZN(
        n8255) );
  OAI22_X1 U4133 ( .A1(n10755), .A2(n12100), .B1(n10090), .B2(n12105), .ZN(
        n8254) );
  OAI22_X1 U4134 ( .A1(n10748), .A2(n12100), .B1(n10058), .B2(n12105), .ZN(
        n8253) );
  OAI22_X1 U4135 ( .A1(n10741), .A2(n12100), .B1(n10026), .B2(n12105), .ZN(
        n8252) );
  OAI22_X1 U4136 ( .A1(n10734), .A2(n12100), .B1(n9696), .B2(n12106), .ZN(
        n8251) );
  OAI22_X1 U4137 ( .A1(n10727), .A2(n12100), .B1(n9632), .B2(n12106), .ZN(
        n8250) );
  OAI22_X1 U4138 ( .A1(n10720), .A2(n12100), .B1(n9600), .B2(n12106), .ZN(
        n8249) );
  OAI22_X1 U4139 ( .A1(n10713), .A2(n12100), .B1(n9568), .B2(n12106), .ZN(
        n8248) );
  OAI22_X1 U4140 ( .A1(n10706), .A2(n12099), .B1(n9202), .B2(n12107), .ZN(
        n8247) );
  OAI22_X1 U4141 ( .A1(n10699), .A2(n12099), .B1(n9170), .B2(n12107), .ZN(
        n8246) );
  OAI22_X1 U4142 ( .A1(n10692), .A2(n12099), .B1(n9138), .B2(n12107), .ZN(
        n8245) );
  OAI22_X1 U4143 ( .A1(n10685), .A2(n12099), .B1(n6003), .B2(n12107), .ZN(
        n8244) );
  OAI22_X1 U4144 ( .A1(n10678), .A2(n12099), .B1(n5939), .B2(n12108), .ZN(
        n8243) );
  OAI22_X1 U4145 ( .A1(n10671), .A2(n12099), .B1(n5907), .B2(n12108), .ZN(
        n8242) );
  OAI22_X1 U4146 ( .A1(n10664), .A2(n12099), .B1(n5875), .B2(n12108), .ZN(
        n8241) );
  OAI22_X1 U4147 ( .A1(n10657), .A2(n12099), .B1(n5843), .B2(n12108), .ZN(
        n8240) );
  OAI22_X1 U4148 ( .A1(n10650), .A2(n12099), .B1(n5811), .B2(n12109), .ZN(
        n8239) );
  OAI22_X1 U4149 ( .A1(n10643), .A2(n12099), .B1(n5779), .B2(n12109), .ZN(
        n8238) );
  OAI22_X1 U4150 ( .A1(n10636), .A2(n12099), .B1(n5747), .B2(n12109), .ZN(
        n8237) );
  OAI22_X1 U4151 ( .A1(n10629), .A2(n12099), .B1(n5715), .B2(n12109), .ZN(
        n8236) );
  OAI22_X1 U4152 ( .A1(n10846), .A2(n12065), .B1(n10517), .B2(n12066), .ZN(
        n8171) );
  OAI22_X1 U4153 ( .A1(n10839), .A2(n12065), .B1(n10485), .B2(n12066), .ZN(
        n8170) );
  OAI22_X1 U4154 ( .A1(n10832), .A2(n12065), .B1(n10453), .B2(n12066), .ZN(
        n8169) );
  OAI22_X1 U4155 ( .A1(n10825), .A2(n12065), .B1(n10421), .B2(n12066), .ZN(
        n8168) );
  OAI22_X1 U4156 ( .A1(n10818), .A2(n12065), .B1(n10386), .B2(n12067), .ZN(
        n8167) );
  OAI22_X1 U4157 ( .A1(n10811), .A2(n12065), .B1(n10354), .B2(n12067), .ZN(
        n8166) );
  OAI22_X1 U4158 ( .A1(n10804), .A2(n12065), .B1(n10322), .B2(n12067), .ZN(
        n8165) );
  OAI22_X1 U4159 ( .A1(n10797), .A2(n12065), .B1(n10287), .B2(n12067), .ZN(
        n8164) );
  OAI22_X1 U4160 ( .A1(n10790), .A2(n12064), .B1(n10255), .B2(n12068), .ZN(
        n8163) );
  OAI22_X1 U4161 ( .A1(n10783), .A2(n12064), .B1(n10223), .B2(n12068), .ZN(
        n8162) );
  OAI22_X1 U4162 ( .A1(n10776), .A2(n12064), .B1(n10189), .B2(n12068), .ZN(
        n8161) );
  OAI22_X1 U4163 ( .A1(n10769), .A2(n12064), .B1(n10157), .B2(n12068), .ZN(
        n8160) );
  OAI22_X1 U4164 ( .A1(n10762), .A2(n12064), .B1(n10125), .B2(n12069), .ZN(
        n8159) );
  OAI22_X1 U4165 ( .A1(n10755), .A2(n12064), .B1(n10093), .B2(n12069), .ZN(
        n8158) );
  OAI22_X1 U4166 ( .A1(n10748), .A2(n12064), .B1(n10061), .B2(n12069), .ZN(
        n8157) );
  OAI22_X1 U4167 ( .A1(n10741), .A2(n12064), .B1(n10029), .B2(n12069), .ZN(
        n8156) );
  OAI22_X1 U4168 ( .A1(n10734), .A2(n12064), .B1(n9699), .B2(n12070), .ZN(
        n8155) );
  OAI22_X1 U4169 ( .A1(n10727), .A2(n12064), .B1(n9635), .B2(n12070), .ZN(
        n8154) );
  OAI22_X1 U4170 ( .A1(n10720), .A2(n12064), .B1(n9603), .B2(n12070), .ZN(
        n8153) );
  OAI22_X1 U4171 ( .A1(n10713), .A2(n12064), .B1(n9571), .B2(n12070), .ZN(
        n8152) );
  OAI22_X1 U4172 ( .A1(n10706), .A2(n12063), .B1(n9205), .B2(n12071), .ZN(
        n8151) );
  OAI22_X1 U4173 ( .A1(n10699), .A2(n12063), .B1(n9173), .B2(n12071), .ZN(
        n8150) );
  OAI22_X1 U4174 ( .A1(n10692), .A2(n12063), .B1(n9141), .B2(n12071), .ZN(
        n8149) );
  OAI22_X1 U4175 ( .A1(n10685), .A2(n12063), .B1(n6006), .B2(n12071), .ZN(
        n8148) );
  OAI22_X1 U4176 ( .A1(n10678), .A2(n12063), .B1(n5942), .B2(n12072), .ZN(
        n8147) );
  OAI22_X1 U4177 ( .A1(n10671), .A2(n12063), .B1(n5910), .B2(n12072), .ZN(
        n8146) );
  OAI22_X1 U4178 ( .A1(n10664), .A2(n12063), .B1(n5878), .B2(n12072), .ZN(
        n8145) );
  OAI22_X1 U4179 ( .A1(n10657), .A2(n12063), .B1(n5846), .B2(n12072), .ZN(
        n8144) );
  OAI22_X1 U4180 ( .A1(n10650), .A2(n12063), .B1(n5814), .B2(n12073), .ZN(
        n8143) );
  OAI22_X1 U4181 ( .A1(n10643), .A2(n12063), .B1(n5782), .B2(n12073), .ZN(
        n8142) );
  OAI22_X1 U4182 ( .A1(n10636), .A2(n12063), .B1(n5750), .B2(n12073), .ZN(
        n8141) );
  OAI22_X1 U4183 ( .A1(n10629), .A2(n12063), .B1(n5718), .B2(n12073), .ZN(
        n8140) );
  OAI22_X1 U4184 ( .A1(n10847), .A2(n11837), .B1(n10522), .B2(n11838), .ZN(
        n7563) );
  OAI22_X1 U4185 ( .A1(n10840), .A2(n11837), .B1(n10490), .B2(n11838), .ZN(
        n7562) );
  OAI22_X1 U4186 ( .A1(n10833), .A2(n11837), .B1(n10458), .B2(n11838), .ZN(
        n7561) );
  OAI22_X1 U4187 ( .A1(n10826), .A2(n11837), .B1(n10426), .B2(n11838), .ZN(
        n7560) );
  OAI22_X1 U4188 ( .A1(n10819), .A2(n11837), .B1(n10391), .B2(n11839), .ZN(
        n7559) );
  OAI22_X1 U4189 ( .A1(n10812), .A2(n11837), .B1(n10359), .B2(n11839), .ZN(
        n7558) );
  OAI22_X1 U4190 ( .A1(n10805), .A2(n11837), .B1(n10327), .B2(n11839), .ZN(
        n7557) );
  OAI22_X1 U4191 ( .A1(n10798), .A2(n11837), .B1(n10292), .B2(n11839), .ZN(
        n7556) );
  OAI22_X1 U4192 ( .A1(n10791), .A2(n11836), .B1(n10260), .B2(n11840), .ZN(
        n7555) );
  OAI22_X1 U4193 ( .A1(n10784), .A2(n11836), .B1(n10228), .B2(n11840), .ZN(
        n7554) );
  OAI22_X1 U4194 ( .A1(n10777), .A2(n11836), .B1(n10194), .B2(n11840), .ZN(
        n7553) );
  OAI22_X1 U4195 ( .A1(n10770), .A2(n11836), .B1(n10162), .B2(n11840), .ZN(
        n7552) );
  OAI22_X1 U4196 ( .A1(n10763), .A2(n11836), .B1(n10130), .B2(n11841), .ZN(
        n7551) );
  OAI22_X1 U4197 ( .A1(n10756), .A2(n11836), .B1(n10098), .B2(n11841), .ZN(
        n7550) );
  OAI22_X1 U4198 ( .A1(n10749), .A2(n11836), .B1(n10066), .B2(n11841), .ZN(
        n7549) );
  OAI22_X1 U4199 ( .A1(n10742), .A2(n11836), .B1(n10034), .B2(n11841), .ZN(
        n7548) );
  OAI22_X1 U4200 ( .A1(n10735), .A2(n11836), .B1(n10002), .B2(n11842), .ZN(
        n7547) );
  OAI22_X1 U4201 ( .A1(n10728), .A2(n11836), .B1(n9640), .B2(n11842), .ZN(
        n7546) );
  OAI22_X1 U4202 ( .A1(n10721), .A2(n11836), .B1(n9608), .B2(n11842), .ZN(
        n7545) );
  OAI22_X1 U4203 ( .A1(n10714), .A2(n11836), .B1(n9576), .B2(n11842), .ZN(
        n7544) );
  OAI22_X1 U4204 ( .A1(n10707), .A2(n11835), .B1(n9210), .B2(n11843), .ZN(
        n7543) );
  OAI22_X1 U4205 ( .A1(n10700), .A2(n11835), .B1(n9178), .B2(n11843), .ZN(
        n7542) );
  OAI22_X1 U4206 ( .A1(n10693), .A2(n11835), .B1(n9146), .B2(n11843), .ZN(
        n7541) );
  OAI22_X1 U4207 ( .A1(n10686), .A2(n11835), .B1(n6011), .B2(n11843), .ZN(
        n7540) );
  OAI22_X1 U4208 ( .A1(n10679), .A2(n11835), .B1(n5947), .B2(n11844), .ZN(
        n7539) );
  OAI22_X1 U4209 ( .A1(n10672), .A2(n11835), .B1(n5915), .B2(n11844), .ZN(
        n7538) );
  OAI22_X1 U4210 ( .A1(n10665), .A2(n11835), .B1(n5883), .B2(n11844), .ZN(
        n7537) );
  OAI22_X1 U4211 ( .A1(n10658), .A2(n11835), .B1(n5851), .B2(n11844), .ZN(
        n7536) );
  OAI22_X1 U4212 ( .A1(n10651), .A2(n11835), .B1(n5819), .B2(n11845), .ZN(
        n7535) );
  OAI22_X1 U4213 ( .A1(n10644), .A2(n11835), .B1(n5787), .B2(n11845), .ZN(
        n7534) );
  OAI22_X1 U4214 ( .A1(n10637), .A2(n11835), .B1(n5755), .B2(n11845), .ZN(
        n7533) );
  OAI22_X1 U4215 ( .A1(n10630), .A2(n11835), .B1(n5723), .B2(n11845), .ZN(
        n7532) );
  OAI22_X1 U4216 ( .A1(n10848), .A2(n11801), .B1(n10525), .B2(n11802), .ZN(
        n7467) );
  OAI22_X1 U4217 ( .A1(n10841), .A2(n11801), .B1(n10493), .B2(n11802), .ZN(
        n7466) );
  OAI22_X1 U4218 ( .A1(n10834), .A2(n11801), .B1(n10461), .B2(n11802), .ZN(
        n7465) );
  OAI22_X1 U4219 ( .A1(n10827), .A2(n11801), .B1(n10429), .B2(n11802), .ZN(
        n7464) );
  OAI22_X1 U4220 ( .A1(n10820), .A2(n11801), .B1(n10394), .B2(n11803), .ZN(
        n7463) );
  OAI22_X1 U4221 ( .A1(n10813), .A2(n11801), .B1(n10362), .B2(n11803), .ZN(
        n7462) );
  OAI22_X1 U4222 ( .A1(n10806), .A2(n11801), .B1(n10330), .B2(n11803), .ZN(
        n7461) );
  OAI22_X1 U4223 ( .A1(n10799), .A2(n11801), .B1(n10295), .B2(n11803), .ZN(
        n7460) );
  OAI22_X1 U4224 ( .A1(n10792), .A2(n11800), .B1(n10263), .B2(n11804), .ZN(
        n7459) );
  OAI22_X1 U4225 ( .A1(n10785), .A2(n11800), .B1(n10231), .B2(n11804), .ZN(
        n7458) );
  OAI22_X1 U4226 ( .A1(n10778), .A2(n11800), .B1(n10197), .B2(n11804), .ZN(
        n7457) );
  OAI22_X1 U4227 ( .A1(n10771), .A2(n11800), .B1(n10165), .B2(n11804), .ZN(
        n7456) );
  OAI22_X1 U4228 ( .A1(n10764), .A2(n11800), .B1(n10133), .B2(n11805), .ZN(
        n7455) );
  OAI22_X1 U4229 ( .A1(n10757), .A2(n11800), .B1(n10101), .B2(n11805), .ZN(
        n7454) );
  OAI22_X1 U4230 ( .A1(n10750), .A2(n11800), .B1(n10069), .B2(n11805), .ZN(
        n7453) );
  OAI22_X1 U4231 ( .A1(n10743), .A2(n11800), .B1(n10037), .B2(n11805), .ZN(
        n7452) );
  OAI22_X1 U4232 ( .A1(n10736), .A2(n11800), .B1(n10005), .B2(n11806), .ZN(
        n7451) );
  OAI22_X1 U4233 ( .A1(n10729), .A2(n11800), .B1(n9643), .B2(n11806), .ZN(
        n7450) );
  OAI22_X1 U4234 ( .A1(n10722), .A2(n11800), .B1(n9611), .B2(n11806), .ZN(
        n7449) );
  OAI22_X1 U4235 ( .A1(n10715), .A2(n11800), .B1(n9579), .B2(n11806), .ZN(
        n7448) );
  OAI22_X1 U4236 ( .A1(n10708), .A2(n11799), .B1(n9213), .B2(n11807), .ZN(
        n7447) );
  OAI22_X1 U4237 ( .A1(n10701), .A2(n11799), .B1(n9181), .B2(n11807), .ZN(
        n7446) );
  OAI22_X1 U4238 ( .A1(n10694), .A2(n11799), .B1(n9149), .B2(n11807), .ZN(
        n7445) );
  OAI22_X1 U4239 ( .A1(n10687), .A2(n11799), .B1(n6140), .B2(n11807), .ZN(
        n7444) );
  OAI22_X1 U4240 ( .A1(n10680), .A2(n11799), .B1(n5982), .B2(n11808), .ZN(
        n7443) );
  OAI22_X1 U4241 ( .A1(n10673), .A2(n11799), .B1(n5918), .B2(n11808), .ZN(
        n7442) );
  OAI22_X1 U4242 ( .A1(n10666), .A2(n11799), .B1(n5886), .B2(n11808), .ZN(
        n7441) );
  OAI22_X1 U4243 ( .A1(n10659), .A2(n11799), .B1(n5854), .B2(n11808), .ZN(
        n7440) );
  OAI22_X1 U4244 ( .A1(n10652), .A2(n11799), .B1(n5822), .B2(n11809), .ZN(
        n7439) );
  OAI22_X1 U4245 ( .A1(n10645), .A2(n11799), .B1(n5790), .B2(n11809), .ZN(
        n7438) );
  OAI22_X1 U4246 ( .A1(n10638), .A2(n11799), .B1(n5758), .B2(n11809), .ZN(
        n7437) );
  OAI22_X1 U4247 ( .A1(n10631), .A2(n11799), .B1(n5726), .B2(n11809), .ZN(
        n7436) );
  OAI22_X1 U4248 ( .A1(n10849), .A2(n11537), .B1(n10533), .B2(n11538), .ZN(
        n6763) );
  OAI22_X1 U4249 ( .A1(n10842), .A2(n11537), .B1(n10501), .B2(n11538), .ZN(
        n6762) );
  OAI22_X1 U4250 ( .A1(n10835), .A2(n11537), .B1(n10469), .B2(n11538), .ZN(
        n6761) );
  OAI22_X1 U4251 ( .A1(n10828), .A2(n11537), .B1(n10437), .B2(n11538), .ZN(
        n6760) );
  OAI22_X1 U4252 ( .A1(n10821), .A2(n11537), .B1(n10405), .B2(n11539), .ZN(
        n6759) );
  OAI22_X1 U4253 ( .A1(n10814), .A2(n11537), .B1(n10370), .B2(n11539), .ZN(
        n6758) );
  OAI22_X1 U4254 ( .A1(n10807), .A2(n11537), .B1(n10338), .B2(n11539), .ZN(
        n6757) );
  OAI22_X1 U4255 ( .A1(n10800), .A2(n11537), .B1(n10306), .B2(n11539), .ZN(
        n6756) );
  OAI22_X1 U4256 ( .A1(n10793), .A2(n11536), .B1(n10271), .B2(n11540), .ZN(
        n6755) );
  OAI22_X1 U4257 ( .A1(n10786), .A2(n11536), .B1(n10239), .B2(n11540), .ZN(
        n6754) );
  OAI22_X1 U4258 ( .A1(n10779), .A2(n11536), .B1(n10205), .B2(n11540), .ZN(
        n6753) );
  OAI22_X1 U4259 ( .A1(n10772), .A2(n11536), .B1(n10173), .B2(n11540), .ZN(
        n6752) );
  OAI22_X1 U4260 ( .A1(n10765), .A2(n11536), .B1(n10141), .B2(n11541), .ZN(
        n6751) );
  OAI22_X1 U4261 ( .A1(n10758), .A2(n11536), .B1(n10109), .B2(n11541), .ZN(
        n6750) );
  OAI22_X1 U4262 ( .A1(n10751), .A2(n11536), .B1(n10077), .B2(n11541), .ZN(
        n6749) );
  OAI22_X1 U4263 ( .A1(n10744), .A2(n11536), .B1(n10045), .B2(n11541), .ZN(
        n6748) );
  OAI22_X1 U4264 ( .A1(n10737), .A2(n11536), .B1(n10013), .B2(n11542), .ZN(
        n6747) );
  OAI22_X1 U4265 ( .A1(n10730), .A2(n11536), .B1(n9651), .B2(n11542), .ZN(
        n6746) );
  OAI22_X1 U4266 ( .A1(n10723), .A2(n11536), .B1(n9619), .B2(n11542), .ZN(
        n6745) );
  OAI22_X1 U4267 ( .A1(n10716), .A2(n11536), .B1(n9587), .B2(n11542), .ZN(
        n6744) );
  OAI22_X1 U4268 ( .A1(n10709), .A2(n11535), .B1(n9253), .B2(n11543), .ZN(
        n6743) );
  OAI22_X1 U4269 ( .A1(n10702), .A2(n11535), .B1(n9189), .B2(n11543), .ZN(
        n6742) );
  OAI22_X1 U4270 ( .A1(n10695), .A2(n11535), .B1(n9157), .B2(n11543), .ZN(
        n6741) );
  OAI22_X1 U4271 ( .A1(n10688), .A2(n11535), .B1(n6307), .B2(n11543), .ZN(
        n6740) );
  OAI22_X1 U4272 ( .A1(n10681), .A2(n11535), .B1(n5990), .B2(n11544), .ZN(
        n6739) );
  OAI22_X1 U4273 ( .A1(n10674), .A2(n11535), .B1(n5926), .B2(n11544), .ZN(
        n6738) );
  OAI22_X1 U4274 ( .A1(n10667), .A2(n11535), .B1(n5894), .B2(n11544), .ZN(
        n6737) );
  OAI22_X1 U4275 ( .A1(n10660), .A2(n11535), .B1(n5862), .B2(n11544), .ZN(
        n6736) );
  OAI22_X1 U4276 ( .A1(n10653), .A2(n11535), .B1(n5830), .B2(n11545), .ZN(
        n6735) );
  OAI22_X1 U4277 ( .A1(n10646), .A2(n11535), .B1(n5798), .B2(n11545), .ZN(
        n6734) );
  OAI22_X1 U4278 ( .A1(n10639), .A2(n11535), .B1(n5766), .B2(n11545), .ZN(
        n6733) );
  OAI22_X1 U4279 ( .A1(n10632), .A2(n11535), .B1(n5734), .B2(n11545), .ZN(
        n6732) );
  OAI22_X1 U4280 ( .A1(n10849), .A2(n11501), .B1(n1859), .B2(n11502), .ZN(
        n6667) );
  OAI22_X1 U4281 ( .A1(n10842), .A2(n11501), .B1(n1855), .B2(n11502), .ZN(
        n6666) );
  OAI22_X1 U4282 ( .A1(n10835), .A2(n11501), .B1(n1851), .B2(n11502), .ZN(
        n6665) );
  OAI22_X1 U4283 ( .A1(n10828), .A2(n11501), .B1(n1847), .B2(n11502), .ZN(
        n6664) );
  OAI22_X1 U4284 ( .A1(n10821), .A2(n11501), .B1(n1843), .B2(n11503), .ZN(
        n6663) );
  OAI22_X1 U4285 ( .A1(n10814), .A2(n11501), .B1(n1839), .B2(n11503), .ZN(
        n6662) );
  OAI22_X1 U4286 ( .A1(n10807), .A2(n11501), .B1(n1835), .B2(n11503), .ZN(
        n6661) );
  OAI22_X1 U4287 ( .A1(n10800), .A2(n11501), .B1(n1831), .B2(n11503), .ZN(
        n6660) );
  OAI22_X1 U4288 ( .A1(n10793), .A2(n11500), .B1(n1827), .B2(n11504), .ZN(
        n6659) );
  OAI22_X1 U4289 ( .A1(n10786), .A2(n11500), .B1(n1823), .B2(n11504), .ZN(
        n6658) );
  OAI22_X1 U4290 ( .A1(n10779), .A2(n11500), .B1(n1819), .B2(n11504), .ZN(
        n6657) );
  OAI22_X1 U4291 ( .A1(n10772), .A2(n11500), .B1(n1815), .B2(n11504), .ZN(
        n6656) );
  OAI22_X1 U4292 ( .A1(n10765), .A2(n11500), .B1(n1811), .B2(n11505), .ZN(
        n6655) );
  OAI22_X1 U4293 ( .A1(n10758), .A2(n11500), .B1(n1807), .B2(n11505), .ZN(
        n6654) );
  OAI22_X1 U4294 ( .A1(n10751), .A2(n11500), .B1(n1803), .B2(n11505), .ZN(
        n6653) );
  OAI22_X1 U4295 ( .A1(n10744), .A2(n11500), .B1(n1799), .B2(n11505), .ZN(
        n6652) );
  OAI22_X1 U4296 ( .A1(n10737), .A2(n11500), .B1(n1795), .B2(n11506), .ZN(
        n6651) );
  OAI22_X1 U4297 ( .A1(n10730), .A2(n11500), .B1(n1791), .B2(n11506), .ZN(
        n6650) );
  OAI22_X1 U4298 ( .A1(n10723), .A2(n11500), .B1(n1787), .B2(n11506), .ZN(
        n6649) );
  OAI22_X1 U4299 ( .A1(n10716), .A2(n11500), .B1(n1783), .B2(n11506), .ZN(
        n6648) );
  OAI22_X1 U4300 ( .A1(n10709), .A2(n11499), .B1(n1779), .B2(n11507), .ZN(
        n6647) );
  OAI22_X1 U4301 ( .A1(n10702), .A2(n11499), .B1(n1775), .B2(n11507), .ZN(
        n6646) );
  OAI22_X1 U4302 ( .A1(n10695), .A2(n11499), .B1(n1771), .B2(n11507), .ZN(
        n6645) );
  OAI22_X1 U4303 ( .A1(n10688), .A2(n11499), .B1(n1767), .B2(n11507), .ZN(
        n6644) );
  OAI22_X1 U4304 ( .A1(n10681), .A2(n11499), .B1(n1763), .B2(n11508), .ZN(
        n6643) );
  OAI22_X1 U4305 ( .A1(n10674), .A2(n11499), .B1(n1759), .B2(n11508), .ZN(
        n6642) );
  OAI22_X1 U4306 ( .A1(n10667), .A2(n11499), .B1(n1755), .B2(n11508), .ZN(
        n6641) );
  OAI22_X1 U4307 ( .A1(n10660), .A2(n11499), .B1(n1751), .B2(n11508), .ZN(
        n6640) );
  OAI22_X1 U4308 ( .A1(n10653), .A2(n11499), .B1(n1747), .B2(n11509), .ZN(
        n6639) );
  OAI22_X1 U4309 ( .A1(n10646), .A2(n11499), .B1(n1743), .B2(n11509), .ZN(
        n6638) );
  OAI22_X1 U4310 ( .A1(n10639), .A2(n11499), .B1(n1739), .B2(n11509), .ZN(
        n6637) );
  OAI22_X1 U4311 ( .A1(n10632), .A2(n11499), .B1(n1735), .B2(n11509), .ZN(
        n6636) );
  OAI22_X1 U4312 ( .A1(n10850), .A2(n11465), .B1(n513), .B2(n11466), .ZN(n6571) );
  OAI22_X1 U4313 ( .A1(n10843), .A2(n11465), .B1(n501), .B2(n11466), .ZN(n6570) );
  OAI22_X1 U4314 ( .A1(n10836), .A2(n11465), .B1(n489), .B2(n11466), .ZN(n6569) );
  OAI22_X1 U4315 ( .A1(n10829), .A2(n11465), .B1(n477), .B2(n11466), .ZN(n6568) );
  OAI22_X1 U4316 ( .A1(n10822), .A2(n11465), .B1(n465), .B2(n11467), .ZN(n6567) );
  OAI22_X1 U4317 ( .A1(n10815), .A2(n11465), .B1(n453), .B2(n11467), .ZN(n6566) );
  OAI22_X1 U4318 ( .A1(n10808), .A2(n11465), .B1(n441), .B2(n11467), .ZN(n6565) );
  OAI22_X1 U4319 ( .A1(n10801), .A2(n11465), .B1(n429), .B2(n11467), .ZN(n6564) );
  OAI22_X1 U4320 ( .A1(n10794), .A2(n11464), .B1(n417), .B2(n11468), .ZN(n6563) );
  OAI22_X1 U4321 ( .A1(n10787), .A2(n11464), .B1(n405), .B2(n11468), .ZN(n6562) );
  OAI22_X1 U4322 ( .A1(n10780), .A2(n11464), .B1(n393), .B2(n11468), .ZN(n6561) );
  OAI22_X1 U4323 ( .A1(n10773), .A2(n11464), .B1(n381), .B2(n11468), .ZN(n6560) );
  OAI22_X1 U4324 ( .A1(n10766), .A2(n11464), .B1(n369), .B2(n11469), .ZN(n6559) );
  OAI22_X1 U4325 ( .A1(n10759), .A2(n11464), .B1(n357), .B2(n11469), .ZN(n6558) );
  OAI22_X1 U4326 ( .A1(n10752), .A2(n11464), .B1(n345), .B2(n11469), .ZN(n6557) );
  OAI22_X1 U4327 ( .A1(n10745), .A2(n11464), .B1(n333), .B2(n11469), .ZN(n6556) );
  OAI22_X1 U4328 ( .A1(n10738), .A2(n11464), .B1(n321), .B2(n11470), .ZN(n6555) );
  OAI22_X1 U4329 ( .A1(n10731), .A2(n11464), .B1(n309), .B2(n11470), .ZN(n6554) );
  OAI22_X1 U4330 ( .A1(n10724), .A2(n11464), .B1(n297), .B2(n11470), .ZN(n6553) );
  OAI22_X1 U4331 ( .A1(n10717), .A2(n11464), .B1(n285), .B2(n11470), .ZN(n6552) );
  OAI22_X1 U4332 ( .A1(n10710), .A2(n11463), .B1(n273), .B2(n11471), .ZN(n6551) );
  OAI22_X1 U4333 ( .A1(n10703), .A2(n11463), .B1(n261), .B2(n11471), .ZN(n6550) );
  OAI22_X1 U4334 ( .A1(n10696), .A2(n11463), .B1(n249), .B2(n11471), .ZN(n6549) );
  OAI22_X1 U4335 ( .A1(n10689), .A2(n11463), .B1(n237), .B2(n11471), .ZN(n6548) );
  OAI22_X1 U4336 ( .A1(n10682), .A2(n11463), .B1(n225), .B2(n11472), .ZN(n6547) );
  OAI22_X1 U4337 ( .A1(n10675), .A2(n11463), .B1(n213), .B2(n11472), .ZN(n6546) );
  OAI22_X1 U4338 ( .A1(n10668), .A2(n11463), .B1(n201), .B2(n11472), .ZN(n6545) );
  OAI22_X1 U4339 ( .A1(n10661), .A2(n11463), .B1(n189), .B2(n11472), .ZN(n6544) );
  OAI22_X1 U4340 ( .A1(n10654), .A2(n11463), .B1(n177), .B2(n11473), .ZN(n6543) );
  OAI22_X1 U4341 ( .A1(n10647), .A2(n11463), .B1(n165), .B2(n11473), .ZN(n6542) );
  OAI22_X1 U4342 ( .A1(n10640), .A2(n11463), .B1(n153), .B2(n11473), .ZN(n6541) );
  OAI22_X1 U4343 ( .A1(n10633), .A2(n11463), .B1(n141), .B2(n11473), .ZN(n6540) );
  OAI22_X1 U4344 ( .A1(n10850), .A2(n11429), .B1(n514), .B2(n11430), .ZN(n6475) );
  OAI22_X1 U4345 ( .A1(n10843), .A2(n11429), .B1(n502), .B2(n11430), .ZN(n6474) );
  OAI22_X1 U4346 ( .A1(n10836), .A2(n11429), .B1(n490), .B2(n11430), .ZN(n6473) );
  OAI22_X1 U4347 ( .A1(n10829), .A2(n11429), .B1(n478), .B2(n11430), .ZN(n6472) );
  OAI22_X1 U4348 ( .A1(n10822), .A2(n11429), .B1(n466), .B2(n11431), .ZN(n6471) );
  OAI22_X1 U4349 ( .A1(n10815), .A2(n11429), .B1(n454), .B2(n11431), .ZN(n6470) );
  OAI22_X1 U4350 ( .A1(n10808), .A2(n11429), .B1(n442), .B2(n11431), .ZN(n6469) );
  OAI22_X1 U4351 ( .A1(n10801), .A2(n11429), .B1(n430), .B2(n11431), .ZN(n6468) );
  OAI22_X1 U4352 ( .A1(n10794), .A2(n11428), .B1(n418), .B2(n11432), .ZN(n6467) );
  OAI22_X1 U4353 ( .A1(n10787), .A2(n11428), .B1(n406), .B2(n11432), .ZN(n6466) );
  OAI22_X1 U4354 ( .A1(n10780), .A2(n11428), .B1(n394), .B2(n11432), .ZN(n6465) );
  OAI22_X1 U4355 ( .A1(n10773), .A2(n11428), .B1(n382), .B2(n11432), .ZN(n6464) );
  OAI22_X1 U4356 ( .A1(n10766), .A2(n11428), .B1(n370), .B2(n11433), .ZN(n6463) );
  OAI22_X1 U4357 ( .A1(n10759), .A2(n11428), .B1(n358), .B2(n11433), .ZN(n6462) );
  OAI22_X1 U4358 ( .A1(n10752), .A2(n11428), .B1(n346), .B2(n11433), .ZN(n6461) );
  OAI22_X1 U4360 ( .A1(n10745), .A2(n11428), .B1(n334), .B2(n11433), .ZN(n6460) );
  OAI22_X1 U4361 ( .A1(n10738), .A2(n11428), .B1(n322), .B2(n11434), .ZN(n6459) );
  OAI22_X1 U4362 ( .A1(n10731), .A2(n11428), .B1(n310), .B2(n11434), .ZN(n6458) );
  OAI22_X1 U4363 ( .A1(n10724), .A2(n11428), .B1(n298), .B2(n11434), .ZN(n6457) );
  OAI22_X1 U4364 ( .A1(n10717), .A2(n11428), .B1(n286), .B2(n11434), .ZN(n6456) );
  OAI22_X1 U4365 ( .A1(n10710), .A2(n11427), .B1(n274), .B2(n11435), .ZN(n6455) );
  OAI22_X1 U4366 ( .A1(n10703), .A2(n11427), .B1(n262), .B2(n11435), .ZN(n6454) );
  OAI22_X1 U4367 ( .A1(n10696), .A2(n11427), .B1(n250), .B2(n11435), .ZN(n6453) );
  OAI22_X1 U4368 ( .A1(n10689), .A2(n11427), .B1(n238), .B2(n11435), .ZN(n6452) );
  OAI22_X1 U4369 ( .A1(n10682), .A2(n11427), .B1(n226), .B2(n11436), .ZN(n6451) );
  OAI22_X1 U4370 ( .A1(n10675), .A2(n11427), .B1(n214), .B2(n11436), .ZN(n6450) );
  OAI22_X1 U4371 ( .A1(n10668), .A2(n11427), .B1(n202), .B2(n11436), .ZN(n6449) );
  OAI22_X1 U4372 ( .A1(n10661), .A2(n11427), .B1(n190), .B2(n11436), .ZN(n6448) );
  OAI22_X1 U4373 ( .A1(n10654), .A2(n11427), .B1(n178), .B2(n11437), .ZN(n6447) );
  OAI22_X1 U4374 ( .A1(n10647), .A2(n11427), .B1(n166), .B2(n11437), .ZN(n6446) );
  OAI22_X1 U4375 ( .A1(n10640), .A2(n11427), .B1(n154), .B2(n11437), .ZN(n6445) );
  OAI22_X1 U4376 ( .A1(n10633), .A2(n11427), .B1(n142), .B2(n11437), .ZN(n6444) );
  OAI22_X1 U4377 ( .A1(n10844), .A2(n12340), .B1(n10510), .B2(n12341), .ZN(
        n8907) );
  OAI22_X1 U4378 ( .A1(n10837), .A2(n12339), .B1(n10478), .B2(n12341), .ZN(
        n8906) );
  OAI22_X1 U4379 ( .A1(n10830), .A2(n12340), .B1(n10446), .B2(n12341), .ZN(
        n8905) );
  OAI22_X1 U4380 ( .A1(n10823), .A2(n12339), .B1(n10414), .B2(n12341), .ZN(
        n8904) );
  OAI22_X1 U4381 ( .A1(n10816), .A2(n12340), .B1(n10379), .B2(n12342), .ZN(
        n8903) );
  OAI22_X1 U4382 ( .A1(n10809), .A2(n12339), .B1(n10347), .B2(n12342), .ZN(
        n8902) );
  OAI22_X1 U4383 ( .A1(n10802), .A2(n12340), .B1(n10315), .B2(n12342), .ZN(
        n8901) );
  OAI22_X1 U4384 ( .A1(n10795), .A2(n12339), .B1(n10280), .B2(n12342), .ZN(
        n8900) );
  OAI22_X1 U4385 ( .A1(n10788), .A2(n12340), .B1(n10248), .B2(n12343), .ZN(
        n8899) );
  OAI22_X1 U4386 ( .A1(n10781), .A2(n12340), .B1(n10216), .B2(n12343), .ZN(
        n8898) );
  OAI22_X1 U4387 ( .A1(n10774), .A2(n12340), .B1(n10182), .B2(n12343), .ZN(
        n8897) );
  OAI22_X1 U4388 ( .A1(n10767), .A2(n12340), .B1(n10150), .B2(n12343), .ZN(
        n8896) );
  OAI22_X1 U4389 ( .A1(n10760), .A2(n12340), .B1(n10118), .B2(n12344), .ZN(
        n8895) );
  OAI22_X1 U4390 ( .A1(n10753), .A2(n12340), .B1(n10086), .B2(n12344), .ZN(
        n8894) );
  OAI22_X1 U4391 ( .A1(n10746), .A2(n12340), .B1(n10054), .B2(n12344), .ZN(
        n8893) );
  OAI22_X1 U4392 ( .A1(n10739), .A2(n12340), .B1(n10022), .B2(n12344), .ZN(
        n8892) );
  OAI22_X1 U4393 ( .A1(n10732), .A2(n12340), .B1(n9660), .B2(n12345), .ZN(
        n8891) );
  OAI22_X1 U4394 ( .A1(n10725), .A2(n12340), .B1(n9628), .B2(n12345), .ZN(
        n8890) );
  OAI22_X1 U4395 ( .A1(n10718), .A2(n12340), .B1(n9596), .B2(n12345), .ZN(
        n8889) );
  OAI22_X1 U4396 ( .A1(n10711), .A2(n12340), .B1(n9262), .B2(n12345), .ZN(
        n8888) );
  OAI22_X1 U4397 ( .A1(n10704), .A2(n12339), .B1(n9198), .B2(n12346), .ZN(
        n8887) );
  OAI22_X1 U4398 ( .A1(n10697), .A2(n12339), .B1(n9166), .B2(n12346), .ZN(
        n8886) );
  OAI22_X1 U4399 ( .A1(n10690), .A2(n12339), .B1(n9134), .B2(n12346), .ZN(
        n8885) );
  OAI22_X1 U4400 ( .A1(n10683), .A2(n12339), .B1(n5999), .B2(n12346), .ZN(
        n8884) );
  OAI22_X1 U4401 ( .A1(n10676), .A2(n12339), .B1(n5935), .B2(n12347), .ZN(
        n8883) );
  OAI22_X1 U4402 ( .A1(n10669), .A2(n12339), .B1(n5903), .B2(n12347), .ZN(
        n8882) );
  OAI22_X1 U4403 ( .A1(n10662), .A2(n12339), .B1(n5871), .B2(n12347), .ZN(
        n8881) );
  OAI22_X1 U4404 ( .A1(n10655), .A2(n12339), .B1(n5839), .B2(n12347), .ZN(
        n8880) );
  OAI22_X1 U4405 ( .A1(n10648), .A2(n12339), .B1(n5807), .B2(n12348), .ZN(
        n8879) );
  OAI22_X1 U4406 ( .A1(n10641), .A2(n12339), .B1(n5775), .B2(n12348), .ZN(
        n8878) );
  OAI22_X1 U4407 ( .A1(n10634), .A2(n12339), .B1(n5743), .B2(n12348), .ZN(
        n8877) );
  OAI22_X1 U4408 ( .A1(n10627), .A2(n12339), .B1(n5711), .B2(n12348), .ZN(
        n8876) );
  OAI22_X1 U4409 ( .A1(n10844), .A2(n12281), .B1(n992), .B2(n12282), .ZN(n8747) );
  OAI22_X1 U4410 ( .A1(n10837), .A2(n12281), .B1(n988), .B2(n12282), .ZN(n8746) );
  OAI22_X1 U4411 ( .A1(n10830), .A2(n12281), .B1(n984), .B2(n12282), .ZN(n8745) );
  OAI22_X1 U4412 ( .A1(n10823), .A2(n12281), .B1(n980), .B2(n12282), .ZN(n8744) );
  OAI22_X1 U4413 ( .A1(n10816), .A2(n12281), .B1(n976), .B2(n12283), .ZN(n8743) );
  OAI22_X1 U4414 ( .A1(n10809), .A2(n12281), .B1(n972), .B2(n12283), .ZN(n8742) );
  OAI22_X1 U4415 ( .A1(n10802), .A2(n12281), .B1(n968), .B2(n12283), .ZN(n8741) );
  OAI22_X1 U4416 ( .A1(n10795), .A2(n12281), .B1(n964), .B2(n12283), .ZN(n8740) );
  OAI22_X1 U4417 ( .A1(n10788), .A2(n12280), .B1(n960), .B2(n12284), .ZN(n8739) );
  OAI22_X1 U4418 ( .A1(n10781), .A2(n12280), .B1(n956), .B2(n12284), .ZN(n8738) );
  OAI22_X1 U4419 ( .A1(n10774), .A2(n12280), .B1(n952), .B2(n12284), .ZN(n8737) );
  OAI22_X1 U4420 ( .A1(n10767), .A2(n12280), .B1(n948), .B2(n12284), .ZN(n8736) );
  OAI22_X1 U4421 ( .A1(n10760), .A2(n12280), .B1(n944), .B2(n12285), .ZN(n8735) );
  OAI22_X1 U4422 ( .A1(n10753), .A2(n12280), .B1(n940), .B2(n12285), .ZN(n8734) );
  OAI22_X1 U4423 ( .A1(n10746), .A2(n12280), .B1(n936), .B2(n12285), .ZN(n8733) );
  OAI22_X1 U4424 ( .A1(n10739), .A2(n12280), .B1(n932), .B2(n12285), .ZN(n8732) );
  OAI22_X1 U4425 ( .A1(n10732), .A2(n12280), .B1(n928), .B2(n12286), .ZN(n8731) );
  OAI22_X1 U4426 ( .A1(n10725), .A2(n12280), .B1(n924), .B2(n12286), .ZN(n8730) );
  OAI22_X1 U4427 ( .A1(n10718), .A2(n12280), .B1(n920), .B2(n12286), .ZN(n8729) );
  OAI22_X1 U4428 ( .A1(n10711), .A2(n12280), .B1(n916), .B2(n12286), .ZN(n8728) );
  OAI22_X1 U4429 ( .A1(n10704), .A2(n12279), .B1(n912), .B2(n12287), .ZN(n8727) );
  OAI22_X1 U4430 ( .A1(n10697), .A2(n12279), .B1(n908), .B2(n12287), .ZN(n8726) );
  OAI22_X1 U4431 ( .A1(n10690), .A2(n12279), .B1(n904), .B2(n12287), .ZN(n8725) );
  OAI22_X1 U4432 ( .A1(n10683), .A2(n12279), .B1(n900), .B2(n12287), .ZN(n8724) );
  OAI22_X1 U4433 ( .A1(n10676), .A2(n12279), .B1(n896), .B2(n12288), .ZN(n8723) );
  OAI22_X1 U4434 ( .A1(n10669), .A2(n12279), .B1(n892), .B2(n12288), .ZN(n8722) );
  OAI22_X1 U4435 ( .A1(n10662), .A2(n12279), .B1(n888), .B2(n12288), .ZN(n8721) );
  OAI22_X1 U4436 ( .A1(n10655), .A2(n12279), .B1(n884), .B2(n12288), .ZN(n8720) );
  OAI22_X1 U4437 ( .A1(n10648), .A2(n12279), .B1(n880), .B2(n12289), .ZN(n8719) );
  OAI22_X1 U4438 ( .A1(n10641), .A2(n12279), .B1(n876), .B2(n12289), .ZN(n8718) );
  OAI22_X1 U4439 ( .A1(n10634), .A2(n12279), .B1(n872), .B2(n12289), .ZN(n8717) );
  OAI22_X1 U4440 ( .A1(n10627), .A2(n12279), .B1(n868), .B2(n12289), .ZN(n8716) );
  OAI22_X1 U4441 ( .A1(n10845), .A2(n12125), .B1(n10515), .B2(n12126), .ZN(
        n8331) );
  OAI22_X1 U4442 ( .A1(n10838), .A2(n12125), .B1(n10483), .B2(n12126), .ZN(
        n8330) );
  OAI22_X1 U4443 ( .A1(n10831), .A2(n12125), .B1(n10451), .B2(n12126), .ZN(
        n8329) );
  OAI22_X1 U4444 ( .A1(n10824), .A2(n12125), .B1(n10419), .B2(n12126), .ZN(
        n8328) );
  OAI22_X1 U4445 ( .A1(n10817), .A2(n12125), .B1(n10384), .B2(n12127), .ZN(
        n8327) );
  OAI22_X1 U4446 ( .A1(n10810), .A2(n12125), .B1(n10352), .B2(n12127), .ZN(
        n8326) );
  OAI22_X1 U4447 ( .A1(n10803), .A2(n12125), .B1(n10320), .B2(n12127), .ZN(
        n8325) );
  OAI22_X1 U4448 ( .A1(n10796), .A2(n12125), .B1(n10285), .B2(n12127), .ZN(
        n8324) );
  OAI22_X1 U4449 ( .A1(n10789), .A2(n12124), .B1(n10253), .B2(n12128), .ZN(
        n8323) );
  OAI22_X1 U4450 ( .A1(n10782), .A2(n12124), .B1(n10221), .B2(n12128), .ZN(
        n8322) );
  OAI22_X1 U4451 ( .A1(n10775), .A2(n12124), .B1(n10187), .B2(n12128), .ZN(
        n8321) );
  OAI22_X1 U4452 ( .A1(n10768), .A2(n12124), .B1(n10155), .B2(n12128), .ZN(
        n8320) );
  OAI22_X1 U4453 ( .A1(n10761), .A2(n12124), .B1(n10123), .B2(n12129), .ZN(
        n8319) );
  OAI22_X1 U4454 ( .A1(n10754), .A2(n12124), .B1(n10091), .B2(n12129), .ZN(
        n8318) );
  OAI22_X1 U4455 ( .A1(n10747), .A2(n12124), .B1(n10059), .B2(n12129), .ZN(
        n8317) );
  OAI22_X1 U4456 ( .A1(n10740), .A2(n12124), .B1(n10027), .B2(n12129), .ZN(
        n8316) );
  OAI22_X1 U4457 ( .A1(n10733), .A2(n12124), .B1(n9697), .B2(n12130), .ZN(
        n8315) );
  OAI22_X1 U4458 ( .A1(n10726), .A2(n12124), .B1(n9633), .B2(n12130), .ZN(
        n8314) );
  OAI22_X1 U4459 ( .A1(n10719), .A2(n12124), .B1(n9601), .B2(n12130), .ZN(
        n8313) );
  OAI22_X1 U4460 ( .A1(n10712), .A2(n12124), .B1(n9569), .B2(n12130), .ZN(
        n8312) );
  OAI22_X1 U4461 ( .A1(n10705), .A2(n12123), .B1(n9203), .B2(n12131), .ZN(
        n8311) );
  OAI22_X1 U4462 ( .A1(n10698), .A2(n12123), .B1(n9171), .B2(n12131), .ZN(
        n8310) );
  OAI22_X1 U4463 ( .A1(n10691), .A2(n12123), .B1(n9139), .B2(n12131), .ZN(
        n8309) );
  OAI22_X1 U4464 ( .A1(n10684), .A2(n12123), .B1(n6004), .B2(n12131), .ZN(
        n8308) );
  OAI22_X1 U4465 ( .A1(n10677), .A2(n12123), .B1(n5940), .B2(n12132), .ZN(
        n8307) );
  OAI22_X1 U4466 ( .A1(n10670), .A2(n12123), .B1(n5908), .B2(n12132), .ZN(
        n8306) );
  OAI22_X1 U4467 ( .A1(n10663), .A2(n12123), .B1(n5876), .B2(n12132), .ZN(
        n8305) );
  OAI22_X1 U4468 ( .A1(n10656), .A2(n12123), .B1(n5844), .B2(n12132), .ZN(
        n8304) );
  OAI22_X1 U4469 ( .A1(n10649), .A2(n12123), .B1(n5812), .B2(n12133), .ZN(
        n8303) );
  OAI22_X1 U4470 ( .A1(n10642), .A2(n12123), .B1(n5780), .B2(n12133), .ZN(
        n8302) );
  OAI22_X1 U4471 ( .A1(n10635), .A2(n12123), .B1(n5748), .B2(n12133), .ZN(
        n8301) );
  OAI22_X1 U4472 ( .A1(n10628), .A2(n12123), .B1(n5716), .B2(n12133), .ZN(
        n8300) );
  OAI22_X1 U4473 ( .A1(n10846), .A2(n12077), .B1(n10518), .B2(n12078), .ZN(
        n8203) );
  OAI22_X1 U4474 ( .A1(n10839), .A2(n12077), .B1(n10486), .B2(n12078), .ZN(
        n8202) );
  OAI22_X1 U4475 ( .A1(n10832), .A2(n12077), .B1(n10454), .B2(n12078), .ZN(
        n8201) );
  OAI22_X1 U4476 ( .A1(n10825), .A2(n12077), .B1(n10422), .B2(n12078), .ZN(
        n8200) );
  OAI22_X1 U4477 ( .A1(n10818), .A2(n12077), .B1(n10387), .B2(n12079), .ZN(
        n8199) );
  OAI22_X1 U4478 ( .A1(n10811), .A2(n12077), .B1(n10355), .B2(n12079), .ZN(
        n8198) );
  OAI22_X1 U4479 ( .A1(n10804), .A2(n12077), .B1(n10323), .B2(n12079), .ZN(
        n8197) );
  OAI22_X1 U4480 ( .A1(n10797), .A2(n12077), .B1(n10288), .B2(n12079), .ZN(
        n8196) );
  OAI22_X1 U4481 ( .A1(n10790), .A2(n12076), .B1(n10256), .B2(n12080), .ZN(
        n8195) );
  OAI22_X1 U4482 ( .A1(n10783), .A2(n12076), .B1(n10224), .B2(n12080), .ZN(
        n8194) );
  OAI22_X1 U4483 ( .A1(n10776), .A2(n12076), .B1(n10190), .B2(n12080), .ZN(
        n8193) );
  OAI22_X1 U4484 ( .A1(n10769), .A2(n12076), .B1(n10158), .B2(n12080), .ZN(
        n8192) );
  OAI22_X1 U4485 ( .A1(n10762), .A2(n12076), .B1(n10126), .B2(n12081), .ZN(
        n8191) );
  OAI22_X1 U4486 ( .A1(n10755), .A2(n12076), .B1(n10094), .B2(n12081), .ZN(
        n8190) );
  OAI22_X1 U4487 ( .A1(n10748), .A2(n12076), .B1(n10062), .B2(n12081), .ZN(
        n8189) );
  OAI22_X1 U4488 ( .A1(n10741), .A2(n12076), .B1(n10030), .B2(n12081), .ZN(
        n8188) );
  OAI22_X1 U4489 ( .A1(n10734), .A2(n12076), .B1(n9700), .B2(n12082), .ZN(
        n8187) );
  OAI22_X1 U4490 ( .A1(n10727), .A2(n12076), .B1(n9636), .B2(n12082), .ZN(
        n8186) );
  OAI22_X1 U4491 ( .A1(n10720), .A2(n12076), .B1(n9604), .B2(n12082), .ZN(
        n8185) );
  OAI22_X1 U4492 ( .A1(n10713), .A2(n12076), .B1(n9572), .B2(n12082), .ZN(
        n8184) );
  OAI22_X1 U4493 ( .A1(n10706), .A2(n12075), .B1(n9206), .B2(n12083), .ZN(
        n8183) );
  OAI22_X1 U4494 ( .A1(n10699), .A2(n12075), .B1(n9174), .B2(n12083), .ZN(
        n8182) );
  OAI22_X1 U4495 ( .A1(n10692), .A2(n12075), .B1(n9142), .B2(n12083), .ZN(
        n8181) );
  OAI22_X1 U4496 ( .A1(n10685), .A2(n12075), .B1(n6007), .B2(n12083), .ZN(
        n8180) );
  OAI22_X1 U4497 ( .A1(n10678), .A2(n12075), .B1(n5943), .B2(n12084), .ZN(
        n8179) );
  OAI22_X1 U4498 ( .A1(n10671), .A2(n12075), .B1(n5911), .B2(n12084), .ZN(
        n8178) );
  OAI22_X1 U4499 ( .A1(n10664), .A2(n12075), .B1(n5879), .B2(n12084), .ZN(
        n8177) );
  OAI22_X1 U4500 ( .A1(n10657), .A2(n12075), .B1(n5847), .B2(n12084), .ZN(
        n8176) );
  OAI22_X1 U4501 ( .A1(n10650), .A2(n12075), .B1(n5815), .B2(n12085), .ZN(
        n8175) );
  OAI22_X1 U4502 ( .A1(n10643), .A2(n12075), .B1(n5783), .B2(n12085), .ZN(
        n8174) );
  OAI22_X1 U4503 ( .A1(n10636), .A2(n12075), .B1(n5751), .B2(n12085), .ZN(
        n8173) );
  OAI22_X1 U4504 ( .A1(n10629), .A2(n12075), .B1(n5719), .B2(n12085), .ZN(
        n8172) );
  OAI22_X1 U4505 ( .A1(n10847), .A2(n11861), .B1(n10523), .B2(n11862), .ZN(
        n7627) );
  OAI22_X1 U4506 ( .A1(n10840), .A2(n11861), .B1(n10491), .B2(n11862), .ZN(
        n7626) );
  OAI22_X1 U4507 ( .A1(n10833), .A2(n11861), .B1(n10459), .B2(n11862), .ZN(
        n7625) );
  OAI22_X1 U4508 ( .A1(n10826), .A2(n11861), .B1(n10427), .B2(n11862), .ZN(
        n7624) );
  OAI22_X1 U4509 ( .A1(n10819), .A2(n11861), .B1(n10392), .B2(n11863), .ZN(
        n7623) );
  OAI22_X1 U4510 ( .A1(n10812), .A2(n11861), .B1(n10360), .B2(n11863), .ZN(
        n7622) );
  OAI22_X1 U4511 ( .A1(n10805), .A2(n11861), .B1(n10328), .B2(n11863), .ZN(
        n7621) );
  OAI22_X1 U4512 ( .A1(n10798), .A2(n11861), .B1(n10293), .B2(n11863), .ZN(
        n7620) );
  OAI22_X1 U4513 ( .A1(n10791), .A2(n11860), .B1(n10261), .B2(n11864), .ZN(
        n7619) );
  OAI22_X1 U4514 ( .A1(n10784), .A2(n11860), .B1(n10229), .B2(n11864), .ZN(
        n7618) );
  OAI22_X1 U4515 ( .A1(n10777), .A2(n11860), .B1(n10195), .B2(n11864), .ZN(
        n7617) );
  OAI22_X1 U4516 ( .A1(n10770), .A2(n11860), .B1(n10163), .B2(n11864), .ZN(
        n7616) );
  OAI22_X1 U4517 ( .A1(n10763), .A2(n11860), .B1(n10131), .B2(n11865), .ZN(
        n7615) );
  OAI22_X1 U4518 ( .A1(n10756), .A2(n11860), .B1(n10099), .B2(n11865), .ZN(
        n7614) );
  OAI22_X1 U4519 ( .A1(n10749), .A2(n11860), .B1(n10067), .B2(n11865), .ZN(
        n7613) );
  OAI22_X1 U4520 ( .A1(n10742), .A2(n11860), .B1(n10035), .B2(n11865), .ZN(
        n7612) );
  OAI22_X1 U4521 ( .A1(n10735), .A2(n11860), .B1(n10003), .B2(n11866), .ZN(
        n7611) );
  OAI22_X1 U4522 ( .A1(n10728), .A2(n11860), .B1(n9641), .B2(n11866), .ZN(
        n7610) );
  OAI22_X1 U4523 ( .A1(n10721), .A2(n11860), .B1(n9609), .B2(n11866), .ZN(
        n7609) );
  OAI22_X1 U4524 ( .A1(n10714), .A2(n11860), .B1(n9577), .B2(n11866), .ZN(
        n7608) );
  OAI22_X1 U4525 ( .A1(n10707), .A2(n11859), .B1(n9211), .B2(n11867), .ZN(
        n7607) );
  OAI22_X1 U4526 ( .A1(n10700), .A2(n11859), .B1(n9179), .B2(n11867), .ZN(
        n7606) );
  OAI22_X1 U4527 ( .A1(n10693), .A2(n11859), .B1(n9147), .B2(n11867), .ZN(
        n7605) );
  OAI22_X1 U4528 ( .A1(n10686), .A2(n11859), .B1(n6012), .B2(n11867), .ZN(
        n7604) );
  OAI22_X1 U4529 ( .A1(n10679), .A2(n11859), .B1(n5948), .B2(n11868), .ZN(
        n7603) );
  OAI22_X1 U4530 ( .A1(n10672), .A2(n11859), .B1(n5916), .B2(n11868), .ZN(
        n7602) );
  OAI22_X1 U4531 ( .A1(n10665), .A2(n11859), .B1(n5884), .B2(n11868), .ZN(
        n7601) );
  OAI22_X1 U4532 ( .A1(n10658), .A2(n11859), .B1(n5852), .B2(n11868), .ZN(
        n7600) );
  OAI22_X1 U4533 ( .A1(n10651), .A2(n11859), .B1(n5820), .B2(n11869), .ZN(
        n7599) );
  OAI22_X1 U4534 ( .A1(n10644), .A2(n11859), .B1(n5788), .B2(n11869), .ZN(
        n7598) );
  OAI22_X1 U4535 ( .A1(n10637), .A2(n11859), .B1(n5756), .B2(n11869), .ZN(
        n7597) );
  OAI22_X1 U4536 ( .A1(n10630), .A2(n11859), .B1(n5724), .B2(n11869), .ZN(
        n7596) );
  OAI22_X1 U4537 ( .A1(n10847), .A2(n11813), .B1(n10526), .B2(n11814), .ZN(
        n7499) );
  OAI22_X1 U4538 ( .A1(n10840), .A2(n11813), .B1(n10494), .B2(n11814), .ZN(
        n7498) );
  OAI22_X1 U4539 ( .A1(n10833), .A2(n11813), .B1(n10462), .B2(n11814), .ZN(
        n7497) );
  OAI22_X1 U4540 ( .A1(n10826), .A2(n11813), .B1(n10430), .B2(n11814), .ZN(
        n7496) );
  OAI22_X1 U4541 ( .A1(n10819), .A2(n11813), .B1(n10395), .B2(n11815), .ZN(
        n7495) );
  OAI22_X1 U4542 ( .A1(n10812), .A2(n11813), .B1(n10363), .B2(n11815), .ZN(
        n7494) );
  OAI22_X1 U4543 ( .A1(n10805), .A2(n11813), .B1(n10331), .B2(n11815), .ZN(
        n7493) );
  OAI22_X1 U4544 ( .A1(n10798), .A2(n11813), .B1(n10296), .B2(n11815), .ZN(
        n7492) );
  OAI22_X1 U4545 ( .A1(n10791), .A2(n11812), .B1(n10264), .B2(n11816), .ZN(
        n7491) );
  OAI22_X1 U4546 ( .A1(n10784), .A2(n11812), .B1(n10232), .B2(n11816), .ZN(
        n7490) );
  OAI22_X1 U4547 ( .A1(n10777), .A2(n11812), .B1(n10198), .B2(n11816), .ZN(
        n7489) );
  OAI22_X1 U4548 ( .A1(n10770), .A2(n11812), .B1(n10166), .B2(n11816), .ZN(
        n7488) );
  OAI22_X1 U4549 ( .A1(n10763), .A2(n11812), .B1(n10134), .B2(n11817), .ZN(
        n7487) );
  OAI22_X1 U4550 ( .A1(n10756), .A2(n11812), .B1(n10102), .B2(n11817), .ZN(
        n7486) );
  OAI22_X1 U4551 ( .A1(n10749), .A2(n11812), .B1(n10070), .B2(n11817), .ZN(
        n7485) );
  OAI22_X1 U4552 ( .A1(n10742), .A2(n11812), .B1(n10038), .B2(n11817), .ZN(
        n7484) );
  OAI22_X1 U4553 ( .A1(n10735), .A2(n11812), .B1(n10006), .B2(n11818), .ZN(
        n7483) );
  OAI22_X1 U4554 ( .A1(n10728), .A2(n11812), .B1(n9644), .B2(n11818), .ZN(
        n7482) );
  OAI22_X1 U4555 ( .A1(n10721), .A2(n11812), .B1(n9612), .B2(n11818), .ZN(
        n7481) );
  OAI22_X1 U4556 ( .A1(n10714), .A2(n11812), .B1(n9580), .B2(n11818), .ZN(
        n7480) );
  OAI22_X1 U4557 ( .A1(n10707), .A2(n11811), .B1(n9214), .B2(n11819), .ZN(
        n7479) );
  OAI22_X1 U4558 ( .A1(n10700), .A2(n11811), .B1(n9182), .B2(n11819), .ZN(
        n7478) );
  OAI22_X1 U4559 ( .A1(n10693), .A2(n11811), .B1(n9150), .B2(n11819), .ZN(
        n7477) );
  OAI22_X1 U4560 ( .A1(n10686), .A2(n11811), .B1(n6236), .B2(n11819), .ZN(
        n7476) );
  OAI22_X1 U4561 ( .A1(n10679), .A2(n11811), .B1(n5983), .B2(n11820), .ZN(
        n7475) );
  OAI22_X1 U4562 ( .A1(n10672), .A2(n11811), .B1(n5919), .B2(n11820), .ZN(
        n7474) );
  OAI22_X1 U4563 ( .A1(n10665), .A2(n11811), .B1(n5887), .B2(n11820), .ZN(
        n7473) );
  OAI22_X1 U4564 ( .A1(n10658), .A2(n11811), .B1(n5855), .B2(n11820), .ZN(
        n7472) );
  OAI22_X1 U4565 ( .A1(n10651), .A2(n11811), .B1(n5823), .B2(n11821), .ZN(
        n7471) );
  OAI22_X1 U4566 ( .A1(n10644), .A2(n11811), .B1(n5791), .B2(n11821), .ZN(
        n7470) );
  OAI22_X1 U4567 ( .A1(n10637), .A2(n11811), .B1(n5759), .B2(n11821), .ZN(
        n7469) );
  OAI22_X1 U4568 ( .A1(n10630), .A2(n11811), .B1(n5727), .B2(n11821), .ZN(
        n7468) );
  OAI22_X1 U4569 ( .A1(n10849), .A2(n11549), .B1(n10534), .B2(n11550), .ZN(
        n6795) );
  OAI22_X1 U4570 ( .A1(n10842), .A2(n11549), .B1(n10502), .B2(n11550), .ZN(
        n6794) );
  OAI22_X1 U4571 ( .A1(n10835), .A2(n11549), .B1(n10470), .B2(n11550), .ZN(
        n6793) );
  OAI22_X1 U4572 ( .A1(n10828), .A2(n11549), .B1(n10438), .B2(n11550), .ZN(
        n6792) );
  OAI22_X1 U4573 ( .A1(n10821), .A2(n11549), .B1(n10406), .B2(n11551), .ZN(
        n6791) );
  OAI22_X1 U4574 ( .A1(n10814), .A2(n11549), .B1(n10371), .B2(n11551), .ZN(
        n6790) );
  OAI22_X1 U4575 ( .A1(n10807), .A2(n11549), .B1(n10339), .B2(n11551), .ZN(
        n6789) );
  OAI22_X1 U4576 ( .A1(n10800), .A2(n11549), .B1(n10307), .B2(n11551), .ZN(
        n6788) );
  OAI22_X1 U4577 ( .A1(n10793), .A2(n11548), .B1(n10272), .B2(n11552), .ZN(
        n6787) );
  OAI22_X1 U4578 ( .A1(n10786), .A2(n11548), .B1(n10240), .B2(n11552), .ZN(
        n6786) );
  OAI22_X1 U4579 ( .A1(n10779), .A2(n11548), .B1(n10208), .B2(n11552), .ZN(
        n6785) );
  OAI22_X1 U4580 ( .A1(n10772), .A2(n11548), .B1(n10174), .B2(n11552), .ZN(
        n6784) );
  OAI22_X1 U4581 ( .A1(n10765), .A2(n11548), .B1(n10142), .B2(n11553), .ZN(
        n6783) );
  OAI22_X1 U4582 ( .A1(n10758), .A2(n11548), .B1(n10110), .B2(n11553), .ZN(
        n6782) );
  OAI22_X1 U4583 ( .A1(n10751), .A2(n11548), .B1(n10078), .B2(n11553), .ZN(
        n6781) );
  OAI22_X1 U4584 ( .A1(n10744), .A2(n11548), .B1(n10046), .B2(n11553), .ZN(
        n6780) );
  OAI22_X1 U4585 ( .A1(n10737), .A2(n11548), .B1(n10014), .B2(n11554), .ZN(
        n6779) );
  OAI22_X1 U4586 ( .A1(n10730), .A2(n11548), .B1(n9652), .B2(n11554), .ZN(
        n6778) );
  OAI22_X1 U4587 ( .A1(n10723), .A2(n11548), .B1(n9620), .B2(n11554), .ZN(
        n6777) );
  OAI22_X1 U4588 ( .A1(n10716), .A2(n11548), .B1(n9588), .B2(n11554), .ZN(
        n6776) );
  OAI22_X1 U4589 ( .A1(n10709), .A2(n11547), .B1(n9254), .B2(n11555), .ZN(
        n6775) );
  OAI22_X1 U4590 ( .A1(n10702), .A2(n11547), .B1(n9190), .B2(n11555), .ZN(
        n6774) );
  OAI22_X1 U4591 ( .A1(n10695), .A2(n11547), .B1(n9158), .B2(n11555), .ZN(
        n6773) );
  OAI22_X1 U4592 ( .A1(n10688), .A2(n11547), .B1(n6308), .B2(n11555), .ZN(
        n6772) );
  OAI22_X1 U4593 ( .A1(n10681), .A2(n11547), .B1(n5991), .B2(n11556), .ZN(
        n6771) );
  OAI22_X1 U4594 ( .A1(n10674), .A2(n11547), .B1(n5927), .B2(n11556), .ZN(
        n6770) );
  OAI22_X1 U4595 ( .A1(n10667), .A2(n11547), .B1(n5895), .B2(n11556), .ZN(
        n6769) );
  OAI22_X1 U4596 ( .A1(n10660), .A2(n11547), .B1(n5863), .B2(n11556), .ZN(
        n6768) );
  OAI22_X1 U4597 ( .A1(n10653), .A2(n11547), .B1(n5831), .B2(n11557), .ZN(
        n6767) );
  OAI22_X1 U4598 ( .A1(n10646), .A2(n11547), .B1(n5799), .B2(n11557), .ZN(
        n6766) );
  OAI22_X1 U4599 ( .A1(n10639), .A2(n11547), .B1(n5767), .B2(n11557), .ZN(
        n6765) );
  OAI22_X1 U4600 ( .A1(n10632), .A2(n11547), .B1(n5735), .B2(n11557), .ZN(
        n6764) );
  OAI22_X1 U4601 ( .A1(n10850), .A2(n11489), .B1(n995), .B2(n11490), .ZN(n6635) );
  OAI22_X1 U4602 ( .A1(n10843), .A2(n11489), .B1(n991), .B2(n11490), .ZN(n6634) );
  OAI22_X1 U4603 ( .A1(n10836), .A2(n11489), .B1(n987), .B2(n11490), .ZN(n6633) );
  OAI22_X1 U4604 ( .A1(n10829), .A2(n11489), .B1(n983), .B2(n11490), .ZN(n6632) );
  OAI22_X1 U4605 ( .A1(n10822), .A2(n11489), .B1(n979), .B2(n11491), .ZN(n6631) );
  OAI22_X1 U4606 ( .A1(n10815), .A2(n11489), .B1(n975), .B2(n11491), .ZN(n6630) );
  OAI22_X1 U4607 ( .A1(n10808), .A2(n11489), .B1(n971), .B2(n11491), .ZN(n6629) );
  OAI22_X1 U4608 ( .A1(n10801), .A2(n11489), .B1(n967), .B2(n11491), .ZN(n6628) );
  OAI22_X1 U4609 ( .A1(n10794), .A2(n11488), .B1(n963), .B2(n11492), .ZN(n6627) );
  OAI22_X1 U4610 ( .A1(n10787), .A2(n11488), .B1(n959), .B2(n11492), .ZN(n6626) );
  OAI22_X1 U4611 ( .A1(n10780), .A2(n11488), .B1(n955), .B2(n11492), .ZN(n6625) );
  OAI22_X1 U4612 ( .A1(n10773), .A2(n11488), .B1(n951), .B2(n11492), .ZN(n6624) );
  OAI22_X1 U4613 ( .A1(n10766), .A2(n11488), .B1(n947), .B2(n11493), .ZN(n6623) );
  OAI22_X1 U4614 ( .A1(n10759), .A2(n11488), .B1(n943), .B2(n11493), .ZN(n6622) );
  OAI22_X1 U4615 ( .A1(n10752), .A2(n11488), .B1(n939), .B2(n11493), .ZN(n6621) );
  OAI22_X1 U4616 ( .A1(n10745), .A2(n11488), .B1(n935), .B2(n11493), .ZN(n6620) );
  OAI22_X1 U4617 ( .A1(n10738), .A2(n11488), .B1(n931), .B2(n11494), .ZN(n6619) );
  OAI22_X1 U4618 ( .A1(n10731), .A2(n11488), .B1(n927), .B2(n11494), .ZN(n6618) );
  OAI22_X1 U4619 ( .A1(n10724), .A2(n11488), .B1(n923), .B2(n11494), .ZN(n6617) );
  OAI22_X1 U4620 ( .A1(n10717), .A2(n11488), .B1(n919), .B2(n11494), .ZN(n6616) );
  OAI22_X1 U4621 ( .A1(n10710), .A2(n11487), .B1(n915), .B2(n11495), .ZN(n6615) );
  OAI22_X1 U4622 ( .A1(n10703), .A2(n11487), .B1(n911), .B2(n11495), .ZN(n6614) );
  OAI22_X1 U4623 ( .A1(n10696), .A2(n11487), .B1(n907), .B2(n11495), .ZN(n6613) );
  OAI22_X1 U4624 ( .A1(n10689), .A2(n11487), .B1(n903), .B2(n11495), .ZN(n6612) );
  OAI22_X1 U4625 ( .A1(n10682), .A2(n11487), .B1(n899), .B2(n11496), .ZN(n6611) );
  OAI22_X1 U4626 ( .A1(n10675), .A2(n11487), .B1(n895), .B2(n11496), .ZN(n6610) );
  OAI22_X1 U4627 ( .A1(n10668), .A2(n11487), .B1(n891), .B2(n11496), .ZN(n6609) );
  OAI22_X1 U4628 ( .A1(n10661), .A2(n11487), .B1(n887), .B2(n11496), .ZN(n6608) );
  OAI22_X1 U4629 ( .A1(n10654), .A2(n11487), .B1(n883), .B2(n11497), .ZN(n6607) );
  OAI22_X1 U4630 ( .A1(n10647), .A2(n11487), .B1(n879), .B2(n11497), .ZN(n6606) );
  OAI22_X1 U4631 ( .A1(n10640), .A2(n11487), .B1(n875), .B2(n11497), .ZN(n6605) );
  OAI22_X1 U4632 ( .A1(n10633), .A2(n11487), .B1(n871), .B2(n11497), .ZN(n6604) );
  OAI22_X1 U4633 ( .A1(n10850), .A2(n11453), .B1(n2337), .B2(n11454), .ZN(
        n6539) );
  OAI22_X1 U4634 ( .A1(n10843), .A2(n11453), .B1(n2325), .B2(n11454), .ZN(
        n6538) );
  OAI22_X1 U4635 ( .A1(n10836), .A2(n11453), .B1(n2313), .B2(n11454), .ZN(
        n6537) );
  OAI22_X1 U4636 ( .A1(n10829), .A2(n11453), .B1(n2301), .B2(n11454), .ZN(
        n6536) );
  OAI22_X1 U4637 ( .A1(n10822), .A2(n11453), .B1(n2289), .B2(n11455), .ZN(
        n6535) );
  OAI22_X1 U4638 ( .A1(n10815), .A2(n11453), .B1(n2277), .B2(n11455), .ZN(
        n6534) );
  OAI22_X1 U4639 ( .A1(n10808), .A2(n11453), .B1(n2265), .B2(n11455), .ZN(
        n6533) );
  OAI22_X1 U4640 ( .A1(n10801), .A2(n11453), .B1(n2253), .B2(n11455), .ZN(
        n6532) );
  OAI22_X1 U4641 ( .A1(n10794), .A2(n11452), .B1(n2241), .B2(n11456), .ZN(
        n6531) );
  OAI22_X1 U4642 ( .A1(n10787), .A2(n11452), .B1(n2229), .B2(n11456), .ZN(
        n6530) );
  OAI22_X1 U4643 ( .A1(n10780), .A2(n11452), .B1(n2217), .B2(n11456), .ZN(
        n6529) );
  OAI22_X1 U4644 ( .A1(n10773), .A2(n11452), .B1(n2173), .B2(n11456), .ZN(
        n6528) );
  OAI22_X1 U4645 ( .A1(n10766), .A2(n11452), .B1(n2161), .B2(n11457), .ZN(
        n6527) );
  OAI22_X1 U4646 ( .A1(n10759), .A2(n11452), .B1(n2149), .B2(n11457), .ZN(
        n6526) );
  OAI22_X1 U4647 ( .A1(n10752), .A2(n11452), .B1(n2105), .B2(n11457), .ZN(
        n6525) );
  OAI22_X1 U4648 ( .A1(n10745), .A2(n11452), .B1(n2093), .B2(n11457), .ZN(
        n6524) );
  OAI22_X1 U4649 ( .A1(n10738), .A2(n11452), .B1(n2049), .B2(n11458), .ZN(
        n6523) );
  OAI22_X1 U4650 ( .A1(n10731), .A2(n11452), .B1(n2037), .B2(n11458), .ZN(
        n6522) );
  OAI22_X1 U4651 ( .A1(n10724), .A2(n11452), .B1(n2025), .B2(n11458), .ZN(
        n6521) );
  OAI22_X1 U4652 ( .A1(n10717), .A2(n11452), .B1(n2013), .B2(n11458), .ZN(
        n6520) );
  OAI22_X1 U4653 ( .A1(n10710), .A2(n11451), .B1(n2001), .B2(n11459), .ZN(
        n6519) );
  OAI22_X1 U4654 ( .A1(n10703), .A2(n11451), .B1(n1989), .B2(n11459), .ZN(
        n6518) );
  OAI22_X1 U4655 ( .A1(n10696), .A2(n11451), .B1(n1977), .B2(n11459), .ZN(
        n6517) );
  OAI22_X1 U4656 ( .A1(n10689), .A2(n11451), .B1(n1965), .B2(n11459), .ZN(
        n6516) );
  OAI22_X1 U4657 ( .A1(n10682), .A2(n11451), .B1(n1953), .B2(n11460), .ZN(
        n6515) );
  OAI22_X1 U4658 ( .A1(n10675), .A2(n11451), .B1(n1941), .B2(n11460), .ZN(
        n6514) );
  OAI22_X1 U4659 ( .A1(n10668), .A2(n11451), .B1(n1929), .B2(n11460), .ZN(
        n6513) );
  OAI22_X1 U4660 ( .A1(n10661), .A2(n11451), .B1(n1917), .B2(n11460), .ZN(
        n6512) );
  OAI22_X1 U4661 ( .A1(n10654), .A2(n11451), .B1(n1905), .B2(n11461), .ZN(
        n6511) );
  OAI22_X1 U4662 ( .A1(n10647), .A2(n11451), .B1(n1893), .B2(n11461), .ZN(
        n6510) );
  OAI22_X1 U4663 ( .A1(n10640), .A2(n11451), .B1(n1881), .B2(n11461), .ZN(
        n6509) );
  OAI22_X1 U4664 ( .A1(n10633), .A2(n11451), .B1(n1869), .B2(n11461), .ZN(
        n6508) );
  OAI22_X1 U4665 ( .A1(n10850), .A2(n11417), .B1(n2338), .B2(n11418), .ZN(
        n6443) );
  OAI22_X1 U4666 ( .A1(n10843), .A2(n11417), .B1(n2326), .B2(n11418), .ZN(
        n6442) );
  OAI22_X1 U4667 ( .A1(n10836), .A2(n11417), .B1(n2314), .B2(n11418), .ZN(
        n6441) );
  OAI22_X1 U4668 ( .A1(n10829), .A2(n11417), .B1(n2302), .B2(n11418), .ZN(
        n6440) );
  OAI22_X1 U4669 ( .A1(n10822), .A2(n11417), .B1(n2290), .B2(n11419), .ZN(
        n6439) );
  OAI22_X1 U4670 ( .A1(n10815), .A2(n11417), .B1(n2278), .B2(n11419), .ZN(
        n6438) );
  OAI22_X1 U4671 ( .A1(n10808), .A2(n11417), .B1(n2266), .B2(n11419), .ZN(
        n6437) );
  OAI22_X1 U4672 ( .A1(n10801), .A2(n11417), .B1(n2254), .B2(n11419), .ZN(
        n6436) );
  OAI22_X1 U4673 ( .A1(n10794), .A2(n11416), .B1(n2242), .B2(n11420), .ZN(
        n6435) );
  OAI22_X1 U4674 ( .A1(n10787), .A2(n11416), .B1(n2230), .B2(n11420), .ZN(
        n6434) );
  OAI22_X1 U4675 ( .A1(n10780), .A2(n11416), .B1(n2218), .B2(n11420), .ZN(
        n6433) );
  OAI22_X1 U4676 ( .A1(n10773), .A2(n11416), .B1(n2174), .B2(n11420), .ZN(
        n6432) );
  OAI22_X1 U4677 ( .A1(n10766), .A2(n11416), .B1(n2162), .B2(n11421), .ZN(
        n6431) );
  OAI22_X1 U4678 ( .A1(n10759), .A2(n11416), .B1(n2150), .B2(n11421), .ZN(
        n6430) );
  OAI22_X1 U4679 ( .A1(n10752), .A2(n11416), .B1(n2106), .B2(n11421), .ZN(
        n6429) );
  OAI22_X1 U4680 ( .A1(n10745), .A2(n11416), .B1(n2094), .B2(n11421), .ZN(
        n6428) );
  OAI22_X1 U4681 ( .A1(n10738), .A2(n11416), .B1(n2082), .B2(n11422), .ZN(
        n6427) );
  OAI22_X1 U4682 ( .A1(n10731), .A2(n11416), .B1(n2038), .B2(n11422), .ZN(
        n6426) );
  OAI22_X1 U4683 ( .A1(n10724), .A2(n11416), .B1(n2026), .B2(n11422), .ZN(
        n6425) );
  OAI22_X1 U4684 ( .A1(n10717), .A2(n11416), .B1(n2014), .B2(n11422), .ZN(
        n6424) );
  OAI22_X1 U4685 ( .A1(n10710), .A2(n11415), .B1(n2002), .B2(n11423), .ZN(
        n6423) );
  OAI22_X1 U4686 ( .A1(n10703), .A2(n11415), .B1(n1990), .B2(n11423), .ZN(
        n6422) );
  OAI22_X1 U4687 ( .A1(n10696), .A2(n11415), .B1(n1978), .B2(n11423), .ZN(
        n6421) );
  OAI22_X1 U4688 ( .A1(n10689), .A2(n11415), .B1(n1966), .B2(n11423), .ZN(
        n6420) );
  OAI22_X1 U4689 ( .A1(n10682), .A2(n11415), .B1(n1954), .B2(n11424), .ZN(
        n6419) );
  OAI22_X1 U4690 ( .A1(n10675), .A2(n11415), .B1(n1942), .B2(n11424), .ZN(
        n6418) );
  OAI22_X1 U4691 ( .A1(n10668), .A2(n11415), .B1(n1930), .B2(n11424), .ZN(
        n6417) );
  OAI22_X1 U4692 ( .A1(n10661), .A2(n11415), .B1(n1918), .B2(n11424), .ZN(
        n6416) );
  OAI22_X1 U4693 ( .A1(n10654), .A2(n11415), .B1(n1906), .B2(n11425), .ZN(
        n6415) );
  OAI22_X1 U4694 ( .A1(n10647), .A2(n11415), .B1(n1894), .B2(n11425), .ZN(
        n6414) );
  OAI22_X1 U4695 ( .A1(n10640), .A2(n11415), .B1(n1882), .B2(n11425), .ZN(
        n6413) );
  OAI22_X1 U4696 ( .A1(n10633), .A2(n11415), .B1(n1870), .B2(n11425), .ZN(
        n6412) );
  OAI22_X1 U4697 ( .A1(n10846), .A2(n12041), .B1(n10520), .B2(n12042), .ZN(
        n8107) );
  OAI22_X1 U4698 ( .A1(n10839), .A2(n12041), .B1(n10488), .B2(n12042), .ZN(
        n8106) );
  OAI22_X1 U4699 ( .A1(n10832), .A2(n12041), .B1(n10456), .B2(n12042), .ZN(
        n8105) );
  OAI22_X1 U4700 ( .A1(n10825), .A2(n12041), .B1(n10424), .B2(n12042), .ZN(
        n8104) );
  OAI22_X1 U4701 ( .A1(n10818), .A2(n12041), .B1(n10389), .B2(n12043), .ZN(
        n8103) );
  OAI22_X1 U4702 ( .A1(n10811), .A2(n12041), .B1(n10357), .B2(n12043), .ZN(
        n8102) );
  OAI22_X1 U4703 ( .A1(n10804), .A2(n12041), .B1(n10325), .B2(n12043), .ZN(
        n8101) );
  OAI22_X1 U4704 ( .A1(n10797), .A2(n12041), .B1(n10290), .B2(n12043), .ZN(
        n8100) );
  OAI22_X1 U4705 ( .A1(n10790), .A2(n12040), .B1(n10258), .B2(n12044), .ZN(
        n8099) );
  OAI22_X1 U4706 ( .A1(n10783), .A2(n12040), .B1(n10226), .B2(n12044), .ZN(
        n8098) );
  OAI22_X1 U4707 ( .A1(n10776), .A2(n12040), .B1(n10192), .B2(n12044), .ZN(
        n8097) );
  OAI22_X1 U4708 ( .A1(n10769), .A2(n12040), .B1(n10160), .B2(n12044), .ZN(
        n8096) );
  OAI22_X1 U4709 ( .A1(n10762), .A2(n12040), .B1(n10128), .B2(n12045), .ZN(
        n8095) );
  OAI22_X1 U4710 ( .A1(n10755), .A2(n12040), .B1(n10096), .B2(n12045), .ZN(
        n8094) );
  OAI22_X1 U4711 ( .A1(n10748), .A2(n12040), .B1(n10064), .B2(n12045), .ZN(
        n8093) );
  OAI22_X1 U4712 ( .A1(n10741), .A2(n12040), .B1(n10032), .B2(n12045), .ZN(
        n8092) );
  OAI22_X1 U4713 ( .A1(n10734), .A2(n12040), .B1(n10000), .B2(n12046), .ZN(
        n8091) );
  OAI22_X1 U4714 ( .A1(n10727), .A2(n12040), .B1(n9638), .B2(n12046), .ZN(
        n8090) );
  OAI22_X1 U4715 ( .A1(n10720), .A2(n12040), .B1(n9606), .B2(n12046), .ZN(
        n8089) );
  OAI22_X1 U4716 ( .A1(n10713), .A2(n12040), .B1(n9574), .B2(n12046), .ZN(
        n8088) );
  OAI22_X1 U4717 ( .A1(n10706), .A2(n12039), .B1(n9208), .B2(n12047), .ZN(
        n8087) );
  OAI22_X1 U4718 ( .A1(n10699), .A2(n12039), .B1(n9176), .B2(n12047), .ZN(
        n8086) );
  OAI22_X1 U4719 ( .A1(n10692), .A2(n12039), .B1(n9144), .B2(n12047), .ZN(
        n8085) );
  OAI22_X1 U4720 ( .A1(n10685), .A2(n12039), .B1(n6009), .B2(n12047), .ZN(
        n8084) );
  OAI22_X1 U4721 ( .A1(n10678), .A2(n12039), .B1(n5945), .B2(n12048), .ZN(
        n8083) );
  OAI22_X1 U4722 ( .A1(n10671), .A2(n12039), .B1(n5913), .B2(n12048), .ZN(
        n8082) );
  OAI22_X1 U4723 ( .A1(n10664), .A2(n12039), .B1(n5881), .B2(n12048), .ZN(
        n8081) );
  OAI22_X1 U4724 ( .A1(n10657), .A2(n12039), .B1(n5849), .B2(n12048), .ZN(
        n8080) );
  OAI22_X1 U4725 ( .A1(n10650), .A2(n12039), .B1(n5817), .B2(n12049), .ZN(
        n8079) );
  OAI22_X1 U4726 ( .A1(n10643), .A2(n12039), .B1(n5785), .B2(n12049), .ZN(
        n8078) );
  OAI22_X1 U4727 ( .A1(n10636), .A2(n12039), .B1(n5753), .B2(n12049), .ZN(
        n8077) );
  OAI22_X1 U4728 ( .A1(n10629), .A2(n12039), .B1(n5721), .B2(n12049), .ZN(
        n8076) );
  OAI22_X1 U4729 ( .A1(n10848), .A2(n11777), .B1(n10528), .B2(n11778), .ZN(
        n7403) );
  OAI22_X1 U4730 ( .A1(n10841), .A2(n11777), .B1(n10496), .B2(n11778), .ZN(
        n7402) );
  OAI22_X1 U4731 ( .A1(n10834), .A2(n11777), .B1(n10464), .B2(n11778), .ZN(
        n7401) );
  OAI22_X1 U4732 ( .A1(n10827), .A2(n11777), .B1(n10432), .B2(n11778), .ZN(
        n7400) );
  OAI22_X1 U4733 ( .A1(n10820), .A2(n11777), .B1(n10400), .B2(n11779), .ZN(
        n7399) );
  OAI22_X1 U4734 ( .A1(n10813), .A2(n11777), .B1(n10365), .B2(n11779), .ZN(
        n7398) );
  OAI22_X1 U4735 ( .A1(n10806), .A2(n11777), .B1(n10333), .B2(n11779), .ZN(
        n7397) );
  OAI22_X1 U4736 ( .A1(n10799), .A2(n11777), .B1(n10298), .B2(n11779), .ZN(
        n7396) );
  OAI22_X1 U4737 ( .A1(n10792), .A2(n11776), .B1(n10266), .B2(n11780), .ZN(
        n7395) );
  OAI22_X1 U4738 ( .A1(n10785), .A2(n11776), .B1(n10234), .B2(n11780), .ZN(
        n7394) );
  OAI22_X1 U4739 ( .A1(n10778), .A2(n11776), .B1(n10200), .B2(n11780), .ZN(
        n7393) );
  OAI22_X1 U4740 ( .A1(n10771), .A2(n11776), .B1(n10168), .B2(n11780), .ZN(
        n7392) );
  OAI22_X1 U4741 ( .A1(n10764), .A2(n11776), .B1(n10136), .B2(n11781), .ZN(
        n7391) );
  OAI22_X1 U4742 ( .A1(n10757), .A2(n11776), .B1(n10104), .B2(n11781), .ZN(
        n7390) );
  OAI22_X1 U4743 ( .A1(n10750), .A2(n11776), .B1(n10072), .B2(n11781), .ZN(
        n7389) );
  OAI22_X1 U4744 ( .A1(n10743), .A2(n11776), .B1(n10040), .B2(n11781), .ZN(
        n7388) );
  OAI22_X1 U4745 ( .A1(n10736), .A2(n11776), .B1(n10008), .B2(n11782), .ZN(
        n7387) );
  OAI22_X1 U4746 ( .A1(n10729), .A2(n11776), .B1(n9646), .B2(n11782), .ZN(
        n7386) );
  OAI22_X1 U4747 ( .A1(n10722), .A2(n11776), .B1(n9614), .B2(n11782), .ZN(
        n7385) );
  OAI22_X1 U4748 ( .A1(n10715), .A2(n11776), .B1(n9582), .B2(n11782), .ZN(
        n7384) );
  OAI22_X1 U4749 ( .A1(n10708), .A2(n11775), .B1(n9248), .B2(n11783), .ZN(
        n7383) );
  OAI22_X1 U4750 ( .A1(n10701), .A2(n11775), .B1(n9184), .B2(n11783), .ZN(
        n7382) );
  OAI22_X1 U4751 ( .A1(n10694), .A2(n11775), .B1(n9152), .B2(n11783), .ZN(
        n7381) );
  OAI22_X1 U4752 ( .A1(n10687), .A2(n11775), .B1(n6302), .B2(n11783), .ZN(
        n7380) );
  OAI22_X1 U4753 ( .A1(n10680), .A2(n11775), .B1(n5985), .B2(n11784), .ZN(
        n7379) );
  OAI22_X1 U4754 ( .A1(n10673), .A2(n11775), .B1(n5921), .B2(n11784), .ZN(
        n7378) );
  OAI22_X1 U4755 ( .A1(n10666), .A2(n11775), .B1(n5889), .B2(n11784), .ZN(
        n7377) );
  OAI22_X1 U4756 ( .A1(n10659), .A2(n11775), .B1(n5857), .B2(n11784), .ZN(
        n7376) );
  OAI22_X1 U4757 ( .A1(n10652), .A2(n11775), .B1(n5825), .B2(n11785), .ZN(
        n7375) );
  OAI22_X1 U4758 ( .A1(n10645), .A2(n11775), .B1(n5793), .B2(n11785), .ZN(
        n7374) );
  OAI22_X1 U4759 ( .A1(n10638), .A2(n11775), .B1(n5761), .B2(n11785), .ZN(
        n7373) );
  OAI22_X1 U4760 ( .A1(n10631), .A2(n11775), .B1(n5729), .B2(n11785), .ZN(
        n7372) );
  OAI22_X1 U4761 ( .A1(n10850), .A2(n11393), .B1(n515), .B2(n11394), .ZN(n6379) );
  OAI22_X1 U4762 ( .A1(n10843), .A2(n11393), .B1(n503), .B2(n11394), .ZN(n6378) );
  OAI22_X1 U4763 ( .A1(n10836), .A2(n11393), .B1(n491), .B2(n11394), .ZN(n6377) );
  OAI22_X1 U4764 ( .A1(n10829), .A2(n11393), .B1(n479), .B2(n11394), .ZN(n6376) );
  OAI22_X1 U4765 ( .A1(n10822), .A2(n11393), .B1(n467), .B2(n11395), .ZN(n6375) );
  OAI22_X1 U4766 ( .A1(n10815), .A2(n11393), .B1(n455), .B2(n11395), .ZN(n6374) );
  OAI22_X1 U4767 ( .A1(n10808), .A2(n11393), .B1(n443), .B2(n11395), .ZN(n6373) );
  OAI22_X1 U4768 ( .A1(n10801), .A2(n11393), .B1(n431), .B2(n11395), .ZN(n6372) );
  OAI22_X1 U4769 ( .A1(n10794), .A2(n11392), .B1(n419), .B2(n11396), .ZN(n6371) );
  OAI22_X1 U4770 ( .A1(n10787), .A2(n11392), .B1(n407), .B2(n11396), .ZN(n6370) );
  OAI22_X1 U4771 ( .A1(n10780), .A2(n11392), .B1(n395), .B2(n11396), .ZN(n6369) );
  OAI22_X1 U4772 ( .A1(n10773), .A2(n11392), .B1(n383), .B2(n11396), .ZN(n6368) );
  OAI22_X1 U4773 ( .A1(n10766), .A2(n11392), .B1(n371), .B2(n11397), .ZN(n6367) );
  OAI22_X1 U4774 ( .A1(n10759), .A2(n11392), .B1(n359), .B2(n11397), .ZN(n6366) );
  OAI22_X1 U4775 ( .A1(n10752), .A2(n11392), .B1(n347), .B2(n11397), .ZN(n6365) );
  OAI22_X1 U4776 ( .A1(n10745), .A2(n11392), .B1(n335), .B2(n11397), .ZN(n6364) );
  OAI22_X1 U4777 ( .A1(n10738), .A2(n11392), .B1(n323), .B2(n11398), .ZN(n6363) );
  OAI22_X1 U4778 ( .A1(n10731), .A2(n11392), .B1(n311), .B2(n11398), .ZN(n6362) );
  OAI22_X1 U4779 ( .A1(n10724), .A2(n11392), .B1(n299), .B2(n11398), .ZN(n6361) );
  OAI22_X1 U4780 ( .A1(n10717), .A2(n11392), .B1(n287), .B2(n11398), .ZN(n6360) );
  OAI22_X1 U4781 ( .A1(n10710), .A2(n11391), .B1(n275), .B2(n11399), .ZN(n6359) );
  OAI22_X1 U4782 ( .A1(n10703), .A2(n11391), .B1(n263), .B2(n11399), .ZN(n6358) );
  OAI22_X1 U4783 ( .A1(n10696), .A2(n11391), .B1(n251), .B2(n11399), .ZN(n6357) );
  OAI22_X1 U4784 ( .A1(n10689), .A2(n11391), .B1(n239), .B2(n11399), .ZN(n6356) );
  OAI22_X1 U4785 ( .A1(n10682), .A2(n11391), .B1(n227), .B2(n11400), .ZN(n6355) );
  OAI22_X1 U4786 ( .A1(n10675), .A2(n11391), .B1(n215), .B2(n11400), .ZN(n6354) );
  OAI22_X1 U4787 ( .A1(n10668), .A2(n11391), .B1(n203), .B2(n11400), .ZN(n6353) );
  OAI22_X1 U4788 ( .A1(n10661), .A2(n11391), .B1(n191), .B2(n11400), .ZN(n6352) );
  OAI22_X1 U4789 ( .A1(n10654), .A2(n11391), .B1(n179), .B2(n11401), .ZN(n6351) );
  OAI22_X1 U4790 ( .A1(n10647), .A2(n11391), .B1(n167), .B2(n11401), .ZN(n6350) );
  OAI22_X1 U4791 ( .A1(n10640), .A2(n11391), .B1(n155), .B2(n11401), .ZN(n6349) );
  OAI22_X1 U4792 ( .A1(n10633), .A2(n11391), .B1(n143), .B2(n11401), .ZN(n6348) );
  OAI22_X1 U4793 ( .A1(n10845), .A2(n12149), .B1(n10521), .B2(n12150), .ZN(
        n8395) );
  OAI22_X1 U4794 ( .A1(n10838), .A2(n12149), .B1(n10489), .B2(n12150), .ZN(
        n8394) );
  OAI22_X1 U4795 ( .A1(n10831), .A2(n12149), .B1(n10457), .B2(n12150), .ZN(
        n8393) );
  OAI22_X1 U4796 ( .A1(n10824), .A2(n12149), .B1(n10425), .B2(n12150), .ZN(
        n8392) );
  OAI22_X1 U4797 ( .A1(n10817), .A2(n12149), .B1(n10390), .B2(n12151), .ZN(
        n8391) );
  OAI22_X1 U4798 ( .A1(n10810), .A2(n12149), .B1(n10358), .B2(n12151), .ZN(
        n8390) );
  OAI22_X1 U4799 ( .A1(n10803), .A2(n12149), .B1(n10326), .B2(n12151), .ZN(
        n8389) );
  OAI22_X1 U4800 ( .A1(n10796), .A2(n12149), .B1(n10291), .B2(n12151), .ZN(
        n8388) );
  OAI22_X1 U4801 ( .A1(n10789), .A2(n12148), .B1(n10259), .B2(n12152), .ZN(
        n8387) );
  OAI22_X1 U4802 ( .A1(n10782), .A2(n12148), .B1(n10227), .B2(n12152), .ZN(
        n8386) );
  OAI22_X1 U4803 ( .A1(n10775), .A2(n12148), .B1(n10193), .B2(n12152), .ZN(
        n8385) );
  OAI22_X1 U4804 ( .A1(n10768), .A2(n12148), .B1(n10161), .B2(n12152), .ZN(
        n8384) );
  OAI22_X1 U4805 ( .A1(n10761), .A2(n12148), .B1(n10129), .B2(n12153), .ZN(
        n8383) );
  OAI22_X1 U4806 ( .A1(n10754), .A2(n12148), .B1(n10097), .B2(n12153), .ZN(
        n8382) );
  OAI22_X1 U4807 ( .A1(n10747), .A2(n12148), .B1(n10065), .B2(n12153), .ZN(
        n8381) );
  OAI22_X1 U4808 ( .A1(n10740), .A2(n12148), .B1(n10033), .B2(n12153), .ZN(
        n8380) );
  OAI22_X1 U4809 ( .A1(n10733), .A2(n12148), .B1(n10001), .B2(n12154), .ZN(
        n8379) );
  OAI22_X1 U4810 ( .A1(n10726), .A2(n12148), .B1(n9639), .B2(n12154), .ZN(
        n8378) );
  OAI22_X1 U4811 ( .A1(n10719), .A2(n12148), .B1(n9607), .B2(n12154), .ZN(
        n8377) );
  OAI22_X1 U4812 ( .A1(n10712), .A2(n12148), .B1(n9575), .B2(n12154), .ZN(
        n8376) );
  OAI22_X1 U4813 ( .A1(n10705), .A2(n12147), .B1(n9209), .B2(n12155), .ZN(
        n8375) );
  OAI22_X1 U4814 ( .A1(n10698), .A2(n12147), .B1(n9177), .B2(n12155), .ZN(
        n8374) );
  OAI22_X1 U4815 ( .A1(n10691), .A2(n12147), .B1(n9145), .B2(n12155), .ZN(
        n8373) );
  OAI22_X1 U4816 ( .A1(n10684), .A2(n12147), .B1(n6010), .B2(n12155), .ZN(
        n8372) );
  OAI22_X1 U4817 ( .A1(n10677), .A2(n12147), .B1(n5946), .B2(n12156), .ZN(
        n8371) );
  OAI22_X1 U4818 ( .A1(n10670), .A2(n12147), .B1(n5914), .B2(n12156), .ZN(
        n8370) );
  OAI22_X1 U4819 ( .A1(n10663), .A2(n12147), .B1(n5882), .B2(n12156), .ZN(
        n8369) );
  OAI22_X1 U4820 ( .A1(n10656), .A2(n12147), .B1(n5850), .B2(n12156), .ZN(
        n8368) );
  OAI22_X1 U4821 ( .A1(n10649), .A2(n12147), .B1(n5818), .B2(n12157), .ZN(
        n8367) );
  OAI22_X1 U4822 ( .A1(n10642), .A2(n12147), .B1(n5786), .B2(n12157), .ZN(
        n8366) );
  OAI22_X1 U4823 ( .A1(n10635), .A2(n12147), .B1(n5754), .B2(n12157), .ZN(
        n8365) );
  OAI22_X1 U4824 ( .A1(n10628), .A2(n12147), .B1(n5722), .B2(n12157), .ZN(
        n8364) );
  OAI22_X1 U4825 ( .A1(n10847), .A2(n11885), .B1(n10529), .B2(n11886), .ZN(
        n7691) );
  OAI22_X1 U4826 ( .A1(n10840), .A2(n11885), .B1(n10497), .B2(n11886), .ZN(
        n7690) );
  OAI22_X1 U4827 ( .A1(n10833), .A2(n11885), .B1(n10465), .B2(n11886), .ZN(
        n7689) );
  OAI22_X1 U4828 ( .A1(n10826), .A2(n11885), .B1(n10433), .B2(n11886), .ZN(
        n7688) );
  OAI22_X1 U4829 ( .A1(n10819), .A2(n11885), .B1(n10401), .B2(n11887), .ZN(
        n7687) );
  OAI22_X1 U4830 ( .A1(n10812), .A2(n11885), .B1(n10366), .B2(n11887), .ZN(
        n7686) );
  OAI22_X1 U4831 ( .A1(n10805), .A2(n11885), .B1(n10334), .B2(n11887), .ZN(
        n7685) );
  OAI22_X1 U4832 ( .A1(n10798), .A2(n11885), .B1(n10299), .B2(n11887), .ZN(
        n7684) );
  OAI22_X1 U4833 ( .A1(n10791), .A2(n11884), .B1(n10267), .B2(n11888), .ZN(
        n7683) );
  OAI22_X1 U4834 ( .A1(n10784), .A2(n11884), .B1(n10235), .B2(n11888), .ZN(
        n7682) );
  OAI22_X1 U4835 ( .A1(n10777), .A2(n11884), .B1(n10201), .B2(n11888), .ZN(
        n7681) );
  OAI22_X1 U4836 ( .A1(n10770), .A2(n11884), .B1(n10169), .B2(n11888), .ZN(
        n7680) );
  OAI22_X1 U4837 ( .A1(n10763), .A2(n11884), .B1(n10137), .B2(n11889), .ZN(
        n7679) );
  OAI22_X1 U4838 ( .A1(n10756), .A2(n11884), .B1(n10105), .B2(n11889), .ZN(
        n7678) );
  OAI22_X1 U4839 ( .A1(n10749), .A2(n11884), .B1(n10073), .B2(n11889), .ZN(
        n7677) );
  OAI22_X1 U4840 ( .A1(n10742), .A2(n11884), .B1(n10041), .B2(n11889), .ZN(
        n7676) );
  OAI22_X1 U4841 ( .A1(n10735), .A2(n11884), .B1(n10009), .B2(n11890), .ZN(
        n7675) );
  OAI22_X1 U4842 ( .A1(n10728), .A2(n11884), .B1(n9647), .B2(n11890), .ZN(
        n7674) );
  OAI22_X1 U4843 ( .A1(n10721), .A2(n11884), .B1(n9615), .B2(n11890), .ZN(
        n7673) );
  OAI22_X1 U4844 ( .A1(n10714), .A2(n11884), .B1(n9583), .B2(n11890), .ZN(
        n7672) );
  OAI22_X1 U4845 ( .A1(n10707), .A2(n11883), .B1(n9249), .B2(n11891), .ZN(
        n7671) );
  OAI22_X1 U4846 ( .A1(n10700), .A2(n11883), .B1(n9185), .B2(n11891), .ZN(
        n7670) );
  OAI22_X1 U4847 ( .A1(n10693), .A2(n11883), .B1(n9153), .B2(n11891), .ZN(
        n7669) );
  OAI22_X1 U4848 ( .A1(n10686), .A2(n11883), .B1(n6303), .B2(n11891), .ZN(
        n7668) );
  OAI22_X1 U4849 ( .A1(n10679), .A2(n11883), .B1(n5986), .B2(n11892), .ZN(
        n7667) );
  OAI22_X1 U4850 ( .A1(n10672), .A2(n11883), .B1(n5922), .B2(n11892), .ZN(
        n7666) );
  OAI22_X1 U4851 ( .A1(n10665), .A2(n11883), .B1(n5890), .B2(n11892), .ZN(
        n7665) );
  OAI22_X1 U4852 ( .A1(n10658), .A2(n11883), .B1(n5858), .B2(n11892), .ZN(
        n7664) );
  OAI22_X1 U4853 ( .A1(n10651), .A2(n11883), .B1(n5826), .B2(n11893), .ZN(
        n7663) );
  OAI22_X1 U4854 ( .A1(n10644), .A2(n11883), .B1(n5794), .B2(n11893), .ZN(
        n7662) );
  OAI22_X1 U4855 ( .A1(n10637), .A2(n11883), .B1(n5762), .B2(n11893), .ZN(
        n7661) );
  OAI22_X1 U4856 ( .A1(n10630), .A2(n11883), .B1(n5730), .B2(n11893), .ZN(
        n7660) );
  OAI22_X1 U4857 ( .A1(n10850), .A2(n11381), .B1(n2339), .B2(n11382), .ZN(
        n6347) );
  OAI22_X1 U4858 ( .A1(n10843), .A2(n11381), .B1(n2327), .B2(n11382), .ZN(
        n6346) );
  OAI22_X1 U4859 ( .A1(n10836), .A2(n11381), .B1(n2315), .B2(n11382), .ZN(
        n6345) );
  OAI22_X1 U4860 ( .A1(n10829), .A2(n11381), .B1(n2303), .B2(n11382), .ZN(
        n6344) );
  OAI22_X1 U4861 ( .A1(n10822), .A2(n11381), .B1(n2291), .B2(n11383), .ZN(
        n6343) );
  OAI22_X1 U4862 ( .A1(n10815), .A2(n11381), .B1(n2279), .B2(n11383), .ZN(
        n6342) );
  OAI22_X1 U4863 ( .A1(n10808), .A2(n11381), .B1(n2267), .B2(n11383), .ZN(
        n6341) );
  OAI22_X1 U4864 ( .A1(n10801), .A2(n11381), .B1(n2255), .B2(n11383), .ZN(
        n6340) );
  OAI22_X1 U4865 ( .A1(n10794), .A2(n11380), .B1(n2243), .B2(n11384), .ZN(
        n6339) );
  OAI22_X1 U4866 ( .A1(n10787), .A2(n11380), .B1(n2231), .B2(n11384), .ZN(
        n6338) );
  OAI22_X1 U4867 ( .A1(n10780), .A2(n11380), .B1(n2219), .B2(n11384), .ZN(
        n6337) );
  OAI22_X1 U4868 ( .A1(n10773), .A2(n11380), .B1(n2175), .B2(n11384), .ZN(
        n6336) );
  OAI22_X1 U4869 ( .A1(n10766), .A2(n11380), .B1(n2163), .B2(n11385), .ZN(
        n6335) );
  OAI22_X1 U4870 ( .A1(n10759), .A2(n11380), .B1(n2151), .B2(n11385), .ZN(
        n6334) );
  OAI22_X1 U4871 ( .A1(n10752), .A2(n11380), .B1(n2107), .B2(n11385), .ZN(
        n6333) );
  OAI22_X1 U4872 ( .A1(n10745), .A2(n11380), .B1(n2095), .B2(n11385), .ZN(
        n6332) );
  OAI22_X1 U4873 ( .A1(n10738), .A2(n11380), .B1(n2083), .B2(n11386), .ZN(
        n6331) );
  OAI22_X1 U4874 ( .A1(n10731), .A2(n11380), .B1(n2039), .B2(n11386), .ZN(
        n6330) );
  OAI22_X1 U4875 ( .A1(n10724), .A2(n11380), .B1(n2027), .B2(n11386), .ZN(
        n6329) );
  OAI22_X1 U4876 ( .A1(n10717), .A2(n11380), .B1(n2015), .B2(n11386), .ZN(
        n6328) );
  OAI22_X1 U4877 ( .A1(n10710), .A2(n11379), .B1(n2003), .B2(n11387), .ZN(
        n6327) );
  OAI22_X1 U4878 ( .A1(n10703), .A2(n11379), .B1(n1991), .B2(n11387), .ZN(
        n6326) );
  OAI22_X1 U4879 ( .A1(n10696), .A2(n11379), .B1(n1979), .B2(n11387), .ZN(
        n6325) );
  OAI22_X1 U4880 ( .A1(n10689), .A2(n11379), .B1(n1967), .B2(n11387), .ZN(
        n6324) );
  OAI22_X1 U4881 ( .A1(n10682), .A2(n11379), .B1(n1955), .B2(n11388), .ZN(
        n6323) );
  OAI22_X1 U4882 ( .A1(n10675), .A2(n11379), .B1(n1943), .B2(n11388), .ZN(
        n6322) );
  OAI22_X1 U4883 ( .A1(n10668), .A2(n11379), .B1(n1931), .B2(n11388), .ZN(
        n6321) );
  OAI22_X1 U4884 ( .A1(n10661), .A2(n11379), .B1(n1919), .B2(n11388), .ZN(
        n6320) );
  OAI22_X1 U4885 ( .A1(n10654), .A2(n11379), .B1(n1907), .B2(n11389), .ZN(
        n6319) );
  OAI22_X1 U4886 ( .A1(n10647), .A2(n11379), .B1(n1895), .B2(n11389), .ZN(
        n6318) );
  OAI22_X1 U4887 ( .A1(n10640), .A2(n11379), .B1(n1883), .B2(n11389), .ZN(
        n6317) );
  OAI22_X1 U4888 ( .A1(n10633), .A2(n11379), .B1(n1871), .B2(n11389), .ZN(
        n6316) );
  OAI22_X1 U4889 ( .A1(n10844), .A2(n12406), .B1(n10513), .B2(n12407), .ZN(
        n9099) );
  OAI22_X1 U4890 ( .A1(n10837), .A2(n12405), .B1(n10481), .B2(n12407), .ZN(
        n9098) );
  OAI22_X1 U4891 ( .A1(n10830), .A2(n12406), .B1(n10449), .B2(n12407), .ZN(
        n9097) );
  OAI22_X1 U4892 ( .A1(n10823), .A2(n12405), .B1(n10417), .B2(n12407), .ZN(
        n9096) );
  OAI22_X1 U4893 ( .A1(n10816), .A2(n12406), .B1(n10382), .B2(n12408), .ZN(
        n9095) );
  OAI22_X1 U4894 ( .A1(n10809), .A2(n12405), .B1(n10350), .B2(n12408), .ZN(
        n9094) );
  OAI22_X1 U4895 ( .A1(n10802), .A2(n12406), .B1(n10318), .B2(n12408), .ZN(
        n9093) );
  OAI22_X1 U4896 ( .A1(n10795), .A2(n12405), .B1(n10283), .B2(n12408), .ZN(
        n9092) );
  OAI22_X1 U4897 ( .A1(n10788), .A2(n12406), .B1(n10251), .B2(n12409), .ZN(
        n9091) );
  OAI22_X1 U4898 ( .A1(n10781), .A2(n12406), .B1(n10219), .B2(n12409), .ZN(
        n9090) );
  OAI22_X1 U4899 ( .A1(n10774), .A2(n12406), .B1(n10185), .B2(n12409), .ZN(
        n9089) );
  OAI22_X1 U4900 ( .A1(n10767), .A2(n12406), .B1(n10153), .B2(n12409), .ZN(
        n9088) );
  OAI22_X1 U4901 ( .A1(n10760), .A2(n12406), .B1(n10121), .B2(n12410), .ZN(
        n9087) );
  OAI22_X1 U4902 ( .A1(n10753), .A2(n12406), .B1(n10089), .B2(n12410), .ZN(
        n9086) );
  OAI22_X1 U4903 ( .A1(n10746), .A2(n12406), .B1(n10057), .B2(n12410), .ZN(
        n9085) );
  OAI22_X1 U4904 ( .A1(n10739), .A2(n12406), .B1(n10025), .B2(n12410), .ZN(
        n9084) );
  OAI22_X1 U4905 ( .A1(n10732), .A2(n12406), .B1(n9663), .B2(n12411), .ZN(
        n9083) );
  OAI22_X1 U4906 ( .A1(n10725), .A2(n12406), .B1(n9631), .B2(n12411), .ZN(
        n9082) );
  OAI22_X1 U4907 ( .A1(n10718), .A2(n12406), .B1(n9599), .B2(n12411), .ZN(
        n9081) );
  OAI22_X1 U4908 ( .A1(n10711), .A2(n12406), .B1(n9311), .B2(n12411), .ZN(
        n9080) );
  OAI22_X1 U4909 ( .A1(n10704), .A2(n12405), .B1(n9201), .B2(n12412), .ZN(
        n9079) );
  OAI22_X1 U4910 ( .A1(n10697), .A2(n12405), .B1(n9169), .B2(n12412), .ZN(
        n9078) );
  OAI22_X1 U4911 ( .A1(n10690), .A2(n12405), .B1(n9137), .B2(n12412), .ZN(
        n9077) );
  OAI22_X1 U4912 ( .A1(n10683), .A2(n12405), .B1(n6002), .B2(n12412), .ZN(
        n9076) );
  OAI22_X1 U4913 ( .A1(n10676), .A2(n12405), .B1(n5938), .B2(n12413), .ZN(
        n9075) );
  OAI22_X1 U4914 ( .A1(n10669), .A2(n12405), .B1(n5906), .B2(n12413), .ZN(
        n9074) );
  OAI22_X1 U4915 ( .A1(n10662), .A2(n12405), .B1(n5874), .B2(n12413), .ZN(
        n9073) );
  OAI22_X1 U4916 ( .A1(n10655), .A2(n12405), .B1(n5842), .B2(n12413), .ZN(
        n9072) );
  OAI22_X1 U4917 ( .A1(n10648), .A2(n12405), .B1(n5810), .B2(n12414), .ZN(
        n9071) );
  OAI22_X1 U4918 ( .A1(n10641), .A2(n12405), .B1(n5778), .B2(n12414), .ZN(
        n9070) );
  OAI22_X1 U4919 ( .A1(n10634), .A2(n12405), .B1(n5746), .B2(n12414), .ZN(
        n9069) );
  OAI22_X1 U4920 ( .A1(n10627), .A2(n12405), .B1(n5714), .B2(n12414), .ZN(
        n9068) );
  OAI22_X1 U4921 ( .A1(n10844), .A2(n12395), .B1(n2849), .B2(n12396), .ZN(
        n9067) );
  OAI22_X1 U4922 ( .A1(n10837), .A2(n12394), .B1(n2848), .B2(n12396), .ZN(
        n9066) );
  OAI22_X1 U4923 ( .A1(n10830), .A2(n12395), .B1(n2847), .B2(n12396), .ZN(
        n9065) );
  OAI22_X1 U4924 ( .A1(n10823), .A2(n12394), .B1(n2846), .B2(n12396), .ZN(
        n9064) );
  OAI22_X1 U4925 ( .A1(n10816), .A2(n12395), .B1(n2845), .B2(n12397), .ZN(
        n9063) );
  OAI22_X1 U4926 ( .A1(n10809), .A2(n12394), .B1(n2844), .B2(n12397), .ZN(
        n9062) );
  OAI22_X1 U4927 ( .A1(n10802), .A2(n12395), .B1(n2843), .B2(n12397), .ZN(
        n9061) );
  OAI22_X1 U4928 ( .A1(n10795), .A2(n12394), .B1(n2842), .B2(n12397), .ZN(
        n9060) );
  OAI22_X1 U4929 ( .A1(n10788), .A2(n12395), .B1(n2841), .B2(n12398), .ZN(
        n9059) );
  OAI22_X1 U4930 ( .A1(n10781), .A2(n12395), .B1(n2840), .B2(n12398), .ZN(
        n9058) );
  OAI22_X1 U4931 ( .A1(n10774), .A2(n12395), .B1(n2839), .B2(n12398), .ZN(
        n9057) );
  OAI22_X1 U4932 ( .A1(n10767), .A2(n12395), .B1(n2838), .B2(n12398), .ZN(
        n9056) );
  OAI22_X1 U4933 ( .A1(n10760), .A2(n12395), .B1(n2837), .B2(n12399), .ZN(
        n9055) );
  OAI22_X1 U4934 ( .A1(n10753), .A2(n12395), .B1(n2836), .B2(n12399), .ZN(
        n9054) );
  OAI22_X1 U4935 ( .A1(n10746), .A2(n12395), .B1(n2835), .B2(n12399), .ZN(
        n9053) );
  OAI22_X1 U4936 ( .A1(n10739), .A2(n12395), .B1(n2834), .B2(n12399), .ZN(
        n9052) );
  OAI22_X1 U4937 ( .A1(n10732), .A2(n12395), .B1(n2833), .B2(n12400), .ZN(
        n9051) );
  OAI22_X1 U4938 ( .A1(n10725), .A2(n12395), .B1(n2832), .B2(n12400), .ZN(
        n9050) );
  OAI22_X1 U4939 ( .A1(n10718), .A2(n12395), .B1(n2831), .B2(n12400), .ZN(
        n9049) );
  OAI22_X1 U4940 ( .A1(n10711), .A2(n12395), .B1(n2830), .B2(n12400), .ZN(
        n9048) );
  OAI22_X1 U4941 ( .A1(n10704), .A2(n12394), .B1(n2829), .B2(n12401), .ZN(
        n9047) );
  OAI22_X1 U4942 ( .A1(n10697), .A2(n12394), .B1(n2828), .B2(n12401), .ZN(
        n9046) );
  OAI22_X1 U4943 ( .A1(n10690), .A2(n12394), .B1(n2827), .B2(n12401), .ZN(
        n9045) );
  OAI22_X1 U4944 ( .A1(n10683), .A2(n12394), .B1(n2826), .B2(n12401), .ZN(
        n9044) );
  OAI22_X1 U4945 ( .A1(n10676), .A2(n12394), .B1(n2825), .B2(n12402), .ZN(
        n9043) );
  OAI22_X1 U4946 ( .A1(n10669), .A2(n12394), .B1(n2824), .B2(n12402), .ZN(
        n9042) );
  OAI22_X1 U4947 ( .A1(n10662), .A2(n12394), .B1(n2823), .B2(n12402), .ZN(
        n9041) );
  OAI22_X1 U4948 ( .A1(n10655), .A2(n12394), .B1(n2822), .B2(n12402), .ZN(
        n9040) );
  OAI22_X1 U4949 ( .A1(n10648), .A2(n12394), .B1(n2821), .B2(n12403), .ZN(
        n9039) );
  OAI22_X1 U4950 ( .A1(n10641), .A2(n12394), .B1(n2820), .B2(n12403), .ZN(
        n9038) );
  OAI22_X1 U4951 ( .A1(n10634), .A2(n12394), .B1(n2819), .B2(n12403), .ZN(
        n9037) );
  OAI22_X1 U4952 ( .A1(n10627), .A2(n12394), .B1(n2818), .B2(n12403), .ZN(
        n9036) );
  OAI22_X1 U4953 ( .A1(n10844), .A2(n12384), .B1(n10507), .B2(n12385), .ZN(
        n9035) );
  OAI22_X1 U4954 ( .A1(n10837), .A2(n12383), .B1(n10475), .B2(n12385), .ZN(
        n9034) );
  OAI22_X1 U4955 ( .A1(n10830), .A2(n12384), .B1(n10443), .B2(n12385), .ZN(
        n9033) );
  OAI22_X1 U4956 ( .A1(n10823), .A2(n12383), .B1(n10411), .B2(n12385), .ZN(
        n9032) );
  OAI22_X1 U4957 ( .A1(n10816), .A2(n12384), .B1(n10376), .B2(n12386), .ZN(
        n9031) );
  OAI22_X1 U4958 ( .A1(n10809), .A2(n12383), .B1(n10344), .B2(n12386), .ZN(
        n9030) );
  OAI22_X1 U4959 ( .A1(n10802), .A2(n12384), .B1(n10312), .B2(n12386), .ZN(
        n9029) );
  OAI22_X1 U4960 ( .A1(n10795), .A2(n12383), .B1(n10277), .B2(n12386), .ZN(
        n9028) );
  OAI22_X1 U4961 ( .A1(n10788), .A2(n12384), .B1(n10245), .B2(n12387), .ZN(
        n9027) );
  OAI22_X1 U4962 ( .A1(n10781), .A2(n12384), .B1(n10213), .B2(n12387), .ZN(
        n9026) );
  OAI22_X1 U4963 ( .A1(n10774), .A2(n12384), .B1(n10179), .B2(n12387), .ZN(
        n9025) );
  OAI22_X1 U4964 ( .A1(n10767), .A2(n12384), .B1(n10147), .B2(n12387), .ZN(
        n9024) );
  OAI22_X1 U4965 ( .A1(n10760), .A2(n12384), .B1(n10115), .B2(n12388), .ZN(
        n9023) );
  OAI22_X1 U4966 ( .A1(n10753), .A2(n12384), .B1(n10083), .B2(n12388), .ZN(
        n9022) );
  OAI22_X1 U4967 ( .A1(n10746), .A2(n12384), .B1(n10051), .B2(n12388), .ZN(
        n9021) );
  OAI22_X1 U4968 ( .A1(n10739), .A2(n12384), .B1(n10019), .B2(n12388), .ZN(
        n9020) );
  OAI22_X1 U4969 ( .A1(n10732), .A2(n12384), .B1(n9657), .B2(n12389), .ZN(
        n9019) );
  OAI22_X1 U4970 ( .A1(n10725), .A2(n12384), .B1(n9625), .B2(n12389), .ZN(
        n9018) );
  OAI22_X1 U4971 ( .A1(n10718), .A2(n12384), .B1(n9593), .B2(n12389), .ZN(
        n9017) );
  OAI22_X1 U4972 ( .A1(n10711), .A2(n12384), .B1(n9259), .B2(n12389), .ZN(
        n9016) );
  OAI22_X1 U4973 ( .A1(n10704), .A2(n12383), .B1(n9195), .B2(n12390), .ZN(
        n9015) );
  OAI22_X1 U4974 ( .A1(n10697), .A2(n12383), .B1(n9163), .B2(n12390), .ZN(
        n9014) );
  OAI22_X1 U4975 ( .A1(n10690), .A2(n12383), .B1(n6313), .B2(n12390), .ZN(
        n9013) );
  OAI22_X1 U4976 ( .A1(n10683), .A2(n12383), .B1(n5996), .B2(n12390), .ZN(
        n9012) );
  OAI22_X1 U4977 ( .A1(n10676), .A2(n12383), .B1(n5932), .B2(n12391), .ZN(
        n9011) );
  OAI22_X1 U4978 ( .A1(n10669), .A2(n12383), .B1(n5900), .B2(n12391), .ZN(
        n9010) );
  OAI22_X1 U4979 ( .A1(n10662), .A2(n12383), .B1(n5868), .B2(n12391), .ZN(
        n9009) );
  OAI22_X1 U4980 ( .A1(n10655), .A2(n12383), .B1(n5836), .B2(n12391), .ZN(
        n9008) );
  OAI22_X1 U4981 ( .A1(n10648), .A2(n12383), .B1(n5804), .B2(n12392), .ZN(
        n9007) );
  OAI22_X1 U4982 ( .A1(n10641), .A2(n12383), .B1(n5772), .B2(n12392), .ZN(
        n9006) );
  OAI22_X1 U4983 ( .A1(n10634), .A2(n12383), .B1(n5740), .B2(n12392), .ZN(
        n9005) );
  OAI22_X1 U4984 ( .A1(n10627), .A2(n12383), .B1(n5708), .B2(n12392), .ZN(
        n9004) );
  OAI22_X1 U4985 ( .A1(n10844), .A2(n12373), .B1(n2785), .B2(n12374), .ZN(
        n9003) );
  OAI22_X1 U4986 ( .A1(n10837), .A2(n12372), .B1(n2784), .B2(n12374), .ZN(
        n9002) );
  OAI22_X1 U4987 ( .A1(n10830), .A2(n12373), .B1(n2783), .B2(n12374), .ZN(
        n9001) );
  OAI22_X1 U4988 ( .A1(n10823), .A2(n12372), .B1(n2782), .B2(n12374), .ZN(
        n9000) );
  OAI22_X1 U4989 ( .A1(n10816), .A2(n12373), .B1(n2781), .B2(n12375), .ZN(
        n8999) );
  OAI22_X1 U4990 ( .A1(n10809), .A2(n12372), .B1(n2780), .B2(n12375), .ZN(
        n8998) );
  OAI22_X1 U4991 ( .A1(n10802), .A2(n12373), .B1(n2779), .B2(n12375), .ZN(
        n8997) );
  OAI22_X1 U4992 ( .A1(n10795), .A2(n12372), .B1(n2778), .B2(n12375), .ZN(
        n8996) );
  OAI22_X1 U4993 ( .A1(n10788), .A2(n12373), .B1(n2777), .B2(n12376), .ZN(
        n8995) );
  OAI22_X1 U4994 ( .A1(n10781), .A2(n12373), .B1(n2776), .B2(n12376), .ZN(
        n8994) );
  OAI22_X1 U4995 ( .A1(n10774), .A2(n12373), .B1(n2775), .B2(n12376), .ZN(
        n8993) );
  OAI22_X1 U4996 ( .A1(n10767), .A2(n12373), .B1(n2774), .B2(n12376), .ZN(
        n8992) );
  OAI22_X1 U4997 ( .A1(n10760), .A2(n12373), .B1(n2773), .B2(n12377), .ZN(
        n8991) );
  OAI22_X1 U4998 ( .A1(n10753), .A2(n12373), .B1(n2772), .B2(n12377), .ZN(
        n8990) );
  OAI22_X1 U4999 ( .A1(n10746), .A2(n12373), .B1(n2771), .B2(n12377), .ZN(
        n8989) );
  OAI22_X1 U5000 ( .A1(n10739), .A2(n12373), .B1(n2770), .B2(n12377), .ZN(
        n8988) );
  OAI22_X1 U5001 ( .A1(n10732), .A2(n12373), .B1(n2769), .B2(n12378), .ZN(
        n8987) );
  OAI22_X1 U5002 ( .A1(n10725), .A2(n12373), .B1(n2768), .B2(n12378), .ZN(
        n8986) );
  OAI22_X1 U5003 ( .A1(n10718), .A2(n12373), .B1(n2767), .B2(n12378), .ZN(
        n8985) );
  OAI22_X1 U5004 ( .A1(n10711), .A2(n12373), .B1(n2766), .B2(n12378), .ZN(
        n8984) );
  OAI22_X1 U5005 ( .A1(n10704), .A2(n12372), .B1(n2765), .B2(n12379), .ZN(
        n8983) );
  OAI22_X1 U5006 ( .A1(n10697), .A2(n12372), .B1(n2764), .B2(n12379), .ZN(
        n8982) );
  OAI22_X1 U5007 ( .A1(n10690), .A2(n12372), .B1(n2763), .B2(n12379), .ZN(
        n8981) );
  OAI22_X1 U5008 ( .A1(n10683), .A2(n12372), .B1(n2762), .B2(n12379), .ZN(
        n8980) );
  OAI22_X1 U5009 ( .A1(n10676), .A2(n12372), .B1(n2761), .B2(n12380), .ZN(
        n8979) );
  OAI22_X1 U5010 ( .A1(n10669), .A2(n12372), .B1(n2760), .B2(n12380), .ZN(
        n8978) );
  OAI22_X1 U5011 ( .A1(n10662), .A2(n12372), .B1(n2759), .B2(n12380), .ZN(
        n8977) );
  OAI22_X1 U5012 ( .A1(n10655), .A2(n12372), .B1(n2758), .B2(n12380), .ZN(
        n8976) );
  OAI22_X1 U5013 ( .A1(n10648), .A2(n12372), .B1(n2757), .B2(n12381), .ZN(
        n8975) );
  OAI22_X1 U5014 ( .A1(n10641), .A2(n12372), .B1(n2756), .B2(n12381), .ZN(
        n8974) );
  OAI22_X1 U5015 ( .A1(n10634), .A2(n12372), .B1(n2755), .B2(n12381), .ZN(
        n8973) );
  OAI22_X1 U5016 ( .A1(n10627), .A2(n12372), .B1(n2754), .B2(n12381), .ZN(
        n8972) );
  OAI22_X1 U5017 ( .A1(n10844), .A2(n12362), .B1(n10506), .B2(n12363), .ZN(
        n8971) );
  OAI22_X1 U5018 ( .A1(n10837), .A2(n12361), .B1(n10474), .B2(n12363), .ZN(
        n8970) );
  OAI22_X1 U5019 ( .A1(n10830), .A2(n12362), .B1(n10442), .B2(n12363), .ZN(
        n8969) );
  OAI22_X1 U5020 ( .A1(n10823), .A2(n12361), .B1(n10410), .B2(n12363), .ZN(
        n8968) );
  OAI22_X1 U5021 ( .A1(n10816), .A2(n12362), .B1(n10375), .B2(n12364), .ZN(
        n8967) );
  OAI22_X1 U5022 ( .A1(n10809), .A2(n12361), .B1(n10343), .B2(n12364), .ZN(
        n8966) );
  OAI22_X1 U5023 ( .A1(n10802), .A2(n12362), .B1(n10311), .B2(n12364), .ZN(
        n8965) );
  OAI22_X1 U5024 ( .A1(n10795), .A2(n12361), .B1(n10276), .B2(n12364), .ZN(
        n8964) );
  OAI22_X1 U5025 ( .A1(n10788), .A2(n12362), .B1(n10244), .B2(n12365), .ZN(
        n8963) );
  OAI22_X1 U5026 ( .A1(n10781), .A2(n12362), .B1(n10212), .B2(n12365), .ZN(
        n8962) );
  OAI22_X1 U5027 ( .A1(n10774), .A2(n12362), .B1(n10178), .B2(n12365), .ZN(
        n8961) );
  OAI22_X1 U5028 ( .A1(n10767), .A2(n12362), .B1(n10146), .B2(n12365), .ZN(
        n8960) );
  OAI22_X1 U5029 ( .A1(n10760), .A2(n12362), .B1(n10114), .B2(n12366), .ZN(
        n8959) );
  OAI22_X1 U5030 ( .A1(n10753), .A2(n12362), .B1(n10082), .B2(n12366), .ZN(
        n8958) );
  OAI22_X1 U5031 ( .A1(n10746), .A2(n12362), .B1(n10050), .B2(n12366), .ZN(
        n8957) );
  OAI22_X1 U5032 ( .A1(n10739), .A2(n12362), .B1(n10018), .B2(n12366), .ZN(
        n8956) );
  OAI22_X1 U5033 ( .A1(n10732), .A2(n12362), .B1(n9656), .B2(n12367), .ZN(
        n8955) );
  OAI22_X1 U5034 ( .A1(n10725), .A2(n12362), .B1(n9624), .B2(n12367), .ZN(
        n8954) );
  OAI22_X1 U5035 ( .A1(n10718), .A2(n12362), .B1(n9592), .B2(n12367), .ZN(
        n8953) );
  OAI22_X1 U5036 ( .A1(n10711), .A2(n12362), .B1(n9258), .B2(n12367), .ZN(
        n8952) );
  OAI22_X1 U5037 ( .A1(n10704), .A2(n12361), .B1(n9194), .B2(n12368), .ZN(
        n8951) );
  OAI22_X1 U5038 ( .A1(n10697), .A2(n12361), .B1(n9162), .B2(n12368), .ZN(
        n8950) );
  OAI22_X1 U5039 ( .A1(n10690), .A2(n12361), .B1(n6312), .B2(n12368), .ZN(
        n8949) );
  OAI22_X1 U5040 ( .A1(n10683), .A2(n12361), .B1(n5995), .B2(n12368), .ZN(
        n8948) );
  OAI22_X1 U5041 ( .A1(n10676), .A2(n12361), .B1(n5931), .B2(n12369), .ZN(
        n8947) );
  OAI22_X1 U5042 ( .A1(n10669), .A2(n12361), .B1(n5899), .B2(n12369), .ZN(
        n8946) );
  OAI22_X1 U5043 ( .A1(n10662), .A2(n12361), .B1(n5867), .B2(n12369), .ZN(
        n8945) );
  OAI22_X1 U5044 ( .A1(n10655), .A2(n12361), .B1(n5835), .B2(n12369), .ZN(
        n8944) );
  OAI22_X1 U5045 ( .A1(n10648), .A2(n12361), .B1(n5803), .B2(n12370), .ZN(
        n8943) );
  OAI22_X1 U5046 ( .A1(n10641), .A2(n12361), .B1(n5771), .B2(n12370), .ZN(
        n8942) );
  OAI22_X1 U5047 ( .A1(n10634), .A2(n12361), .B1(n5739), .B2(n12370), .ZN(
        n8941) );
  OAI22_X1 U5048 ( .A1(n10627), .A2(n12361), .B1(n5707), .B2(n12370), .ZN(
        n8940) );
  OAI22_X1 U5049 ( .A1(n10844), .A2(n12351), .B1(n10508), .B2(n12352), .ZN(
        n8939) );
  OAI22_X1 U5050 ( .A1(n10837), .A2(n12350), .B1(n10476), .B2(n12352), .ZN(
        n8938) );
  OAI22_X1 U5051 ( .A1(n10830), .A2(n12351), .B1(n10444), .B2(n12352), .ZN(
        n8937) );
  OAI22_X1 U5052 ( .A1(n10823), .A2(n12350), .B1(n10412), .B2(n12352), .ZN(
        n8936) );
  OAI22_X1 U5053 ( .A1(n10816), .A2(n12351), .B1(n10377), .B2(n12353), .ZN(
        n8935) );
  OAI22_X1 U5054 ( .A1(n10809), .A2(n12350), .B1(n10345), .B2(n12353), .ZN(
        n8934) );
  OAI22_X1 U5055 ( .A1(n10802), .A2(n12351), .B1(n10313), .B2(n12353), .ZN(
        n8933) );
  OAI22_X1 U5056 ( .A1(n10795), .A2(n12350), .B1(n10278), .B2(n12353), .ZN(
        n8932) );
  OAI22_X1 U5057 ( .A1(n10788), .A2(n12351), .B1(n10246), .B2(n12354), .ZN(
        n8931) );
  OAI22_X1 U5058 ( .A1(n10781), .A2(n12351), .B1(n10214), .B2(n12354), .ZN(
        n8930) );
  OAI22_X1 U5059 ( .A1(n10774), .A2(n12351), .B1(n10180), .B2(n12354), .ZN(
        n8929) );
  OAI22_X1 U5060 ( .A1(n10767), .A2(n12351), .B1(n10148), .B2(n12354), .ZN(
        n8928) );
  OAI22_X1 U5061 ( .A1(n10760), .A2(n12351), .B1(n10116), .B2(n12355), .ZN(
        n8927) );
  OAI22_X1 U5062 ( .A1(n10753), .A2(n12351), .B1(n10084), .B2(n12355), .ZN(
        n8926) );
  OAI22_X1 U5063 ( .A1(n10746), .A2(n12351), .B1(n10052), .B2(n12355), .ZN(
        n8925) );
  OAI22_X1 U5064 ( .A1(n10739), .A2(n12351), .B1(n10020), .B2(n12355), .ZN(
        n8924) );
  OAI22_X1 U5065 ( .A1(n10732), .A2(n12351), .B1(n9658), .B2(n12356), .ZN(
        n8923) );
  OAI22_X1 U5066 ( .A1(n10725), .A2(n12351), .B1(n9626), .B2(n12356), .ZN(
        n8922) );
  OAI22_X1 U5067 ( .A1(n10718), .A2(n12351), .B1(n9594), .B2(n12356), .ZN(
        n8921) );
  OAI22_X1 U5068 ( .A1(n10711), .A2(n12351), .B1(n9260), .B2(n12356), .ZN(
        n8920) );
  OAI22_X1 U5069 ( .A1(n10704), .A2(n12350), .B1(n9196), .B2(n12357), .ZN(
        n8919) );
  OAI22_X1 U5070 ( .A1(n10697), .A2(n12350), .B1(n9164), .B2(n12357), .ZN(
        n8918) );
  OAI22_X1 U5071 ( .A1(n10690), .A2(n12350), .B1(n6314), .B2(n12357), .ZN(
        n8917) );
  OAI22_X1 U5072 ( .A1(n10683), .A2(n12350), .B1(n5997), .B2(n12357), .ZN(
        n8916) );
  OAI22_X1 U5073 ( .A1(n10676), .A2(n12350), .B1(n5933), .B2(n12358), .ZN(
        n8915) );
  OAI22_X1 U5074 ( .A1(n10669), .A2(n12350), .B1(n5901), .B2(n12358), .ZN(
        n8914) );
  OAI22_X1 U5075 ( .A1(n10662), .A2(n12350), .B1(n5869), .B2(n12358), .ZN(
        n8913) );
  OAI22_X1 U5076 ( .A1(n10655), .A2(n12350), .B1(n5837), .B2(n12358), .ZN(
        n8912) );
  OAI22_X1 U5077 ( .A1(n10648), .A2(n12350), .B1(n5805), .B2(n12359), .ZN(
        n8911) );
  OAI22_X1 U5078 ( .A1(n10641), .A2(n12350), .B1(n5773), .B2(n12359), .ZN(
        n8910) );
  OAI22_X1 U5079 ( .A1(n10634), .A2(n12350), .B1(n5741), .B2(n12359), .ZN(
        n8909) );
  OAI22_X1 U5080 ( .A1(n10627), .A2(n12350), .B1(n5709), .B2(n12359), .ZN(
        n8908) );
  OAI22_X1 U5081 ( .A1(n10844), .A2(n12305), .B1(n10512), .B2(n12306), .ZN(
        n8811) );
  OAI22_X1 U5082 ( .A1(n10837), .A2(n12305), .B1(n10480), .B2(n12306), .ZN(
        n8810) );
  OAI22_X1 U5083 ( .A1(n10830), .A2(n12305), .B1(n10448), .B2(n12306), .ZN(
        n8809) );
  OAI22_X1 U5084 ( .A1(n10823), .A2(n12305), .B1(n10416), .B2(n12306), .ZN(
        n8808) );
  OAI22_X1 U5085 ( .A1(n10816), .A2(n12305), .B1(n10381), .B2(n12307), .ZN(
        n8807) );
  OAI22_X1 U5086 ( .A1(n10809), .A2(n12305), .B1(n10349), .B2(n12307), .ZN(
        n8806) );
  OAI22_X1 U5087 ( .A1(n10802), .A2(n12305), .B1(n10317), .B2(n12307), .ZN(
        n8805) );
  OAI22_X1 U5088 ( .A1(n10795), .A2(n12305), .B1(n10282), .B2(n12307), .ZN(
        n8804) );
  OAI22_X1 U5089 ( .A1(n10788), .A2(n12304), .B1(n10250), .B2(n12308), .ZN(
        n8803) );
  OAI22_X1 U5090 ( .A1(n10781), .A2(n12304), .B1(n10218), .B2(n12308), .ZN(
        n8802) );
  OAI22_X1 U5091 ( .A1(n10774), .A2(n12304), .B1(n10184), .B2(n12308), .ZN(
        n8801) );
  OAI22_X1 U5092 ( .A1(n10767), .A2(n12304), .B1(n10152), .B2(n12308), .ZN(
        n8800) );
  OAI22_X1 U5093 ( .A1(n10760), .A2(n12304), .B1(n10120), .B2(n12309), .ZN(
        n8799) );
  OAI22_X1 U5094 ( .A1(n10753), .A2(n12304), .B1(n10088), .B2(n12309), .ZN(
        n8798) );
  OAI22_X1 U5095 ( .A1(n10746), .A2(n12304), .B1(n10056), .B2(n12309), .ZN(
        n8797) );
  OAI22_X1 U5096 ( .A1(n10739), .A2(n12304), .B1(n10024), .B2(n12309), .ZN(
        n8796) );
  OAI22_X1 U5097 ( .A1(n10732), .A2(n12304), .B1(n9662), .B2(n12310), .ZN(
        n8795) );
  OAI22_X1 U5098 ( .A1(n10725), .A2(n12304), .B1(n9630), .B2(n12310), .ZN(
        n8794) );
  OAI22_X1 U5099 ( .A1(n10718), .A2(n12304), .B1(n9598), .B2(n12310), .ZN(
        n8793) );
  OAI22_X1 U5100 ( .A1(n10711), .A2(n12304), .B1(n9264), .B2(n12310), .ZN(
        n8792) );
  OAI22_X1 U5101 ( .A1(n10704), .A2(n12303), .B1(n9200), .B2(n12311), .ZN(
        n8791) );
  OAI22_X1 U5102 ( .A1(n10697), .A2(n12303), .B1(n9168), .B2(n12311), .ZN(
        n8790) );
  OAI22_X1 U5103 ( .A1(n10690), .A2(n12303), .B1(n9136), .B2(n12311), .ZN(
        n8789) );
  OAI22_X1 U5104 ( .A1(n10683), .A2(n12303), .B1(n6001), .B2(n12311), .ZN(
        n8788) );
  OAI22_X1 U5105 ( .A1(n10676), .A2(n12303), .B1(n5937), .B2(n12312), .ZN(
        n8787) );
  OAI22_X1 U5106 ( .A1(n10669), .A2(n12303), .B1(n5905), .B2(n12312), .ZN(
        n8786) );
  OAI22_X1 U5107 ( .A1(n10662), .A2(n12303), .B1(n5873), .B2(n12312), .ZN(
        n8785) );
  OAI22_X1 U5108 ( .A1(n10655), .A2(n12303), .B1(n5841), .B2(n12312), .ZN(
        n8784) );
  OAI22_X1 U5109 ( .A1(n10648), .A2(n12303), .B1(n5809), .B2(n12313), .ZN(
        n8783) );
  OAI22_X1 U5110 ( .A1(n10641), .A2(n12303), .B1(n5777), .B2(n12313), .ZN(
        n8782) );
  OAI22_X1 U5111 ( .A1(n10634), .A2(n12303), .B1(n5745), .B2(n12313), .ZN(
        n8781) );
  OAI22_X1 U5112 ( .A1(n10627), .A2(n12303), .B1(n5713), .B2(n12313), .ZN(
        n8780) );
  OAI22_X1 U5113 ( .A1(n10846), .A2(n12017), .B1(n993), .B2(n12018), .ZN(n8043) );
  OAI22_X1 U5114 ( .A1(n10839), .A2(n12017), .B1(n989), .B2(n12018), .ZN(n8042) );
  OAI22_X1 U5115 ( .A1(n10832), .A2(n12017), .B1(n985), .B2(n12018), .ZN(n8041) );
  OAI22_X1 U5116 ( .A1(n10825), .A2(n12017), .B1(n981), .B2(n12018), .ZN(n8040) );
  OAI22_X1 U5117 ( .A1(n10818), .A2(n12017), .B1(n977), .B2(n12019), .ZN(n8039) );
  OAI22_X1 U5118 ( .A1(n10811), .A2(n12017), .B1(n973), .B2(n12019), .ZN(n8038) );
  OAI22_X1 U5119 ( .A1(n10804), .A2(n12017), .B1(n969), .B2(n12019), .ZN(n8037) );
  OAI22_X1 U5120 ( .A1(n10797), .A2(n12017), .B1(n965), .B2(n12019), .ZN(n8036) );
  OAI22_X1 U5121 ( .A1(n10790), .A2(n12016), .B1(n961), .B2(n12020), .ZN(n8035) );
  OAI22_X1 U5122 ( .A1(n10783), .A2(n12016), .B1(n957), .B2(n12020), .ZN(n8034) );
  OAI22_X1 U5123 ( .A1(n10776), .A2(n12016), .B1(n953), .B2(n12020), .ZN(n8033) );
  OAI22_X1 U5124 ( .A1(n10769), .A2(n12016), .B1(n949), .B2(n12020), .ZN(n8032) );
  OAI22_X1 U5125 ( .A1(n10762), .A2(n12016), .B1(n945), .B2(n12021), .ZN(n8031) );
  OAI22_X1 U5126 ( .A1(n10755), .A2(n12016), .B1(n941), .B2(n12021), .ZN(n8030) );
  OAI22_X1 U5127 ( .A1(n10748), .A2(n12016), .B1(n937), .B2(n12021), .ZN(n8029) );
  OAI22_X1 U5128 ( .A1(n10741), .A2(n12016), .B1(n933), .B2(n12021), .ZN(n8028) );
  OAI22_X1 U5129 ( .A1(n10734), .A2(n12016), .B1(n929), .B2(n12022), .ZN(n8027) );
  OAI22_X1 U5130 ( .A1(n10629), .A2(n12003), .B1(n999), .B2(n12006), .ZN(n7980) );
  OAI22_X1 U5131 ( .A1(n10848), .A2(n11753), .B1(n994), .B2(n11754), .ZN(n7339) );
  OAI22_X1 U5132 ( .A1(n10841), .A2(n11753), .B1(n990), .B2(n11754), .ZN(n7338) );
  OAI22_X1 U5133 ( .A1(n10834), .A2(n11753), .B1(n986), .B2(n11754), .ZN(n7337) );
  OAI22_X1 U5134 ( .A1(n10827), .A2(n11753), .B1(n982), .B2(n11754), .ZN(n7336) );
  OAI22_X1 U5135 ( .A1(n10820), .A2(n11753), .B1(n978), .B2(n11755), .ZN(n7335) );
  OAI22_X1 U5136 ( .A1(n10813), .A2(n11753), .B1(n974), .B2(n11755), .ZN(n7334) );
  OAI22_X1 U5137 ( .A1(n10737), .A2(n11644), .B1(n2048), .B2(n11646), .ZN(
        n7035) );
  OAI22_X1 U5138 ( .A1(n10730), .A2(n11644), .B1(n2036), .B2(n11646), .ZN(
        n7034) );
  OAI22_X1 U5139 ( .A1(n10723), .A2(n11644), .B1(n2024), .B2(n11646), .ZN(
        n7033) );
  OAI22_X1 U5140 ( .A1(n10716), .A2(n11644), .B1(n2012), .B2(n11646), .ZN(
        n7032) );
  OAI22_X1 U5141 ( .A1(n10709), .A2(n11643), .B1(n2000), .B2(n11647), .ZN(
        n7031) );
  OAI22_X1 U5142 ( .A1(n10702), .A2(n11643), .B1(n1988), .B2(n11647), .ZN(
        n7030) );
  OAI22_X1 U5143 ( .A1(n10695), .A2(n11643), .B1(n1976), .B2(n11647), .ZN(
        n7029) );
  OAI22_X1 U5144 ( .A1(n10688), .A2(n11643), .B1(n1964), .B2(n11647), .ZN(
        n7028) );
  OAI22_X1 U5145 ( .A1(n10681), .A2(n11643), .B1(n1952), .B2(n11648), .ZN(
        n7027) );
  OAI22_X1 U5146 ( .A1(n10674), .A2(n11643), .B1(n1940), .B2(n11648), .ZN(
        n7026) );
  OAI22_X1 U5147 ( .A1(n10667), .A2(n11643), .B1(n1928), .B2(n11648), .ZN(
        n7025) );
  OAI22_X1 U5148 ( .A1(n10660), .A2(n11643), .B1(n1916), .B2(n11648), .ZN(
        n7024) );
  OAI22_X1 U5149 ( .A1(n10653), .A2(n11643), .B1(n1904), .B2(n11649), .ZN(
        n7023) );
  OAI22_X1 U5150 ( .A1(n10646), .A2(n11643), .B1(n1892), .B2(n11649), .ZN(
        n7022) );
  OAI22_X1 U5151 ( .A1(n10639), .A2(n11643), .B1(n1880), .B2(n11649), .ZN(
        n7021) );
  OAI22_X1 U5152 ( .A1(n10632), .A2(n11643), .B1(n1868), .B2(n11649), .ZN(
        n7020) );
  OAI22_X1 U5153 ( .A1(n10849), .A2(n11633), .B1(n801), .B2(n11634), .ZN(n7019) );
  OAI22_X1 U5154 ( .A1(n10842), .A2(n11633), .B1(n800), .B2(n11634), .ZN(n7018) );
  OAI22_X1 U5155 ( .A1(n10835), .A2(n11633), .B1(n799), .B2(n11634), .ZN(n7017) );
  OAI22_X1 U5156 ( .A1(n10828), .A2(n11633), .B1(n798), .B2(n11634), .ZN(n7016) );
  OAI22_X1 U5157 ( .A1(n10821), .A2(n11633), .B1(n797), .B2(n11635), .ZN(n7015) );
  OAI22_X1 U5158 ( .A1(n10814), .A2(n11633), .B1(n796), .B2(n11635), .ZN(n7014) );
  OAI22_X1 U5159 ( .A1(n10807), .A2(n11633), .B1(n795), .B2(n11635), .ZN(n7013) );
  OAI22_X1 U5160 ( .A1(n10800), .A2(n11633), .B1(n794), .B2(n11635), .ZN(n7012) );
  OAI22_X1 U5161 ( .A1(n10793), .A2(n11632), .B1(n793), .B2(n11636), .ZN(n7011) );
  OAI22_X1 U5162 ( .A1(n10786), .A2(n11632), .B1(n792), .B2(n11636), .ZN(n7010) );
  OAI22_X1 U5163 ( .A1(n10779), .A2(n11632), .B1(n791), .B2(n11636), .ZN(n7009) );
  OAI22_X1 U5164 ( .A1(n10772), .A2(n11632), .B1(n790), .B2(n11636), .ZN(n7008) );
  OAI22_X1 U5165 ( .A1(n10765), .A2(n11632), .B1(n789), .B2(n11637), .ZN(n7007) );
  OAI22_X1 U5166 ( .A1(n10758), .A2(n11632), .B1(n788), .B2(n11637), .ZN(n7006) );
  OAI22_X1 U5167 ( .A1(n10751), .A2(n11632), .B1(n787), .B2(n11637), .ZN(n7005) );
  OAI22_X1 U5168 ( .A1(n10744), .A2(n11632), .B1(n786), .B2(n11637), .ZN(n7004) );
  OAI22_X1 U5169 ( .A1(n10737), .A2(n11632), .B1(n785), .B2(n11638), .ZN(n7003) );
  OAI22_X1 U5170 ( .A1(n10730), .A2(n11632), .B1(n784), .B2(n11638), .ZN(n7002) );
  OAI22_X1 U5171 ( .A1(n10723), .A2(n11632), .B1(n783), .B2(n11638), .ZN(n7001) );
  OAI22_X1 U5172 ( .A1(n10716), .A2(n11632), .B1(n782), .B2(n11638), .ZN(n7000) );
  OAI22_X1 U5173 ( .A1(n10709), .A2(n11631), .B1(n781), .B2(n11639), .ZN(n6999) );
  OAI22_X1 U5174 ( .A1(n10702), .A2(n11631), .B1(n780), .B2(n11639), .ZN(n6998) );
  OAI22_X1 U5175 ( .A1(n10695), .A2(n11631), .B1(n779), .B2(n11639), .ZN(n6997) );
  OAI22_X1 U5176 ( .A1(n10688), .A2(n11631), .B1(n778), .B2(n11639), .ZN(n6996) );
  OAI22_X1 U5177 ( .A1(n10681), .A2(n11631), .B1(n777), .B2(n11640), .ZN(n6995) );
  OAI22_X1 U5178 ( .A1(n10674), .A2(n11631), .B1(n776), .B2(n11640), .ZN(n6994) );
  OAI22_X1 U5179 ( .A1(n10667), .A2(n11631), .B1(n775), .B2(n11640), .ZN(n6993) );
  OAI22_X1 U5180 ( .A1(n10660), .A2(n11631), .B1(n774), .B2(n11640), .ZN(n6992) );
  OAI22_X1 U5181 ( .A1(n10653), .A2(n11631), .B1(n773), .B2(n11641), .ZN(n6991) );
  OAI22_X1 U5182 ( .A1(n10646), .A2(n11631), .B1(n772), .B2(n11641), .ZN(n6990) );
  OAI22_X1 U5183 ( .A1(n10639), .A2(n11631), .B1(n771), .B2(n11641), .ZN(n6989) );
  OAI22_X1 U5184 ( .A1(n10632), .A2(n11631), .B1(n770), .B2(n11641), .ZN(n6988) );
  OAI22_X1 U5185 ( .A1(n10849), .A2(n11621), .B1(n10537), .B2(n11622), .ZN(
        n6987) );
  OAI22_X1 U5186 ( .A1(n10842), .A2(n11621), .B1(n10505), .B2(n11622), .ZN(
        n6986) );
  OAI22_X1 U5187 ( .A1(n10835), .A2(n11621), .B1(n10473), .B2(n11622), .ZN(
        n6985) );
  OAI22_X1 U5188 ( .A1(n10828), .A2(n11621), .B1(n10441), .B2(n11622), .ZN(
        n6984) );
  OAI22_X1 U5189 ( .A1(n10821), .A2(n11621), .B1(n10409), .B2(n11623), .ZN(
        n6983) );
  OAI22_X1 U5190 ( .A1(n10814), .A2(n11621), .B1(n10374), .B2(n11623), .ZN(
        n6982) );
  OAI22_X1 U5191 ( .A1(n10807), .A2(n11621), .B1(n10342), .B2(n11623), .ZN(
        n6981) );
  OAI22_X1 U5192 ( .A1(n10800), .A2(n11621), .B1(n10310), .B2(n11623), .ZN(
        n6980) );
  OAI22_X1 U5193 ( .A1(n10793), .A2(n11620), .B1(n10275), .B2(n11624), .ZN(
        n6979) );
  OAI22_X1 U5194 ( .A1(n10786), .A2(n11620), .B1(n10243), .B2(n11624), .ZN(
        n6978) );
  OAI22_X1 U5195 ( .A1(n10779), .A2(n11620), .B1(n10211), .B2(n11624), .ZN(
        n6977) );
  OAI22_X1 U5196 ( .A1(n10772), .A2(n11620), .B1(n10177), .B2(n11624), .ZN(
        n6976) );
  OAI22_X1 U5197 ( .A1(n10765), .A2(n11620), .B1(n10145), .B2(n11625), .ZN(
        n6975) );
  OAI22_X1 U5198 ( .A1(n10758), .A2(n11620), .B1(n10113), .B2(n11625), .ZN(
        n6974) );
  OAI22_X1 U5199 ( .A1(n10751), .A2(n11620), .B1(n10081), .B2(n11625), .ZN(
        n6973) );
  OAI22_X1 U5200 ( .A1(n10744), .A2(n11620), .B1(n10049), .B2(n11625), .ZN(
        n6972) );
  OAI22_X1 U5201 ( .A1(n10737), .A2(n11620), .B1(n10017), .B2(n11626), .ZN(
        n6971) );
  OAI22_X1 U5202 ( .A1(n10730), .A2(n11620), .B1(n9655), .B2(n11626), .ZN(
        n6970) );
  OAI22_X1 U5203 ( .A1(n10723), .A2(n11620), .B1(n9623), .B2(n11626), .ZN(
        n6969) );
  OAI22_X1 U5204 ( .A1(n10716), .A2(n11620), .B1(n9591), .B2(n11626), .ZN(
        n6968) );
  OAI22_X1 U5205 ( .A1(n10709), .A2(n11619), .B1(n9257), .B2(n11627), .ZN(
        n6967) );
  OAI22_X1 U5206 ( .A1(n10702), .A2(n11619), .B1(n9193), .B2(n11627), .ZN(
        n6966) );
  OAI22_X1 U5207 ( .A1(n10695), .A2(n11619), .B1(n9161), .B2(n11627), .ZN(
        n6965) );
  OAI22_X1 U5208 ( .A1(n10688), .A2(n11619), .B1(n6311), .B2(n11627), .ZN(
        n6964) );
  OAI22_X1 U5209 ( .A1(n10681), .A2(n11619), .B1(n5994), .B2(n11628), .ZN(
        n6963) );
  OAI22_X1 U5210 ( .A1(n10674), .A2(n11619), .B1(n5930), .B2(n11628), .ZN(
        n6962) );
  OAI22_X1 U5211 ( .A1(n10667), .A2(n11619), .B1(n5898), .B2(n11628), .ZN(
        n6961) );
  OAI22_X1 U5212 ( .A1(n10660), .A2(n11619), .B1(n5866), .B2(n11628), .ZN(
        n6960) );
  OAI22_X1 U5213 ( .A1(n10653), .A2(n11619), .B1(n5834), .B2(n11629), .ZN(
        n6959) );
  OAI22_X1 U5214 ( .A1(n10646), .A2(n11619), .B1(n5802), .B2(n11629), .ZN(
        n6958) );
  OAI22_X1 U5215 ( .A1(n10639), .A2(n11619), .B1(n5770), .B2(n11629), .ZN(
        n6957) );
  OAI22_X1 U5216 ( .A1(n10632), .A2(n11619), .B1(n5738), .B2(n11629), .ZN(
        n6956) );
  OAI22_X1 U5217 ( .A1(n10849), .A2(n11609), .B1(n737), .B2(n11610), .ZN(n6955) );
  OAI22_X1 U5218 ( .A1(n10842), .A2(n11609), .B1(n736), .B2(n11610), .ZN(n6954) );
  OAI22_X1 U5219 ( .A1(n10835), .A2(n11609), .B1(n735), .B2(n11610), .ZN(n6953) );
  OAI22_X1 U5220 ( .A1(n10828), .A2(n11609), .B1(n734), .B2(n11610), .ZN(n6952) );
  OAI22_X1 U5221 ( .A1(n10821), .A2(n11609), .B1(n733), .B2(n11611), .ZN(n6951) );
  OAI22_X1 U5222 ( .A1(n10814), .A2(n11609), .B1(n732), .B2(n11611), .ZN(n6950) );
  OAI22_X1 U5223 ( .A1(n10807), .A2(n11609), .B1(n731), .B2(n11611), .ZN(n6949) );
  OAI22_X1 U5224 ( .A1(n10800), .A2(n11609), .B1(n730), .B2(n11611), .ZN(n6948) );
  OAI22_X1 U5225 ( .A1(n10793), .A2(n11608), .B1(n729), .B2(n11612), .ZN(n6947) );
  OAI22_X1 U5226 ( .A1(n10786), .A2(n11608), .B1(n728), .B2(n11612), .ZN(n6946) );
  OAI22_X1 U5227 ( .A1(n10779), .A2(n11608), .B1(n727), .B2(n11612), .ZN(n6945) );
  OAI22_X1 U5228 ( .A1(n10772), .A2(n11608), .B1(n726), .B2(n11612), .ZN(n6944) );
  OAI22_X1 U5229 ( .A1(n10765), .A2(n11608), .B1(n725), .B2(n11613), .ZN(n6943) );
  OAI22_X1 U5230 ( .A1(n10758), .A2(n11608), .B1(n724), .B2(n11613), .ZN(n6942) );
  OAI22_X1 U5231 ( .A1(n10751), .A2(n11608), .B1(n723), .B2(n11613), .ZN(n6941) );
  OAI22_X1 U5232 ( .A1(n10744), .A2(n11608), .B1(n722), .B2(n11613), .ZN(n6940) );
  OAI22_X1 U5233 ( .A1(n10737), .A2(n11608), .B1(n721), .B2(n11614), .ZN(n6939) );
  OAI22_X1 U5234 ( .A1(n10730), .A2(n11608), .B1(n720), .B2(n11614), .ZN(n6938) );
  OAI22_X1 U5235 ( .A1(n10723), .A2(n11608), .B1(n719), .B2(n11614), .ZN(n6937) );
  OAI22_X1 U5236 ( .A1(n10716), .A2(n11608), .B1(n718), .B2(n11614), .ZN(n6936) );
  OAI22_X1 U5237 ( .A1(n10709), .A2(n11607), .B1(n717), .B2(n11615), .ZN(n6935) );
  OAI22_X1 U5238 ( .A1(n10702), .A2(n11607), .B1(n716), .B2(n11615), .ZN(n6934) );
  OAI22_X1 U5239 ( .A1(n10695), .A2(n11607), .B1(n715), .B2(n11615), .ZN(n6933) );
  OAI22_X1 U5240 ( .A1(n10688), .A2(n11607), .B1(n714), .B2(n11615), .ZN(n6932) );
  OAI22_X1 U5241 ( .A1(n10681), .A2(n11607), .B1(n713), .B2(n11616), .ZN(n6931) );
  OAI22_X1 U5242 ( .A1(n10674), .A2(n11607), .B1(n712), .B2(n11616), .ZN(n6930) );
  OAI22_X1 U5243 ( .A1(n10667), .A2(n11607), .B1(n711), .B2(n11616), .ZN(n6929) );
  OAI22_X1 U5244 ( .A1(n10660), .A2(n11607), .B1(n710), .B2(n11616), .ZN(n6928) );
  OAI22_X1 U5245 ( .A1(n10653), .A2(n11607), .B1(n709), .B2(n11617), .ZN(n6927) );
  OAI22_X1 U5246 ( .A1(n10646), .A2(n11607), .B1(n708), .B2(n11617), .ZN(n6926) );
  OAI22_X1 U5247 ( .A1(n10639), .A2(n11607), .B1(n707), .B2(n11617), .ZN(n6925) );
  OAI22_X1 U5248 ( .A1(n10632), .A2(n11607), .B1(n706), .B2(n11617), .ZN(n6924) );
  OAI22_X1 U5249 ( .A1(n10849), .A2(n11597), .B1(n10531), .B2(n11598), .ZN(
        n6923) );
  OAI22_X1 U5250 ( .A1(n10842), .A2(n11597), .B1(n10499), .B2(n11598), .ZN(
        n6922) );
  OAI22_X1 U5251 ( .A1(n10835), .A2(n11597), .B1(n10467), .B2(n11598), .ZN(
        n6921) );
  OAI22_X1 U5252 ( .A1(n10828), .A2(n11597), .B1(n10435), .B2(n11598), .ZN(
        n6920) );
  OAI22_X1 U5253 ( .A1(n10821), .A2(n11597), .B1(n10403), .B2(n11599), .ZN(
        n6919) );
  OAI22_X1 U5254 ( .A1(n10814), .A2(n11597), .B1(n10368), .B2(n11599), .ZN(
        n6918) );
  OAI22_X1 U5255 ( .A1(n10807), .A2(n11597), .B1(n10336), .B2(n11599), .ZN(
        n6917) );
  OAI22_X1 U5256 ( .A1(n10800), .A2(n11597), .B1(n10304), .B2(n11599), .ZN(
        n6916) );
  OAI22_X1 U5257 ( .A1(n10793), .A2(n11596), .B1(n10269), .B2(n11600), .ZN(
        n6915) );
  OAI22_X1 U5258 ( .A1(n10786), .A2(n11596), .B1(n10237), .B2(n11600), .ZN(
        n6914) );
  OAI22_X1 U5259 ( .A1(n10779), .A2(n11596), .B1(n10203), .B2(n11600), .ZN(
        n6913) );
  OAI22_X1 U5260 ( .A1(n10772), .A2(n11596), .B1(n10171), .B2(n11600), .ZN(
        n6912) );
  OAI22_X1 U5261 ( .A1(n10765), .A2(n11596), .B1(n10139), .B2(n11601), .ZN(
        n6911) );
  OAI22_X1 U5262 ( .A1(n10758), .A2(n11596), .B1(n10107), .B2(n11601), .ZN(
        n6910) );
  OAI22_X1 U5263 ( .A1(n10751), .A2(n11596), .B1(n10075), .B2(n11601), .ZN(
        n6909) );
  OAI22_X1 U5264 ( .A1(n10744), .A2(n11596), .B1(n10043), .B2(n11601), .ZN(
        n6908) );
  OAI22_X1 U5265 ( .A1(n10737), .A2(n11596), .B1(n10011), .B2(n11602), .ZN(
        n6907) );
  OAI22_X1 U5266 ( .A1(n10730), .A2(n11596), .B1(n9649), .B2(n11602), .ZN(
        n6906) );
  OAI22_X1 U5267 ( .A1(n10723), .A2(n11596), .B1(n9617), .B2(n11602), .ZN(
        n6905) );
  OAI22_X1 U5268 ( .A1(n10716), .A2(n11596), .B1(n9585), .B2(n11602), .ZN(
        n6904) );
  OAI22_X1 U5269 ( .A1(n10709), .A2(n11595), .B1(n9251), .B2(n11603), .ZN(
        n6903) );
  OAI22_X1 U5270 ( .A1(n10702), .A2(n11595), .B1(n9187), .B2(n11603), .ZN(
        n6902) );
  OAI22_X1 U5271 ( .A1(n10695), .A2(n11595), .B1(n9155), .B2(n11603), .ZN(
        n6901) );
  OAI22_X1 U5272 ( .A1(n10688), .A2(n11595), .B1(n6305), .B2(n11603), .ZN(
        n6900) );
  OAI22_X1 U5273 ( .A1(n10681), .A2(n11595), .B1(n5988), .B2(n11604), .ZN(
        n6899) );
  OAI22_X1 U5274 ( .A1(n10674), .A2(n11595), .B1(n5924), .B2(n11604), .ZN(
        n6898) );
  OAI22_X1 U5275 ( .A1(n10667), .A2(n11595), .B1(n5892), .B2(n11604), .ZN(
        n6897) );
  OAI22_X1 U5276 ( .A1(n10660), .A2(n11595), .B1(n5860), .B2(n11604), .ZN(
        n6896) );
  OAI22_X1 U5277 ( .A1(n10653), .A2(n11595), .B1(n5828), .B2(n11605), .ZN(
        n6895) );
  OAI22_X1 U5278 ( .A1(n10646), .A2(n11595), .B1(n5796), .B2(n11605), .ZN(
        n6894) );
  OAI22_X1 U5279 ( .A1(n10639), .A2(n11595), .B1(n5764), .B2(n11605), .ZN(
        n6893) );
  OAI22_X1 U5280 ( .A1(n10632), .A2(n11595), .B1(n5732), .B2(n11605), .ZN(
        n6892) );
  OAI22_X1 U5281 ( .A1(n10849), .A2(n11585), .B1(n673), .B2(n11586), .ZN(n6891) );
  OAI22_X1 U5282 ( .A1(n10842), .A2(n11585), .B1(n672), .B2(n11586), .ZN(n6890) );
  OAI22_X1 U5283 ( .A1(n10835), .A2(n11585), .B1(n671), .B2(n11586), .ZN(n6889) );
  OAI22_X1 U5284 ( .A1(n10828), .A2(n11585), .B1(n670), .B2(n11586), .ZN(n6888) );
  OAI22_X1 U5285 ( .A1(n10821), .A2(n11585), .B1(n669), .B2(n11587), .ZN(n6887) );
  OAI22_X1 U5286 ( .A1(n10814), .A2(n11585), .B1(n668), .B2(n11587), .ZN(n6886) );
  OAI22_X1 U5287 ( .A1(n10807), .A2(n11585), .B1(n667), .B2(n11587), .ZN(n6885) );
  OAI22_X1 U5288 ( .A1(n10800), .A2(n11585), .B1(n666), .B2(n11587), .ZN(n6884) );
  OAI22_X1 U5289 ( .A1(n10793), .A2(n11584), .B1(n665), .B2(n11588), .ZN(n6883) );
  OAI22_X1 U5290 ( .A1(n10786), .A2(n11584), .B1(n664), .B2(n11588), .ZN(n6882) );
  OAI22_X1 U5291 ( .A1(n10779), .A2(n11584), .B1(n663), .B2(n11588), .ZN(n6881) );
  OAI22_X1 U5292 ( .A1(n10772), .A2(n11584), .B1(n662), .B2(n11588), .ZN(n6880) );
  OAI22_X1 U5293 ( .A1(n10765), .A2(n11584), .B1(n661), .B2(n11589), .ZN(n6879) );
  OAI22_X1 U5294 ( .A1(n10758), .A2(n11584), .B1(n660), .B2(n11589), .ZN(n6878) );
  OAI22_X1 U5295 ( .A1(n10751), .A2(n11584), .B1(n659), .B2(n11589), .ZN(n6877) );
  OAI22_X1 U5296 ( .A1(n10744), .A2(n11584), .B1(n658), .B2(n11589), .ZN(n6876) );
  OAI22_X1 U5297 ( .A1(n10737), .A2(n11584), .B1(n657), .B2(n11590), .ZN(n6875) );
  OAI22_X1 U5298 ( .A1(n10730), .A2(n11584), .B1(n656), .B2(n11590), .ZN(n6874) );
  OAI22_X1 U5299 ( .A1(n10723), .A2(n11584), .B1(n655), .B2(n11590), .ZN(n6873) );
  OAI22_X1 U5300 ( .A1(n10716), .A2(n11584), .B1(n654), .B2(n11590), .ZN(n6872) );
  OAI22_X1 U5301 ( .A1(n10709), .A2(n11583), .B1(n653), .B2(n11591), .ZN(n6871) );
  OAI22_X1 U5302 ( .A1(n10702), .A2(n11583), .B1(n652), .B2(n11591), .ZN(n6870) );
  OAI22_X1 U5303 ( .A1(n10695), .A2(n11583), .B1(n651), .B2(n11591), .ZN(n6869) );
  OAI22_X1 U5304 ( .A1(n10688), .A2(n11583), .B1(n650), .B2(n11591), .ZN(n6868) );
  OAI22_X1 U5305 ( .A1(n10681), .A2(n11583), .B1(n649), .B2(n11592), .ZN(n6867) );
  OAI22_X1 U5306 ( .A1(n10674), .A2(n11583), .B1(n648), .B2(n11592), .ZN(n6866) );
  OAI22_X1 U5307 ( .A1(n10667), .A2(n11583), .B1(n647), .B2(n11592), .ZN(n6865) );
  OAI22_X1 U5308 ( .A1(n10660), .A2(n11583), .B1(n646), .B2(n11592), .ZN(n6864) );
  OAI22_X1 U5309 ( .A1(n10653), .A2(n11583), .B1(n645), .B2(n11593), .ZN(n6863) );
  OAI22_X1 U5310 ( .A1(n10646), .A2(n11583), .B1(n644), .B2(n11593), .ZN(n6862) );
  OAI22_X1 U5311 ( .A1(n10639), .A2(n11583), .B1(n643), .B2(n11593), .ZN(n6861) );
  OAI22_X1 U5312 ( .A1(n10632), .A2(n11583), .B1(n642), .B2(n11593), .ZN(n6860) );
  OAI22_X1 U5313 ( .A1(n10849), .A2(n11573), .B1(n10530), .B2(n11574), .ZN(
        n6859) );
  OAI22_X1 U5314 ( .A1(n10842), .A2(n11573), .B1(n10498), .B2(n11574), .ZN(
        n6858) );
  OAI22_X1 U5315 ( .A1(n10835), .A2(n11573), .B1(n10466), .B2(n11574), .ZN(
        n6857) );
  OAI22_X1 U5316 ( .A1(n10828), .A2(n11573), .B1(n10434), .B2(n11574), .ZN(
        n6856) );
  OAI22_X1 U5317 ( .A1(n10821), .A2(n11573), .B1(n10402), .B2(n11575), .ZN(
        n6855) );
  OAI22_X1 U5318 ( .A1(n10814), .A2(n11573), .B1(n10367), .B2(n11575), .ZN(
        n6854) );
  OAI22_X1 U5319 ( .A1(n10807), .A2(n11573), .B1(n10335), .B2(n11575), .ZN(
        n6853) );
  OAI22_X1 U5320 ( .A1(n10800), .A2(n11573), .B1(n10300), .B2(n11575), .ZN(
        n6852) );
  OAI22_X1 U5321 ( .A1(n10793), .A2(n11572), .B1(n10268), .B2(n11576), .ZN(
        n6851) );
  OAI22_X1 U5322 ( .A1(n10786), .A2(n11572), .B1(n10236), .B2(n11576), .ZN(
        n6850) );
  OAI22_X1 U5323 ( .A1(n10779), .A2(n11572), .B1(n10202), .B2(n11576), .ZN(
        n6849) );
  OAI22_X1 U5324 ( .A1(n10772), .A2(n11572), .B1(n10170), .B2(n11576), .ZN(
        n6848) );
  OAI22_X1 U5325 ( .A1(n10765), .A2(n11572), .B1(n10138), .B2(n11577), .ZN(
        n6847) );
  OAI22_X1 U5326 ( .A1(n10758), .A2(n11572), .B1(n10106), .B2(n11577), .ZN(
        n6846) );
  OAI22_X1 U5327 ( .A1(n10751), .A2(n11572), .B1(n10074), .B2(n11577), .ZN(
        n6845) );
  OAI22_X1 U5328 ( .A1(n10744), .A2(n11572), .B1(n10042), .B2(n11577), .ZN(
        n6844) );
  OAI22_X1 U5329 ( .A1(n10737), .A2(n11572), .B1(n10010), .B2(n11578), .ZN(
        n6843) );
  OAI22_X1 U5330 ( .A1(n10730), .A2(n11572), .B1(n9648), .B2(n11578), .ZN(
        n6842) );
  OAI22_X1 U5331 ( .A1(n10723), .A2(n11572), .B1(n9616), .B2(n11578), .ZN(
        n6841) );
  OAI22_X1 U5332 ( .A1(n10716), .A2(n11572), .B1(n9584), .B2(n11578), .ZN(
        n6840) );
  OAI22_X1 U5333 ( .A1(n10709), .A2(n11571), .B1(n9250), .B2(n11579), .ZN(
        n6839) );
  OAI22_X1 U5334 ( .A1(n10702), .A2(n11571), .B1(n9186), .B2(n11579), .ZN(
        n6838) );
  OAI22_X1 U5335 ( .A1(n10695), .A2(n11571), .B1(n9154), .B2(n11579), .ZN(
        n6837) );
  OAI22_X1 U5336 ( .A1(n10688), .A2(n11571), .B1(n6304), .B2(n11579), .ZN(
        n6836) );
  OAI22_X1 U5337 ( .A1(n10681), .A2(n11571), .B1(n5987), .B2(n11580), .ZN(
        n6835) );
  OAI22_X1 U5338 ( .A1(n10674), .A2(n11571), .B1(n5923), .B2(n11580), .ZN(
        n6834) );
  OAI22_X1 U5339 ( .A1(n10667), .A2(n11571), .B1(n5891), .B2(n11580), .ZN(
        n6833) );
  OAI22_X1 U5340 ( .A1(n10660), .A2(n11571), .B1(n5859), .B2(n11580), .ZN(
        n6832) );
  OAI22_X1 U5341 ( .A1(n10653), .A2(n11571), .B1(n5827), .B2(n11581), .ZN(
        n6831) );
  OAI22_X1 U5342 ( .A1(n10646), .A2(n11571), .B1(n5795), .B2(n11581), .ZN(
        n6830) );
  OAI22_X1 U5343 ( .A1(n10639), .A2(n11571), .B1(n5763), .B2(n11581), .ZN(
        n6829) );
  OAI22_X1 U5344 ( .A1(n10632), .A2(n11571), .B1(n5731), .B2(n11581), .ZN(
        n6828) );
  OAI22_X1 U5345 ( .A1(n10849), .A2(n11561), .B1(n10532), .B2(n11562), .ZN(
        n6827) );
  OAI22_X1 U5346 ( .A1(n10842), .A2(n11561), .B1(n10500), .B2(n11562), .ZN(
        n6826) );
  OAI22_X1 U5347 ( .A1(n10835), .A2(n11561), .B1(n10468), .B2(n11562), .ZN(
        n6825) );
  OAI22_X1 U5348 ( .A1(n10828), .A2(n11561), .B1(n10436), .B2(n11562), .ZN(
        n6824) );
  OAI22_X1 U5349 ( .A1(n10821), .A2(n11561), .B1(n10404), .B2(n11563), .ZN(
        n6823) );
  OAI22_X1 U5350 ( .A1(n10814), .A2(n11561), .B1(n10369), .B2(n11563), .ZN(
        n6822) );
  OAI22_X1 U5351 ( .A1(n10807), .A2(n11561), .B1(n10337), .B2(n11563), .ZN(
        n6821) );
  OAI22_X1 U5352 ( .A1(n10800), .A2(n11561), .B1(n10305), .B2(n11563), .ZN(
        n6820) );
  OAI22_X1 U5353 ( .A1(n10793), .A2(n11560), .B1(n10270), .B2(n11564), .ZN(
        n6819) );
  OAI22_X1 U5354 ( .A1(n10786), .A2(n11560), .B1(n10238), .B2(n11564), .ZN(
        n6818) );
  OAI22_X1 U5355 ( .A1(n10779), .A2(n11560), .B1(n10204), .B2(n11564), .ZN(
        n6817) );
  OAI22_X1 U5356 ( .A1(n10772), .A2(n11560), .B1(n10172), .B2(n11564), .ZN(
        n6816) );
  OAI22_X1 U5357 ( .A1(n10765), .A2(n11560), .B1(n10140), .B2(n11565), .ZN(
        n6815) );
  OAI22_X1 U5358 ( .A1(n10758), .A2(n11560), .B1(n10108), .B2(n11565), .ZN(
        n6814) );
  OAI22_X1 U5359 ( .A1(n10751), .A2(n11560), .B1(n10076), .B2(n11565), .ZN(
        n6813) );
  OAI22_X1 U5360 ( .A1(n10744), .A2(n11560), .B1(n10044), .B2(n11565), .ZN(
        n6812) );
  OAI22_X1 U5361 ( .A1(n10737), .A2(n11560), .B1(n10012), .B2(n11566), .ZN(
        n6811) );
  OAI22_X1 U5362 ( .A1(n10730), .A2(n11560), .B1(n9650), .B2(n11566), .ZN(
        n6810) );
  OAI22_X1 U5363 ( .A1(n10723), .A2(n11560), .B1(n9618), .B2(n11566), .ZN(
        n6809) );
  OAI22_X1 U5364 ( .A1(n10716), .A2(n11560), .B1(n9586), .B2(n11566), .ZN(
        n6808) );
  OAI22_X1 U5365 ( .A1(n10709), .A2(n11559), .B1(n9252), .B2(n11567), .ZN(
        n6807) );
  OAI22_X1 U5366 ( .A1(n10702), .A2(n11559), .B1(n9188), .B2(n11567), .ZN(
        n6806) );
  OAI22_X1 U5367 ( .A1(n10695), .A2(n11559), .B1(n9156), .B2(n11567), .ZN(
        n6805) );
  OAI22_X1 U5368 ( .A1(n10688), .A2(n11559), .B1(n6306), .B2(n11567), .ZN(
        n6804) );
  OAI22_X1 U5369 ( .A1(n10681), .A2(n11559), .B1(n5989), .B2(n11568), .ZN(
        n6803) );
  OAI22_X1 U5370 ( .A1(n10674), .A2(n11559), .B1(n5925), .B2(n11568), .ZN(
        n6802) );
  OAI22_X1 U5371 ( .A1(n10667), .A2(n11559), .B1(n5893), .B2(n11568), .ZN(
        n6801) );
  OAI22_X1 U5372 ( .A1(n10660), .A2(n11559), .B1(n5861), .B2(n11568), .ZN(
        n6800) );
  OAI22_X1 U5373 ( .A1(n10653), .A2(n11559), .B1(n5829), .B2(n11569), .ZN(
        n6799) );
  OAI22_X1 U5374 ( .A1(n10646), .A2(n11559), .B1(n5797), .B2(n11569), .ZN(
        n6798) );
  OAI22_X1 U5375 ( .A1(n10639), .A2(n11559), .B1(n5765), .B2(n11569), .ZN(
        n6797) );
  OAI22_X1 U5376 ( .A1(n10632), .A2(n11559), .B1(n5733), .B2(n11569), .ZN(
        n6796) );
  OAI22_X1 U5377 ( .A1(n10849), .A2(n11513), .B1(n10536), .B2(n11514), .ZN(
        n6699) );
  OAI22_X1 U5378 ( .A1(n10842), .A2(n11513), .B1(n10504), .B2(n11514), .ZN(
        n6698) );
  OAI22_X1 U5379 ( .A1(n10835), .A2(n11513), .B1(n10472), .B2(n11514), .ZN(
        n6697) );
  OAI22_X1 U5380 ( .A1(n10828), .A2(n11513), .B1(n10440), .B2(n11514), .ZN(
        n6696) );
  OAI22_X1 U5381 ( .A1(n10821), .A2(n11513), .B1(n10408), .B2(n11515), .ZN(
        n6695) );
  OAI22_X1 U5382 ( .A1(n10814), .A2(n11513), .B1(n10373), .B2(n11515), .ZN(
        n6694) );
  OAI22_X1 U5383 ( .A1(n10807), .A2(n11513), .B1(n10341), .B2(n11515), .ZN(
        n6693) );
  OAI22_X1 U5384 ( .A1(n10800), .A2(n11513), .B1(n10309), .B2(n11515), .ZN(
        n6692) );
  OAI22_X1 U5385 ( .A1(n10793), .A2(n11512), .B1(n10274), .B2(n11516), .ZN(
        n6691) );
  OAI22_X1 U5386 ( .A1(n10786), .A2(n11512), .B1(n10242), .B2(n11516), .ZN(
        n6690) );
  OAI22_X1 U5387 ( .A1(n10779), .A2(n11512), .B1(n10210), .B2(n11516), .ZN(
        n6689) );
  OAI22_X1 U5388 ( .A1(n10772), .A2(n11512), .B1(n10176), .B2(n11516), .ZN(
        n6688) );
  OAI22_X1 U5389 ( .A1(n10765), .A2(n11512), .B1(n10144), .B2(n11517), .ZN(
        n6687) );
  OAI22_X1 U5390 ( .A1(n10758), .A2(n11512), .B1(n10112), .B2(n11517), .ZN(
        n6686) );
  OAI22_X1 U5391 ( .A1(n10751), .A2(n11512), .B1(n10080), .B2(n11517), .ZN(
        n6685) );
  OAI22_X1 U5392 ( .A1(n10744), .A2(n11512), .B1(n10048), .B2(n11517), .ZN(
        n6684) );
  OAI22_X1 U5393 ( .A1(n10737), .A2(n11512), .B1(n10016), .B2(n11518), .ZN(
        n6683) );
  OAI22_X1 U5394 ( .A1(n10730), .A2(n11512), .B1(n9654), .B2(n11518), .ZN(
        n6682) );
  OAI22_X1 U5395 ( .A1(n10723), .A2(n11512), .B1(n9622), .B2(n11518), .ZN(
        n6681) );
  OAI22_X1 U5396 ( .A1(n10716), .A2(n11512), .B1(n9590), .B2(n11518), .ZN(
        n6680) );
  OAI22_X1 U5397 ( .A1(n10709), .A2(n11511), .B1(n9256), .B2(n11519), .ZN(
        n6679) );
  OAI22_X1 U5398 ( .A1(n10702), .A2(n11511), .B1(n9192), .B2(n11519), .ZN(
        n6678) );
  OAI22_X1 U5399 ( .A1(n10695), .A2(n11511), .B1(n9160), .B2(n11519), .ZN(
        n6677) );
  OAI22_X1 U5400 ( .A1(n10688), .A2(n11511), .B1(n6310), .B2(n11519), .ZN(
        n6676) );
  OAI22_X1 U5401 ( .A1(n10681), .A2(n11511), .B1(n5993), .B2(n11520), .ZN(
        n6675) );
  OAI22_X1 U5402 ( .A1(n10674), .A2(n11511), .B1(n5929), .B2(n11520), .ZN(
        n6674) );
  OAI22_X1 U5403 ( .A1(n10667), .A2(n11511), .B1(n5897), .B2(n11520), .ZN(
        n6673) );
  OAI22_X1 U5404 ( .A1(n10660), .A2(n11511), .B1(n5865), .B2(n11520), .ZN(
        n6672) );
  OAI22_X1 U5405 ( .A1(n10653), .A2(n11511), .B1(n5833), .B2(n11521), .ZN(
        n6671) );
  OAI22_X1 U5406 ( .A1(n10646), .A2(n11511), .B1(n5801), .B2(n11521), .ZN(
        n6670) );
  OAI22_X1 U5407 ( .A1(n10639), .A2(n11511), .B1(n5769), .B2(n11521), .ZN(
        n6669) );
  OAI22_X1 U5408 ( .A1(n10632), .A2(n11511), .B1(n5737), .B2(n11521), .ZN(
        n6668) );
  OAI22_X1 U5409 ( .A1(n10846), .A2(n12029), .B1(n12030), .B2(n13843), .ZN(
        n8075) );
  OAI22_X1 U5410 ( .A1(n10839), .A2(n12029), .B1(n12030), .B2(n13842), .ZN(
        n8074) );
  OAI22_X1 U5411 ( .A1(n10832), .A2(n12029), .B1(n12030), .B2(n13841), .ZN(
        n8073) );
  OAI22_X1 U5412 ( .A1(n10825), .A2(n12029), .B1(n12030), .B2(n13840), .ZN(
        n8072) );
  OAI22_X1 U5413 ( .A1(n10818), .A2(n12029), .B1(n12031), .B2(n13839), .ZN(
        n8071) );
  OAI22_X1 U5414 ( .A1(n10811), .A2(n12029), .B1(n12031), .B2(n13838), .ZN(
        n8070) );
  OAI22_X1 U5415 ( .A1(n10804), .A2(n12029), .B1(n12031), .B2(n13837), .ZN(
        n8069) );
  OAI22_X1 U5416 ( .A1(n10797), .A2(n12029), .B1(n12031), .B2(n13836), .ZN(
        n8068) );
  OAI22_X1 U5417 ( .A1(n10790), .A2(n12028), .B1(n12032), .B2(n13835), .ZN(
        n8067) );
  OAI22_X1 U5418 ( .A1(n10783), .A2(n12028), .B1(n12032), .B2(n13834), .ZN(
        n8066) );
  OAI22_X1 U5419 ( .A1(n10776), .A2(n12028), .B1(n12032), .B2(n13833), .ZN(
        n8065) );
  OAI22_X1 U5420 ( .A1(n10769), .A2(n12028), .B1(n12032), .B2(n13832), .ZN(
        n8064) );
  OAI22_X1 U5421 ( .A1(n10762), .A2(n12028), .B1(n12033), .B2(n13831), .ZN(
        n8063) );
  OAI22_X1 U5422 ( .A1(n10755), .A2(n12028), .B1(n12033), .B2(n13830), .ZN(
        n8062) );
  OAI22_X1 U5423 ( .A1(n10748), .A2(n12028), .B1(n12033), .B2(n13829), .ZN(
        n8061) );
  OAI22_X1 U5424 ( .A1(n10741), .A2(n12028), .B1(n12033), .B2(n13828), .ZN(
        n8060) );
  OAI22_X1 U5425 ( .A1(n10734), .A2(n12028), .B1(n12034), .B2(n13827), .ZN(
        n8059) );
  OAI22_X1 U5426 ( .A1(n10727), .A2(n12028), .B1(n12034), .B2(n13826), .ZN(
        n8058) );
  OAI22_X1 U5427 ( .A1(n10720), .A2(n12028), .B1(n12034), .B2(n13825), .ZN(
        n8057) );
  OAI22_X1 U5428 ( .A1(n10713), .A2(n12028), .B1(n12034), .B2(n13824), .ZN(
        n8056) );
  OAI22_X1 U5429 ( .A1(n10706), .A2(n12027), .B1(n12035), .B2(n13823), .ZN(
        n8055) );
  OAI22_X1 U5430 ( .A1(n10699), .A2(n12027), .B1(n12035), .B2(n13822), .ZN(
        n8054) );
  OAI22_X1 U5431 ( .A1(n10692), .A2(n12027), .B1(n12035), .B2(n13821), .ZN(
        n8053) );
  OAI22_X1 U5432 ( .A1(n10685), .A2(n12027), .B1(n12035), .B2(n13820), .ZN(
        n8052) );
  OAI22_X1 U5433 ( .A1(n10678), .A2(n12027), .B1(n12036), .B2(n13819), .ZN(
        n8051) );
  OAI22_X1 U5434 ( .A1(n10671), .A2(n12027), .B1(n12036), .B2(n13818), .ZN(
        n8050) );
  OAI22_X1 U5435 ( .A1(n10664), .A2(n12027), .B1(n12036), .B2(n13817), .ZN(
        n8049) );
  OAI22_X1 U5436 ( .A1(n10657), .A2(n12027), .B1(n12036), .B2(n13816), .ZN(
        n8048) );
  OAI22_X1 U5437 ( .A1(n10650), .A2(n12027), .B1(n12037), .B2(n13815), .ZN(
        n8047) );
  OAI22_X1 U5438 ( .A1(n10643), .A2(n12027), .B1(n12037), .B2(n13814), .ZN(
        n8046) );
  OAI22_X1 U5439 ( .A1(n10636), .A2(n12027), .B1(n12037), .B2(n13813), .ZN(
        n8045) );
  OAI22_X1 U5440 ( .A1(n10629), .A2(n12027), .B1(n12037), .B2(n13812), .ZN(
        n8044) );
  OAI22_X1 U5441 ( .A1(n10727), .A2(n12016), .B1(n12022), .B2(n13794), .ZN(
        n8026) );
  OAI22_X1 U5442 ( .A1(n10720), .A2(n12016), .B1(n12022), .B2(n13793), .ZN(
        n8025) );
  OAI22_X1 U5443 ( .A1(n10713), .A2(n12016), .B1(n12022), .B2(n13792), .ZN(
        n8024) );
  OAI22_X1 U5444 ( .A1(n10706), .A2(n12015), .B1(n12023), .B2(n13791), .ZN(
        n8023) );
  OAI22_X1 U5445 ( .A1(n10699), .A2(n12015), .B1(n12023), .B2(n13790), .ZN(
        n8022) );
  OAI22_X1 U5446 ( .A1(n10692), .A2(n12015), .B1(n12023), .B2(n13789), .ZN(
        n8021) );
  OAI22_X1 U5447 ( .A1(n10685), .A2(n12015), .B1(n12023), .B2(n13788), .ZN(
        n8020) );
  OAI22_X1 U5448 ( .A1(n10678), .A2(n12015), .B1(n12024), .B2(n13787), .ZN(
        n8019) );
  OAI22_X1 U5449 ( .A1(n10671), .A2(n12015), .B1(n12024), .B2(n13786), .ZN(
        n8018) );
  OAI22_X1 U5450 ( .A1(n10664), .A2(n12015), .B1(n12024), .B2(n13785), .ZN(
        n8017) );
  OAI22_X1 U5451 ( .A1(n10657), .A2(n12015), .B1(n12024), .B2(n13784), .ZN(
        n8016) );
  OAI22_X1 U5452 ( .A1(n10650), .A2(n12015), .B1(n12025), .B2(n13783), .ZN(
        n8015) );
  OAI22_X1 U5453 ( .A1(n10643), .A2(n12015), .B1(n12025), .B2(n13782), .ZN(
        n8014) );
  OAI22_X1 U5454 ( .A1(n10636), .A2(n12015), .B1(n12025), .B2(n13781), .ZN(
        n8013) );
  OAI22_X1 U5455 ( .A1(n10629), .A2(n12015), .B1(n12025), .B2(n13780), .ZN(
        n8012) );
  OAI22_X1 U5456 ( .A1(n10846), .A2(n12005), .B1(n12010), .B2(n13779), .ZN(
        n8011) );
  OAI22_X1 U5457 ( .A1(n10839), .A2(n12005), .B1(n12006), .B2(n13778), .ZN(
        n8010) );
  OAI22_X1 U5458 ( .A1(n10832), .A2(n12005), .B1(n12006), .B2(n13777), .ZN(
        n8009) );
  OAI22_X1 U5459 ( .A1(n10825), .A2(n12005), .B1(n12006), .B2(n13776), .ZN(
        n8008) );
  OAI22_X1 U5460 ( .A1(n10818), .A2(n12005), .B1(n12007), .B2(n13775), .ZN(
        n8007) );
  OAI22_X1 U5461 ( .A1(n10811), .A2(n12005), .B1(n12007), .B2(n13774), .ZN(
        n8006) );
  OAI22_X1 U5462 ( .A1(n10804), .A2(n12005), .B1(n12007), .B2(n13773), .ZN(
        n8005) );
  OAI22_X1 U5463 ( .A1(n10797), .A2(n12005), .B1(n12007), .B2(n13772), .ZN(
        n8004) );
  OAI22_X1 U5464 ( .A1(n10790), .A2(n12004), .B1(n12008), .B2(n13771), .ZN(
        n8003) );
  OAI22_X1 U5465 ( .A1(n10783), .A2(n12004), .B1(n12008), .B2(n13770), .ZN(
        n8002) );
  OAI22_X1 U5466 ( .A1(n10776), .A2(n12004), .B1(n12008), .B2(n13769), .ZN(
        n8001) );
  OAI22_X1 U5467 ( .A1(n10769), .A2(n12004), .B1(n12008), .B2(n13768), .ZN(
        n8000) );
  OAI22_X1 U5468 ( .A1(n10762), .A2(n12004), .B1(n12009), .B2(n13767), .ZN(
        n7999) );
  OAI22_X1 U5469 ( .A1(n10755), .A2(n12004), .B1(n12009), .B2(n13766), .ZN(
        n7998) );
  OAI22_X1 U5470 ( .A1(n10748), .A2(n12004), .B1(n12009), .B2(n13765), .ZN(
        n7997) );
  OAI22_X1 U5471 ( .A1(n10741), .A2(n12004), .B1(n12009), .B2(n13764), .ZN(
        n7996) );
  OAI22_X1 U5472 ( .A1(n10734), .A2(n12004), .B1(n12010), .B2(n13763), .ZN(
        n7995) );
  OAI22_X1 U5473 ( .A1(n10727), .A2(n12004), .B1(n12010), .B2(n13762), .ZN(
        n7994) );
  OAI22_X1 U5474 ( .A1(n10720), .A2(n12004), .B1(n12010), .B2(n13761), .ZN(
        n7993) );
  OAI22_X1 U5475 ( .A1(n10713), .A2(n12004), .B1(n12011), .B2(n13760), .ZN(
        n7992) );
  OAI22_X1 U5476 ( .A1(n10706), .A2(n12003), .B1(n12011), .B2(n13759), .ZN(
        n7991) );
  OAI22_X1 U5477 ( .A1(n10699), .A2(n12003), .B1(n12011), .B2(n13758), .ZN(
        n7990) );
  OAI22_X1 U5478 ( .A1(n10692), .A2(n12003), .B1(n12011), .B2(n13757), .ZN(
        n7989) );
  OAI22_X1 U5479 ( .A1(n10685), .A2(n12003), .B1(n12012), .B2(n13756), .ZN(
        n7988) );
  OAI22_X1 U5480 ( .A1(n10678), .A2(n12003), .B1(n12012), .B2(n13755), .ZN(
        n7987) );
  OAI22_X1 U5481 ( .A1(n10671), .A2(n12003), .B1(n12012), .B2(n13754), .ZN(
        n7986) );
  OAI22_X1 U5482 ( .A1(n10664), .A2(n12003), .B1(n12012), .B2(n13753), .ZN(
        n7985) );
  OAI22_X1 U5483 ( .A1(n10657), .A2(n12003), .B1(n12013), .B2(n13752), .ZN(
        n7984) );
  OAI22_X1 U5484 ( .A1(n10650), .A2(n12003), .B1(n12013), .B2(n13751), .ZN(
        n7983) );
  OAI22_X1 U5485 ( .A1(n10643), .A2(n12003), .B1(n12013), .B2(n13750), .ZN(
        n7982) );
  OAI22_X1 U5486 ( .A1(n10636), .A2(n12003), .B1(n12013), .B2(n13749), .ZN(
        n7981) );
  OAI22_X1 U5487 ( .A1(n10846), .A2(n11993), .B1(n11994), .B2(n13747), .ZN(
        n7979) );
  OAI22_X1 U5488 ( .A1(n10839), .A2(n11993), .B1(n11994), .B2(n13746), .ZN(
        n7978) );
  OAI22_X1 U5489 ( .A1(n10832), .A2(n11993), .B1(n11994), .B2(n13745), .ZN(
        n7977) );
  OAI22_X1 U5490 ( .A1(n10825), .A2(n11993), .B1(n11994), .B2(n13744), .ZN(
        n7976) );
  OAI22_X1 U5491 ( .A1(n10818), .A2(n11993), .B1(n11995), .B2(n13743), .ZN(
        n7975) );
  OAI22_X1 U5492 ( .A1(n10811), .A2(n11993), .B1(n11995), .B2(n13742), .ZN(
        n7974) );
  OAI22_X1 U5493 ( .A1(n10804), .A2(n11993), .B1(n11995), .B2(n13741), .ZN(
        n7973) );
  OAI22_X1 U5494 ( .A1(n10797), .A2(n11993), .B1(n11995), .B2(n13740), .ZN(
        n7972) );
  OAI22_X1 U5495 ( .A1(n10790), .A2(n11992), .B1(n11996), .B2(n13739), .ZN(
        n7971) );
  OAI22_X1 U5496 ( .A1(n10783), .A2(n11992), .B1(n11996), .B2(n13738), .ZN(
        n7970) );
  OAI22_X1 U5497 ( .A1(n10776), .A2(n11992), .B1(n11996), .B2(n13737), .ZN(
        n7969) );
  OAI22_X1 U5498 ( .A1(n10769), .A2(n11992), .B1(n11996), .B2(n13736), .ZN(
        n7968) );
  OAI22_X1 U5499 ( .A1(n10762), .A2(n11992), .B1(n11997), .B2(n13735), .ZN(
        n7967) );
  OAI22_X1 U5500 ( .A1(n10755), .A2(n11992), .B1(n11997), .B2(n13734), .ZN(
        n7966) );
  OAI22_X1 U5501 ( .A1(n10748), .A2(n11992), .B1(n11997), .B2(n13733), .ZN(
        n7965) );
  OAI22_X1 U5502 ( .A1(n10741), .A2(n11992), .B1(n11997), .B2(n13732), .ZN(
        n7964) );
  OAI22_X1 U5503 ( .A1(n10734), .A2(n11992), .B1(n11998), .B2(n13731), .ZN(
        n7963) );
  OAI22_X1 U5504 ( .A1(n10727), .A2(n11992), .B1(n11998), .B2(n13730), .ZN(
        n7962) );
  OAI22_X1 U5505 ( .A1(n10720), .A2(n11992), .B1(n11998), .B2(n13729), .ZN(
        n7961) );
  OAI22_X1 U5506 ( .A1(n10713), .A2(n11992), .B1(n11998), .B2(n13728), .ZN(
        n7960) );
  OAI22_X1 U5507 ( .A1(n10706), .A2(n11991), .B1(n11999), .B2(n13727), .ZN(
        n7959) );
  OAI22_X1 U5508 ( .A1(n10699), .A2(n11991), .B1(n11999), .B2(n13726), .ZN(
        n7958) );
  OAI22_X1 U5509 ( .A1(n10692), .A2(n11991), .B1(n11999), .B2(n13725), .ZN(
        n7957) );
  OAI22_X1 U5510 ( .A1(n10685), .A2(n11991), .B1(n11999), .B2(n13724), .ZN(
        n7956) );
  OAI22_X1 U5511 ( .A1(n10678), .A2(n11991), .B1(n12000), .B2(n13723), .ZN(
        n7955) );
  OAI22_X1 U5512 ( .A1(n10671), .A2(n11991), .B1(n12000), .B2(n13722), .ZN(
        n7954) );
  OAI22_X1 U5513 ( .A1(n10664), .A2(n11991), .B1(n12000), .B2(n13721), .ZN(
        n7953) );
  OAI22_X1 U5514 ( .A1(n10657), .A2(n11991), .B1(n12000), .B2(n13720), .ZN(
        n7952) );
  OAI22_X1 U5515 ( .A1(n10650), .A2(n11991), .B1(n12001), .B2(n13719), .ZN(
        n7951) );
  OAI22_X1 U5516 ( .A1(n10643), .A2(n11991), .B1(n12001), .B2(n13718), .ZN(
        n7950) );
  OAI22_X1 U5517 ( .A1(n10636), .A2(n11991), .B1(n12001), .B2(n13717), .ZN(
        n7949) );
  OAI22_X1 U5518 ( .A1(n10629), .A2(n11991), .B1(n12001), .B2(n13716), .ZN(
        n7948) );
  OAI22_X1 U5519 ( .A1(n10846), .A2(n11981), .B1(n11982), .B2(n13715), .ZN(
        n7947) );
  OAI22_X1 U5520 ( .A1(n10839), .A2(n11981), .B1(n11982), .B2(n13714), .ZN(
        n7946) );
  OAI22_X1 U5521 ( .A1(n10832), .A2(n11981), .B1(n11982), .B2(n13713), .ZN(
        n7945) );
  OAI22_X1 U5522 ( .A1(n10825), .A2(n11981), .B1(n11982), .B2(n13712), .ZN(
        n7944) );
  OAI22_X1 U5523 ( .A1(n10818), .A2(n11981), .B1(n11983), .B2(n13711), .ZN(
        n7943) );
  OAI22_X1 U5524 ( .A1(n10811), .A2(n11981), .B1(n11983), .B2(n13710), .ZN(
        n7942) );
  OAI22_X1 U5525 ( .A1(n10804), .A2(n11981), .B1(n11983), .B2(n13709), .ZN(
        n7941) );
  OAI22_X1 U5526 ( .A1(n10797), .A2(n11981), .B1(n11983), .B2(n13708), .ZN(
        n7940) );
  OAI22_X1 U5527 ( .A1(n10790), .A2(n11980), .B1(n11984), .B2(n13707), .ZN(
        n7939) );
  OAI22_X1 U5528 ( .A1(n10783), .A2(n11980), .B1(n11984), .B2(n13706), .ZN(
        n7938) );
  OAI22_X1 U5529 ( .A1(n10776), .A2(n11980), .B1(n11984), .B2(n13705), .ZN(
        n7937) );
  OAI22_X1 U5530 ( .A1(n10769), .A2(n11980), .B1(n11984), .B2(n13704), .ZN(
        n7936) );
  OAI22_X1 U5531 ( .A1(n10762), .A2(n11980), .B1(n11985), .B2(n13703), .ZN(
        n7935) );
  OAI22_X1 U5532 ( .A1(n10755), .A2(n11980), .B1(n11985), .B2(n13702), .ZN(
        n7934) );
  OAI22_X1 U5533 ( .A1(n10748), .A2(n11980), .B1(n11985), .B2(n13701), .ZN(
        n7933) );
  OAI22_X1 U5534 ( .A1(n10741), .A2(n11980), .B1(n11985), .B2(n13700), .ZN(
        n7932) );
  OAI22_X1 U5535 ( .A1(n10734), .A2(n11980), .B1(n11986), .B2(n13699), .ZN(
        n7931) );
  OAI22_X1 U5536 ( .A1(n10727), .A2(n11980), .B1(n11986), .B2(n13698), .ZN(
        n7930) );
  OAI22_X1 U5537 ( .A1(n10720), .A2(n11980), .B1(n11986), .B2(n13697), .ZN(
        n7929) );
  OAI22_X1 U5538 ( .A1(n10713), .A2(n11980), .B1(n11986), .B2(n13696), .ZN(
        n7928) );
  OAI22_X1 U5539 ( .A1(n10706), .A2(n11979), .B1(n11987), .B2(n13695), .ZN(
        n7927) );
  OAI22_X1 U5540 ( .A1(n10699), .A2(n11979), .B1(n11987), .B2(n13694), .ZN(
        n7926) );
  OAI22_X1 U5541 ( .A1(n10692), .A2(n11979), .B1(n11987), .B2(n13693), .ZN(
        n7925) );
  OAI22_X1 U5542 ( .A1(n10685), .A2(n11979), .B1(n11987), .B2(n13692), .ZN(
        n7924) );
  OAI22_X1 U5543 ( .A1(n10678), .A2(n11979), .B1(n11988), .B2(n13691), .ZN(
        n7923) );
  OAI22_X1 U5544 ( .A1(n10671), .A2(n11979), .B1(n11988), .B2(n13690), .ZN(
        n7922) );
  OAI22_X1 U5545 ( .A1(n10664), .A2(n11979), .B1(n11988), .B2(n13689), .ZN(
        n7921) );
  OAI22_X1 U5546 ( .A1(n10657), .A2(n11979), .B1(n11988), .B2(n13688), .ZN(
        n7920) );
  OAI22_X1 U5547 ( .A1(n10650), .A2(n11979), .B1(n11989), .B2(n13687), .ZN(
        n7919) );
  OAI22_X1 U5548 ( .A1(n10643), .A2(n11979), .B1(n11989), .B2(n13686), .ZN(
        n7918) );
  OAI22_X1 U5549 ( .A1(n10636), .A2(n11979), .B1(n11989), .B2(n13685), .ZN(
        n7917) );
  OAI22_X1 U5550 ( .A1(n10629), .A2(n11979), .B1(n11989), .B2(n13684), .ZN(
        n7916) );
  OAI22_X1 U5551 ( .A1(n10846), .A2(n11969), .B1(n11970), .B2(n13683), .ZN(
        n7915) );
  OAI22_X1 U5552 ( .A1(n10839), .A2(n11969), .B1(n11970), .B2(n13682), .ZN(
        n7914) );
  OAI22_X1 U5553 ( .A1(n10832), .A2(n11969), .B1(n11970), .B2(n13681), .ZN(
        n7913) );
  OAI22_X1 U5554 ( .A1(n10825), .A2(n11969), .B1(n11970), .B2(n13680), .ZN(
        n7912) );
  OAI22_X1 U5555 ( .A1(n10818), .A2(n11969), .B1(n11971), .B2(n13679), .ZN(
        n7911) );
  OAI22_X1 U5556 ( .A1(n10811), .A2(n11969), .B1(n11971), .B2(n13678), .ZN(
        n7910) );
  OAI22_X1 U5557 ( .A1(n10804), .A2(n11969), .B1(n11971), .B2(n13677), .ZN(
        n7909) );
  OAI22_X1 U5558 ( .A1(n10797), .A2(n11969), .B1(n11971), .B2(n13676), .ZN(
        n7908) );
  OAI22_X1 U5559 ( .A1(n10790), .A2(n11968), .B1(n11972), .B2(n13675), .ZN(
        n7907) );
  OAI22_X1 U5560 ( .A1(n10783), .A2(n11968), .B1(n11972), .B2(n13674), .ZN(
        n7906) );
  OAI22_X1 U5561 ( .A1(n10776), .A2(n11968), .B1(n11972), .B2(n13673), .ZN(
        n7905) );
  OAI22_X1 U5562 ( .A1(n10769), .A2(n11968), .B1(n11972), .B2(n13672), .ZN(
        n7904) );
  OAI22_X1 U5563 ( .A1(n10762), .A2(n11968), .B1(n11973), .B2(n13671), .ZN(
        n7903) );
  OAI22_X1 U5564 ( .A1(n10755), .A2(n11968), .B1(n11973), .B2(n13670), .ZN(
        n7902) );
  OAI22_X1 U5565 ( .A1(n10748), .A2(n11968), .B1(n11973), .B2(n13669), .ZN(
        n7901) );
  OAI22_X1 U5566 ( .A1(n10741), .A2(n11968), .B1(n11973), .B2(n13668), .ZN(
        n7900) );
  OAI22_X1 U5567 ( .A1(n10734), .A2(n11968), .B1(n11974), .B2(n13667), .ZN(
        n7899) );
  OAI22_X1 U5568 ( .A1(n10727), .A2(n11968), .B1(n11974), .B2(n13666), .ZN(
        n7898) );
  OAI22_X1 U5569 ( .A1(n10720), .A2(n11968), .B1(n11974), .B2(n13665), .ZN(
        n7897) );
  OAI22_X1 U5570 ( .A1(n10713), .A2(n11968), .B1(n11974), .B2(n13664), .ZN(
        n7896) );
  OAI22_X1 U5571 ( .A1(n10706), .A2(n11967), .B1(n11975), .B2(n13663), .ZN(
        n7895) );
  OAI22_X1 U5572 ( .A1(n10699), .A2(n11967), .B1(n11975), .B2(n13662), .ZN(
        n7894) );
  OAI22_X1 U5573 ( .A1(n10692), .A2(n11967), .B1(n11975), .B2(n13661), .ZN(
        n7893) );
  OAI22_X1 U5574 ( .A1(n10685), .A2(n11967), .B1(n11975), .B2(n13660), .ZN(
        n7892) );
  OAI22_X1 U5575 ( .A1(n10678), .A2(n11967), .B1(n11976), .B2(n13659), .ZN(
        n7891) );
  OAI22_X1 U5576 ( .A1(n10671), .A2(n11967), .B1(n11976), .B2(n13658), .ZN(
        n7890) );
  OAI22_X1 U5577 ( .A1(n10664), .A2(n11967), .B1(n11976), .B2(n13657), .ZN(
        n7889) );
  OAI22_X1 U5578 ( .A1(n10657), .A2(n11967), .B1(n11976), .B2(n13656), .ZN(
        n7888) );
  OAI22_X1 U5579 ( .A1(n10650), .A2(n11967), .B1(n11977), .B2(n13655), .ZN(
        n7887) );
  OAI22_X1 U5580 ( .A1(n10643), .A2(n11967), .B1(n11977), .B2(n13654), .ZN(
        n7886) );
  OAI22_X1 U5581 ( .A1(n10636), .A2(n11967), .B1(n11977), .B2(n13653), .ZN(
        n7885) );
  OAI22_X1 U5582 ( .A1(n10629), .A2(n11967), .B1(n11977), .B2(n13652), .ZN(
        n7884) );
  OAI22_X1 U5583 ( .A1(n10847), .A2(n11921), .B1(n11922), .B2(n13555), .ZN(
        n7787) );
  OAI22_X1 U5584 ( .A1(n10840), .A2(n11921), .B1(n11922), .B2(n13554), .ZN(
        n7786) );
  OAI22_X1 U5585 ( .A1(n10833), .A2(n11921), .B1(n11922), .B2(n13553), .ZN(
        n7785) );
  OAI22_X1 U5586 ( .A1(n10826), .A2(n11921), .B1(n11922), .B2(n13552), .ZN(
        n7784) );
  OAI22_X1 U5587 ( .A1(n10819), .A2(n11921), .B1(n11923), .B2(n13551), .ZN(
        n7783) );
  OAI22_X1 U5588 ( .A1(n10812), .A2(n11921), .B1(n11923), .B2(n13550), .ZN(
        n7782) );
  OAI22_X1 U5589 ( .A1(n10805), .A2(n11921), .B1(n11923), .B2(n13549), .ZN(
        n7781) );
  OAI22_X1 U5590 ( .A1(n10798), .A2(n11921), .B1(n11923), .B2(n13548), .ZN(
        n7780) );
  OAI22_X1 U5591 ( .A1(n10791), .A2(n11920), .B1(n11924), .B2(n13547), .ZN(
        n7779) );
  OAI22_X1 U5592 ( .A1(n10784), .A2(n11920), .B1(n11924), .B2(n13546), .ZN(
        n7778) );
  OAI22_X1 U5593 ( .A1(n10777), .A2(n11920), .B1(n11924), .B2(n13545), .ZN(
        n7777) );
  OAI22_X1 U5594 ( .A1(n10770), .A2(n11920), .B1(n11924), .B2(n13544), .ZN(
        n7776) );
  OAI22_X1 U5595 ( .A1(n10763), .A2(n11920), .B1(n11925), .B2(n13543), .ZN(
        n7775) );
  OAI22_X1 U5596 ( .A1(n10756), .A2(n11920), .B1(n11925), .B2(n13542), .ZN(
        n7774) );
  OAI22_X1 U5597 ( .A1(n10749), .A2(n11920), .B1(n11925), .B2(n13541), .ZN(
        n7773) );
  OAI22_X1 U5598 ( .A1(n10742), .A2(n11920), .B1(n11925), .B2(n13540), .ZN(
        n7772) );
  OAI22_X1 U5599 ( .A1(n10735), .A2(n11920), .B1(n11926), .B2(n13539), .ZN(
        n7771) );
  OAI22_X1 U5600 ( .A1(n10728), .A2(n11920), .B1(n11926), .B2(n13538), .ZN(
        n7770) );
  OAI22_X1 U5601 ( .A1(n10721), .A2(n11920), .B1(n11926), .B2(n13537), .ZN(
        n7769) );
  OAI22_X1 U5602 ( .A1(n10714), .A2(n11920), .B1(n11926), .B2(n13536), .ZN(
        n7768) );
  OAI22_X1 U5603 ( .A1(n10707), .A2(n11919), .B1(n11927), .B2(n13535), .ZN(
        n7767) );
  OAI22_X1 U5604 ( .A1(n10700), .A2(n11919), .B1(n11927), .B2(n13534), .ZN(
        n7766) );
  OAI22_X1 U5605 ( .A1(n10693), .A2(n11919), .B1(n11927), .B2(n13533), .ZN(
        n7765) );
  OAI22_X1 U5606 ( .A1(n10686), .A2(n11919), .B1(n11927), .B2(n13532), .ZN(
        n7764) );
  OAI22_X1 U5607 ( .A1(n10679), .A2(n11919), .B1(n11928), .B2(n13531), .ZN(
        n7763) );
  OAI22_X1 U5608 ( .A1(n10672), .A2(n11919), .B1(n11928), .B2(n13530), .ZN(
        n7762) );
  OAI22_X1 U5609 ( .A1(n10665), .A2(n11919), .B1(n11928), .B2(n13529), .ZN(
        n7761) );
  OAI22_X1 U5610 ( .A1(n10658), .A2(n11919), .B1(n11928), .B2(n13528), .ZN(
        n7760) );
  OAI22_X1 U5611 ( .A1(n10651), .A2(n11919), .B1(n11929), .B2(n13527), .ZN(
        n7759) );
  OAI22_X1 U5612 ( .A1(n10644), .A2(n11919), .B1(n11929), .B2(n13526), .ZN(
        n7758) );
  OAI22_X1 U5613 ( .A1(n10637), .A2(n11919), .B1(n11929), .B2(n13525), .ZN(
        n7757) );
  OAI22_X1 U5614 ( .A1(n10630), .A2(n11919), .B1(n11929), .B2(n13524), .ZN(
        n7756) );
  OAI22_X1 U5615 ( .A1(n10847), .A2(n11909), .B1(n11910), .B2(n13523), .ZN(
        n7755) );
  OAI22_X1 U5616 ( .A1(n10840), .A2(n11909), .B1(n11910), .B2(n13522), .ZN(
        n7754) );
  OAI22_X1 U5617 ( .A1(n10833), .A2(n11909), .B1(n11910), .B2(n13521), .ZN(
        n7753) );
  OAI22_X1 U5618 ( .A1(n10826), .A2(n11909), .B1(n11910), .B2(n13520), .ZN(
        n7752) );
  OAI22_X1 U5619 ( .A1(n10819), .A2(n11909), .B1(n11911), .B2(n13519), .ZN(
        n7751) );
  OAI22_X1 U5620 ( .A1(n10812), .A2(n11909), .B1(n11911), .B2(n13518), .ZN(
        n7750) );
  OAI22_X1 U5621 ( .A1(n10805), .A2(n11909), .B1(n11911), .B2(n13517), .ZN(
        n7749) );
  OAI22_X1 U5622 ( .A1(n10798), .A2(n11909), .B1(n11911), .B2(n13516), .ZN(
        n7748) );
  OAI22_X1 U5623 ( .A1(n10791), .A2(n11908), .B1(n11912), .B2(n13515), .ZN(
        n7747) );
  OAI22_X1 U5624 ( .A1(n10784), .A2(n11908), .B1(n11912), .B2(n13514), .ZN(
        n7746) );
  OAI22_X1 U5625 ( .A1(n10777), .A2(n11908), .B1(n11912), .B2(n13513), .ZN(
        n7745) );
  OAI22_X1 U5626 ( .A1(n10770), .A2(n11908), .B1(n11912), .B2(n13512), .ZN(
        n7744) );
  OAI22_X1 U5627 ( .A1(n10763), .A2(n11908), .B1(n11913), .B2(n13511), .ZN(
        n7743) );
  OAI22_X1 U5628 ( .A1(n10756), .A2(n11908), .B1(n11913), .B2(n13510), .ZN(
        n7742) );
  OAI22_X1 U5629 ( .A1(n10749), .A2(n11908), .B1(n11913), .B2(n13509), .ZN(
        n7741) );
  OAI22_X1 U5630 ( .A1(n10742), .A2(n11908), .B1(n11913), .B2(n13508), .ZN(
        n7740) );
  OAI22_X1 U5631 ( .A1(n10735), .A2(n11908), .B1(n11914), .B2(n13507), .ZN(
        n7739) );
  OAI22_X1 U5632 ( .A1(n10728), .A2(n11908), .B1(n11914), .B2(n13506), .ZN(
        n7738) );
  OAI22_X1 U5633 ( .A1(n10721), .A2(n11908), .B1(n11914), .B2(n13505), .ZN(
        n7737) );
  OAI22_X1 U5634 ( .A1(n10714), .A2(n11908), .B1(n11914), .B2(n13504), .ZN(
        n7736) );
  OAI22_X1 U5635 ( .A1(n10707), .A2(n11907), .B1(n11915), .B2(n13503), .ZN(
        n7735) );
  OAI22_X1 U5636 ( .A1(n10700), .A2(n11907), .B1(n11915), .B2(n13502), .ZN(
        n7734) );
  OAI22_X1 U5637 ( .A1(n10693), .A2(n11907), .B1(n11915), .B2(n13501), .ZN(
        n7733) );
  OAI22_X1 U5638 ( .A1(n10686), .A2(n11907), .B1(n11915), .B2(n13500), .ZN(
        n7732) );
  OAI22_X1 U5639 ( .A1(n10679), .A2(n11907), .B1(n11916), .B2(n13499), .ZN(
        n7731) );
  OAI22_X1 U5640 ( .A1(n10672), .A2(n11907), .B1(n11916), .B2(n13498), .ZN(
        n7730) );
  OAI22_X1 U5641 ( .A1(n10665), .A2(n11907), .B1(n11916), .B2(n13497), .ZN(
        n7729) );
  OAI22_X1 U5642 ( .A1(n10658), .A2(n11907), .B1(n11916), .B2(n13496), .ZN(
        n7728) );
  OAI22_X1 U5643 ( .A1(n10651), .A2(n11907), .B1(n11917), .B2(n13495), .ZN(
        n7727) );
  OAI22_X1 U5644 ( .A1(n10644), .A2(n11907), .B1(n11917), .B2(n13494), .ZN(
        n7726) );
  OAI22_X1 U5645 ( .A1(n10637), .A2(n11907), .B1(n11917), .B2(n13493), .ZN(
        n7725) );
  OAI22_X1 U5646 ( .A1(n10630), .A2(n11907), .B1(n11917), .B2(n13492), .ZN(
        n7724) );
  OAI22_X1 U5647 ( .A1(n10848), .A2(n11765), .B1(n11766), .B2(n13395), .ZN(
        n7371) );
  OAI22_X1 U5648 ( .A1(n10841), .A2(n11765), .B1(n11766), .B2(n13394), .ZN(
        n7370) );
  OAI22_X1 U5649 ( .A1(n10834), .A2(n11765), .B1(n11766), .B2(n13393), .ZN(
        n7369) );
  OAI22_X1 U5650 ( .A1(n10827), .A2(n11765), .B1(n11766), .B2(n13392), .ZN(
        n7368) );
  OAI22_X1 U5651 ( .A1(n10820), .A2(n11765), .B1(n11767), .B2(n13391), .ZN(
        n7367) );
  OAI22_X1 U5652 ( .A1(n10813), .A2(n11765), .B1(n11767), .B2(n13390), .ZN(
        n7366) );
  OAI22_X1 U5653 ( .A1(n10806), .A2(n11765), .B1(n11767), .B2(n13389), .ZN(
        n7365) );
  OAI22_X1 U5654 ( .A1(n10799), .A2(n11765), .B1(n11767), .B2(n13388), .ZN(
        n7364) );
  OAI22_X1 U5655 ( .A1(n10792), .A2(n11764), .B1(n11768), .B2(n13387), .ZN(
        n7363) );
  OAI22_X1 U5656 ( .A1(n10785), .A2(n11764), .B1(n11768), .B2(n13386), .ZN(
        n7362) );
  OAI22_X1 U5657 ( .A1(n10778), .A2(n11764), .B1(n11768), .B2(n13385), .ZN(
        n7361) );
  OAI22_X1 U5658 ( .A1(n10771), .A2(n11764), .B1(n11768), .B2(n13384), .ZN(
        n7360) );
  OAI22_X1 U5659 ( .A1(n10764), .A2(n11764), .B1(n11769), .B2(n13383), .ZN(
        n7359) );
  OAI22_X1 U5660 ( .A1(n10757), .A2(n11764), .B1(n11769), .B2(n13382), .ZN(
        n7358) );
  OAI22_X1 U5661 ( .A1(n10750), .A2(n11764), .B1(n11769), .B2(n13381), .ZN(
        n7357) );
  OAI22_X1 U5662 ( .A1(n10743), .A2(n11764), .B1(n11769), .B2(n13380), .ZN(
        n7356) );
  OAI22_X1 U5663 ( .A1(n10736), .A2(n11764), .B1(n11770), .B2(n13379), .ZN(
        n7355) );
  OAI22_X1 U5664 ( .A1(n10729), .A2(n11764), .B1(n11770), .B2(n13378), .ZN(
        n7354) );
  OAI22_X1 U5665 ( .A1(n10722), .A2(n11764), .B1(n11770), .B2(n13377), .ZN(
        n7353) );
  OAI22_X1 U5666 ( .A1(n10715), .A2(n11764), .B1(n11770), .B2(n13376), .ZN(
        n7352) );
  OAI22_X1 U5667 ( .A1(n10708), .A2(n11763), .B1(n11771), .B2(n13375), .ZN(
        n7351) );
  OAI22_X1 U5668 ( .A1(n10701), .A2(n11763), .B1(n11771), .B2(n13374), .ZN(
        n7350) );
  OAI22_X1 U5669 ( .A1(n10694), .A2(n11763), .B1(n11771), .B2(n13373), .ZN(
        n7349) );
  OAI22_X1 U5670 ( .A1(n10687), .A2(n11763), .B1(n11771), .B2(n13372), .ZN(
        n7348) );
  OAI22_X1 U5671 ( .A1(n10680), .A2(n11763), .B1(n11772), .B2(n13371), .ZN(
        n7347) );
  OAI22_X1 U5672 ( .A1(n10673), .A2(n11763), .B1(n11772), .B2(n13370), .ZN(
        n7346) );
  OAI22_X1 U5673 ( .A1(n10666), .A2(n11763), .B1(n11772), .B2(n13369), .ZN(
        n7345) );
  OAI22_X1 U5674 ( .A1(n10659), .A2(n11763), .B1(n11772), .B2(n13368), .ZN(
        n7344) );
  OAI22_X1 U5675 ( .A1(n10652), .A2(n11763), .B1(n11773), .B2(n13367), .ZN(
        n7343) );
  OAI22_X1 U5676 ( .A1(n10645), .A2(n11763), .B1(n11773), .B2(n13366), .ZN(
        n7342) );
  OAI22_X1 U5677 ( .A1(n10638), .A2(n11763), .B1(n11773), .B2(n13365), .ZN(
        n7341) );
  OAI22_X1 U5678 ( .A1(n10631), .A2(n11763), .B1(n11773), .B2(n13364), .ZN(
        n7340) );
  OAI22_X1 U5679 ( .A1(n10806), .A2(n11753), .B1(n11755), .B2(n13357), .ZN(
        n7333) );
  OAI22_X1 U5680 ( .A1(n10799), .A2(n11753), .B1(n11755), .B2(n13356), .ZN(
        n7332) );
  OAI22_X1 U5681 ( .A1(n10792), .A2(n11752), .B1(n11756), .B2(n13355), .ZN(
        n7331) );
  OAI22_X1 U5682 ( .A1(n10785), .A2(n11752), .B1(n11756), .B2(n13354), .ZN(
        n7330) );
  OAI22_X1 U5683 ( .A1(n10778), .A2(n11752), .B1(n11756), .B2(n13353), .ZN(
        n7329) );
  OAI22_X1 U5684 ( .A1(n10771), .A2(n11752), .B1(n11756), .B2(n13352), .ZN(
        n7328) );
  OAI22_X1 U5685 ( .A1(n10764), .A2(n11752), .B1(n11757), .B2(n13351), .ZN(
        n7327) );
  OAI22_X1 U5686 ( .A1(n10757), .A2(n11752), .B1(n11757), .B2(n13350), .ZN(
        n7326) );
  OAI22_X1 U5687 ( .A1(n10750), .A2(n11752), .B1(n11757), .B2(n13349), .ZN(
        n7325) );
  OAI22_X1 U5688 ( .A1(n10743), .A2(n11752), .B1(n11757), .B2(n13348), .ZN(
        n7324) );
  OAI22_X1 U5689 ( .A1(n10736), .A2(n11752), .B1(n11758), .B2(n13347), .ZN(
        n7323) );
  OAI22_X1 U5690 ( .A1(n10729), .A2(n11752), .B1(n11758), .B2(n13346), .ZN(
        n7322) );
  OAI22_X1 U5691 ( .A1(n10722), .A2(n11752), .B1(n11758), .B2(n13345), .ZN(
        n7321) );
  OAI22_X1 U5692 ( .A1(n10715), .A2(n11752), .B1(n11758), .B2(n13344), .ZN(
        n7320) );
  OAI22_X1 U5693 ( .A1(n10708), .A2(n11751), .B1(n11759), .B2(n13343), .ZN(
        n7319) );
  OAI22_X1 U5694 ( .A1(n10701), .A2(n11751), .B1(n11759), .B2(n13342), .ZN(
        n7318) );
  OAI22_X1 U5695 ( .A1(n10694), .A2(n11751), .B1(n11759), .B2(n13341), .ZN(
        n7317) );
  OAI22_X1 U5696 ( .A1(n10687), .A2(n11751), .B1(n11759), .B2(n13340), .ZN(
        n7316) );
  OAI22_X1 U5697 ( .A1(n10680), .A2(n11751), .B1(n11760), .B2(n13339), .ZN(
        n7315) );
  OAI22_X1 U5698 ( .A1(n10673), .A2(n11751), .B1(n11760), .B2(n13338), .ZN(
        n7314) );
  OAI22_X1 U5699 ( .A1(n10666), .A2(n11751), .B1(n11760), .B2(n13337), .ZN(
        n7313) );
  OAI22_X1 U5700 ( .A1(n10659), .A2(n11751), .B1(n11760), .B2(n13336), .ZN(
        n7312) );
  OAI22_X1 U5701 ( .A1(n10652), .A2(n11751), .B1(n11761), .B2(n13335), .ZN(
        n7311) );
  OAI22_X1 U5702 ( .A1(n10645), .A2(n11751), .B1(n11761), .B2(n13334), .ZN(
        n7310) );
  OAI22_X1 U5703 ( .A1(n10638), .A2(n11751), .B1(n11761), .B2(n13333), .ZN(
        n7309) );
  OAI22_X1 U5704 ( .A1(n10631), .A2(n11751), .B1(n11761), .B2(n13332), .ZN(
        n7308) );
  OAI22_X1 U5705 ( .A1(n10848), .A2(n11741), .B1(n11742), .B2(n13331), .ZN(
        n7307) );
  OAI22_X1 U5706 ( .A1(n10841), .A2(n11741), .B1(n11742), .B2(n13330), .ZN(
        n7306) );
  OAI22_X1 U5707 ( .A1(n10834), .A2(n11741), .B1(n11742), .B2(n13329), .ZN(
        n7305) );
  OAI22_X1 U5708 ( .A1(n10827), .A2(n11741), .B1(n11742), .B2(n13328), .ZN(
        n7304) );
  OAI22_X1 U5709 ( .A1(n10820), .A2(n11741), .B1(n11743), .B2(n13327), .ZN(
        n7303) );
  OAI22_X1 U5710 ( .A1(n10813), .A2(n11741), .B1(n11743), .B2(n13326), .ZN(
        n7302) );
  OAI22_X1 U5711 ( .A1(n10806), .A2(n11741), .B1(n11743), .B2(n13325), .ZN(
        n7301) );
  OAI22_X1 U5712 ( .A1(n10799), .A2(n11741), .B1(n11743), .B2(n13324), .ZN(
        n7300) );
  OAI22_X1 U5713 ( .A1(n10792), .A2(n11740), .B1(n11744), .B2(n13323), .ZN(
        n7299) );
  OAI22_X1 U5714 ( .A1(n10785), .A2(n11740), .B1(n11744), .B2(n13322), .ZN(
        n7298) );
  OAI22_X1 U5715 ( .A1(n10778), .A2(n11740), .B1(n11744), .B2(n13321), .ZN(
        n7297) );
  OAI22_X1 U5716 ( .A1(n10771), .A2(n11740), .B1(n11744), .B2(n13320), .ZN(
        n7296) );
  OAI22_X1 U5717 ( .A1(n10764), .A2(n11740), .B1(n11745), .B2(n13319), .ZN(
        n7295) );
  OAI22_X1 U5718 ( .A1(n10757), .A2(n11740), .B1(n11745), .B2(n13318), .ZN(
        n7294) );
  OAI22_X1 U5719 ( .A1(n10750), .A2(n11740), .B1(n11745), .B2(n13317), .ZN(
        n7293) );
  OAI22_X1 U5720 ( .A1(n10743), .A2(n11740), .B1(n11745), .B2(n13316), .ZN(
        n7292) );
  OAI22_X1 U5721 ( .A1(n10736), .A2(n11740), .B1(n11746), .B2(n13315), .ZN(
        n7291) );
  OAI22_X1 U5722 ( .A1(n10729), .A2(n11740), .B1(n11746), .B2(n13314), .ZN(
        n7290) );
  OAI22_X1 U5723 ( .A1(n10722), .A2(n11740), .B1(n11746), .B2(n13313), .ZN(
        n7289) );
  OAI22_X1 U5724 ( .A1(n10715), .A2(n11740), .B1(n11746), .B2(n13312), .ZN(
        n7288) );
  OAI22_X1 U5725 ( .A1(n10708), .A2(n11739), .B1(n11747), .B2(n13311), .ZN(
        n7287) );
  OAI22_X1 U5726 ( .A1(n10701), .A2(n11739), .B1(n11747), .B2(n13310), .ZN(
        n7286) );
  OAI22_X1 U5727 ( .A1(n10694), .A2(n11739), .B1(n11747), .B2(n13309), .ZN(
        n7285) );
  OAI22_X1 U5728 ( .A1(n10687), .A2(n11739), .B1(n11747), .B2(n13308), .ZN(
        n7284) );
  OAI22_X1 U5729 ( .A1(n10680), .A2(n11739), .B1(n11748), .B2(n13307), .ZN(
        n7283) );
  OAI22_X1 U5730 ( .A1(n10673), .A2(n11739), .B1(n11748), .B2(n13306), .ZN(
        n7282) );
  OAI22_X1 U5731 ( .A1(n10666), .A2(n11739), .B1(n11748), .B2(n13305), .ZN(
        n7281) );
  OAI22_X1 U5732 ( .A1(n10659), .A2(n11739), .B1(n11748), .B2(n13304), .ZN(
        n7280) );
  OAI22_X1 U5733 ( .A1(n10652), .A2(n11739), .B1(n11749), .B2(n13303), .ZN(
        n7279) );
  OAI22_X1 U5734 ( .A1(n10645), .A2(n11739), .B1(n11749), .B2(n13302), .ZN(
        n7278) );
  OAI22_X1 U5735 ( .A1(n10638), .A2(n11739), .B1(n11749), .B2(n13301), .ZN(
        n7277) );
  OAI22_X1 U5736 ( .A1(n10631), .A2(n11739), .B1(n11749), .B2(n13300), .ZN(
        n7276) );
  OAI22_X1 U5737 ( .A1(n10848), .A2(n11729), .B1(n11730), .B2(n13299), .ZN(
        n7275) );
  OAI22_X1 U5738 ( .A1(n10841), .A2(n11729), .B1(n11730), .B2(n13298), .ZN(
        n7274) );
  OAI22_X1 U5739 ( .A1(n10834), .A2(n11729), .B1(n11730), .B2(n13297), .ZN(
        n7273) );
  OAI22_X1 U5740 ( .A1(n10827), .A2(n11729), .B1(n11730), .B2(n13296), .ZN(
        n7272) );
  OAI22_X1 U5741 ( .A1(n10820), .A2(n11729), .B1(n11731), .B2(n13295), .ZN(
        n7271) );
  OAI22_X1 U5742 ( .A1(n10813), .A2(n11729), .B1(n11731), .B2(n13294), .ZN(
        n7270) );
  OAI22_X1 U5743 ( .A1(n10806), .A2(n11729), .B1(n11731), .B2(n13293), .ZN(
        n7269) );
  OAI22_X1 U5744 ( .A1(n10799), .A2(n11729), .B1(n11731), .B2(n13292), .ZN(
        n7268) );
  OAI22_X1 U5745 ( .A1(n10792), .A2(n11728), .B1(n11732), .B2(n13291), .ZN(
        n7267) );
  OAI22_X1 U5746 ( .A1(n10785), .A2(n11728), .B1(n11732), .B2(n13290), .ZN(
        n7266) );
  OAI22_X1 U5747 ( .A1(n10778), .A2(n11728), .B1(n11732), .B2(n13289), .ZN(
        n7265) );
  OAI22_X1 U5748 ( .A1(n10771), .A2(n11728), .B1(n11732), .B2(n13288), .ZN(
        n7264) );
  OAI22_X1 U5749 ( .A1(n10764), .A2(n11728), .B1(n11733), .B2(n13287), .ZN(
        n7263) );
  OAI22_X1 U5750 ( .A1(n10757), .A2(n11728), .B1(n11733), .B2(n13286), .ZN(
        n7262) );
  OAI22_X1 U5751 ( .A1(n10750), .A2(n11728), .B1(n11733), .B2(n13285), .ZN(
        n7261) );
  OAI22_X1 U5752 ( .A1(n10743), .A2(n11728), .B1(n11733), .B2(n13284), .ZN(
        n7260) );
  OAI22_X1 U5753 ( .A1(n10736), .A2(n11728), .B1(n11734), .B2(n13283), .ZN(
        n7259) );
  OAI22_X1 U5754 ( .A1(n10729), .A2(n11728), .B1(n11734), .B2(n13282), .ZN(
        n7258) );
  OAI22_X1 U5755 ( .A1(n10722), .A2(n11728), .B1(n11734), .B2(n13281), .ZN(
        n7257) );
  OAI22_X1 U5756 ( .A1(n10715), .A2(n11728), .B1(n11734), .B2(n13280), .ZN(
        n7256) );
  OAI22_X1 U5757 ( .A1(n10708), .A2(n11727), .B1(n11735), .B2(n13279), .ZN(
        n7255) );
  OAI22_X1 U5758 ( .A1(n10701), .A2(n11727), .B1(n11735), .B2(n13278), .ZN(
        n7254) );
  OAI22_X1 U5759 ( .A1(n10694), .A2(n11727), .B1(n11735), .B2(n13277), .ZN(
        n7253) );
  OAI22_X1 U5760 ( .A1(n10687), .A2(n11727), .B1(n11735), .B2(n13276), .ZN(
        n7252) );
  OAI22_X1 U5761 ( .A1(n10680), .A2(n11727), .B1(n11736), .B2(n13275), .ZN(
        n7251) );
  OAI22_X1 U5762 ( .A1(n10673), .A2(n11727), .B1(n11736), .B2(n13274), .ZN(
        n7250) );
  OAI22_X1 U5763 ( .A1(n10666), .A2(n11727), .B1(n11736), .B2(n13273), .ZN(
        n7249) );
  OAI22_X1 U5764 ( .A1(n10659), .A2(n11727), .B1(n11736), .B2(n13272), .ZN(
        n7248) );
  OAI22_X1 U5765 ( .A1(n10652), .A2(n11727), .B1(n11737), .B2(n13271), .ZN(
        n7247) );
  OAI22_X1 U5766 ( .A1(n10645), .A2(n11727), .B1(n11737), .B2(n13270), .ZN(
        n7246) );
  OAI22_X1 U5767 ( .A1(n10638), .A2(n11727), .B1(n11737), .B2(n13269), .ZN(
        n7245) );
  OAI22_X1 U5768 ( .A1(n10631), .A2(n11727), .B1(n11737), .B2(n13268), .ZN(
        n7244) );
  OAI22_X1 U5769 ( .A1(n10848), .A2(n11717), .B1(n11718), .B2(n13267), .ZN(
        n7243) );
  OAI22_X1 U5770 ( .A1(n10841), .A2(n11717), .B1(n11718), .B2(n13266), .ZN(
        n7242) );
  OAI22_X1 U5771 ( .A1(n10834), .A2(n11717), .B1(n11718), .B2(n13265), .ZN(
        n7241) );
  OAI22_X1 U5772 ( .A1(n10827), .A2(n11717), .B1(n11718), .B2(n13264), .ZN(
        n7240) );
  OAI22_X1 U5773 ( .A1(n10820), .A2(n11717), .B1(n11719), .B2(n13263), .ZN(
        n7239) );
  OAI22_X1 U5774 ( .A1(n10813), .A2(n11717), .B1(n11719), .B2(n13262), .ZN(
        n7238) );
  OAI22_X1 U5775 ( .A1(n10806), .A2(n11717), .B1(n11719), .B2(n13261), .ZN(
        n7237) );
  OAI22_X1 U5776 ( .A1(n10799), .A2(n11717), .B1(n11719), .B2(n13260), .ZN(
        n7236) );
  OAI22_X1 U5777 ( .A1(n10792), .A2(n11716), .B1(n11720), .B2(n13259), .ZN(
        n7235) );
  OAI22_X1 U5778 ( .A1(n10785), .A2(n11716), .B1(n11720), .B2(n13258), .ZN(
        n7234) );
  OAI22_X1 U5779 ( .A1(n10778), .A2(n11716), .B1(n11720), .B2(n13257), .ZN(
        n7233) );
  OAI22_X1 U5780 ( .A1(n10771), .A2(n11716), .B1(n11720), .B2(n13256), .ZN(
        n7232) );
  OAI22_X1 U5781 ( .A1(n10764), .A2(n11716), .B1(n11721), .B2(n13255), .ZN(
        n7231) );
  OAI22_X1 U5782 ( .A1(n10757), .A2(n11716), .B1(n11721), .B2(n13254), .ZN(
        n7230) );
  OAI22_X1 U5783 ( .A1(n10750), .A2(n11716), .B1(n11721), .B2(n13253), .ZN(
        n7229) );
  OAI22_X1 U5784 ( .A1(n10743), .A2(n11716), .B1(n11721), .B2(n13252), .ZN(
        n7228) );
  OAI22_X1 U5785 ( .A1(n10736), .A2(n11716), .B1(n11722), .B2(n13251), .ZN(
        n7227) );
  OAI22_X1 U5786 ( .A1(n10729), .A2(n11716), .B1(n11722), .B2(n13250), .ZN(
        n7226) );
  OAI22_X1 U5787 ( .A1(n10722), .A2(n11716), .B1(n11722), .B2(n13249), .ZN(
        n7225) );
  OAI22_X1 U5788 ( .A1(n10715), .A2(n11716), .B1(n11722), .B2(n13248), .ZN(
        n7224) );
  OAI22_X1 U5789 ( .A1(n10708), .A2(n11715), .B1(n11723), .B2(n13247), .ZN(
        n7223) );
  OAI22_X1 U5790 ( .A1(n10701), .A2(n11715), .B1(n11723), .B2(n13246), .ZN(
        n7222) );
  OAI22_X1 U5791 ( .A1(n10694), .A2(n11715), .B1(n11723), .B2(n13245), .ZN(
        n7221) );
  OAI22_X1 U5792 ( .A1(n10687), .A2(n11715), .B1(n11723), .B2(n13244), .ZN(
        n7220) );
  OAI22_X1 U5793 ( .A1(n10680), .A2(n11715), .B1(n11724), .B2(n13243), .ZN(
        n7219) );
  OAI22_X1 U5794 ( .A1(n10673), .A2(n11715), .B1(n11724), .B2(n13242), .ZN(
        n7218) );
  OAI22_X1 U5795 ( .A1(n10666), .A2(n11715), .B1(n11724), .B2(n13241), .ZN(
        n7217) );
  OAI22_X1 U5796 ( .A1(n10659), .A2(n11715), .B1(n11724), .B2(n13240), .ZN(
        n7216) );
  OAI22_X1 U5797 ( .A1(n10652), .A2(n11715), .B1(n11725), .B2(n13239), .ZN(
        n7215) );
  OAI22_X1 U5798 ( .A1(n10645), .A2(n11715), .B1(n11725), .B2(n13238), .ZN(
        n7214) );
  OAI22_X1 U5799 ( .A1(n10638), .A2(n11715), .B1(n11725), .B2(n13237), .ZN(
        n7213) );
  OAI22_X1 U5800 ( .A1(n10631), .A2(n11715), .B1(n11725), .B2(n13236), .ZN(
        n7212) );
  OAI22_X1 U5801 ( .A1(n10848), .A2(n11705), .B1(n11706), .B2(n13235), .ZN(
        n7211) );
  OAI22_X1 U5802 ( .A1(n10841), .A2(n11705), .B1(n11706), .B2(n13234), .ZN(
        n7210) );
  OAI22_X1 U5803 ( .A1(n10834), .A2(n11705), .B1(n11706), .B2(n13233), .ZN(
        n7209) );
  OAI22_X1 U5804 ( .A1(n10827), .A2(n11705), .B1(n11706), .B2(n13232), .ZN(
        n7208) );
  OAI22_X1 U5805 ( .A1(n10820), .A2(n11705), .B1(n11707), .B2(n13231), .ZN(
        n7207) );
  OAI22_X1 U5806 ( .A1(n10813), .A2(n11705), .B1(n11707), .B2(n13230), .ZN(
        n7206) );
  OAI22_X1 U5807 ( .A1(n10806), .A2(n11705), .B1(n11707), .B2(n13229), .ZN(
        n7205) );
  OAI22_X1 U5808 ( .A1(n10799), .A2(n11705), .B1(n11707), .B2(n13228), .ZN(
        n7204) );
  OAI22_X1 U5809 ( .A1(n10792), .A2(n11704), .B1(n11708), .B2(n13227), .ZN(
        n7203) );
  OAI22_X1 U5810 ( .A1(n10785), .A2(n11704), .B1(n11708), .B2(n13226), .ZN(
        n7202) );
  OAI22_X1 U5811 ( .A1(n10778), .A2(n11704), .B1(n11708), .B2(n13225), .ZN(
        n7201) );
  OAI22_X1 U5812 ( .A1(n10771), .A2(n11704), .B1(n11708), .B2(n13224), .ZN(
        n7200) );
  OAI22_X1 U5813 ( .A1(n10764), .A2(n11704), .B1(n11709), .B2(n13223), .ZN(
        n7199) );
  OAI22_X1 U5814 ( .A1(n10757), .A2(n11704), .B1(n11709), .B2(n13222), .ZN(
        n7198) );
  OAI22_X1 U5815 ( .A1(n10750), .A2(n11704), .B1(n11709), .B2(n13221), .ZN(
        n7197) );
  OAI22_X1 U5816 ( .A1(n10743), .A2(n11704), .B1(n11709), .B2(n13220), .ZN(
        n7196) );
  OAI22_X1 U5817 ( .A1(n10736), .A2(n11704), .B1(n11710), .B2(n13219), .ZN(
        n7195) );
  OAI22_X1 U5818 ( .A1(n10729), .A2(n11704), .B1(n11710), .B2(n13218), .ZN(
        n7194) );
  OAI22_X1 U5819 ( .A1(n10722), .A2(n11704), .B1(n11710), .B2(n13217), .ZN(
        n7193) );
  OAI22_X1 U5820 ( .A1(n10715), .A2(n11704), .B1(n11710), .B2(n13216), .ZN(
        n7192) );
  OAI22_X1 U5821 ( .A1(n10708), .A2(n11703), .B1(n11711), .B2(n13215), .ZN(
        n7191) );
  OAI22_X1 U5822 ( .A1(n10701), .A2(n11703), .B1(n11711), .B2(n13214), .ZN(
        n7190) );
  OAI22_X1 U5823 ( .A1(n10694), .A2(n11703), .B1(n11711), .B2(n13213), .ZN(
        n7189) );
  OAI22_X1 U5824 ( .A1(n10687), .A2(n11703), .B1(n11711), .B2(n13212), .ZN(
        n7188) );
  OAI22_X1 U5826 ( .A1(n10680), .A2(n11703), .B1(n11712), .B2(n13211), .ZN(
        n7187) );
  OAI22_X1 U5827 ( .A1(n10673), .A2(n11703), .B1(n11712), .B2(n13210), .ZN(
        n7186) );
  OAI22_X1 U5828 ( .A1(n10666), .A2(n11703), .B1(n11712), .B2(n13209), .ZN(
        n7185) );
  OAI22_X1 U5829 ( .A1(n10659), .A2(n11703), .B1(n11712), .B2(n13208), .ZN(
        n7184) );
  OAI22_X1 U5830 ( .A1(n10652), .A2(n11703), .B1(n11713), .B2(n13207), .ZN(
        n7183) );
  OAI22_X1 U5831 ( .A1(n10645), .A2(n11703), .B1(n11713), .B2(n13206), .ZN(
        n7182) );
  OAI22_X1 U5832 ( .A1(n10638), .A2(n11703), .B1(n11713), .B2(n13205), .ZN(
        n7181) );
  OAI22_X1 U5833 ( .A1(n10631), .A2(n11703), .B1(n11713), .B2(n13204), .ZN(
        n7180) );
  OAI22_X1 U5834 ( .A1(n10848), .A2(n11657), .B1(n11658), .B2(n13107), .ZN(
        n7083) );
  OAI22_X1 U5835 ( .A1(n10841), .A2(n11657), .B1(n11658), .B2(n13106), .ZN(
        n7082) );
  OAI22_X1 U5836 ( .A1(n10834), .A2(n11657), .B1(n11658), .B2(n13105), .ZN(
        n7081) );
  OAI22_X1 U5837 ( .A1(n10827), .A2(n11657), .B1(n11658), .B2(n13104), .ZN(
        n7080) );
  OAI22_X1 U5838 ( .A1(n10820), .A2(n11657), .B1(n11659), .B2(n13103), .ZN(
        n7079) );
  OAI22_X1 U5839 ( .A1(n10813), .A2(n11657), .B1(n11659), .B2(n13102), .ZN(
        n7078) );
  OAI22_X1 U5840 ( .A1(n10806), .A2(n11657), .B1(n11659), .B2(n13101), .ZN(
        n7077) );
  OAI22_X1 U5841 ( .A1(n10799), .A2(n11657), .B1(n11659), .B2(n13100), .ZN(
        n7076) );
  OAI22_X1 U5842 ( .A1(n10792), .A2(n11656), .B1(n11660), .B2(n13099), .ZN(
        n7075) );
  OAI22_X1 U5843 ( .A1(n10785), .A2(n11656), .B1(n11660), .B2(n13098), .ZN(
        n7074) );
  OAI22_X1 U5844 ( .A1(n10778), .A2(n11656), .B1(n11660), .B2(n13097), .ZN(
        n7073) );
  OAI22_X1 U5845 ( .A1(n10771), .A2(n11656), .B1(n11660), .B2(n13096), .ZN(
        n7072) );
  OAI22_X1 U5846 ( .A1(n10764), .A2(n11656), .B1(n11661), .B2(n13095), .ZN(
        n7071) );
  OAI22_X1 U5847 ( .A1(n10757), .A2(n11656), .B1(n11661), .B2(n13094), .ZN(
        n7070) );
  OAI22_X1 U5848 ( .A1(n10750), .A2(n11656), .B1(n11661), .B2(n13093), .ZN(
        n7069) );
  OAI22_X1 U5849 ( .A1(n10743), .A2(n11656), .B1(n11661), .B2(n13092), .ZN(
        n7068) );
  OAI22_X1 U5850 ( .A1(n10736), .A2(n11656), .B1(n11662), .B2(n13091), .ZN(
        n7067) );
  OAI22_X1 U5851 ( .A1(n10729), .A2(n11656), .B1(n11662), .B2(n13090), .ZN(
        n7066) );
  OAI22_X1 U5852 ( .A1(n10722), .A2(n11656), .B1(n11662), .B2(n13089), .ZN(
        n7065) );
  OAI22_X1 U5853 ( .A1(n10715), .A2(n11656), .B1(n11662), .B2(n13088), .ZN(
        n7064) );
  OAI22_X1 U5854 ( .A1(n10708), .A2(n11655), .B1(n11663), .B2(n13087), .ZN(
        n7063) );
  OAI22_X1 U5855 ( .A1(n10701), .A2(n11655), .B1(n11663), .B2(n13086), .ZN(
        n7062) );
  OAI22_X1 U5856 ( .A1(n10694), .A2(n11655), .B1(n11663), .B2(n13085), .ZN(
        n7061) );
  OAI22_X1 U5857 ( .A1(n10687), .A2(n11655), .B1(n11663), .B2(n13084), .ZN(
        n7060) );
  OAI22_X1 U5858 ( .A1(n10680), .A2(n11655), .B1(n11664), .B2(n13083), .ZN(
        n7059) );
  OAI22_X1 U5859 ( .A1(n10673), .A2(n11655), .B1(n11664), .B2(n13082), .ZN(
        n7058) );
  OAI22_X1 U5860 ( .A1(n10666), .A2(n11655), .B1(n11664), .B2(n13081), .ZN(
        n7057) );
  OAI22_X1 U5861 ( .A1(n10659), .A2(n11655), .B1(n11664), .B2(n13080), .ZN(
        n7056) );
  OAI22_X1 U5862 ( .A1(n10652), .A2(n11655), .B1(n11665), .B2(n13079), .ZN(
        n7055) );
  OAI22_X1 U5863 ( .A1(n10645), .A2(n11655), .B1(n11665), .B2(n13078), .ZN(
        n7054) );
  OAI22_X1 U5864 ( .A1(n10638), .A2(n11655), .B1(n11665), .B2(n13077), .ZN(
        n7053) );
  OAI22_X1 U5865 ( .A1(n10631), .A2(n11655), .B1(n11665), .B2(n13076), .ZN(
        n7052) );
  OAI22_X1 U5866 ( .A1(n10849), .A2(n11645), .B1(n11650), .B2(n13075), .ZN(
        n7051) );
  OAI22_X1 U5867 ( .A1(n10842), .A2(n11645), .B1(n11653), .B2(n13074), .ZN(
        n7050) );
  OAI22_X1 U5868 ( .A1(n10835), .A2(n11645), .B1(n11653), .B2(n13073), .ZN(
        n7049) );
  OAI22_X1 U5869 ( .A1(n10828), .A2(n11645), .B1(n11653), .B2(n13072), .ZN(
        n7048) );
  OAI22_X1 U5870 ( .A1(n10821), .A2(n11645), .B1(n11652), .B2(n13071), .ZN(
        n7047) );
  OAI22_X1 U5871 ( .A1(n10814), .A2(n11645), .B1(n11653), .B2(n13070), .ZN(
        n7046) );
  OAI22_X1 U5872 ( .A1(n10807), .A2(n11645), .B1(n11652), .B2(n13069), .ZN(
        n7045) );
  OAI22_X1 U5873 ( .A1(n10800), .A2(n11645), .B1(n11652), .B2(n13068), .ZN(
        n7044) );
  OAI22_X1 U5874 ( .A1(n10793), .A2(n11644), .B1(n11651), .B2(n13067), .ZN(
        n7043) );
  OAI22_X1 U5875 ( .A1(n10786), .A2(n11644), .B1(n11652), .B2(n13066), .ZN(
        n7042) );
  OAI22_X1 U5876 ( .A1(n10779), .A2(n11644), .B1(n11651), .B2(n13065), .ZN(
        n7041) );
  OAI22_X1 U5877 ( .A1(n10772), .A2(n11644), .B1(n11651), .B2(n13064), .ZN(
        n7040) );
  OAI22_X1 U5878 ( .A1(n10765), .A2(n11644), .B1(n11650), .B2(n13063), .ZN(
        n7039) );
  OAI22_X1 U5879 ( .A1(n10758), .A2(n11644), .B1(n11651), .B2(n13062), .ZN(
        n7038) );
  OAI22_X1 U5880 ( .A1(n10751), .A2(n11644), .B1(n11650), .B2(n13061), .ZN(
        n7037) );
  OAI22_X1 U5881 ( .A1(n10744), .A2(n11644), .B1(n11650), .B2(n13060), .ZN(
        n7036) );
  AOI21_X1 U5882 ( .B1(n2937), .B2(n2936), .A(n14518), .ZN(n2488) );
  OAI22_X1 U5883 ( .A1(n12419), .A2(n10844), .B1(n2913), .B2(n12418), .ZN(
        n9131) );
  OAI22_X1 U5884 ( .A1(n12419), .A2(n10837), .B1(n2912), .B2(n12418), .ZN(
        n9130) );
  OAI22_X1 U5885 ( .A1(n12419), .A2(n10830), .B1(n2911), .B2(n12418), .ZN(
        n9129) );
  OAI22_X1 U5886 ( .A1(n12419), .A2(n10823), .B1(n2910), .B2(n12418), .ZN(
        n9128) );
  OAI22_X1 U5887 ( .A1(n12419), .A2(n10816), .B1(n2909), .B2(n12418), .ZN(
        n9127) );
  OAI22_X1 U5888 ( .A1(n12420), .A2(n10809), .B1(n2908), .B2(n12418), .ZN(
        n9126) );
  OAI22_X1 U5889 ( .A1(n12420), .A2(n10802), .B1(n2907), .B2(n12418), .ZN(
        n9125) );
  OAI22_X1 U5890 ( .A1(n12420), .A2(n10795), .B1(n2906), .B2(n12418), .ZN(
        n9124) );
  OAI22_X1 U5891 ( .A1(n12420), .A2(n10788), .B1(n2905), .B2(n12417), .ZN(
        n9123) );
  OAI22_X1 U5892 ( .A1(n12420), .A2(n10781), .B1(n2904), .B2(n12417), .ZN(
        n9122) );
  OAI22_X1 U5893 ( .A1(n12421), .A2(n10774), .B1(n2903), .B2(n12417), .ZN(
        n9121) );
  OAI22_X1 U5894 ( .A1(n12421), .A2(n10767), .B1(n2902), .B2(n12417), .ZN(
        n9120) );
  OAI22_X1 U5895 ( .A1(n12421), .A2(n10760), .B1(n2901), .B2(n12417), .ZN(
        n9119) );
  OAI22_X1 U5896 ( .A1(n12421), .A2(n10753), .B1(n2900), .B2(n12417), .ZN(
        n9118) );
  OAI22_X1 U5897 ( .A1(n12421), .A2(n10746), .B1(n2899), .B2(n12417), .ZN(
        n9117) );
  OAI22_X1 U5898 ( .A1(n12422), .A2(n10739), .B1(n2898), .B2(n12417), .ZN(
        n9116) );
  OAI22_X1 U5899 ( .A1(n12422), .A2(n10732), .B1(n2897), .B2(n12417), .ZN(
        n9115) );
  OAI22_X1 U5900 ( .A1(n12422), .A2(n10725), .B1(n2896), .B2(n12417), .ZN(
        n9114) );
  OAI22_X1 U5901 ( .A1(n12422), .A2(n10718), .B1(n2895), .B2(n12417), .ZN(
        n9113) );
  OAI22_X1 U5902 ( .A1(n12422), .A2(n10711), .B1(n2894), .B2(n12417), .ZN(
        n9112) );
  OAI22_X1 U5903 ( .A1(n12423), .A2(n10704), .B1(n2893), .B2(n12416), .ZN(
        n9111) );
  OAI22_X1 U5904 ( .A1(n12423), .A2(n10697), .B1(n2892), .B2(n12416), .ZN(
        n9110) );
  OAI22_X1 U5905 ( .A1(n12423), .A2(n10690), .B1(n2891), .B2(n12416), .ZN(
        n9109) );
  OAI22_X1 U5906 ( .A1(n12423), .A2(n10683), .B1(n2890), .B2(n12416), .ZN(
        n9108) );
  OAI22_X1 U5907 ( .A1(n12423), .A2(n10676), .B1(n2889), .B2(n12416), .ZN(
        n9107) );
  OAI22_X1 U5908 ( .A1(n12424), .A2(n10669), .B1(n2888), .B2(n12416), .ZN(
        n9106) );
  OAI22_X1 U5909 ( .A1(n12424), .A2(n10662), .B1(n2887), .B2(n12416), .ZN(
        n9105) );
  OAI22_X1 U5910 ( .A1(n12424), .A2(n10655), .B1(n2886), .B2(n12416), .ZN(
        n9104) );
  OAI22_X1 U5911 ( .A1(n12424), .A2(n10648), .B1(n2885), .B2(n12416), .ZN(
        n9103) );
  OAI22_X1 U5912 ( .A1(n12424), .A2(n10641), .B1(n2884), .B2(n12416), .ZN(
        n9102) );
  OAI22_X1 U5913 ( .A1(n12425), .A2(n10634), .B1(n2883), .B2(n12416), .ZN(
        n9101) );
  OAI22_X1 U5914 ( .A1(n12425), .A2(n10627), .B1(n2882), .B2(n12416), .ZN(
        n9100) );
  INV_X1 U5915 ( .A(RETRN), .ZN(n14518) );
  NAND2_X1 U5916 ( .A1(\U3/U98/Z_5 ), .A2(\r480/carry[5] ), .ZN(\r480/n4 ) );
  NOR2_X1 U5917 ( .A1(n2935), .A2(\r480/A[3] ), .ZN(\U3/U98/Z_6 ) );
  NAND2_X1 U5918 ( .A1(\U3/U99/Z_5 ), .A2(\r486/carry[5] ), .ZN(\r486/n4 ) );
  NOR2_X1 U5919 ( .A1(n2935), .A2(\r486/A[3] ), .ZN(\U3/U99/Z_6 ) );
  NOR2_X2 U5920 ( .A1(N8432), .A2(N8433), .ZN(n5647) );
  NOR2_X2 U5921 ( .A1(N8576), .A2(N8577), .ZN(n4214) );
  NOR2_X2 U5922 ( .A1(n14513), .A2(N8433), .ZN(n5649) );
  NOR2_X2 U5923 ( .A1(n14515), .A2(N8577), .ZN(n4216) );
  NOR3_X1 U5924 ( .A1(n12769), .A2(N8431), .A3(n12771), .ZN(n5705) );
  NOR3_X1 U5925 ( .A1(n12773), .A2(N8575), .A3(n12775), .ZN(n4272) );
  AOI222_X1 U5926 ( .A1(n10998), .A2(n9728), .B1(n10995), .B2(n9664), .C1(
        n10992), .C2(n13363), .ZN(n5667) );
  AOI222_X1 U5927 ( .A1(n10932), .A2(n9280), .B1(n10929), .B2(n9216), .C1(
        n10926), .C2(n13811), .ZN(n5680) );
  AOI222_X1 U5928 ( .A1(n11262), .A2(n9728), .B1(n11259), .B2(n9664), .C1(
        n11256), .C2(n13363), .ZN(n4234) );
  AOI222_X1 U5929 ( .A1(n11196), .A2(n9280), .B1(n11193), .B2(n9216), .C1(
        n11190), .C2(n13811), .ZN(n4247) );
  AOI222_X1 U5930 ( .A1(n10998), .A2(n9729), .B1(n10995), .B2(n9665), .C1(
        n10992), .C2(n13362), .ZN(n5607) );
  AOI222_X1 U5931 ( .A1(n10932), .A2(n9281), .B1(n10929), .B2(n9217), .C1(
        n10926), .C2(n13810), .ZN(n5616) );
  AOI222_X1 U5932 ( .A1(n11262), .A2(n9729), .B1(n11259), .B2(n9665), .C1(
        n11256), .C2(n13362), .ZN(n4174) );
  AOI222_X1 U5933 ( .A1(n11196), .A2(n9281), .B1(n11193), .B2(n9217), .C1(
        n11190), .C2(n13810), .ZN(n4183) );
  AOI222_X1 U5934 ( .A1(n10998), .A2(n9730), .B1(n10995), .B2(n9666), .C1(
        n10992), .C2(n13361), .ZN(n5566) );
  AOI222_X1 U5935 ( .A1(n10932), .A2(n9282), .B1(n10929), .B2(n9218), .C1(
        n10926), .C2(n13809), .ZN(n5575) );
  AOI222_X1 U5936 ( .A1(n11262), .A2(n9730), .B1(n11259), .B2(n9666), .C1(
        n11256), .C2(n13361), .ZN(n4133) );
  AOI222_X1 U5937 ( .A1(n11196), .A2(n9282), .B1(n11193), .B2(n9218), .C1(
        n11190), .C2(n13809), .ZN(n4142) );
  AOI222_X1 U5938 ( .A1(n10998), .A2(n9731), .B1(n10995), .B2(n9667), .C1(
        n10992), .C2(n13360), .ZN(n5525) );
  AOI222_X1 U5939 ( .A1(n10932), .A2(n9283), .B1(n10929), .B2(n9219), .C1(
        n10926), .C2(n13808), .ZN(n5534) );
  AOI222_X1 U5940 ( .A1(n11262), .A2(n9731), .B1(n11259), .B2(n9667), .C1(
        n11256), .C2(n13360), .ZN(n4092) );
  AOI222_X1 U5941 ( .A1(n11196), .A2(n9283), .B1(n11193), .B2(n9219), .C1(
        n11190), .C2(n13808), .ZN(n4101) );
  AOI222_X1 U5942 ( .A1(n10998), .A2(n9732), .B1(n10995), .B2(n9668), .C1(
        n10992), .C2(n13359), .ZN(n5484) );
  AOI222_X1 U5943 ( .A1(n10932), .A2(n9284), .B1(n10929), .B2(n9220), .C1(
        n10926), .C2(n13807), .ZN(n5493) );
  AOI222_X1 U5944 ( .A1(n11262), .A2(n9732), .B1(n11259), .B2(n9668), .C1(
        n11256), .C2(n13359), .ZN(n4051) );
  AOI222_X1 U5945 ( .A1(n11196), .A2(n9284), .B1(n11193), .B2(n9220), .C1(
        n11190), .C2(n13807), .ZN(n4060) );
  AOI222_X1 U5946 ( .A1(n10998), .A2(n9733), .B1(n10995), .B2(n9669), .C1(
        n10992), .C2(n13358), .ZN(n5443) );
  AOI222_X1 U5947 ( .A1(n10932), .A2(n9285), .B1(n10929), .B2(n9221), .C1(
        n10926), .C2(n13806), .ZN(n5452) );
  AOI222_X1 U5948 ( .A1(n11262), .A2(n9733), .B1(n11259), .B2(n9669), .C1(
        n11256), .C2(n13358), .ZN(n4010) );
  AOI222_X1 U5949 ( .A1(n11196), .A2(n9285), .B1(n11193), .B2(n9221), .C1(
        n11190), .C2(n13806), .ZN(n4019) );
  AOI222_X1 U5950 ( .A1(n10998), .A2(n9734), .B1(n10995), .B2(n9670), .C1(
        n10992), .C2(n9702), .ZN(n5402) );
  AOI222_X1 U5951 ( .A1(n10932), .A2(n9286), .B1(n10929), .B2(n9222), .C1(
        n10926), .C2(n13805), .ZN(n5411) );
  AOI222_X1 U5952 ( .A1(n11262), .A2(n9734), .B1(n11259), .B2(n9670), .C1(
        n11256), .C2(n9702), .ZN(n3969) );
  AOI222_X1 U5953 ( .A1(n11196), .A2(n9286), .B1(n11193), .B2(n9222), .C1(
        n11190), .C2(n13805), .ZN(n3978) );
  AOI222_X1 U5954 ( .A1(n10998), .A2(n9735), .B1(n10995), .B2(n9671), .C1(
        n10992), .C2(n9703), .ZN(n5361) );
  AOI222_X1 U5955 ( .A1(n10932), .A2(n9287), .B1(n10929), .B2(n9223), .C1(
        n10926), .C2(n13804), .ZN(n5370) );
  AOI222_X1 U5956 ( .A1(n11262), .A2(n9735), .B1(n11259), .B2(n9671), .C1(
        n11256), .C2(n9703), .ZN(n3928) );
  AOI222_X1 U5957 ( .A1(n11196), .A2(n9287), .B1(n11193), .B2(n9223), .C1(
        n11190), .C2(n13804), .ZN(n3937) );
  AOI222_X1 U5958 ( .A1(n10998), .A2(n9736), .B1(n10995), .B2(n9672), .C1(
        n10992), .C2(n9704), .ZN(n5320) );
  AOI222_X1 U5959 ( .A1(n10932), .A2(n9288), .B1(n10929), .B2(n9224), .C1(
        n10926), .C2(n13803), .ZN(n5329) );
  AOI222_X1 U5960 ( .A1(n11262), .A2(n9736), .B1(n11259), .B2(n9672), .C1(
        n11256), .C2(n9704), .ZN(n3887) );
  AOI222_X1 U5961 ( .A1(n11196), .A2(n9288), .B1(n11193), .B2(n9224), .C1(
        n11190), .C2(n13803), .ZN(n3896) );
  AOI222_X1 U5962 ( .A1(n10998), .A2(n9737), .B1(n10995), .B2(n9673), .C1(
        n10992), .C2(n9705), .ZN(n5279) );
  AOI222_X1 U5963 ( .A1(n10932), .A2(n9289), .B1(n10929), .B2(n9225), .C1(
        n10926), .C2(n13802), .ZN(n5288) );
  AOI222_X1 U5964 ( .A1(n11262), .A2(n9737), .B1(n11259), .B2(n9673), .C1(
        n11256), .C2(n9705), .ZN(n3846) );
  AOI222_X1 U5965 ( .A1(n11196), .A2(n9289), .B1(n11193), .B2(n9225), .C1(
        n11190), .C2(n13802), .ZN(n3855) );
  AOI222_X1 U5966 ( .A1(n10998), .A2(n9738), .B1(n10995), .B2(n9674), .C1(
        n10992), .C2(n9706), .ZN(n5238) );
  AOI222_X1 U5967 ( .A1(n10932), .A2(n9290), .B1(n10929), .B2(n9226), .C1(
        n10926), .C2(n13801), .ZN(n5247) );
  AOI222_X1 U5968 ( .A1(n11262), .A2(n9738), .B1(n11259), .B2(n9674), .C1(
        n11256), .C2(n9706), .ZN(n3805) );
  AOI222_X1 U5969 ( .A1(n11196), .A2(n9290), .B1(n11193), .B2(n9226), .C1(
        n11190), .C2(n13801), .ZN(n3814) );
  AOI222_X1 U5970 ( .A1(n10998), .A2(n9739), .B1(n10995), .B2(n9675), .C1(
        n10992), .C2(n9707), .ZN(n5197) );
  AOI222_X1 U5971 ( .A1(n10932), .A2(n9291), .B1(n10929), .B2(n9227), .C1(
        n10926), .C2(n13800), .ZN(n5206) );
  AOI222_X1 U5972 ( .A1(n11262), .A2(n9739), .B1(n11259), .B2(n9675), .C1(
        n11256), .C2(n9707), .ZN(n3764) );
  AOI222_X1 U5973 ( .A1(n11196), .A2(n9291), .B1(n11193), .B2(n9227), .C1(
        n11190), .C2(n13800), .ZN(n3773) );
  AOI222_X1 U5974 ( .A1(n10999), .A2(n9740), .B1(n10996), .B2(n9676), .C1(
        n10993), .C2(n9708), .ZN(n5156) );
  AOI222_X1 U5975 ( .A1(n10933), .A2(n9292), .B1(n10930), .B2(n9228), .C1(
        n10927), .C2(n13799), .ZN(n5165) );
  AOI222_X1 U5976 ( .A1(n11263), .A2(n9740), .B1(n11260), .B2(n9676), .C1(
        n11257), .C2(n9708), .ZN(n3723) );
  AOI222_X1 U5977 ( .A1(n11197), .A2(n9292), .B1(n11194), .B2(n9228), .C1(
        n11191), .C2(n13799), .ZN(n3732) );
  AOI222_X1 U5978 ( .A1(n10999), .A2(n9741), .B1(n10996), .B2(n9677), .C1(
        n10993), .C2(n9709), .ZN(n5115) );
  AOI222_X1 U5979 ( .A1(n10933), .A2(n9293), .B1(n10930), .B2(n9229), .C1(
        n10927), .C2(n13798), .ZN(n5124) );
  AOI222_X1 U5980 ( .A1(n11263), .A2(n9741), .B1(n11260), .B2(n9677), .C1(
        n11257), .C2(n9709), .ZN(n3682) );
  AOI222_X1 U5981 ( .A1(n11197), .A2(n9293), .B1(n11194), .B2(n9229), .C1(
        n11191), .C2(n13798), .ZN(n3691) );
  AOI222_X1 U5982 ( .A1(n10999), .A2(n9742), .B1(n10996), .B2(n9678), .C1(
        n10993), .C2(n9710), .ZN(n5074) );
  AOI222_X1 U5983 ( .A1(n10933), .A2(n9294), .B1(n10930), .B2(n9230), .C1(
        n10927), .C2(n13797), .ZN(n5083) );
  AOI222_X1 U5984 ( .A1(n11263), .A2(n9742), .B1(n11260), .B2(n9678), .C1(
        n11257), .C2(n9710), .ZN(n3641) );
  AOI222_X1 U5985 ( .A1(n11197), .A2(n9294), .B1(n11194), .B2(n9230), .C1(
        n11191), .C2(n13797), .ZN(n3650) );
  AOI222_X1 U5986 ( .A1(n10999), .A2(n9743), .B1(n10996), .B2(n9679), .C1(
        n10993), .C2(n9711), .ZN(n5033) );
  AOI222_X1 U5987 ( .A1(n10933), .A2(n9295), .B1(n10930), .B2(n9231), .C1(
        n10927), .C2(n13796), .ZN(n5042) );
  AOI222_X1 U5988 ( .A1(n11263), .A2(n9743), .B1(n11260), .B2(n9679), .C1(
        n11257), .C2(n9711), .ZN(n3600) );
  AOI222_X1 U5989 ( .A1(n11197), .A2(n9295), .B1(n11194), .B2(n9231), .C1(
        n11191), .C2(n13796), .ZN(n3609) );
  AOI222_X1 U5990 ( .A1(n10999), .A2(n9744), .B1(n10996), .B2(n9680), .C1(
        n10993), .C2(n9712), .ZN(n4992) );
  AOI222_X1 U5991 ( .A1(n10933), .A2(n9296), .B1(n10930), .B2(n9232), .C1(
        n10927), .C2(n13795), .ZN(n5001) );
  AOI222_X1 U5992 ( .A1(n11263), .A2(n9744), .B1(n11260), .B2(n9680), .C1(
        n11257), .C2(n9712), .ZN(n3559) );
  AOI222_X1 U5993 ( .A1(n11197), .A2(n9296), .B1(n11194), .B2(n9232), .C1(
        n11191), .C2(n13795), .ZN(n3568) );
  AOI222_X1 U5994 ( .A1(n10999), .A2(n9745), .B1(n10996), .B2(n9681), .C1(
        n10993), .C2(n9713), .ZN(n4951) );
  AOI222_X1 U5995 ( .A1(n10933), .A2(n9297), .B1(n10930), .B2(n9233), .C1(
        n10927), .C2(n9265), .ZN(n4960) );
  AOI222_X1 U5996 ( .A1(n11263), .A2(n9745), .B1(n11260), .B2(n9681), .C1(
        n11257), .C2(n9713), .ZN(n3518) );
  AOI222_X1 U5997 ( .A1(n11197), .A2(n9297), .B1(n11194), .B2(n9233), .C1(
        n11191), .C2(n9265), .ZN(n3527) );
  AOI222_X1 U5998 ( .A1(n10999), .A2(n9746), .B1(n10996), .B2(n9682), .C1(
        n10993), .C2(n9714), .ZN(n4910) );
  AOI222_X1 U5999 ( .A1(n10933), .A2(n9298), .B1(n10930), .B2(n9234), .C1(
        n10927), .C2(n9266), .ZN(n4919) );
  AOI222_X1 U6000 ( .A1(n11263), .A2(n9746), .B1(n11260), .B2(n9682), .C1(
        n11257), .C2(n9714), .ZN(n3477) );
  AOI222_X1 U6001 ( .A1(n11197), .A2(n9298), .B1(n11194), .B2(n9234), .C1(
        n11191), .C2(n9266), .ZN(n3486) );
  AOI222_X1 U6002 ( .A1(n10999), .A2(n9747), .B1(n10996), .B2(n9683), .C1(
        n10993), .C2(n9715), .ZN(n4869) );
  AOI222_X1 U6003 ( .A1(n10933), .A2(n9299), .B1(n10930), .B2(n9235), .C1(
        n10927), .C2(n9267), .ZN(n4878) );
  AOI222_X1 U6004 ( .A1(n11263), .A2(n9747), .B1(n11260), .B2(n9683), .C1(
        n11257), .C2(n9715), .ZN(n3436) );
  AOI222_X1 U6005 ( .A1(n11197), .A2(n9299), .B1(n11194), .B2(n9235), .C1(
        n11191), .C2(n9267), .ZN(n3445) );
  AOI222_X1 U6006 ( .A1(n10999), .A2(n9748), .B1(n10996), .B2(n9684), .C1(
        n10993), .C2(n9716), .ZN(n4828) );
  AOI222_X1 U6007 ( .A1(n10933), .A2(n9300), .B1(n10930), .B2(n9236), .C1(
        n10927), .C2(n9268), .ZN(n4837) );
  AOI222_X1 U6008 ( .A1(n11263), .A2(n9748), .B1(n11260), .B2(n9684), .C1(
        n11257), .C2(n9716), .ZN(n3395) );
  AOI222_X1 U6009 ( .A1(n11197), .A2(n9300), .B1(n11194), .B2(n9236), .C1(
        n11191), .C2(n9268), .ZN(n3404) );
  AOI222_X1 U6010 ( .A1(n10999), .A2(n9749), .B1(n10996), .B2(n9685), .C1(
        n10993), .C2(n9717), .ZN(n4787) );
  AOI222_X1 U6011 ( .A1(n10933), .A2(n9301), .B1(n10930), .B2(n9237), .C1(
        n10927), .C2(n9269), .ZN(n4796) );
  AOI222_X1 U6012 ( .A1(n11263), .A2(n9749), .B1(n11260), .B2(n9685), .C1(
        n11257), .C2(n9717), .ZN(n3354) );
  AOI222_X1 U6013 ( .A1(n11197), .A2(n9301), .B1(n11194), .B2(n9237), .C1(
        n11191), .C2(n9269), .ZN(n3363) );
  AOI222_X1 U6014 ( .A1(n10999), .A2(n9750), .B1(n10996), .B2(n9686), .C1(
        n10993), .C2(n9718), .ZN(n4746) );
  AOI222_X1 U6015 ( .A1(n10933), .A2(n9302), .B1(n10930), .B2(n9238), .C1(
        n10927), .C2(n9270), .ZN(n4755) );
  AOI222_X1 U6016 ( .A1(n11263), .A2(n9750), .B1(n11260), .B2(n9686), .C1(
        n11257), .C2(n9718), .ZN(n3313) );
  AOI222_X1 U6017 ( .A1(n11197), .A2(n9302), .B1(n11194), .B2(n9238), .C1(
        n11191), .C2(n9270), .ZN(n3322) );
  AOI222_X1 U6018 ( .A1(n10999), .A2(n9751), .B1(n10996), .B2(n9687), .C1(
        n10993), .C2(n9719), .ZN(n4705) );
  AOI222_X1 U6019 ( .A1(n10933), .A2(n9303), .B1(n10930), .B2(n9239), .C1(
        n10927), .C2(n9271), .ZN(n4714) );
  AOI222_X1 U6020 ( .A1(n11263), .A2(n9751), .B1(n11260), .B2(n9687), .C1(
        n11257), .C2(n9719), .ZN(n3272) );
  AOI222_X1 U6021 ( .A1(n11197), .A2(n9303), .B1(n11194), .B2(n9239), .C1(
        n11191), .C2(n9271), .ZN(n3281) );
  AOI222_X1 U6022 ( .A1(n11000), .A2(n9752), .B1(n10997), .B2(n9688), .C1(
        n10994), .C2(n9720), .ZN(n4664) );
  AOI222_X1 U6023 ( .A1(n10934), .A2(n9304), .B1(n10931), .B2(n9240), .C1(
        n10928), .C2(n9272), .ZN(n4673) );
  AOI222_X1 U6024 ( .A1(n11264), .A2(n9752), .B1(n11261), .B2(n9688), .C1(
        n11258), .C2(n9720), .ZN(n3231) );
  AOI222_X1 U6025 ( .A1(n11198), .A2(n9304), .B1(n11195), .B2(n9240), .C1(
        n11192), .C2(n9272), .ZN(n3240) );
  AOI222_X1 U6026 ( .A1(n11000), .A2(n9753), .B1(n10997), .B2(n9689), .C1(
        n10994), .C2(n9721), .ZN(n4623) );
  AOI222_X1 U6027 ( .A1(n10934), .A2(n9305), .B1(n10931), .B2(n9241), .C1(
        n10928), .C2(n9273), .ZN(n4632) );
  AOI222_X1 U6028 ( .A1(n11264), .A2(n9753), .B1(n11261), .B2(n9689), .C1(
        n11258), .C2(n9721), .ZN(n3190) );
  AOI222_X1 U6029 ( .A1(n11198), .A2(n9305), .B1(n11195), .B2(n9241), .C1(
        n11192), .C2(n9273), .ZN(n3199) );
  AOI222_X1 U6030 ( .A1(n11000), .A2(n9754), .B1(n10997), .B2(n9690), .C1(
        n10994), .C2(n9722), .ZN(n4582) );
  AOI222_X1 U6031 ( .A1(n10934), .A2(n9306), .B1(n10931), .B2(n9242), .C1(
        n10928), .C2(n9274), .ZN(n4591) );
  AOI222_X1 U6032 ( .A1(n11264), .A2(n9754), .B1(n11261), .B2(n9690), .C1(
        n11258), .C2(n9722), .ZN(n3149) );
  AOI222_X1 U6033 ( .A1(n11198), .A2(n9306), .B1(n11195), .B2(n9242), .C1(
        n11192), .C2(n9274), .ZN(n3158) );
  AOI222_X1 U6034 ( .A1(n11000), .A2(n9755), .B1(n10997), .B2(n9691), .C1(
        n10994), .C2(n9723), .ZN(n4541) );
  AOI222_X1 U6035 ( .A1(n10934), .A2(n9307), .B1(n10931), .B2(n9243), .C1(
        n10928), .C2(n9275), .ZN(n4550) );
  AOI222_X1 U6036 ( .A1(n11264), .A2(n9755), .B1(n11261), .B2(n9691), .C1(
        n11258), .C2(n9723), .ZN(n3108) );
  AOI222_X1 U6037 ( .A1(n11198), .A2(n9307), .B1(n11195), .B2(n9243), .C1(
        n11192), .C2(n9275), .ZN(n3117) );
  AOI222_X1 U6038 ( .A1(n11000), .A2(n9756), .B1(n10997), .B2(n9692), .C1(
        n10994), .C2(n9724), .ZN(n4500) );
  AOI222_X1 U6039 ( .A1(n10934), .A2(n9308), .B1(n10931), .B2(n9244), .C1(
        n10928), .C2(n9276), .ZN(n4509) );
  AOI222_X1 U6040 ( .A1(n11264), .A2(n9756), .B1(n11261), .B2(n9692), .C1(
        n11258), .C2(n9724), .ZN(n3067) );
  AOI222_X1 U6041 ( .A1(n11198), .A2(n9308), .B1(n11195), .B2(n9244), .C1(
        n11192), .C2(n9276), .ZN(n3076) );
  AOI222_X1 U6042 ( .A1(n11000), .A2(n9757), .B1(n10997), .B2(n9693), .C1(
        n10994), .C2(n9725), .ZN(n4459) );
  AOI222_X1 U6043 ( .A1(n10934), .A2(n9309), .B1(n10931), .B2(n9245), .C1(
        n10928), .C2(n9277), .ZN(n4468) );
  AOI222_X1 U6044 ( .A1(n11264), .A2(n9757), .B1(n11261), .B2(n9693), .C1(
        n11258), .C2(n9725), .ZN(n3026) );
  AOI222_X1 U6045 ( .A1(n11198), .A2(n9309), .B1(n11195), .B2(n9245), .C1(
        n11192), .C2(n9277), .ZN(n3035) );
  AOI222_X1 U6046 ( .A1(n11000), .A2(n9758), .B1(n10997), .B2(n9694), .C1(
        n10994), .C2(n9726), .ZN(n4418) );
  AOI222_X1 U6047 ( .A1(n10934), .A2(n9310), .B1(n10931), .B2(n9246), .C1(
        n10928), .C2(n9278), .ZN(n4427) );
  AOI222_X1 U6048 ( .A1(n11264), .A2(n9758), .B1(n11261), .B2(n9694), .C1(
        n11258), .C2(n9726), .ZN(n2985) );
  AOI222_X1 U6049 ( .A1(n11198), .A2(n9310), .B1(n11195), .B2(n9246), .C1(
        n11192), .C2(n9278), .ZN(n2994) );
  AOI222_X1 U6050 ( .A1(n11000), .A2(n9759), .B1(n10997), .B2(n9695), .C1(
        n10994), .C2(n9727), .ZN(n4311) );
  AOI222_X1 U6051 ( .A1(n10934), .A2(n13748), .B1(n10931), .B2(n9247), .C1(
        n10928), .C2(n9279), .ZN(n4342) );
  AOI222_X1 U6052 ( .A1(n11264), .A2(n9759), .B1(n11261), .B2(n9695), .C1(
        n11258), .C2(n9727), .ZN(n2811) );
  AOI222_X1 U6053 ( .A1(n11198), .A2(n13748), .B1(n11195), .B2(n9247), .C1(
        n11192), .C2(n9279), .ZN(n2874) );
  OAI222_X1 U6054 ( .A1(n2338), .A2(n11106), .B1(n514), .B2(n11103), .C1(n1443), .C2(n11100), .ZN(n5644) );
  OAI222_X1 U6055 ( .A1(n10526), .A2(n11040), .B1(n10525), .B2(n11037), .C1(
        n10527), .C2(n11034), .ZN(n5672) );
  OAI222_X1 U6056 ( .A1(n10518), .A2(n10974), .B1(n10517), .B2(n10971), .C1(
        n10519), .C2(n10968), .ZN(n5685) );
  OAI222_X1 U6057 ( .A1(n2338), .A2(n11370), .B1(n514), .B2(n11367), .C1(n1443), .C2(n11364), .ZN(n4211) );
  OAI222_X1 U6058 ( .A1(n10526), .A2(n11304), .B1(n10525), .B2(n11301), .C1(
        n10527), .C2(n11298), .ZN(n4239) );
  OAI222_X1 U6059 ( .A1(n10518), .A2(n11238), .B1(n10517), .B2(n11235), .C1(
        n10519), .C2(n11232), .ZN(n4252) );
  OAI222_X1 U6060 ( .A1(n2326), .A2(n11106), .B1(n502), .B2(n11103), .C1(n1399), .C2(n11100), .ZN(n5603) );
  OAI222_X1 U6061 ( .A1(n10494), .A2(n11040), .B1(n10493), .B2(n11037), .C1(
        n10495), .C2(n11034), .ZN(n5612) );
  OAI222_X1 U6062 ( .A1(n10486), .A2(n10974), .B1(n10485), .B2(n10971), .C1(
        n10487), .C2(n10968), .ZN(n5621) );
  OAI222_X1 U6063 ( .A1(n2326), .A2(n11370), .B1(n502), .B2(n11367), .C1(n1399), .C2(n11364), .ZN(n4170) );
  OAI222_X1 U6064 ( .A1(n10494), .A2(n11304), .B1(n10493), .B2(n11301), .C1(
        n10495), .C2(n11298), .ZN(n4179) );
  OAI222_X1 U6065 ( .A1(n10486), .A2(n11238), .B1(n10485), .B2(n11235), .C1(
        n10487), .C2(n11232), .ZN(n4188) );
  OAI222_X1 U6066 ( .A1(n2314), .A2(n11106), .B1(n490), .B2(n11103), .C1(n1387), .C2(n11100), .ZN(n5562) );
  OAI222_X1 U6067 ( .A1(n10462), .A2(n11040), .B1(n10461), .B2(n11037), .C1(
        n10463), .C2(n11034), .ZN(n5571) );
  OAI222_X1 U6068 ( .A1(n10454), .A2(n10974), .B1(n10453), .B2(n10971), .C1(
        n10455), .C2(n10968), .ZN(n5580) );
  OAI222_X1 U6069 ( .A1(n2314), .A2(n11370), .B1(n490), .B2(n11367), .C1(n1387), .C2(n11364), .ZN(n4129) );
  OAI222_X1 U6070 ( .A1(n10462), .A2(n11304), .B1(n10461), .B2(n11301), .C1(
        n10463), .C2(n11298), .ZN(n4138) );
  OAI222_X1 U6071 ( .A1(n10454), .A2(n11238), .B1(n10453), .B2(n11235), .C1(
        n10455), .C2(n11232), .ZN(n4147) );
  OAI222_X1 U6072 ( .A1(n2302), .A2(n11106), .B1(n478), .B2(n11103), .C1(n1343), .C2(n11100), .ZN(n5521) );
  OAI222_X1 U6073 ( .A1(n10430), .A2(n11040), .B1(n10429), .B2(n11037), .C1(
        n10431), .C2(n11034), .ZN(n5530) );
  OAI222_X1 U6074 ( .A1(n10422), .A2(n10974), .B1(n10421), .B2(n10971), .C1(
        n10423), .C2(n10968), .ZN(n5539) );
  OAI222_X1 U6075 ( .A1(n2302), .A2(n11370), .B1(n478), .B2(n11367), .C1(n1343), .C2(n11364), .ZN(n4088) );
  OAI222_X1 U6076 ( .A1(n10430), .A2(n11304), .B1(n10429), .B2(n11301), .C1(
        n10431), .C2(n11298), .ZN(n4097) );
  OAI222_X1 U6077 ( .A1(n10422), .A2(n11238), .B1(n10421), .B2(n11235), .C1(
        n10423), .C2(n11232), .ZN(n4106) );
  OAI222_X1 U6078 ( .A1(n2290), .A2(n11106), .B1(n466), .B2(n11103), .C1(n1331), .C2(n11100), .ZN(n5480) );
  OAI222_X1 U6079 ( .A1(n10395), .A2(n11040), .B1(n10394), .B2(n11037), .C1(
        n10396), .C2(n11034), .ZN(n5489) );
  OAI222_X1 U6080 ( .A1(n10387), .A2(n10974), .B1(n10386), .B2(n10971), .C1(
        n10388), .C2(n10968), .ZN(n5498) );
  OAI222_X1 U6081 ( .A1(n2290), .A2(n11370), .B1(n466), .B2(n11367), .C1(n1331), .C2(n11364), .ZN(n4047) );
  OAI222_X1 U6082 ( .A1(n10395), .A2(n11304), .B1(n10394), .B2(n11301), .C1(
        n10396), .C2(n11298), .ZN(n4056) );
  OAI222_X1 U6083 ( .A1(n10387), .A2(n11238), .B1(n10386), .B2(n11235), .C1(
        n10388), .C2(n11232), .ZN(n4065) );
  OAI222_X1 U6084 ( .A1(n2278), .A2(n11106), .B1(n454), .B2(n11103), .C1(n1319), .C2(n11100), .ZN(n5439) );
  OAI222_X1 U6085 ( .A1(n10363), .A2(n11040), .B1(n10362), .B2(n11037), .C1(
        n10364), .C2(n11034), .ZN(n5448) );
  OAI222_X1 U6086 ( .A1(n10355), .A2(n10974), .B1(n10354), .B2(n10971), .C1(
        n10356), .C2(n10968), .ZN(n5457) );
  OAI222_X1 U6087 ( .A1(n2278), .A2(n11370), .B1(n454), .B2(n11367), .C1(n1319), .C2(n11364), .ZN(n4006) );
  OAI222_X1 U6088 ( .A1(n10363), .A2(n11304), .B1(n10362), .B2(n11301), .C1(
        n10364), .C2(n11298), .ZN(n4015) );
  OAI222_X1 U6089 ( .A1(n10355), .A2(n11238), .B1(n10354), .B2(n11235), .C1(
        n10356), .C2(n11232), .ZN(n4024) );
  OAI222_X1 U6090 ( .A1(n2266), .A2(n11106), .B1(n442), .B2(n11103), .C1(n1307), .C2(n11100), .ZN(n5398) );
  OAI222_X1 U6091 ( .A1(n10331), .A2(n11040), .B1(n10330), .B2(n11037), .C1(
        n10332), .C2(n11034), .ZN(n5407) );
  OAI222_X1 U6092 ( .A1(n10323), .A2(n10974), .B1(n10322), .B2(n10971), .C1(
        n10324), .C2(n10968), .ZN(n5416) );
  OAI222_X1 U6093 ( .A1(n2266), .A2(n11370), .B1(n442), .B2(n11367), .C1(n1307), .C2(n11364), .ZN(n3965) );
  OAI222_X1 U6094 ( .A1(n10331), .A2(n11304), .B1(n10330), .B2(n11301), .C1(
        n10332), .C2(n11298), .ZN(n3974) );
  OAI222_X1 U6095 ( .A1(n10323), .A2(n11238), .B1(n10322), .B2(n11235), .C1(
        n10324), .C2(n11232), .ZN(n3983) );
  OAI222_X1 U6096 ( .A1(n2254), .A2(n11106), .B1(n430), .B2(n11103), .C1(n1295), .C2(n11100), .ZN(n5357) );
  OAI222_X1 U6097 ( .A1(n10296), .A2(n11040), .B1(n10295), .B2(n11037), .C1(
        n10297), .C2(n11034), .ZN(n5366) );
  OAI222_X1 U6098 ( .A1(n10288), .A2(n10974), .B1(n10287), .B2(n10971), .C1(
        n10289), .C2(n10968), .ZN(n5375) );
  OAI222_X1 U6099 ( .A1(n2254), .A2(n11370), .B1(n430), .B2(n11367), .C1(n1295), .C2(n11364), .ZN(n3924) );
  OAI222_X1 U6100 ( .A1(n10296), .A2(n11304), .B1(n10295), .B2(n11301), .C1(
        n10297), .C2(n11298), .ZN(n3933) );
  OAI222_X1 U6101 ( .A1(n10288), .A2(n11238), .B1(n10287), .B2(n11235), .C1(
        n10289), .C2(n11232), .ZN(n3942) );
  OAI222_X1 U6102 ( .A1(n2242), .A2(n11106), .B1(n418), .B2(n11103), .C1(n1283), .C2(n11100), .ZN(n5316) );
  OAI222_X1 U6103 ( .A1(n10264), .A2(n11040), .B1(n10263), .B2(n11037), .C1(
        n10265), .C2(n11034), .ZN(n5325) );
  OAI222_X1 U6104 ( .A1(n10256), .A2(n10974), .B1(n10255), .B2(n10971), .C1(
        n10257), .C2(n10968), .ZN(n5334) );
  OAI222_X1 U6105 ( .A1(n2242), .A2(n11370), .B1(n418), .B2(n11367), .C1(n1283), .C2(n11364), .ZN(n3883) );
  OAI222_X1 U6106 ( .A1(n10264), .A2(n11304), .B1(n10263), .B2(n11301), .C1(
        n10265), .C2(n11298), .ZN(n3892) );
  OAI222_X1 U6107 ( .A1(n10256), .A2(n11238), .B1(n10255), .B2(n11235), .C1(
        n10257), .C2(n11232), .ZN(n3901) );
  OAI222_X1 U6108 ( .A1(n2230), .A2(n11106), .B1(n406), .B2(n11103), .C1(n1271), .C2(n11100), .ZN(n5275) );
  OAI222_X1 U6109 ( .A1(n10232), .A2(n11040), .B1(n10231), .B2(n11037), .C1(
        n10233), .C2(n11034), .ZN(n5284) );
  OAI222_X1 U6110 ( .A1(n10224), .A2(n10974), .B1(n10223), .B2(n10971), .C1(
        n10225), .C2(n10968), .ZN(n5293) );
  OAI222_X1 U6111 ( .A1(n2230), .A2(n11370), .B1(n406), .B2(n11367), .C1(n1271), .C2(n11364), .ZN(n3842) );
  OAI222_X1 U6112 ( .A1(n10232), .A2(n11304), .B1(n10231), .B2(n11301), .C1(
        n10233), .C2(n11298), .ZN(n3851) );
  OAI222_X1 U6113 ( .A1(n10224), .A2(n11238), .B1(n10223), .B2(n11235), .C1(
        n10225), .C2(n11232), .ZN(n3860) );
  OAI222_X1 U6114 ( .A1(n2218), .A2(n11106), .B1(n394), .B2(n11103), .C1(n1259), .C2(n11100), .ZN(n5234) );
  OAI222_X1 U6115 ( .A1(n10198), .A2(n11040), .B1(n10197), .B2(n11037), .C1(
        n10199), .C2(n11034), .ZN(n5243) );
  OAI222_X1 U6116 ( .A1(n10190), .A2(n10974), .B1(n10189), .B2(n10971), .C1(
        n10191), .C2(n10968), .ZN(n5252) );
  OAI222_X1 U6117 ( .A1(n2218), .A2(n11370), .B1(n394), .B2(n11367), .C1(n1259), .C2(n11364), .ZN(n3801) );
  OAI222_X1 U6118 ( .A1(n10198), .A2(n11304), .B1(n10197), .B2(n11301), .C1(
        n10199), .C2(n11298), .ZN(n3810) );
  OAI222_X1 U6119 ( .A1(n10190), .A2(n11238), .B1(n10189), .B2(n11235), .C1(
        n10191), .C2(n11232), .ZN(n3819) );
  OAI222_X1 U6120 ( .A1(n2174), .A2(n11106), .B1(n382), .B2(n11103), .C1(n1247), .C2(n11100), .ZN(n5193) );
  OAI222_X1 U6121 ( .A1(n10166), .A2(n11040), .B1(n10165), .B2(n11037), .C1(
        n10167), .C2(n11034), .ZN(n5202) );
  OAI222_X1 U6122 ( .A1(n10158), .A2(n10974), .B1(n10157), .B2(n10971), .C1(
        n10159), .C2(n10968), .ZN(n5211) );
  OAI222_X1 U6123 ( .A1(n2174), .A2(n11370), .B1(n382), .B2(n11367), .C1(n1247), .C2(n11364), .ZN(n3760) );
  OAI222_X1 U6124 ( .A1(n10166), .A2(n11304), .B1(n10165), .B2(n11301), .C1(
        n10167), .C2(n11298), .ZN(n3769) );
  OAI222_X1 U6125 ( .A1(n10158), .A2(n11238), .B1(n10157), .B2(n11235), .C1(
        n10159), .C2(n11232), .ZN(n3778) );
  OAI222_X1 U6126 ( .A1(n2162), .A2(n11107), .B1(n370), .B2(n11104), .C1(n1235), .C2(n11101), .ZN(n5152) );
  OAI222_X1 U6127 ( .A1(n10134), .A2(n11041), .B1(n10133), .B2(n11038), .C1(
        n10135), .C2(n11035), .ZN(n5161) );
  OAI222_X1 U6128 ( .A1(n10126), .A2(n10975), .B1(n10125), .B2(n10972), .C1(
        n10127), .C2(n10969), .ZN(n5170) );
  OAI222_X1 U6129 ( .A1(n2162), .A2(n11371), .B1(n370), .B2(n11368), .C1(n1235), .C2(n11365), .ZN(n3719) );
  OAI222_X1 U6130 ( .A1(n10134), .A2(n11305), .B1(n10133), .B2(n11302), .C1(
        n10135), .C2(n11299), .ZN(n3728) );
  OAI222_X1 U6131 ( .A1(n10126), .A2(n11239), .B1(n10125), .B2(n11236), .C1(
        n10127), .C2(n11233), .ZN(n3737) );
  OAI222_X1 U6132 ( .A1(n2150), .A2(n11107), .B1(n358), .B2(n11104), .C1(n1223), .C2(n11101), .ZN(n5111) );
  OAI222_X1 U6133 ( .A1(n10102), .A2(n11041), .B1(n10101), .B2(n11038), .C1(
        n10103), .C2(n11035), .ZN(n5120) );
  OAI222_X1 U6134 ( .A1(n10094), .A2(n10975), .B1(n10093), .B2(n10972), .C1(
        n10095), .C2(n10969), .ZN(n5129) );
  OAI222_X1 U6135 ( .A1(n2150), .A2(n11371), .B1(n358), .B2(n11368), .C1(n1223), .C2(n11365), .ZN(n3678) );
  OAI222_X1 U6136 ( .A1(n10102), .A2(n11305), .B1(n10101), .B2(n11302), .C1(
        n10103), .C2(n11299), .ZN(n3687) );
  OAI222_X1 U6137 ( .A1(n10094), .A2(n11239), .B1(n10093), .B2(n11236), .C1(
        n10095), .C2(n11233), .ZN(n3696) );
  OAI222_X1 U6138 ( .A1(n2106), .A2(n11107), .B1(n346), .B2(n11104), .C1(n1211), .C2(n11101), .ZN(n5070) );
  OAI222_X1 U6139 ( .A1(n10070), .A2(n11041), .B1(n10069), .B2(n11038), .C1(
        n10071), .C2(n11035), .ZN(n5079) );
  OAI222_X1 U6140 ( .A1(n10062), .A2(n10975), .B1(n10061), .B2(n10972), .C1(
        n10063), .C2(n10969), .ZN(n5088) );
  OAI222_X1 U6141 ( .A1(n2106), .A2(n11371), .B1(n346), .B2(n11368), .C1(n1211), .C2(n11365), .ZN(n3637) );
  OAI222_X1 U6142 ( .A1(n10070), .A2(n11305), .B1(n10069), .B2(n11302), .C1(
        n10071), .C2(n11299), .ZN(n3646) );
  OAI222_X1 U6143 ( .A1(n10062), .A2(n11239), .B1(n10061), .B2(n11236), .C1(
        n10063), .C2(n11233), .ZN(n3655) );
  OAI222_X1 U6144 ( .A1(n2094), .A2(n11107), .B1(n334), .B2(n11104), .C1(n1199), .C2(n11101), .ZN(n5029) );
  OAI222_X1 U6145 ( .A1(n10038), .A2(n11041), .B1(n10037), .B2(n11038), .C1(
        n10039), .C2(n11035), .ZN(n5038) );
  OAI222_X1 U6146 ( .A1(n10030), .A2(n10975), .B1(n10029), .B2(n10972), .C1(
        n10031), .C2(n10969), .ZN(n5047) );
  OAI222_X1 U6147 ( .A1(n2094), .A2(n11371), .B1(n334), .B2(n11368), .C1(n1199), .C2(n11365), .ZN(n3596) );
  OAI222_X1 U6148 ( .A1(n10038), .A2(n11305), .B1(n10037), .B2(n11302), .C1(
        n10039), .C2(n11299), .ZN(n3605) );
  OAI222_X1 U6149 ( .A1(n10030), .A2(n11239), .B1(n10029), .B2(n11236), .C1(
        n10031), .C2(n11233), .ZN(n3614) );
  OAI222_X1 U6150 ( .A1(n2082), .A2(n11107), .B1(n322), .B2(n11104), .C1(n1187), .C2(n11101), .ZN(n4988) );
  OAI222_X1 U6151 ( .A1(n10006), .A2(n11041), .B1(n10005), .B2(n11038), .C1(
        n10007), .C2(n11035), .ZN(n4997) );
  OAI222_X1 U6152 ( .A1(n9700), .A2(n10975), .B1(n9699), .B2(n10972), .C1(
        n9701), .C2(n10969), .ZN(n5006) );
  OAI222_X1 U6153 ( .A1(n2082), .A2(n11371), .B1(n322), .B2(n11368), .C1(n1187), .C2(n11365), .ZN(n3555) );
  OAI222_X1 U6154 ( .A1(n10006), .A2(n11305), .B1(n10005), .B2(n11302), .C1(
        n10007), .C2(n11299), .ZN(n3564) );
  OAI222_X1 U6155 ( .A1(n9700), .A2(n11239), .B1(n9699), .B2(n11236), .C1(
        n9701), .C2(n11233), .ZN(n3573) );
  OAI222_X1 U6156 ( .A1(n2038), .A2(n11107), .B1(n310), .B2(n11104), .C1(n1175), .C2(n11101), .ZN(n4947) );
  OAI222_X1 U6157 ( .A1(n9644), .A2(n11041), .B1(n9643), .B2(n11038), .C1(
        n9645), .C2(n11035), .ZN(n4956) );
  OAI222_X1 U6158 ( .A1(n9636), .A2(n10975), .B1(n9635), .B2(n10972), .C1(
        n9637), .C2(n10969), .ZN(n4965) );
  OAI222_X1 U6159 ( .A1(n2038), .A2(n11371), .B1(n310), .B2(n11368), .C1(n1175), .C2(n11365), .ZN(n3514) );
  OAI222_X1 U6160 ( .A1(n9644), .A2(n11305), .B1(n9643), .B2(n11302), .C1(
        n9645), .C2(n11299), .ZN(n3523) );
  OAI222_X1 U6161 ( .A1(n9636), .A2(n11239), .B1(n9635), .B2(n11236), .C1(
        n9637), .C2(n11233), .ZN(n3532) );
  OAI222_X1 U6162 ( .A1(n2026), .A2(n11107), .B1(n298), .B2(n11104), .C1(n1163), .C2(n11101), .ZN(n4906) );
  OAI222_X1 U6163 ( .A1(n9612), .A2(n11041), .B1(n9611), .B2(n11038), .C1(
        n9613), .C2(n11035), .ZN(n4915) );
  OAI222_X1 U6164 ( .A1(n9604), .A2(n10975), .B1(n9603), .B2(n10972), .C1(
        n9605), .C2(n10969), .ZN(n4924) );
  OAI222_X1 U6165 ( .A1(n2026), .A2(n11371), .B1(n298), .B2(n11368), .C1(n1163), .C2(n11365), .ZN(n3473) );
  OAI222_X1 U6166 ( .A1(n9612), .A2(n11305), .B1(n9611), .B2(n11302), .C1(
        n9613), .C2(n11299), .ZN(n3482) );
  OAI222_X1 U6167 ( .A1(n9604), .A2(n11239), .B1(n9603), .B2(n11236), .C1(
        n9605), .C2(n11233), .ZN(n3491) );
  OAI222_X1 U6168 ( .A1(n2014), .A2(n11107), .B1(n286), .B2(n11104), .C1(n1151), .C2(n11101), .ZN(n4865) );
  OAI222_X1 U6169 ( .A1(n9580), .A2(n11041), .B1(n9579), .B2(n11038), .C1(
        n9581), .C2(n11035), .ZN(n4874) );
  OAI222_X1 U6170 ( .A1(n9572), .A2(n10975), .B1(n9571), .B2(n10972), .C1(
        n9573), .C2(n10969), .ZN(n4883) );
  OAI222_X1 U6171 ( .A1(n2014), .A2(n11371), .B1(n286), .B2(n11368), .C1(n1151), .C2(n11365), .ZN(n3432) );
  OAI222_X1 U6172 ( .A1(n9580), .A2(n11305), .B1(n9579), .B2(n11302), .C1(
        n9581), .C2(n11299), .ZN(n3441) );
  OAI222_X1 U6173 ( .A1(n9572), .A2(n11239), .B1(n9571), .B2(n11236), .C1(
        n9573), .C2(n11233), .ZN(n3450) );
  OAI222_X1 U6174 ( .A1(n2002), .A2(n11107), .B1(n274), .B2(n11104), .C1(n1139), .C2(n11101), .ZN(n4824) );
  OAI222_X1 U6175 ( .A1(n9214), .A2(n11041), .B1(n9213), .B2(n11038), .C1(
        n9215), .C2(n11035), .ZN(n4833) );
  OAI222_X1 U6176 ( .A1(n9206), .A2(n10975), .B1(n9205), .B2(n10972), .C1(
        n9207), .C2(n10969), .ZN(n4842) );
  OAI222_X1 U6177 ( .A1(n2002), .A2(n11371), .B1(n274), .B2(n11368), .C1(n1139), .C2(n11365), .ZN(n3391) );
  OAI222_X1 U6178 ( .A1(n9214), .A2(n11305), .B1(n9213), .B2(n11302), .C1(
        n9215), .C2(n11299), .ZN(n3400) );
  OAI222_X1 U6179 ( .A1(n9206), .A2(n11239), .B1(n9205), .B2(n11236), .C1(
        n9207), .C2(n11233), .ZN(n3409) );
  OAI222_X1 U6180 ( .A1(n1990), .A2(n11107), .B1(n262), .B2(n11104), .C1(n1127), .C2(n11101), .ZN(n4783) );
  OAI222_X1 U6181 ( .A1(n9182), .A2(n11041), .B1(n9181), .B2(n11038), .C1(
        n9183), .C2(n11035), .ZN(n4792) );
  OAI222_X1 U6182 ( .A1(n9174), .A2(n10975), .B1(n9173), .B2(n10972), .C1(
        n9175), .C2(n10969), .ZN(n4801) );
  OAI222_X1 U6183 ( .A1(n1990), .A2(n11371), .B1(n262), .B2(n11368), .C1(n1127), .C2(n11365), .ZN(n3350) );
  OAI222_X1 U6184 ( .A1(n9182), .A2(n11305), .B1(n9181), .B2(n11302), .C1(
        n9183), .C2(n11299), .ZN(n3359) );
  OAI222_X1 U6185 ( .A1(n9174), .A2(n11239), .B1(n9173), .B2(n11236), .C1(
        n9175), .C2(n11233), .ZN(n3368) );
  OAI222_X1 U6186 ( .A1(n1978), .A2(n11107), .B1(n250), .B2(n11104), .C1(n1115), .C2(n11101), .ZN(n4742) );
  OAI222_X1 U6187 ( .A1(n9150), .A2(n11041), .B1(n9149), .B2(n11038), .C1(
        n9151), .C2(n11035), .ZN(n4751) );
  OAI222_X1 U6188 ( .A1(n9142), .A2(n10975), .B1(n9141), .B2(n10972), .C1(
        n9143), .C2(n10969), .ZN(n4760) );
  OAI222_X1 U6189 ( .A1(n1978), .A2(n11371), .B1(n250), .B2(n11368), .C1(n1115), .C2(n11365), .ZN(n3309) );
  OAI222_X1 U6190 ( .A1(n9150), .A2(n11305), .B1(n9149), .B2(n11302), .C1(
        n9151), .C2(n11299), .ZN(n3318) );
  OAI222_X1 U6191 ( .A1(n9142), .A2(n11239), .B1(n9141), .B2(n11236), .C1(
        n9143), .C2(n11233), .ZN(n3327) );
  OAI222_X1 U6192 ( .A1(n1966), .A2(n11107), .B1(n238), .B2(n11104), .C1(n1103), .C2(n11101), .ZN(n4701) );
  OAI222_X1 U6193 ( .A1(n6236), .A2(n11041), .B1(n6140), .B2(n11038), .C1(
        n6301), .C2(n11035), .ZN(n4710) );
  OAI222_X1 U6194 ( .A1(n6007), .A2(n10975), .B1(n6006), .B2(n10972), .C1(
        n6008), .C2(n10969), .ZN(n4719) );
  OAI222_X1 U6195 ( .A1(n1966), .A2(n11371), .B1(n238), .B2(n11368), .C1(n1103), .C2(n11365), .ZN(n3268) );
  OAI222_X1 U6196 ( .A1(n6236), .A2(n11305), .B1(n6140), .B2(n11302), .C1(
        n6301), .C2(n11299), .ZN(n3277) );
  OAI222_X1 U6197 ( .A1(n6007), .A2(n11239), .B1(n6006), .B2(n11236), .C1(
        n6008), .C2(n11233), .ZN(n3286) );
  OAI222_X1 U6198 ( .A1(n1954), .A2(n11108), .B1(n226), .B2(n11105), .C1(n1091), .C2(n11102), .ZN(n4660) );
  OAI222_X1 U6199 ( .A1(n5983), .A2(n11042), .B1(n5982), .B2(n11039), .C1(
        n5984), .C2(n11036), .ZN(n4669) );
  OAI222_X1 U6200 ( .A1(n5943), .A2(n10976), .B1(n5942), .B2(n10973), .C1(
        n5944), .C2(n10970), .ZN(n4678) );
  OAI222_X1 U6201 ( .A1(n1954), .A2(n11372), .B1(n226), .B2(n11369), .C1(n1091), .C2(n11366), .ZN(n3227) );
  OAI222_X1 U6202 ( .A1(n5983), .A2(n11306), .B1(n5982), .B2(n11303), .C1(
        n5984), .C2(n11300), .ZN(n3236) );
  OAI222_X1 U6203 ( .A1(n5943), .A2(n11240), .B1(n5942), .B2(n11237), .C1(
        n5944), .C2(n11234), .ZN(n3245) );
  OAI222_X1 U6204 ( .A1(n1942), .A2(n11108), .B1(n214), .B2(n11105), .C1(n1079), .C2(n11102), .ZN(n4619) );
  OAI222_X1 U6205 ( .A1(n5919), .A2(n11042), .B1(n5918), .B2(n11039), .C1(
        n5920), .C2(n11036), .ZN(n4628) );
  OAI222_X1 U6206 ( .A1(n5911), .A2(n10976), .B1(n5910), .B2(n10973), .C1(
        n5912), .C2(n10970), .ZN(n4637) );
  OAI222_X1 U6207 ( .A1(n1942), .A2(n11372), .B1(n214), .B2(n11369), .C1(n1079), .C2(n11366), .ZN(n3186) );
  OAI222_X1 U6208 ( .A1(n5919), .A2(n11306), .B1(n5918), .B2(n11303), .C1(
        n5920), .C2(n11300), .ZN(n3195) );
  OAI222_X1 U6209 ( .A1(n5911), .A2(n11240), .B1(n5910), .B2(n11237), .C1(
        n5912), .C2(n11234), .ZN(n3204) );
  OAI222_X1 U6210 ( .A1(n1930), .A2(n11108), .B1(n202), .B2(n11105), .C1(n1067), .C2(n11102), .ZN(n4578) );
  OAI222_X1 U6211 ( .A1(n5887), .A2(n11042), .B1(n5886), .B2(n11039), .C1(
        n5888), .C2(n11036), .ZN(n4587) );
  OAI222_X1 U6212 ( .A1(n5879), .A2(n10976), .B1(n5878), .B2(n10973), .C1(
        n5880), .C2(n10970), .ZN(n4596) );
  OAI222_X1 U6213 ( .A1(n1930), .A2(n11372), .B1(n202), .B2(n11369), .C1(n1067), .C2(n11366), .ZN(n3145) );
  OAI222_X1 U6214 ( .A1(n5887), .A2(n11306), .B1(n5886), .B2(n11303), .C1(
        n5888), .C2(n11300), .ZN(n3154) );
  OAI222_X1 U6215 ( .A1(n5879), .A2(n11240), .B1(n5878), .B2(n11237), .C1(
        n5880), .C2(n11234), .ZN(n3163) );
  OAI222_X1 U6216 ( .A1(n1918), .A2(n11108), .B1(n190), .B2(n11105), .C1(n1055), .C2(n11102), .ZN(n4537) );
  OAI222_X1 U6217 ( .A1(n5855), .A2(n11042), .B1(n5854), .B2(n11039), .C1(
        n5856), .C2(n11036), .ZN(n4546) );
  OAI222_X1 U6218 ( .A1(n5847), .A2(n10976), .B1(n5846), .B2(n10973), .C1(
        n5848), .C2(n10970), .ZN(n4555) );
  OAI222_X1 U6219 ( .A1(n1918), .A2(n11372), .B1(n190), .B2(n11369), .C1(n1055), .C2(n11366), .ZN(n3104) );
  OAI222_X1 U6220 ( .A1(n5855), .A2(n11306), .B1(n5854), .B2(n11303), .C1(
        n5856), .C2(n11300), .ZN(n3113) );
  OAI222_X1 U6221 ( .A1(n5847), .A2(n11240), .B1(n5846), .B2(n11237), .C1(
        n5848), .C2(n11234), .ZN(n3122) );
  OAI222_X1 U6222 ( .A1(n1906), .A2(n11108), .B1(n178), .B2(n11105), .C1(n1043), .C2(n11102), .ZN(n4496) );
  OAI222_X1 U6223 ( .A1(n5823), .A2(n11042), .B1(n5822), .B2(n11039), .C1(
        n5824), .C2(n11036), .ZN(n4505) );
  OAI222_X1 U6224 ( .A1(n5815), .A2(n10976), .B1(n5814), .B2(n10973), .C1(
        n5816), .C2(n10970), .ZN(n4514) );
  OAI222_X1 U6225 ( .A1(n1906), .A2(n11372), .B1(n178), .B2(n11369), .C1(n1043), .C2(n11366), .ZN(n3063) );
  OAI222_X1 U6226 ( .A1(n5823), .A2(n11306), .B1(n5822), .B2(n11303), .C1(
        n5824), .C2(n11300), .ZN(n3072) );
  OAI222_X1 U6227 ( .A1(n5815), .A2(n11240), .B1(n5814), .B2(n11237), .C1(
        n5816), .C2(n11234), .ZN(n3081) );
  OAI222_X1 U6228 ( .A1(n5791), .A2(n11042), .B1(n5790), .B2(n11039), .C1(
        n5792), .C2(n11036), .ZN(n4464) );
  OAI222_X1 U6229 ( .A1(n5783), .A2(n10976), .B1(n5782), .B2(n10973), .C1(
        n5784), .C2(n10970), .ZN(n4473) );
  OAI222_X1 U6230 ( .A1(n5791), .A2(n11306), .B1(n5790), .B2(n11303), .C1(
        n5792), .C2(n11300), .ZN(n3031) );
  OAI222_X1 U6231 ( .A1(n5783), .A2(n11240), .B1(n5782), .B2(n11237), .C1(
        n5784), .C2(n11234), .ZN(n3040) );
  OAI222_X1 U6232 ( .A1(n5759), .A2(n11042), .B1(n5758), .B2(n11039), .C1(
        n5760), .C2(n11036), .ZN(n4423) );
  OAI222_X1 U6233 ( .A1(n5751), .A2(n10976), .B1(n5750), .B2(n10973), .C1(
        n5752), .C2(n10970), .ZN(n4432) );
  OAI222_X1 U6234 ( .A1(n5759), .A2(n11306), .B1(n5758), .B2(n11303), .C1(
        n5760), .C2(n11300), .ZN(n2990) );
  OAI222_X1 U6235 ( .A1(n5751), .A2(n11240), .B1(n5750), .B2(n11237), .C1(
        n5752), .C2(n11234), .ZN(n2999) );
  OAI222_X1 U6236 ( .A1(n5727), .A2(n11042), .B1(n5726), .B2(n11039), .C1(
        n5728), .C2(n11036), .ZN(n4316) );
  OAI222_X1 U6237 ( .A1(n5719), .A2(n10976), .B1(n5718), .B2(n10973), .C1(
        n5720), .C2(n10970), .ZN(n4347) );
  OAI222_X1 U6238 ( .A1(n14035), .A2(n10910), .B1(n14067), .B2(n10907), .C1(
        n998), .C2(n10904), .ZN(n4378) );
  OAI222_X1 U6239 ( .A1(n5727), .A2(n11306), .B1(n5726), .B2(n11303), .C1(
        n5728), .C2(n11300), .ZN(n2816) );
  OAI222_X1 U6240 ( .A1(n5719), .A2(n11240), .B1(n5718), .B2(n11237), .C1(
        n5720), .C2(n11234), .ZN(n2879) );
  OAI222_X1 U6241 ( .A1(n14035), .A2(n11174), .B1(n14067), .B2(n11171), .C1(
        n998), .C2(n11168), .ZN(n2945) );
  OAI222_X1 U6242 ( .A1(n1894), .A2(n11108), .B1(n166), .B2(n11105), .C1(
        n12782), .C2(n11102), .ZN(n4455) );
  OAI222_X1 U6243 ( .A1(n1894), .A2(n11372), .B1(n166), .B2(n11369), .C1(
        n12782), .C2(n11366), .ZN(n3022) );
  OAI222_X1 U6244 ( .A1(n1882), .A2(n11108), .B1(n154), .B2(n11105), .C1(
        n12781), .C2(n11102), .ZN(n4414) );
  OAI222_X1 U6245 ( .A1(n1882), .A2(n11372), .B1(n154), .B2(n11369), .C1(
        n12781), .C2(n11366), .ZN(n2981) );
  OAI222_X1 U6246 ( .A1(n1870), .A2(n11108), .B1(n142), .B2(n11105), .C1(
        n12780), .C2(n11102), .ZN(n4285) );
  OAI222_X1 U6247 ( .A1(n1870), .A2(n11372), .B1(n142), .B2(n11369), .C1(
        n12780), .C2(n11366), .ZN(n2753) );
  OAI222_X1 U6248 ( .A1(n10534), .A2(n11073), .B1(n10533), .B2(n11070), .C1(
        n10535), .C2(n11067), .ZN(n5658) );
  OAI222_X1 U6249 ( .A1(n10534), .A2(n11337), .B1(n10533), .B2(n11334), .C1(
        n10535), .C2(n11331), .ZN(n4225) );
  OAI222_X1 U6250 ( .A1(n10502), .A2(n11073), .B1(n10501), .B2(n11070), .C1(
        n10503), .C2(n11067), .ZN(n5605) );
  OAI222_X1 U6251 ( .A1(n10502), .A2(n11337), .B1(n10501), .B2(n11334), .C1(
        n10503), .C2(n11331), .ZN(n4172) );
  OAI222_X1 U6252 ( .A1(n10470), .A2(n11073), .B1(n10469), .B2(n11070), .C1(
        n10471), .C2(n11067), .ZN(n5564) );
  OAI222_X1 U6253 ( .A1(n10470), .A2(n11337), .B1(n10469), .B2(n11334), .C1(
        n10471), .C2(n11331), .ZN(n4131) );
  OAI222_X1 U6254 ( .A1(n10438), .A2(n11073), .B1(n10437), .B2(n11070), .C1(
        n10439), .C2(n11067), .ZN(n5523) );
  OAI222_X1 U6255 ( .A1(n10438), .A2(n11337), .B1(n10437), .B2(n11334), .C1(
        n10439), .C2(n11331), .ZN(n4090) );
  OAI222_X1 U6256 ( .A1(n10406), .A2(n11073), .B1(n10405), .B2(n11070), .C1(
        n10407), .C2(n11067), .ZN(n5482) );
  OAI222_X1 U6257 ( .A1(n10406), .A2(n11337), .B1(n10405), .B2(n11334), .C1(
        n10407), .C2(n11331), .ZN(n4049) );
  OAI222_X1 U6258 ( .A1(n10371), .A2(n11073), .B1(n10370), .B2(n11070), .C1(
        n10372), .C2(n11067), .ZN(n5441) );
  OAI222_X1 U6259 ( .A1(n10371), .A2(n11337), .B1(n10370), .B2(n11334), .C1(
        n10372), .C2(n11331), .ZN(n4008) );
  OAI222_X1 U6260 ( .A1(n10339), .A2(n11073), .B1(n10338), .B2(n11070), .C1(
        n10340), .C2(n11067), .ZN(n5400) );
  OAI222_X1 U6261 ( .A1(n10339), .A2(n11337), .B1(n10338), .B2(n11334), .C1(
        n10340), .C2(n11331), .ZN(n3967) );
  OAI222_X1 U6262 ( .A1(n10307), .A2(n11073), .B1(n10306), .B2(n11070), .C1(
        n10308), .C2(n11067), .ZN(n5359) );
  OAI222_X1 U6263 ( .A1(n10307), .A2(n11337), .B1(n10306), .B2(n11334), .C1(
        n10308), .C2(n11331), .ZN(n3926) );
  OAI222_X1 U6264 ( .A1(n10272), .A2(n11073), .B1(n10271), .B2(n11070), .C1(
        n10273), .C2(n11067), .ZN(n5318) );
  OAI222_X1 U6265 ( .A1(n10272), .A2(n11337), .B1(n10271), .B2(n11334), .C1(
        n10273), .C2(n11331), .ZN(n3885) );
  OAI222_X1 U6266 ( .A1(n10240), .A2(n11073), .B1(n10239), .B2(n11070), .C1(
        n10241), .C2(n11067), .ZN(n5277) );
  OAI222_X1 U6267 ( .A1(n10240), .A2(n11337), .B1(n10239), .B2(n11334), .C1(
        n10241), .C2(n11331), .ZN(n3844) );
  OAI222_X1 U6268 ( .A1(n10208), .A2(n11073), .B1(n10205), .B2(n11070), .C1(
        n10209), .C2(n11067), .ZN(n5236) );
  OAI222_X1 U6269 ( .A1(n10208), .A2(n11337), .B1(n10205), .B2(n11334), .C1(
        n10209), .C2(n11331), .ZN(n3803) );
  OAI222_X1 U6270 ( .A1(n10174), .A2(n11073), .B1(n10173), .B2(n11070), .C1(
        n10175), .C2(n11067), .ZN(n5195) );
  OAI222_X1 U6271 ( .A1(n10174), .A2(n11337), .B1(n10173), .B2(n11334), .C1(
        n10175), .C2(n11331), .ZN(n3762) );
  OAI222_X1 U6272 ( .A1(n10142), .A2(n11074), .B1(n10141), .B2(n11071), .C1(
        n10143), .C2(n11068), .ZN(n5154) );
  OAI222_X1 U6273 ( .A1(n10142), .A2(n11338), .B1(n10141), .B2(n11335), .C1(
        n10143), .C2(n11332), .ZN(n3721) );
  OAI222_X1 U6274 ( .A1(n10110), .A2(n11074), .B1(n10109), .B2(n11071), .C1(
        n10111), .C2(n11068), .ZN(n5113) );
  OAI222_X1 U6275 ( .A1(n10110), .A2(n11338), .B1(n10109), .B2(n11335), .C1(
        n10111), .C2(n11332), .ZN(n3680) );
  OAI222_X1 U6276 ( .A1(n10078), .A2(n11074), .B1(n10077), .B2(n11071), .C1(
        n10079), .C2(n11068), .ZN(n5072) );
  OAI222_X1 U6277 ( .A1(n10078), .A2(n11338), .B1(n10077), .B2(n11335), .C1(
        n10079), .C2(n11332), .ZN(n3639) );
  OAI222_X1 U6278 ( .A1(n10046), .A2(n11074), .B1(n10045), .B2(n11071), .C1(
        n10047), .C2(n11068), .ZN(n5031) );
  OAI222_X1 U6279 ( .A1(n10046), .A2(n11338), .B1(n10045), .B2(n11335), .C1(
        n10047), .C2(n11332), .ZN(n3598) );
  OAI222_X1 U6280 ( .A1(n10014), .A2(n11074), .B1(n10013), .B2(n11071), .C1(
        n10015), .C2(n11068), .ZN(n4990) );
  OAI222_X1 U6281 ( .A1(n10014), .A2(n11338), .B1(n10013), .B2(n11335), .C1(
        n10015), .C2(n11332), .ZN(n3557) );
  OAI222_X1 U6282 ( .A1(n9652), .A2(n11074), .B1(n9651), .B2(n11071), .C1(
        n9653), .C2(n11068), .ZN(n4949) );
  OAI222_X1 U6283 ( .A1(n9652), .A2(n11338), .B1(n9651), .B2(n11335), .C1(
        n9653), .C2(n11332), .ZN(n3516) );
  OAI222_X1 U6284 ( .A1(n9620), .A2(n11074), .B1(n9619), .B2(n11071), .C1(
        n9621), .C2(n11068), .ZN(n4908) );
  OAI222_X1 U6285 ( .A1(n9620), .A2(n11338), .B1(n9619), .B2(n11335), .C1(
        n9621), .C2(n11332), .ZN(n3475) );
  OAI222_X1 U6286 ( .A1(n9588), .A2(n11074), .B1(n9587), .B2(n11071), .C1(
        n9589), .C2(n11068), .ZN(n4867) );
  OAI222_X1 U6287 ( .A1(n9588), .A2(n11338), .B1(n9587), .B2(n11335), .C1(
        n9589), .C2(n11332), .ZN(n3434) );
  OAI222_X1 U6288 ( .A1(n9254), .A2(n11074), .B1(n9253), .B2(n11071), .C1(
        n9255), .C2(n11068), .ZN(n4826) );
  OAI222_X1 U6289 ( .A1(n9254), .A2(n11338), .B1(n9253), .B2(n11335), .C1(
        n9255), .C2(n11332), .ZN(n3393) );
  OAI222_X1 U6290 ( .A1(n9190), .A2(n11074), .B1(n9189), .B2(n11071), .C1(
        n9191), .C2(n11068), .ZN(n4785) );
  OAI222_X1 U6291 ( .A1(n9190), .A2(n11338), .B1(n9189), .B2(n11335), .C1(
        n9191), .C2(n11332), .ZN(n3352) );
  OAI222_X1 U6292 ( .A1(n9158), .A2(n11074), .B1(n9157), .B2(n11071), .C1(
        n9159), .C2(n11068), .ZN(n4744) );
  OAI222_X1 U6293 ( .A1(n9158), .A2(n11338), .B1(n9157), .B2(n11335), .C1(
        n9159), .C2(n11332), .ZN(n3311) );
  OAI222_X1 U6294 ( .A1(n6308), .A2(n11074), .B1(n6307), .B2(n11071), .C1(
        n6309), .C2(n11068), .ZN(n4703) );
  OAI222_X1 U6295 ( .A1(n6308), .A2(n11338), .B1(n6307), .B2(n11335), .C1(
        n6309), .C2(n11332), .ZN(n3270) );
  OAI222_X1 U6296 ( .A1(n5991), .A2(n11075), .B1(n5990), .B2(n11072), .C1(
        n5992), .C2(n11069), .ZN(n4662) );
  OAI222_X1 U6297 ( .A1(n5991), .A2(n11339), .B1(n5990), .B2(n11336), .C1(
        n5992), .C2(n11333), .ZN(n3229) );
  OAI222_X1 U6298 ( .A1(n5927), .A2(n11075), .B1(n5926), .B2(n11072), .C1(
        n5928), .C2(n11069), .ZN(n4621) );
  OAI222_X1 U6299 ( .A1(n5927), .A2(n11339), .B1(n5926), .B2(n11336), .C1(
        n5928), .C2(n11333), .ZN(n3188) );
  OAI222_X1 U6300 ( .A1(n5895), .A2(n11075), .B1(n5894), .B2(n11072), .C1(
        n5896), .C2(n11069), .ZN(n4580) );
  OAI222_X1 U6301 ( .A1(n5895), .A2(n11339), .B1(n5894), .B2(n11336), .C1(
        n5896), .C2(n11333), .ZN(n3147) );
  OAI222_X1 U6302 ( .A1(n5863), .A2(n11075), .B1(n5862), .B2(n11072), .C1(
        n5864), .C2(n11069), .ZN(n4539) );
  OAI222_X1 U6303 ( .A1(n5863), .A2(n11339), .B1(n5862), .B2(n11336), .C1(
        n5864), .C2(n11333), .ZN(n3106) );
  OAI222_X1 U6304 ( .A1(n5831), .A2(n11075), .B1(n5830), .B2(n11072), .C1(
        n5832), .C2(n11069), .ZN(n4498) );
  OAI222_X1 U6305 ( .A1(n5831), .A2(n11339), .B1(n5830), .B2(n11336), .C1(
        n5832), .C2(n11333), .ZN(n3065) );
  OAI222_X1 U6306 ( .A1(n5799), .A2(n11075), .B1(n5798), .B2(n11072), .C1(
        n5800), .C2(n11069), .ZN(n4457) );
  OAI222_X1 U6307 ( .A1(n5799), .A2(n11339), .B1(n5798), .B2(n11336), .C1(
        n5800), .C2(n11333), .ZN(n3024) );
  OAI222_X1 U6308 ( .A1(n5767), .A2(n11075), .B1(n5766), .B2(n11072), .C1(
        n5768), .C2(n11069), .ZN(n4416) );
  OAI222_X1 U6309 ( .A1(n5767), .A2(n11339), .B1(n5766), .B2(n11336), .C1(
        n5768), .C2(n11333), .ZN(n2983) );
  OAI222_X1 U6310 ( .A1(n5735), .A2(n11075), .B1(n5734), .B2(n11072), .C1(
        n5736), .C2(n11069), .ZN(n4300) );
  OAI222_X1 U6311 ( .A1(n5735), .A2(n11339), .B1(n5734), .B2(n11336), .C1(
        n5736), .C2(n11333), .ZN(n2800) );
  OAI222_X1 U6312 ( .A1(n2337), .A2(n11097), .B1(n513), .B2(n11094), .C1(n1442), .C2(n11091), .ZN(n5643) );
  OAI222_X1 U6313 ( .A1(n10523), .A2(n11031), .B1(n10522), .B2(n11028), .C1(
        n10524), .C2(n11025), .ZN(n5671) );
  OAI222_X1 U6314 ( .A1(n2337), .A2(n11361), .B1(n513), .B2(n11358), .C1(n1442), .C2(n11355), .ZN(n4210) );
  OAI222_X1 U6315 ( .A1(n10523), .A2(n11295), .B1(n10522), .B2(n11292), .C1(
        n10524), .C2(n11289), .ZN(n4238) );
  OAI222_X1 U6316 ( .A1(n2325), .A2(n11097), .B1(n501), .B2(n11094), .C1(n1398), .C2(n11091), .ZN(n5602) );
  OAI222_X1 U6317 ( .A1(n10491), .A2(n11031), .B1(n10490), .B2(n11028), .C1(
        n10492), .C2(n11025), .ZN(n5611) );
  OAI222_X1 U6318 ( .A1(n2325), .A2(n11361), .B1(n501), .B2(n11358), .C1(n1398), .C2(n11355), .ZN(n4169) );
  OAI222_X1 U6319 ( .A1(n10491), .A2(n11295), .B1(n10490), .B2(n11292), .C1(
        n10492), .C2(n11289), .ZN(n4178) );
  OAI222_X1 U6320 ( .A1(n2313), .A2(n11097), .B1(n489), .B2(n11094), .C1(n1386), .C2(n11091), .ZN(n5561) );
  OAI222_X1 U6321 ( .A1(n10459), .A2(n11031), .B1(n10458), .B2(n11028), .C1(
        n10460), .C2(n11025), .ZN(n5570) );
  OAI222_X1 U6322 ( .A1(n2313), .A2(n11361), .B1(n489), .B2(n11358), .C1(n1386), .C2(n11355), .ZN(n4128) );
  OAI222_X1 U6323 ( .A1(n10459), .A2(n11295), .B1(n10458), .B2(n11292), .C1(
        n10460), .C2(n11289), .ZN(n4137) );
  OAI222_X1 U6324 ( .A1(n2301), .A2(n11097), .B1(n477), .B2(n11094), .C1(n1342), .C2(n11091), .ZN(n5520) );
  OAI222_X1 U6325 ( .A1(n10427), .A2(n11031), .B1(n10426), .B2(n11028), .C1(
        n10428), .C2(n11025), .ZN(n5529) );
  OAI222_X1 U6326 ( .A1(n2301), .A2(n11361), .B1(n477), .B2(n11358), .C1(n1342), .C2(n11355), .ZN(n4087) );
  OAI222_X1 U6327 ( .A1(n10427), .A2(n11295), .B1(n10426), .B2(n11292), .C1(
        n10428), .C2(n11289), .ZN(n4096) );
  OAI222_X1 U6328 ( .A1(n2289), .A2(n11097), .B1(n465), .B2(n11094), .C1(n1330), .C2(n11091), .ZN(n5479) );
  OAI222_X1 U6329 ( .A1(n10392), .A2(n11031), .B1(n10391), .B2(n11028), .C1(
        n10393), .C2(n11025), .ZN(n5488) );
  OAI222_X1 U6330 ( .A1(n2289), .A2(n11361), .B1(n465), .B2(n11358), .C1(n1330), .C2(n11355), .ZN(n4046) );
  OAI222_X1 U6331 ( .A1(n10392), .A2(n11295), .B1(n10391), .B2(n11292), .C1(
        n10393), .C2(n11289), .ZN(n4055) );
  OAI222_X1 U6332 ( .A1(n2277), .A2(n11097), .B1(n453), .B2(n11094), .C1(n1318), .C2(n11091), .ZN(n5438) );
  OAI222_X1 U6333 ( .A1(n10360), .A2(n11031), .B1(n10359), .B2(n11028), .C1(
        n10361), .C2(n11025), .ZN(n5447) );
  OAI222_X1 U6334 ( .A1(n2277), .A2(n11361), .B1(n453), .B2(n11358), .C1(n1318), .C2(n11355), .ZN(n4005) );
  OAI222_X1 U6335 ( .A1(n10360), .A2(n11295), .B1(n10359), .B2(n11292), .C1(
        n10361), .C2(n11289), .ZN(n4014) );
  OAI222_X1 U6336 ( .A1(n2265), .A2(n11097), .B1(n441), .B2(n11094), .C1(n1306), .C2(n11091), .ZN(n5397) );
  OAI222_X1 U6337 ( .A1(n10328), .A2(n11031), .B1(n10327), .B2(n11028), .C1(
        n10329), .C2(n11025), .ZN(n5406) );
  OAI222_X1 U6338 ( .A1(n2265), .A2(n11361), .B1(n441), .B2(n11358), .C1(n1306), .C2(n11355), .ZN(n3964) );
  OAI222_X1 U6339 ( .A1(n10328), .A2(n11295), .B1(n10327), .B2(n11292), .C1(
        n10329), .C2(n11289), .ZN(n3973) );
  OAI222_X1 U6340 ( .A1(n2253), .A2(n11097), .B1(n429), .B2(n11094), .C1(n1294), .C2(n11091), .ZN(n5356) );
  OAI222_X1 U6341 ( .A1(n10293), .A2(n11031), .B1(n10292), .B2(n11028), .C1(
        n10294), .C2(n11025), .ZN(n5365) );
  OAI222_X1 U6342 ( .A1(n2253), .A2(n11361), .B1(n429), .B2(n11358), .C1(n1294), .C2(n11355), .ZN(n3923) );
  OAI222_X1 U6343 ( .A1(n10293), .A2(n11295), .B1(n10292), .B2(n11292), .C1(
        n10294), .C2(n11289), .ZN(n3932) );
  OAI222_X1 U6344 ( .A1(n2241), .A2(n11097), .B1(n417), .B2(n11094), .C1(n1282), .C2(n11091), .ZN(n5315) );
  OAI222_X1 U6345 ( .A1(n10261), .A2(n11031), .B1(n10260), .B2(n11028), .C1(
        n10262), .C2(n11025), .ZN(n5324) );
  OAI222_X1 U6346 ( .A1(n2241), .A2(n11361), .B1(n417), .B2(n11358), .C1(n1282), .C2(n11355), .ZN(n3882) );
  OAI222_X1 U6347 ( .A1(n10261), .A2(n11295), .B1(n10260), .B2(n11292), .C1(
        n10262), .C2(n11289), .ZN(n3891) );
  OAI222_X1 U6348 ( .A1(n2229), .A2(n11097), .B1(n405), .B2(n11094), .C1(n1270), .C2(n11091), .ZN(n5274) );
  OAI222_X1 U6349 ( .A1(n10229), .A2(n11031), .B1(n10228), .B2(n11028), .C1(
        n10230), .C2(n11025), .ZN(n5283) );
  OAI222_X1 U6350 ( .A1(n2229), .A2(n11361), .B1(n405), .B2(n11358), .C1(n1270), .C2(n11355), .ZN(n3841) );
  OAI222_X1 U6351 ( .A1(n10229), .A2(n11295), .B1(n10228), .B2(n11292), .C1(
        n10230), .C2(n11289), .ZN(n3850) );
  OAI222_X1 U6352 ( .A1(n2217), .A2(n11097), .B1(n393), .B2(n11094), .C1(n1258), .C2(n11091), .ZN(n5233) );
  OAI222_X1 U6353 ( .A1(n10195), .A2(n11031), .B1(n10194), .B2(n11028), .C1(
        n10196), .C2(n11025), .ZN(n5242) );
  OAI222_X1 U6354 ( .A1(n2217), .A2(n11361), .B1(n393), .B2(n11358), .C1(n1258), .C2(n11355), .ZN(n3800) );
  OAI222_X1 U6355 ( .A1(n10195), .A2(n11295), .B1(n10194), .B2(n11292), .C1(
        n10196), .C2(n11289), .ZN(n3809) );
  OAI222_X1 U6356 ( .A1(n2173), .A2(n11097), .B1(n381), .B2(n11094), .C1(n1246), .C2(n11091), .ZN(n5192) );
  OAI222_X1 U6357 ( .A1(n10163), .A2(n11031), .B1(n10162), .B2(n11028), .C1(
        n10164), .C2(n11025), .ZN(n5201) );
  OAI222_X1 U6358 ( .A1(n2173), .A2(n11361), .B1(n381), .B2(n11358), .C1(n1246), .C2(n11355), .ZN(n3759) );
  OAI222_X1 U6359 ( .A1(n10163), .A2(n11295), .B1(n10162), .B2(n11292), .C1(
        n10164), .C2(n11289), .ZN(n3768) );
  OAI222_X1 U6360 ( .A1(n2161), .A2(n11098), .B1(n369), .B2(n11095), .C1(n1234), .C2(n11092), .ZN(n5151) );
  OAI222_X1 U6361 ( .A1(n10131), .A2(n11032), .B1(n10130), .B2(n11029), .C1(
        n10132), .C2(n11026), .ZN(n5160) );
  OAI222_X1 U6362 ( .A1(n2161), .A2(n11362), .B1(n369), .B2(n11359), .C1(n1234), .C2(n11356), .ZN(n3718) );
  OAI222_X1 U6363 ( .A1(n10131), .A2(n11296), .B1(n10130), .B2(n11293), .C1(
        n10132), .C2(n11290), .ZN(n3727) );
  OAI222_X1 U6364 ( .A1(n2149), .A2(n11098), .B1(n357), .B2(n11095), .C1(n1222), .C2(n11092), .ZN(n5110) );
  OAI222_X1 U6365 ( .A1(n10099), .A2(n11032), .B1(n10098), .B2(n11029), .C1(
        n10100), .C2(n11026), .ZN(n5119) );
  OAI222_X1 U6366 ( .A1(n2149), .A2(n11362), .B1(n357), .B2(n11359), .C1(n1222), .C2(n11356), .ZN(n3677) );
  OAI222_X1 U6367 ( .A1(n10099), .A2(n11296), .B1(n10098), .B2(n11293), .C1(
        n10100), .C2(n11290), .ZN(n3686) );
  OAI222_X1 U6368 ( .A1(n2105), .A2(n11098), .B1(n345), .B2(n11095), .C1(n1210), .C2(n11092), .ZN(n5069) );
  OAI222_X1 U6369 ( .A1(n10067), .A2(n11032), .B1(n10066), .B2(n11029), .C1(
        n10068), .C2(n11026), .ZN(n5078) );
  OAI222_X1 U6370 ( .A1(n2105), .A2(n11362), .B1(n345), .B2(n11359), .C1(n1210), .C2(n11356), .ZN(n3636) );
  OAI222_X1 U6371 ( .A1(n10067), .A2(n11296), .B1(n10066), .B2(n11293), .C1(
        n10068), .C2(n11290), .ZN(n3645) );
  OAI222_X1 U6372 ( .A1(n2093), .A2(n11098), .B1(n333), .B2(n11095), .C1(n1198), .C2(n11092), .ZN(n5028) );
  OAI222_X1 U6373 ( .A1(n10035), .A2(n11032), .B1(n10034), .B2(n11029), .C1(
        n10036), .C2(n11026), .ZN(n5037) );
  OAI222_X1 U6374 ( .A1(n2093), .A2(n11362), .B1(n333), .B2(n11359), .C1(n1198), .C2(n11356), .ZN(n3595) );
  OAI222_X1 U6375 ( .A1(n10035), .A2(n11296), .B1(n10034), .B2(n11293), .C1(
        n10036), .C2(n11290), .ZN(n3604) );
  OAI222_X1 U6376 ( .A1(n2049), .A2(n11098), .B1(n321), .B2(n11095), .C1(n1186), .C2(n11092), .ZN(n4987) );
  OAI222_X1 U6377 ( .A1(n10003), .A2(n11032), .B1(n10002), .B2(n11029), .C1(
        n10004), .C2(n11026), .ZN(n4996) );
  OAI222_X1 U6378 ( .A1(n2049), .A2(n11362), .B1(n321), .B2(n11359), .C1(n1186), .C2(n11356), .ZN(n3554) );
  OAI222_X1 U6379 ( .A1(n10003), .A2(n11296), .B1(n10002), .B2(n11293), .C1(
        n10004), .C2(n11290), .ZN(n3563) );
  OAI222_X1 U6380 ( .A1(n2037), .A2(n11098), .B1(n309), .B2(n11095), .C1(n1174), .C2(n11092), .ZN(n4946) );
  OAI222_X1 U6381 ( .A1(n9641), .A2(n11032), .B1(n9640), .B2(n11029), .C1(
        n9642), .C2(n11026), .ZN(n4955) );
  OAI222_X1 U6382 ( .A1(n2037), .A2(n11362), .B1(n309), .B2(n11359), .C1(n1174), .C2(n11356), .ZN(n3513) );
  OAI222_X1 U6383 ( .A1(n9641), .A2(n11296), .B1(n9640), .B2(n11293), .C1(
        n9642), .C2(n11290), .ZN(n3522) );
  OAI222_X1 U6384 ( .A1(n2025), .A2(n11098), .B1(n297), .B2(n11095), .C1(n1162), .C2(n11092), .ZN(n4905) );
  OAI222_X1 U6385 ( .A1(n9609), .A2(n11032), .B1(n9608), .B2(n11029), .C1(
        n9610), .C2(n11026), .ZN(n4914) );
  OAI222_X1 U6386 ( .A1(n2025), .A2(n11362), .B1(n297), .B2(n11359), .C1(n1162), .C2(n11356), .ZN(n3472) );
  OAI222_X1 U6387 ( .A1(n9609), .A2(n11296), .B1(n9608), .B2(n11293), .C1(
        n9610), .C2(n11290), .ZN(n3481) );
  OAI222_X1 U6388 ( .A1(n2013), .A2(n11098), .B1(n285), .B2(n11095), .C1(n1150), .C2(n11092), .ZN(n4864) );
  OAI222_X1 U6389 ( .A1(n9577), .A2(n11032), .B1(n9576), .B2(n11029), .C1(
        n9578), .C2(n11026), .ZN(n4873) );
  OAI222_X1 U6390 ( .A1(n2013), .A2(n11362), .B1(n285), .B2(n11359), .C1(n1150), .C2(n11356), .ZN(n3431) );
  OAI222_X1 U6391 ( .A1(n9577), .A2(n11296), .B1(n9576), .B2(n11293), .C1(
        n9578), .C2(n11290), .ZN(n3440) );
  OAI222_X1 U6392 ( .A1(n2001), .A2(n11098), .B1(n273), .B2(n11095), .C1(n1138), .C2(n11092), .ZN(n4823) );
  OAI222_X1 U6393 ( .A1(n9211), .A2(n11032), .B1(n9210), .B2(n11029), .C1(
        n9212), .C2(n11026), .ZN(n4832) );
  OAI222_X1 U6394 ( .A1(n2001), .A2(n11362), .B1(n273), .B2(n11359), .C1(n1138), .C2(n11356), .ZN(n3390) );
  OAI222_X1 U6395 ( .A1(n9211), .A2(n11296), .B1(n9210), .B2(n11293), .C1(
        n9212), .C2(n11290), .ZN(n3399) );
  OAI222_X1 U6396 ( .A1(n1989), .A2(n11098), .B1(n261), .B2(n11095), .C1(n1126), .C2(n11092), .ZN(n4782) );
  OAI222_X1 U6397 ( .A1(n9179), .A2(n11032), .B1(n9178), .B2(n11029), .C1(
        n9180), .C2(n11026), .ZN(n4791) );
  OAI222_X1 U6398 ( .A1(n1989), .A2(n11362), .B1(n261), .B2(n11359), .C1(n1126), .C2(n11356), .ZN(n3349) );
  OAI222_X1 U6399 ( .A1(n9179), .A2(n11296), .B1(n9178), .B2(n11293), .C1(
        n9180), .C2(n11290), .ZN(n3358) );
  OAI222_X1 U6400 ( .A1(n1977), .A2(n11098), .B1(n249), .B2(n11095), .C1(n1114), .C2(n11092), .ZN(n4741) );
  OAI222_X1 U6401 ( .A1(n9147), .A2(n11032), .B1(n9146), .B2(n11029), .C1(
        n9148), .C2(n11026), .ZN(n4750) );
  OAI222_X1 U6402 ( .A1(n1977), .A2(n11362), .B1(n249), .B2(n11359), .C1(n1114), .C2(n11356), .ZN(n3308) );
  OAI222_X1 U6403 ( .A1(n9147), .A2(n11296), .B1(n9146), .B2(n11293), .C1(
        n9148), .C2(n11290), .ZN(n3317) );
  OAI222_X1 U6404 ( .A1(n1965), .A2(n11098), .B1(n237), .B2(n11095), .C1(n1102), .C2(n11092), .ZN(n4700) );
  OAI222_X1 U6405 ( .A1(n6012), .A2(n11032), .B1(n6011), .B2(n11029), .C1(
        n6044), .C2(n11026), .ZN(n4709) );
  OAI222_X1 U6406 ( .A1(n1965), .A2(n11362), .B1(n237), .B2(n11359), .C1(n1102), .C2(n11356), .ZN(n3267) );
  OAI222_X1 U6407 ( .A1(n6012), .A2(n11296), .B1(n6011), .B2(n11293), .C1(
        n6044), .C2(n11290), .ZN(n3276) );
  OAI222_X1 U6408 ( .A1(n1953), .A2(n11099), .B1(n225), .B2(n11096), .C1(n1090), .C2(n11093), .ZN(n4659) );
  OAI222_X1 U6409 ( .A1(n5948), .A2(n11033), .B1(n5947), .B2(n11030), .C1(
        n5981), .C2(n11027), .ZN(n4668) );
  OAI222_X1 U6410 ( .A1(n1953), .A2(n11363), .B1(n225), .B2(n11360), .C1(n1090), .C2(n11357), .ZN(n3226) );
  OAI222_X1 U6411 ( .A1(n5948), .A2(n11297), .B1(n5947), .B2(n11294), .C1(
        n5981), .C2(n11291), .ZN(n3235) );
  OAI222_X1 U6412 ( .A1(n1941), .A2(n11099), .B1(n213), .B2(n11096), .C1(n1078), .C2(n11093), .ZN(n4618) );
  OAI222_X1 U6413 ( .A1(n5916), .A2(n11033), .B1(n5915), .B2(n11030), .C1(
        n5917), .C2(n11027), .ZN(n4627) );
  OAI222_X1 U6414 ( .A1(n1941), .A2(n11363), .B1(n213), .B2(n11360), .C1(n1078), .C2(n11357), .ZN(n3185) );
  OAI222_X1 U6415 ( .A1(n5916), .A2(n11297), .B1(n5915), .B2(n11294), .C1(
        n5917), .C2(n11291), .ZN(n3194) );
  OAI222_X1 U6416 ( .A1(n1929), .A2(n11099), .B1(n201), .B2(n11096), .C1(n1066), .C2(n11093), .ZN(n4577) );
  OAI222_X1 U6417 ( .A1(n5884), .A2(n11033), .B1(n5883), .B2(n11030), .C1(
        n5885), .C2(n11027), .ZN(n4586) );
  OAI222_X1 U6418 ( .A1(n1929), .A2(n11363), .B1(n201), .B2(n11360), .C1(n1066), .C2(n11357), .ZN(n3144) );
  OAI222_X1 U6419 ( .A1(n5884), .A2(n11297), .B1(n5883), .B2(n11294), .C1(
        n5885), .C2(n11291), .ZN(n3153) );
  OAI222_X1 U6420 ( .A1(n1917), .A2(n11099), .B1(n189), .B2(n11096), .C1(n1054), .C2(n11093), .ZN(n4536) );
  OAI222_X1 U6421 ( .A1(n5852), .A2(n11033), .B1(n5851), .B2(n11030), .C1(
        n5853), .C2(n11027), .ZN(n4545) );
  OAI222_X1 U6422 ( .A1(n1917), .A2(n11363), .B1(n189), .B2(n11360), .C1(n1054), .C2(n11357), .ZN(n3103) );
  OAI222_X1 U6423 ( .A1(n5852), .A2(n11297), .B1(n5851), .B2(n11294), .C1(
        n5853), .C2(n11291), .ZN(n3112) );
  OAI222_X1 U6424 ( .A1(n1905), .A2(n11099), .B1(n177), .B2(n11096), .C1(n1042), .C2(n11093), .ZN(n4495) );
  OAI222_X1 U6425 ( .A1(n5820), .A2(n11033), .B1(n5819), .B2(n11030), .C1(
        n5821), .C2(n11027), .ZN(n4504) );
  OAI222_X1 U6426 ( .A1(n1905), .A2(n11363), .B1(n177), .B2(n11360), .C1(n1042), .C2(n11357), .ZN(n3062) );
  OAI222_X1 U6427 ( .A1(n5820), .A2(n11297), .B1(n5819), .B2(n11294), .C1(
        n5821), .C2(n11291), .ZN(n3071) );
  OAI222_X1 U6428 ( .A1(n5788), .A2(n11033), .B1(n5787), .B2(n11030), .C1(
        n5789), .C2(n11027), .ZN(n4463) );
  OAI222_X1 U6429 ( .A1(n5788), .A2(n11297), .B1(n5787), .B2(n11294), .C1(
        n5789), .C2(n11291), .ZN(n3030) );
  OAI222_X1 U6430 ( .A1(n5756), .A2(n11033), .B1(n5755), .B2(n11030), .C1(
        n5757), .C2(n11027), .ZN(n4422) );
  OAI222_X1 U6431 ( .A1(n5756), .A2(n11297), .B1(n5755), .B2(n11294), .C1(
        n5757), .C2(n11291), .ZN(n2989) );
  OAI222_X1 U6432 ( .A1(n5724), .A2(n11033), .B1(n5723), .B2(n11030), .C1(
        n5725), .C2(n11027), .ZN(n4315) );
  OAI222_X1 U6433 ( .A1(n5724), .A2(n11297), .B1(n5723), .B2(n11294), .C1(
        n5725), .C2(n11291), .ZN(n2815) );
  OAI222_X1 U6434 ( .A1(n1893), .A2(n11099), .B1(n165), .B2(n11096), .C1(
        n12785), .C2(n11093), .ZN(n4454) );
  OAI222_X1 U6435 ( .A1(n1893), .A2(n11363), .B1(n165), .B2(n11360), .C1(
        n12785), .C2(n11357), .ZN(n3021) );
  OAI222_X1 U6436 ( .A1(n1881), .A2(n11099), .B1(n153), .B2(n11096), .C1(
        n12784), .C2(n11093), .ZN(n4413) );
  OAI222_X1 U6437 ( .A1(n1881), .A2(n11363), .B1(n153), .B2(n11360), .C1(
        n12784), .C2(n11357), .ZN(n2980) );
  OAI222_X1 U6438 ( .A1(n1869), .A2(n11099), .B1(n141), .B2(n11096), .C1(
        n12783), .C2(n11093), .ZN(n4284) );
  OAI222_X1 U6439 ( .A1(n1869), .A2(n11363), .B1(n141), .B2(n11360), .C1(
        n12783), .C2(n11357), .ZN(n2752) );
  OAI222_X1 U6440 ( .A1(n995), .A2(n11088), .B1(n1859), .B2(n11085), .C1(n1409), .C2(n11082), .ZN(n5642) );
  OAI222_X1 U6441 ( .A1(n995), .A2(n11352), .B1(n1859), .B2(n11349), .C1(n1409), .C2(n11346), .ZN(n4209) );
  OAI222_X1 U6442 ( .A1(n991), .A2(n11088), .B1(n1855), .B2(n11085), .C1(n1397), .C2(n11082), .ZN(n5601) );
  OAI222_X1 U6443 ( .A1(n991), .A2(n11352), .B1(n1855), .B2(n11349), .C1(n1397), .C2(n11346), .ZN(n4168) );
  OAI222_X1 U6444 ( .A1(n987), .A2(n11088), .B1(n1851), .B2(n11085), .C1(n1385), .C2(n11082), .ZN(n5560) );
  OAI222_X1 U6445 ( .A1(n987), .A2(n11352), .B1(n1851), .B2(n11349), .C1(n1385), .C2(n11346), .ZN(n4127) );
  OAI222_X1 U6446 ( .A1(n983), .A2(n11088), .B1(n1847), .B2(n11085), .C1(n1341), .C2(n11082), .ZN(n5519) );
  OAI222_X1 U6447 ( .A1(n983), .A2(n11352), .B1(n1847), .B2(n11349), .C1(n1341), .C2(n11346), .ZN(n4086) );
  OAI222_X1 U6448 ( .A1(n979), .A2(n11088), .B1(n1843), .B2(n11085), .C1(n1329), .C2(n11082), .ZN(n5478) );
  OAI222_X1 U6449 ( .A1(n979), .A2(n11352), .B1(n1843), .B2(n11349), .C1(n1329), .C2(n11346), .ZN(n4045) );
  OAI222_X1 U6450 ( .A1(n975), .A2(n11088), .B1(n1839), .B2(n11085), .C1(n1317), .C2(n11082), .ZN(n5437) );
  OAI222_X1 U6451 ( .A1(n975), .A2(n11352), .B1(n1839), .B2(n11349), .C1(n1317), .C2(n11346), .ZN(n4004) );
  OAI222_X1 U6452 ( .A1(n971), .A2(n11088), .B1(n1835), .B2(n11085), .C1(n1305), .C2(n11082), .ZN(n5396) );
  OAI222_X1 U6453 ( .A1(n971), .A2(n11352), .B1(n1835), .B2(n11349), .C1(n1305), .C2(n11346), .ZN(n3963) );
  OAI222_X1 U6454 ( .A1(n967), .A2(n11088), .B1(n1831), .B2(n11085), .C1(n1293), .C2(n11082), .ZN(n5355) );
  OAI222_X1 U6455 ( .A1(n967), .A2(n11352), .B1(n1831), .B2(n11349), .C1(n1293), .C2(n11346), .ZN(n3922) );
  OAI222_X1 U6456 ( .A1(n963), .A2(n11088), .B1(n1827), .B2(n11085), .C1(n1281), .C2(n11082), .ZN(n5314) );
  OAI222_X1 U6457 ( .A1(n963), .A2(n11352), .B1(n1827), .B2(n11349), .C1(n1281), .C2(n11346), .ZN(n3881) );
  OAI222_X1 U6458 ( .A1(n959), .A2(n11088), .B1(n1823), .B2(n11085), .C1(n1269), .C2(n11082), .ZN(n5273) );
  OAI222_X1 U6459 ( .A1(n959), .A2(n11352), .B1(n1823), .B2(n11349), .C1(n1269), .C2(n11346), .ZN(n3840) );
  OAI222_X1 U6460 ( .A1(n955), .A2(n11088), .B1(n1819), .B2(n11085), .C1(n1257), .C2(n11082), .ZN(n5232) );
  OAI222_X1 U6461 ( .A1(n955), .A2(n11352), .B1(n1819), .B2(n11349), .C1(n1257), .C2(n11346), .ZN(n3799) );
  OAI222_X1 U6462 ( .A1(n951), .A2(n11088), .B1(n1815), .B2(n11085), .C1(n1245), .C2(n11082), .ZN(n5191) );
  OAI222_X1 U6463 ( .A1(n951), .A2(n11352), .B1(n1815), .B2(n11349), .C1(n1245), .C2(n11346), .ZN(n3758) );
  OAI222_X1 U6464 ( .A1(n947), .A2(n11089), .B1(n1811), .B2(n11086), .C1(n1233), .C2(n11083), .ZN(n5150) );
  OAI222_X1 U6465 ( .A1(n947), .A2(n11353), .B1(n1811), .B2(n11350), .C1(n1233), .C2(n11347), .ZN(n3717) );
  OAI222_X1 U6466 ( .A1(n943), .A2(n11089), .B1(n1807), .B2(n11086), .C1(n1221), .C2(n11083), .ZN(n5109) );
  OAI222_X1 U6467 ( .A1(n943), .A2(n11353), .B1(n1807), .B2(n11350), .C1(n1221), .C2(n11347), .ZN(n3676) );
  OAI222_X1 U6468 ( .A1(n939), .A2(n11089), .B1(n1803), .B2(n11086), .C1(n1209), .C2(n11083), .ZN(n5068) );
  OAI222_X1 U6469 ( .A1(n939), .A2(n11353), .B1(n1803), .B2(n11350), .C1(n1209), .C2(n11347), .ZN(n3635) );
  OAI222_X1 U6470 ( .A1(n935), .A2(n11089), .B1(n1799), .B2(n11086), .C1(n1197), .C2(n11083), .ZN(n5027) );
  OAI222_X1 U6471 ( .A1(n935), .A2(n11353), .B1(n1799), .B2(n11350), .C1(n1197), .C2(n11347), .ZN(n3594) );
  OAI222_X1 U6472 ( .A1(n931), .A2(n11089), .B1(n1795), .B2(n11086), .C1(n1185), .C2(n11083), .ZN(n4986) );
  OAI222_X1 U6473 ( .A1(n931), .A2(n11353), .B1(n1795), .B2(n11350), .C1(n1185), .C2(n11347), .ZN(n3553) );
  OAI222_X1 U6474 ( .A1(n927), .A2(n11089), .B1(n1791), .B2(n11086), .C1(n1173), .C2(n11083), .ZN(n4945) );
  OAI222_X1 U6475 ( .A1(n927), .A2(n11353), .B1(n1791), .B2(n11350), .C1(n1173), .C2(n11347), .ZN(n3512) );
  OAI222_X1 U6476 ( .A1(n923), .A2(n11089), .B1(n1787), .B2(n11086), .C1(n1161), .C2(n11083), .ZN(n4904) );
  OAI222_X1 U6477 ( .A1(n923), .A2(n11353), .B1(n1787), .B2(n11350), .C1(n1161), .C2(n11347), .ZN(n3471) );
  OAI222_X1 U6478 ( .A1(n919), .A2(n11089), .B1(n1783), .B2(n11086), .C1(n1149), .C2(n11083), .ZN(n4863) );
  OAI222_X1 U6479 ( .A1(n919), .A2(n11353), .B1(n1783), .B2(n11350), .C1(n1149), .C2(n11347), .ZN(n3430) );
  OAI222_X1 U6480 ( .A1(n915), .A2(n11089), .B1(n1779), .B2(n11086), .C1(n1137), .C2(n11083), .ZN(n4822) );
  OAI222_X1 U6481 ( .A1(n915), .A2(n11353), .B1(n1779), .B2(n11350), .C1(n1137), .C2(n11347), .ZN(n3389) );
  OAI222_X1 U6482 ( .A1(n911), .A2(n11089), .B1(n1775), .B2(n11086), .C1(n1125), .C2(n11083), .ZN(n4781) );
  OAI222_X1 U6483 ( .A1(n911), .A2(n11353), .B1(n1775), .B2(n11350), .C1(n1125), .C2(n11347), .ZN(n3348) );
  OAI222_X1 U6484 ( .A1(n907), .A2(n11089), .B1(n1771), .B2(n11086), .C1(n1113), .C2(n11083), .ZN(n4740) );
  OAI222_X1 U6485 ( .A1(n907), .A2(n11353), .B1(n1771), .B2(n11350), .C1(n1113), .C2(n11347), .ZN(n3307) );
  OAI222_X1 U6486 ( .A1(n903), .A2(n11089), .B1(n1767), .B2(n11086), .C1(n1101), .C2(n11083), .ZN(n4699) );
  OAI222_X1 U6487 ( .A1(n903), .A2(n11353), .B1(n1767), .B2(n11350), .C1(n1101), .C2(n11347), .ZN(n3266) );
  OAI222_X1 U6488 ( .A1(n899), .A2(n11090), .B1(n1763), .B2(n11087), .C1(n1089), .C2(n11084), .ZN(n4658) );
  OAI222_X1 U6489 ( .A1(n899), .A2(n11354), .B1(n1763), .B2(n11351), .C1(n1089), .C2(n11348), .ZN(n3225) );
  OAI222_X1 U6490 ( .A1(n895), .A2(n11090), .B1(n1759), .B2(n11087), .C1(n1077), .C2(n11084), .ZN(n4617) );
  OAI222_X1 U6491 ( .A1(n895), .A2(n11354), .B1(n1759), .B2(n11351), .C1(n1077), .C2(n11348), .ZN(n3184) );
  OAI222_X1 U6492 ( .A1(n891), .A2(n11090), .B1(n1755), .B2(n11087), .C1(n1065), .C2(n11084), .ZN(n4576) );
  OAI222_X1 U6493 ( .A1(n891), .A2(n11354), .B1(n1755), .B2(n11351), .C1(n1065), .C2(n11348), .ZN(n3143) );
  OAI222_X1 U6494 ( .A1(n887), .A2(n11090), .B1(n1751), .B2(n11087), .C1(n1053), .C2(n11084), .ZN(n4535) );
  OAI222_X1 U6495 ( .A1(n887), .A2(n11354), .B1(n1751), .B2(n11351), .C1(n1053), .C2(n11348), .ZN(n3102) );
  OAI222_X1 U6496 ( .A1(n883), .A2(n11090), .B1(n1747), .B2(n11087), .C1(n1041), .C2(n11084), .ZN(n4494) );
  OAI222_X1 U6497 ( .A1(n883), .A2(n11354), .B1(n1747), .B2(n11351), .C1(n1041), .C2(n11348), .ZN(n3061) );
  OAI222_X1 U6498 ( .A1(n879), .A2(n11090), .B1(n1743), .B2(n11087), .C1(n1029), .C2(n11084), .ZN(n4453) );
  OAI222_X1 U6499 ( .A1(n879), .A2(n11354), .B1(n1743), .B2(n11351), .C1(n1029), .C2(n11348), .ZN(n3020) );
  OAI222_X1 U6500 ( .A1(n875), .A2(n11090), .B1(n1739), .B2(n11087), .C1(
        n12787), .C2(n11084), .ZN(n4412) );
  OAI222_X1 U6501 ( .A1(n875), .A2(n11354), .B1(n1739), .B2(n11351), .C1(
        n12787), .C2(n11348), .ZN(n2979) );
  OAI222_X1 U6502 ( .A1(n871), .A2(n11090), .B1(n1735), .B2(n11087), .C1(
        n12786), .C2(n11084), .ZN(n4283) );
  OAI222_X1 U6503 ( .A1(n871), .A2(n11354), .B1(n1735), .B2(n11351), .C1(
        n12786), .C2(n11348), .ZN(n2751) );
  AOI222_X1 U6504 ( .A1(n10923), .A2(n9376), .B1(n10920), .B2(n9312), .C1(
        n10917), .C2(n9344), .ZN(n5679) );
  AOI222_X1 U6505 ( .A1(n11187), .A2(n9376), .B1(n11184), .B2(n9312), .C1(
        n11181), .C2(n9344), .ZN(n4246) );
  AOI222_X1 U6506 ( .A1(n10923), .A2(n9377), .B1(n10920), .B2(n9313), .C1(
        n10917), .C2(n9345), .ZN(n5615) );
  AOI222_X1 U6507 ( .A1(n11187), .A2(n9377), .B1(n11184), .B2(n9313), .C1(
        n11181), .C2(n9345), .ZN(n4182) );
  AOI222_X1 U6508 ( .A1(n10923), .A2(n9378), .B1(n10920), .B2(n9314), .C1(
        n10917), .C2(n9346), .ZN(n5574) );
  AOI222_X1 U6509 ( .A1(n11187), .A2(n9378), .B1(n11184), .B2(n9314), .C1(
        n11181), .C2(n9346), .ZN(n4141) );
  AOI222_X1 U6510 ( .A1(n10923), .A2(n9379), .B1(n10920), .B2(n9315), .C1(
        n10917), .C2(n9347), .ZN(n5533) );
  AOI222_X1 U6511 ( .A1(n11187), .A2(n9379), .B1(n11184), .B2(n9315), .C1(
        n11181), .C2(n9347), .ZN(n4100) );
  AOI222_X1 U6512 ( .A1(n10923), .A2(n9380), .B1(n10920), .B2(n9316), .C1(
        n10917), .C2(n9348), .ZN(n5492) );
  AOI222_X1 U6513 ( .A1(n11187), .A2(n9380), .B1(n11184), .B2(n9316), .C1(
        n11181), .C2(n9348), .ZN(n4059) );
  AOI222_X1 U6514 ( .A1(n10923), .A2(n9381), .B1(n10920), .B2(n9317), .C1(
        n10917), .C2(n9349), .ZN(n5451) );
  AOI222_X1 U6515 ( .A1(n11187), .A2(n9381), .B1(n11184), .B2(n9317), .C1(
        n11181), .C2(n9349), .ZN(n4018) );
  AOI222_X1 U6516 ( .A1(n10923), .A2(n9382), .B1(n10920), .B2(n9318), .C1(
        n10917), .C2(n9350), .ZN(n5410) );
  AOI222_X1 U6517 ( .A1(n11187), .A2(n9382), .B1(n11184), .B2(n9318), .C1(
        n11181), .C2(n9350), .ZN(n3977) );
  AOI222_X1 U6518 ( .A1(n10923), .A2(n9383), .B1(n10920), .B2(n9319), .C1(
        n10917), .C2(n9351), .ZN(n5369) );
  AOI222_X1 U6519 ( .A1(n11187), .A2(n9383), .B1(n11184), .B2(n9319), .C1(
        n11181), .C2(n9351), .ZN(n3936) );
  AOI222_X1 U6520 ( .A1(n10923), .A2(n9384), .B1(n10920), .B2(n9320), .C1(
        n10917), .C2(n9352), .ZN(n5328) );
  AOI222_X1 U6521 ( .A1(n11187), .A2(n9384), .B1(n11184), .B2(n9320), .C1(
        n11181), .C2(n9352), .ZN(n3895) );
  AOI222_X1 U6522 ( .A1(n10923), .A2(n9385), .B1(n10920), .B2(n9321), .C1(
        n10917), .C2(n9353), .ZN(n5287) );
  AOI222_X1 U6523 ( .A1(n11187), .A2(n9385), .B1(n11184), .B2(n9321), .C1(
        n11181), .C2(n9353), .ZN(n3854) );
  AOI222_X1 U6524 ( .A1(n10923), .A2(n9386), .B1(n10920), .B2(n9322), .C1(
        n10917), .C2(n9354), .ZN(n5246) );
  AOI222_X1 U6525 ( .A1(n11187), .A2(n9386), .B1(n11184), .B2(n9322), .C1(
        n11181), .C2(n9354), .ZN(n3813) );
  AOI222_X1 U6526 ( .A1(n10923), .A2(n9387), .B1(n10920), .B2(n9323), .C1(
        n10917), .C2(n9355), .ZN(n5205) );
  AOI222_X1 U6527 ( .A1(n11187), .A2(n9387), .B1(n11184), .B2(n9323), .C1(
        n11181), .C2(n9355), .ZN(n3772) );
  AOI222_X1 U6528 ( .A1(n10924), .A2(n9388), .B1(n10921), .B2(n9324), .C1(
        n10918), .C2(n9356), .ZN(n5164) );
  AOI222_X1 U6529 ( .A1(n11188), .A2(n9388), .B1(n11185), .B2(n9324), .C1(
        n11182), .C2(n9356), .ZN(n3731) );
  AOI222_X1 U6530 ( .A1(n10924), .A2(n9389), .B1(n10921), .B2(n9325), .C1(
        n10918), .C2(n9357), .ZN(n5123) );
  AOI222_X1 U6531 ( .A1(n11188), .A2(n9389), .B1(n11185), .B2(n9325), .C1(
        n11182), .C2(n9357), .ZN(n3690) );
  AOI222_X1 U6532 ( .A1(n10924), .A2(n9390), .B1(n10921), .B2(n9326), .C1(
        n10918), .C2(n9358), .ZN(n5082) );
  AOI222_X1 U6533 ( .A1(n11188), .A2(n9390), .B1(n11185), .B2(n9326), .C1(
        n11182), .C2(n9358), .ZN(n3649) );
  AOI222_X1 U6534 ( .A1(n10924), .A2(n9391), .B1(n10921), .B2(n9327), .C1(
        n10918), .C2(n9359), .ZN(n5041) );
  AOI222_X1 U6535 ( .A1(n11188), .A2(n9391), .B1(n11185), .B2(n9327), .C1(
        n11182), .C2(n9359), .ZN(n3608) );
  AOI222_X1 U6536 ( .A1(n10924), .A2(n9392), .B1(n10921), .B2(n9328), .C1(
        n10918), .C2(n9360), .ZN(n5000) );
  AOI222_X1 U6537 ( .A1(n11188), .A2(n9392), .B1(n11185), .B2(n9328), .C1(
        n11182), .C2(n9360), .ZN(n3567) );
  AOI222_X1 U6538 ( .A1(n10924), .A2(n9393), .B1(n10921), .B2(n9329), .C1(
        n10918), .C2(n9361), .ZN(n4959) );
  AOI222_X1 U6539 ( .A1(n11188), .A2(n9393), .B1(n11185), .B2(n9329), .C1(
        n11182), .C2(n9361), .ZN(n3526) );
  AOI222_X1 U6540 ( .A1(n10924), .A2(n9394), .B1(n10921), .B2(n9330), .C1(
        n10918), .C2(n9362), .ZN(n4918) );
  AOI222_X1 U6541 ( .A1(n11188), .A2(n9394), .B1(n11185), .B2(n9330), .C1(
        n11182), .C2(n9362), .ZN(n3485) );
  AOI222_X1 U6542 ( .A1(n10924), .A2(n9395), .B1(n10921), .B2(n9331), .C1(
        n10918), .C2(n9363), .ZN(n4877) );
  AOI222_X1 U6543 ( .A1(n11188), .A2(n9395), .B1(n11185), .B2(n9331), .C1(
        n11182), .C2(n9363), .ZN(n3444) );
  AOI222_X1 U6544 ( .A1(n10924), .A2(n9396), .B1(n10921), .B2(n9332), .C1(
        n10918), .C2(n9364), .ZN(n4836) );
  AOI222_X1 U6545 ( .A1(n11188), .A2(n9396), .B1(n11185), .B2(n9332), .C1(
        n11182), .C2(n9364), .ZN(n3403) );
  AOI222_X1 U6546 ( .A1(n10924), .A2(n9397), .B1(n10921), .B2(n9333), .C1(
        n10918), .C2(n9365), .ZN(n4795) );
  AOI222_X1 U6547 ( .A1(n11188), .A2(n9397), .B1(n11185), .B2(n9333), .C1(
        n11182), .C2(n9365), .ZN(n3362) );
  AOI222_X1 U6548 ( .A1(n10924), .A2(n9398), .B1(n10921), .B2(n9334), .C1(
        n10918), .C2(n9366), .ZN(n4754) );
  AOI222_X1 U6549 ( .A1(n11188), .A2(n9398), .B1(n11185), .B2(n9334), .C1(
        n11182), .C2(n9366), .ZN(n3321) );
  AOI222_X1 U6550 ( .A1(n10924), .A2(n9399), .B1(n10921), .B2(n9335), .C1(
        n10918), .C2(n9367), .ZN(n4713) );
  AOI222_X1 U6551 ( .A1(n11188), .A2(n9399), .B1(n11185), .B2(n9335), .C1(
        n11182), .C2(n9367), .ZN(n3280) );
  AOI222_X1 U6552 ( .A1(n10925), .A2(n9400), .B1(n10922), .B2(n9336), .C1(
        n10919), .C2(n9368), .ZN(n4672) );
  AOI222_X1 U6553 ( .A1(n11189), .A2(n9400), .B1(n11186), .B2(n9336), .C1(
        n11183), .C2(n9368), .ZN(n3239) );
  AOI222_X1 U6554 ( .A1(n10925), .A2(n9401), .B1(n10922), .B2(n9337), .C1(
        n10919), .C2(n9369), .ZN(n4631) );
  AOI222_X1 U6555 ( .A1(n11189), .A2(n9401), .B1(n11186), .B2(n9337), .C1(
        n11183), .C2(n9369), .ZN(n3198) );
  AOI222_X1 U6556 ( .A1(n10925), .A2(n9402), .B1(n10922), .B2(n9338), .C1(
        n10919), .C2(n9370), .ZN(n4590) );
  AOI222_X1 U6557 ( .A1(n11189), .A2(n9402), .B1(n11186), .B2(n9338), .C1(
        n11183), .C2(n9370), .ZN(n3157) );
  AOI222_X1 U6558 ( .A1(n10925), .A2(n9403), .B1(n10922), .B2(n9339), .C1(
        n10919), .C2(n9371), .ZN(n4549) );
  AOI222_X1 U6559 ( .A1(n11189), .A2(n9403), .B1(n11186), .B2(n9339), .C1(
        n11183), .C2(n9371), .ZN(n3116) );
  AOI222_X1 U6560 ( .A1(n10925), .A2(n9404), .B1(n10922), .B2(n9340), .C1(
        n10919), .C2(n9372), .ZN(n4508) );
  AOI222_X1 U6561 ( .A1(n11189), .A2(n9404), .B1(n11186), .B2(n9340), .C1(
        n11183), .C2(n9372), .ZN(n3075) );
  AOI222_X1 U6562 ( .A1(n10925), .A2(n9405), .B1(n10922), .B2(n9341), .C1(
        n10919), .C2(n9373), .ZN(n4467) );
  AOI222_X1 U6563 ( .A1(n11189), .A2(n9405), .B1(n11186), .B2(n9341), .C1(
        n11183), .C2(n9373), .ZN(n3034) );
  AOI222_X1 U6564 ( .A1(n10925), .A2(n9406), .B1(n10922), .B2(n9342), .C1(
        n10919), .C2(n9374), .ZN(n4426) );
  AOI222_X1 U6565 ( .A1(n11189), .A2(n9406), .B1(n11186), .B2(n9342), .C1(
        n11183), .C2(n9374), .ZN(n2993) );
  AOI222_X1 U6566 ( .A1(n10925), .A2(n9407), .B1(n10922), .B2(n9343), .C1(
        n10919), .C2(n9375), .ZN(n4341) );
  AOI222_X1 U6567 ( .A1(n11189), .A2(n9407), .B1(n11186), .B2(n9343), .C1(
        n11183), .C2(n9375), .ZN(n2873) );
  NOR4_X1 U6568 ( .A1(n5683), .A2(n5684), .A3(n5685), .A4(n5686), .ZN(n5682)
         );
  OAI22_X1 U6569 ( .A1(n10521), .A2(n10980), .B1(n10520), .B2(n10977), .ZN(
        n5686) );
  OAI222_X1 U6570 ( .A1(n13939), .A2(n10956), .B1(n13875), .B2(n10953), .C1(
        n13907), .C2(n10950), .ZN(n5683) );
  OAI222_X1 U6571 ( .A1(n10515), .A2(n10965), .B1(n10514), .B2(n10962), .C1(
        n10516), .C2(n10959), .ZN(n5684) );
  NOR4_X1 U6572 ( .A1(n5697), .A2(n5698), .A3(n5699), .A4(n5700), .ZN(n5696)
         );
  OAI22_X1 U6573 ( .A1(n13971), .A2(n10914), .B1(n14003), .B2(n10911), .ZN(
        n5700) );
  OAI222_X1 U6574 ( .A1(n992), .A2(n10890), .B1(n14256), .B2(n10887), .C1(
        n14224), .C2(n10884), .ZN(n5697) );
  OAI222_X1 U6575 ( .A1(n14161), .A2(n10899), .B1(n14193), .B2(n10896), .C1(
        n14129), .C2(n10893), .ZN(n5698) );
  NOR4_X1 U6576 ( .A1(n4250), .A2(n4251), .A3(n4252), .A4(n4253), .ZN(n4249)
         );
  OAI22_X1 U6577 ( .A1(n10521), .A2(n11244), .B1(n10520), .B2(n11241), .ZN(
        n4253) );
  OAI222_X1 U6578 ( .A1(n13939), .A2(n11220), .B1(n13875), .B2(n11217), .C1(
        n13907), .C2(n11214), .ZN(n4250) );
  OAI222_X1 U6579 ( .A1(n10515), .A2(n11229), .B1(n10514), .B2(n11226), .C1(
        n10516), .C2(n11223), .ZN(n4251) );
  NOR4_X1 U6580 ( .A1(n4264), .A2(n4265), .A3(n4266), .A4(n4267), .ZN(n4263)
         );
  OAI22_X1 U6581 ( .A1(n13971), .A2(n11178), .B1(n14003), .B2(n11175), .ZN(
        n4267) );
  OAI222_X1 U6582 ( .A1(n992), .A2(n11154), .B1(n14256), .B2(n11151), .C1(
        n14224), .C2(n11148), .ZN(n4264) );
  OAI222_X1 U6583 ( .A1(n14161), .A2(n11163), .B1(n14193), .B2(n11160), .C1(
        n14129), .C2(n11157), .ZN(n4265) );
  NOR4_X1 U6584 ( .A1(n5619), .A2(n5620), .A3(n5621), .A4(n5622), .ZN(n5618)
         );
  OAI22_X1 U6585 ( .A1(n10489), .A2(n10980), .B1(n10488), .B2(n10977), .ZN(
        n5622) );
  OAI222_X1 U6586 ( .A1(n13938), .A2(n10956), .B1(n13874), .B2(n10953), .C1(
        n13906), .C2(n10950), .ZN(n5619) );
  OAI222_X1 U6587 ( .A1(n10483), .A2(n10965), .B1(n10482), .B2(n10962), .C1(
        n10484), .C2(n10959), .ZN(n5620) );
  NOR4_X1 U6588 ( .A1(n5628), .A2(n5629), .A3(n5630), .A4(n5631), .ZN(n5627)
         );
  OAI22_X1 U6589 ( .A1(n13970), .A2(n10914), .B1(n14002), .B2(n10911), .ZN(
        n5631) );
  OAI222_X1 U6590 ( .A1(n988), .A2(n10890), .B1(n14255), .B2(n10887), .C1(
        n14223), .C2(n10884), .ZN(n5628) );
  OAI222_X1 U6591 ( .A1(n14160), .A2(n10899), .B1(n14192), .B2(n10896), .C1(
        n14128), .C2(n10893), .ZN(n5629) );
  NOR4_X1 U6592 ( .A1(n4186), .A2(n4187), .A3(n4188), .A4(n4189), .ZN(n4185)
         );
  OAI22_X1 U6593 ( .A1(n10489), .A2(n11244), .B1(n10488), .B2(n11241), .ZN(
        n4189) );
  OAI222_X1 U6594 ( .A1(n13938), .A2(n11220), .B1(n13874), .B2(n11217), .C1(
        n13906), .C2(n11214), .ZN(n4186) );
  OAI222_X1 U6595 ( .A1(n10483), .A2(n11229), .B1(n10482), .B2(n11226), .C1(
        n10484), .C2(n11223), .ZN(n4187) );
  NOR4_X1 U6596 ( .A1(n4195), .A2(n4196), .A3(n4197), .A4(n4198), .ZN(n4194)
         );
  OAI22_X1 U6597 ( .A1(n13970), .A2(n11178), .B1(n14002), .B2(n11175), .ZN(
        n4198) );
  OAI222_X1 U6598 ( .A1(n988), .A2(n11154), .B1(n14255), .B2(n11151), .C1(
        n14223), .C2(n11148), .ZN(n4195) );
  OAI222_X1 U6599 ( .A1(n14160), .A2(n11163), .B1(n14192), .B2(n11160), .C1(
        n14128), .C2(n11157), .ZN(n4196) );
  NOR4_X1 U6600 ( .A1(n5578), .A2(n5579), .A3(n5580), .A4(n5581), .ZN(n5577)
         );
  OAI22_X1 U6601 ( .A1(n10457), .A2(n10980), .B1(n10456), .B2(n10977), .ZN(
        n5581) );
  OAI222_X1 U6602 ( .A1(n13937), .A2(n10956), .B1(n13873), .B2(n10953), .C1(
        n13905), .C2(n10950), .ZN(n5578) );
  OAI222_X1 U6603 ( .A1(n10451), .A2(n10965), .B1(n10450), .B2(n10962), .C1(
        n10452), .C2(n10959), .ZN(n5579) );
  NOR4_X1 U6604 ( .A1(n5587), .A2(n5588), .A3(n5589), .A4(n5590), .ZN(n5586)
         );
  OAI22_X1 U6605 ( .A1(n13969), .A2(n10914), .B1(n14001), .B2(n10911), .ZN(
        n5590) );
  OAI222_X1 U6606 ( .A1(n984), .A2(n10890), .B1(n14254), .B2(n10887), .C1(
        n14222), .C2(n10884), .ZN(n5587) );
  OAI222_X1 U6607 ( .A1(n14159), .A2(n10899), .B1(n14191), .B2(n10896), .C1(
        n14127), .C2(n10893), .ZN(n5588) );
  NOR4_X1 U6608 ( .A1(n4145), .A2(n4146), .A3(n4147), .A4(n4148), .ZN(n4144)
         );
  OAI22_X1 U6609 ( .A1(n10457), .A2(n11244), .B1(n10456), .B2(n11241), .ZN(
        n4148) );
  OAI222_X1 U6610 ( .A1(n13937), .A2(n11220), .B1(n13873), .B2(n11217), .C1(
        n13905), .C2(n11214), .ZN(n4145) );
  OAI222_X1 U6611 ( .A1(n10451), .A2(n11229), .B1(n10450), .B2(n11226), .C1(
        n10452), .C2(n11223), .ZN(n4146) );
  NOR4_X1 U6612 ( .A1(n4154), .A2(n4155), .A3(n4156), .A4(n4157), .ZN(n4153)
         );
  OAI22_X1 U6613 ( .A1(n13969), .A2(n11178), .B1(n14001), .B2(n11175), .ZN(
        n4157) );
  OAI222_X1 U6614 ( .A1(n984), .A2(n11154), .B1(n14254), .B2(n11151), .C1(
        n14222), .C2(n11148), .ZN(n4154) );
  OAI222_X1 U6615 ( .A1(n14159), .A2(n11163), .B1(n14191), .B2(n11160), .C1(
        n14127), .C2(n11157), .ZN(n4155) );
  NOR4_X1 U6616 ( .A1(n5537), .A2(n5538), .A3(n5539), .A4(n5540), .ZN(n5536)
         );
  OAI22_X1 U6617 ( .A1(n10425), .A2(n10980), .B1(n10424), .B2(n10977), .ZN(
        n5540) );
  OAI222_X1 U6618 ( .A1(n13936), .A2(n10956), .B1(n13872), .B2(n10953), .C1(
        n13904), .C2(n10950), .ZN(n5537) );
  OAI222_X1 U6619 ( .A1(n10419), .A2(n10965), .B1(n10418), .B2(n10962), .C1(
        n10420), .C2(n10959), .ZN(n5538) );
  NOR4_X1 U6620 ( .A1(n5546), .A2(n5547), .A3(n5548), .A4(n5549), .ZN(n5545)
         );
  OAI22_X1 U6621 ( .A1(n13968), .A2(n10914), .B1(n14000), .B2(n10911), .ZN(
        n5549) );
  OAI222_X1 U6622 ( .A1(n980), .A2(n10890), .B1(n14253), .B2(n10887), .C1(
        n14221), .C2(n10884), .ZN(n5546) );
  OAI222_X1 U6623 ( .A1(n14158), .A2(n10899), .B1(n14190), .B2(n10896), .C1(
        n14126), .C2(n10893), .ZN(n5547) );
  NOR4_X1 U6624 ( .A1(n4104), .A2(n4105), .A3(n4106), .A4(n4107), .ZN(n4103)
         );
  OAI22_X1 U6625 ( .A1(n10425), .A2(n11244), .B1(n10424), .B2(n11241), .ZN(
        n4107) );
  OAI222_X1 U6626 ( .A1(n13936), .A2(n11220), .B1(n13872), .B2(n11217), .C1(
        n13904), .C2(n11214), .ZN(n4104) );
  OAI222_X1 U6627 ( .A1(n10419), .A2(n11229), .B1(n10418), .B2(n11226), .C1(
        n10420), .C2(n11223), .ZN(n4105) );
  NOR4_X1 U6628 ( .A1(n4113), .A2(n4114), .A3(n4115), .A4(n4116), .ZN(n4112)
         );
  OAI22_X1 U6629 ( .A1(n13968), .A2(n11178), .B1(n14000), .B2(n11175), .ZN(
        n4116) );
  OAI222_X1 U6630 ( .A1(n980), .A2(n11154), .B1(n14253), .B2(n11151), .C1(
        n14221), .C2(n11148), .ZN(n4113) );
  OAI222_X1 U6631 ( .A1(n14158), .A2(n11163), .B1(n14190), .B2(n11160), .C1(
        n14126), .C2(n11157), .ZN(n4114) );
  NOR4_X1 U6632 ( .A1(n5496), .A2(n5497), .A3(n5498), .A4(n5499), .ZN(n5495)
         );
  OAI22_X1 U6633 ( .A1(n10390), .A2(n10980), .B1(n10389), .B2(n10977), .ZN(
        n5499) );
  OAI222_X1 U6634 ( .A1(n13935), .A2(n10956), .B1(n13871), .B2(n10953), .C1(
        n13903), .C2(n10950), .ZN(n5496) );
  OAI222_X1 U6635 ( .A1(n10384), .A2(n10965), .B1(n10383), .B2(n10962), .C1(
        n10385), .C2(n10959), .ZN(n5497) );
  NOR4_X1 U6636 ( .A1(n5505), .A2(n5506), .A3(n5507), .A4(n5508), .ZN(n5504)
         );
  OAI22_X1 U6637 ( .A1(n13967), .A2(n10914), .B1(n13999), .B2(n10911), .ZN(
        n5508) );
  OAI222_X1 U6638 ( .A1(n976), .A2(n10890), .B1(n14252), .B2(n10887), .C1(
        n14220), .C2(n10884), .ZN(n5505) );
  OAI222_X1 U6639 ( .A1(n14157), .A2(n10899), .B1(n14189), .B2(n10896), .C1(
        n14125), .C2(n10893), .ZN(n5506) );
  NOR4_X1 U6640 ( .A1(n4063), .A2(n4064), .A3(n4065), .A4(n4066), .ZN(n4062)
         );
  OAI22_X1 U6641 ( .A1(n10390), .A2(n11244), .B1(n10389), .B2(n11241), .ZN(
        n4066) );
  OAI222_X1 U6642 ( .A1(n13935), .A2(n11220), .B1(n13871), .B2(n11217), .C1(
        n13903), .C2(n11214), .ZN(n4063) );
  OAI222_X1 U6643 ( .A1(n10384), .A2(n11229), .B1(n10383), .B2(n11226), .C1(
        n10385), .C2(n11223), .ZN(n4064) );
  NOR4_X1 U6644 ( .A1(n4072), .A2(n4073), .A3(n4074), .A4(n4075), .ZN(n4071)
         );
  OAI22_X1 U6645 ( .A1(n13967), .A2(n11178), .B1(n13999), .B2(n11175), .ZN(
        n4075) );
  OAI222_X1 U6646 ( .A1(n976), .A2(n11154), .B1(n14252), .B2(n11151), .C1(
        n14220), .C2(n11148), .ZN(n4072) );
  OAI222_X1 U6647 ( .A1(n14157), .A2(n11163), .B1(n14189), .B2(n11160), .C1(
        n14125), .C2(n11157), .ZN(n4073) );
  NOR4_X1 U6648 ( .A1(n5455), .A2(n5456), .A3(n5457), .A4(n5458), .ZN(n5454)
         );
  OAI22_X1 U6649 ( .A1(n10358), .A2(n10980), .B1(n10357), .B2(n10977), .ZN(
        n5458) );
  OAI222_X1 U6650 ( .A1(n13934), .A2(n10956), .B1(n13870), .B2(n10953), .C1(
        n13902), .C2(n10950), .ZN(n5455) );
  OAI222_X1 U6651 ( .A1(n10352), .A2(n10965), .B1(n10351), .B2(n10962), .C1(
        n10353), .C2(n10959), .ZN(n5456) );
  NOR4_X1 U6652 ( .A1(n5464), .A2(n5465), .A3(n5466), .A4(n5467), .ZN(n5463)
         );
  OAI22_X1 U6653 ( .A1(n13966), .A2(n10914), .B1(n13998), .B2(n10911), .ZN(
        n5467) );
  OAI222_X1 U6654 ( .A1(n972), .A2(n10890), .B1(n14251), .B2(n10887), .C1(
        n14219), .C2(n10884), .ZN(n5464) );
  OAI222_X1 U6655 ( .A1(n14156), .A2(n10899), .B1(n14188), .B2(n10896), .C1(
        n14124), .C2(n10893), .ZN(n5465) );
  NOR4_X1 U6656 ( .A1(n4022), .A2(n4023), .A3(n4024), .A4(n4025), .ZN(n4021)
         );
  OAI22_X1 U6657 ( .A1(n10358), .A2(n11244), .B1(n10357), .B2(n11241), .ZN(
        n4025) );
  OAI222_X1 U6658 ( .A1(n13934), .A2(n11220), .B1(n13870), .B2(n11217), .C1(
        n13902), .C2(n11214), .ZN(n4022) );
  OAI222_X1 U6659 ( .A1(n10352), .A2(n11229), .B1(n10351), .B2(n11226), .C1(
        n10353), .C2(n11223), .ZN(n4023) );
  NOR4_X1 U6660 ( .A1(n4031), .A2(n4032), .A3(n4033), .A4(n4034), .ZN(n4030)
         );
  OAI22_X1 U6661 ( .A1(n13966), .A2(n11178), .B1(n13998), .B2(n11175), .ZN(
        n4034) );
  OAI222_X1 U6662 ( .A1(n972), .A2(n11154), .B1(n14251), .B2(n11151), .C1(
        n14219), .C2(n11148), .ZN(n4031) );
  OAI222_X1 U6663 ( .A1(n14156), .A2(n11163), .B1(n14188), .B2(n11160), .C1(
        n14124), .C2(n11157), .ZN(n4032) );
  NOR4_X1 U6664 ( .A1(n5414), .A2(n5415), .A3(n5416), .A4(n5417), .ZN(n5413)
         );
  OAI22_X1 U6665 ( .A1(n10326), .A2(n10980), .B1(n10325), .B2(n10977), .ZN(
        n5417) );
  OAI222_X1 U6666 ( .A1(n13933), .A2(n10956), .B1(n13869), .B2(n10953), .C1(
        n13901), .C2(n10950), .ZN(n5414) );
  OAI222_X1 U6667 ( .A1(n10320), .A2(n10965), .B1(n10319), .B2(n10962), .C1(
        n10321), .C2(n10959), .ZN(n5415) );
  NOR4_X1 U6668 ( .A1(n5423), .A2(n5424), .A3(n5425), .A4(n5426), .ZN(n5422)
         );
  OAI22_X1 U6669 ( .A1(n13965), .A2(n10914), .B1(n13997), .B2(n10911), .ZN(
        n5426) );
  OAI222_X1 U6670 ( .A1(n968), .A2(n10890), .B1(n14250), .B2(n10887), .C1(
        n14218), .C2(n10884), .ZN(n5423) );
  OAI222_X1 U6671 ( .A1(n14155), .A2(n10899), .B1(n14187), .B2(n10896), .C1(
        n14123), .C2(n10893), .ZN(n5424) );
  NOR4_X1 U6672 ( .A1(n3981), .A2(n3982), .A3(n3983), .A4(n3984), .ZN(n3980)
         );
  OAI22_X1 U6673 ( .A1(n10326), .A2(n11244), .B1(n10325), .B2(n11241), .ZN(
        n3984) );
  OAI222_X1 U6674 ( .A1(n13933), .A2(n11220), .B1(n13869), .B2(n11217), .C1(
        n13901), .C2(n11214), .ZN(n3981) );
  OAI222_X1 U6675 ( .A1(n10320), .A2(n11229), .B1(n10319), .B2(n11226), .C1(
        n10321), .C2(n11223), .ZN(n3982) );
  NOR4_X1 U6676 ( .A1(n3990), .A2(n3991), .A3(n3992), .A4(n3993), .ZN(n3989)
         );
  OAI22_X1 U6677 ( .A1(n13965), .A2(n11178), .B1(n13997), .B2(n11175), .ZN(
        n3993) );
  OAI222_X1 U6678 ( .A1(n968), .A2(n11154), .B1(n14250), .B2(n11151), .C1(
        n14218), .C2(n11148), .ZN(n3990) );
  OAI222_X1 U6679 ( .A1(n14155), .A2(n11163), .B1(n14187), .B2(n11160), .C1(
        n14123), .C2(n11157), .ZN(n3991) );
  NOR4_X1 U6680 ( .A1(n5373), .A2(n5374), .A3(n5375), .A4(n5376), .ZN(n5372)
         );
  OAI22_X1 U6681 ( .A1(n10291), .A2(n10980), .B1(n10290), .B2(n10977), .ZN(
        n5376) );
  OAI222_X1 U6682 ( .A1(n13932), .A2(n10956), .B1(n13868), .B2(n10953), .C1(
        n13900), .C2(n10950), .ZN(n5373) );
  OAI222_X1 U6683 ( .A1(n10285), .A2(n10965), .B1(n10284), .B2(n10962), .C1(
        n10286), .C2(n10959), .ZN(n5374) );
  NOR4_X1 U6684 ( .A1(n5382), .A2(n5383), .A3(n5384), .A4(n5385), .ZN(n5381)
         );
  OAI22_X1 U6685 ( .A1(n13964), .A2(n10914), .B1(n13996), .B2(n10911), .ZN(
        n5385) );
  OAI222_X1 U6686 ( .A1(n964), .A2(n10890), .B1(n14249), .B2(n10887), .C1(
        n14217), .C2(n10884), .ZN(n5382) );
  OAI222_X1 U6687 ( .A1(n14154), .A2(n10899), .B1(n14186), .B2(n10896), .C1(
        n14122), .C2(n10893), .ZN(n5383) );
  NOR4_X1 U6688 ( .A1(n3940), .A2(n3941), .A3(n3942), .A4(n3943), .ZN(n3939)
         );
  OAI22_X1 U6689 ( .A1(n10291), .A2(n11244), .B1(n10290), .B2(n11241), .ZN(
        n3943) );
  OAI222_X1 U6690 ( .A1(n13932), .A2(n11220), .B1(n13868), .B2(n11217), .C1(
        n13900), .C2(n11214), .ZN(n3940) );
  OAI222_X1 U6691 ( .A1(n10285), .A2(n11229), .B1(n10284), .B2(n11226), .C1(
        n10286), .C2(n11223), .ZN(n3941) );
  NOR4_X1 U6692 ( .A1(n3949), .A2(n3950), .A3(n3951), .A4(n3952), .ZN(n3948)
         );
  OAI22_X1 U6693 ( .A1(n13964), .A2(n11178), .B1(n13996), .B2(n11175), .ZN(
        n3952) );
  OAI222_X1 U6694 ( .A1(n964), .A2(n11154), .B1(n14249), .B2(n11151), .C1(
        n14217), .C2(n11148), .ZN(n3949) );
  OAI222_X1 U6695 ( .A1(n14154), .A2(n11163), .B1(n14186), .B2(n11160), .C1(
        n14122), .C2(n11157), .ZN(n3950) );
  NOR4_X1 U6696 ( .A1(n5332), .A2(n5333), .A3(n5334), .A4(n5335), .ZN(n5331)
         );
  OAI22_X1 U6697 ( .A1(n10259), .A2(n10980), .B1(n10258), .B2(n10977), .ZN(
        n5335) );
  OAI222_X1 U6698 ( .A1(n13931), .A2(n10956), .B1(n13867), .B2(n10953), .C1(
        n13899), .C2(n10950), .ZN(n5332) );
  OAI222_X1 U6699 ( .A1(n10253), .A2(n10965), .B1(n10252), .B2(n10962), .C1(
        n10254), .C2(n10959), .ZN(n5333) );
  NOR4_X1 U6700 ( .A1(n5341), .A2(n5342), .A3(n5343), .A4(n5344), .ZN(n5340)
         );
  OAI22_X1 U6701 ( .A1(n13963), .A2(n10914), .B1(n13995), .B2(n10911), .ZN(
        n5344) );
  OAI222_X1 U6702 ( .A1(n960), .A2(n10890), .B1(n14248), .B2(n10887), .C1(
        n14216), .C2(n10884), .ZN(n5341) );
  OAI222_X1 U6703 ( .A1(n14153), .A2(n10899), .B1(n14185), .B2(n10896), .C1(
        n14121), .C2(n10893), .ZN(n5342) );
  NOR4_X1 U6704 ( .A1(n3899), .A2(n3900), .A3(n3901), .A4(n3902), .ZN(n3898)
         );
  OAI22_X1 U6705 ( .A1(n10259), .A2(n11244), .B1(n10258), .B2(n11241), .ZN(
        n3902) );
  OAI222_X1 U6706 ( .A1(n13931), .A2(n11220), .B1(n13867), .B2(n11217), .C1(
        n13899), .C2(n11214), .ZN(n3899) );
  OAI222_X1 U6707 ( .A1(n10253), .A2(n11229), .B1(n10252), .B2(n11226), .C1(
        n10254), .C2(n11223), .ZN(n3900) );
  NOR4_X1 U6708 ( .A1(n3908), .A2(n3909), .A3(n3910), .A4(n3911), .ZN(n3907)
         );
  OAI22_X1 U6709 ( .A1(n13963), .A2(n11178), .B1(n13995), .B2(n11175), .ZN(
        n3911) );
  OAI222_X1 U6710 ( .A1(n960), .A2(n11154), .B1(n14248), .B2(n11151), .C1(
        n14216), .C2(n11148), .ZN(n3908) );
  OAI222_X1 U6711 ( .A1(n14153), .A2(n11163), .B1(n14185), .B2(n11160), .C1(
        n14121), .C2(n11157), .ZN(n3909) );
  NOR4_X1 U6712 ( .A1(n5291), .A2(n5292), .A3(n5293), .A4(n5294), .ZN(n5290)
         );
  OAI22_X1 U6713 ( .A1(n10227), .A2(n10980), .B1(n10226), .B2(n10977), .ZN(
        n5294) );
  OAI222_X1 U6714 ( .A1(n13930), .A2(n10956), .B1(n13866), .B2(n10953), .C1(
        n13898), .C2(n10950), .ZN(n5291) );
  OAI222_X1 U6715 ( .A1(n10221), .A2(n10965), .B1(n10220), .B2(n10962), .C1(
        n10222), .C2(n10959), .ZN(n5292) );
  NOR4_X1 U6716 ( .A1(n5300), .A2(n5301), .A3(n5302), .A4(n5303), .ZN(n5299)
         );
  OAI22_X1 U6717 ( .A1(n13962), .A2(n10914), .B1(n13994), .B2(n10911), .ZN(
        n5303) );
  OAI222_X1 U6718 ( .A1(n956), .A2(n10890), .B1(n14247), .B2(n10887), .C1(
        n14215), .C2(n10884), .ZN(n5300) );
  OAI222_X1 U6719 ( .A1(n14152), .A2(n10899), .B1(n14184), .B2(n10896), .C1(
        n14120), .C2(n10893), .ZN(n5301) );
  NOR4_X1 U6720 ( .A1(n3858), .A2(n3859), .A3(n3860), .A4(n3861), .ZN(n3857)
         );
  OAI22_X1 U6721 ( .A1(n10227), .A2(n11244), .B1(n10226), .B2(n11241), .ZN(
        n3861) );
  OAI222_X1 U6722 ( .A1(n13930), .A2(n11220), .B1(n13866), .B2(n11217), .C1(
        n13898), .C2(n11214), .ZN(n3858) );
  OAI222_X1 U6723 ( .A1(n10221), .A2(n11229), .B1(n10220), .B2(n11226), .C1(
        n10222), .C2(n11223), .ZN(n3859) );
  NOR4_X1 U6724 ( .A1(n3867), .A2(n3868), .A3(n3869), .A4(n3870), .ZN(n3866)
         );
  OAI22_X1 U6725 ( .A1(n13962), .A2(n11178), .B1(n13994), .B2(n11175), .ZN(
        n3870) );
  OAI222_X1 U6726 ( .A1(n956), .A2(n11154), .B1(n14247), .B2(n11151), .C1(
        n14215), .C2(n11148), .ZN(n3867) );
  OAI222_X1 U6727 ( .A1(n14152), .A2(n11163), .B1(n14184), .B2(n11160), .C1(
        n14120), .C2(n11157), .ZN(n3868) );
  NOR4_X1 U6728 ( .A1(n5250), .A2(n5251), .A3(n5252), .A4(n5253), .ZN(n5249)
         );
  OAI22_X1 U6729 ( .A1(n10193), .A2(n10980), .B1(n10192), .B2(n10977), .ZN(
        n5253) );
  OAI222_X1 U6730 ( .A1(n13929), .A2(n10956), .B1(n13865), .B2(n10953), .C1(
        n13897), .C2(n10950), .ZN(n5250) );
  OAI222_X1 U6731 ( .A1(n10187), .A2(n10965), .B1(n10186), .B2(n10962), .C1(
        n10188), .C2(n10959), .ZN(n5251) );
  NOR4_X1 U6732 ( .A1(n5259), .A2(n5260), .A3(n5261), .A4(n5262), .ZN(n5258)
         );
  OAI22_X1 U6733 ( .A1(n13961), .A2(n10914), .B1(n13993), .B2(n10911), .ZN(
        n5262) );
  OAI222_X1 U6734 ( .A1(n952), .A2(n10890), .B1(n14246), .B2(n10887), .C1(
        n14214), .C2(n10884), .ZN(n5259) );
  OAI222_X1 U6735 ( .A1(n14151), .A2(n10899), .B1(n14183), .B2(n10896), .C1(
        n14119), .C2(n10893), .ZN(n5260) );
  NOR4_X1 U6736 ( .A1(n3817), .A2(n3818), .A3(n3819), .A4(n3820), .ZN(n3816)
         );
  OAI22_X1 U6737 ( .A1(n10193), .A2(n11244), .B1(n10192), .B2(n11241), .ZN(
        n3820) );
  OAI222_X1 U6738 ( .A1(n13929), .A2(n11220), .B1(n13865), .B2(n11217), .C1(
        n13897), .C2(n11214), .ZN(n3817) );
  OAI222_X1 U6739 ( .A1(n10187), .A2(n11229), .B1(n10186), .B2(n11226), .C1(
        n10188), .C2(n11223), .ZN(n3818) );
  NOR4_X1 U6740 ( .A1(n3826), .A2(n3827), .A3(n3828), .A4(n3829), .ZN(n3825)
         );
  OAI22_X1 U6741 ( .A1(n13961), .A2(n11178), .B1(n13993), .B2(n11175), .ZN(
        n3829) );
  OAI222_X1 U6742 ( .A1(n952), .A2(n11154), .B1(n14246), .B2(n11151), .C1(
        n14214), .C2(n11148), .ZN(n3826) );
  OAI222_X1 U6743 ( .A1(n14151), .A2(n11163), .B1(n14183), .B2(n11160), .C1(
        n14119), .C2(n11157), .ZN(n3827) );
  NOR4_X1 U6744 ( .A1(n5209), .A2(n5210), .A3(n5211), .A4(n5212), .ZN(n5208)
         );
  OAI22_X1 U6745 ( .A1(n10161), .A2(n10980), .B1(n10160), .B2(n10977), .ZN(
        n5212) );
  OAI222_X1 U6746 ( .A1(n13928), .A2(n10956), .B1(n13864), .B2(n10953), .C1(
        n13896), .C2(n10950), .ZN(n5209) );
  OAI222_X1 U6747 ( .A1(n10155), .A2(n10965), .B1(n10154), .B2(n10962), .C1(
        n10156), .C2(n10959), .ZN(n5210) );
  NOR4_X1 U6748 ( .A1(n5218), .A2(n5219), .A3(n5220), .A4(n5221), .ZN(n5217)
         );
  OAI22_X1 U6749 ( .A1(n13960), .A2(n10914), .B1(n13992), .B2(n10911), .ZN(
        n5221) );
  OAI222_X1 U6750 ( .A1(n948), .A2(n10890), .B1(n14245), .B2(n10887), .C1(
        n14213), .C2(n10884), .ZN(n5218) );
  OAI222_X1 U6751 ( .A1(n14150), .A2(n10899), .B1(n14182), .B2(n10896), .C1(
        n14118), .C2(n10893), .ZN(n5219) );
  NOR4_X1 U6752 ( .A1(n3776), .A2(n3777), .A3(n3778), .A4(n3779), .ZN(n3775)
         );
  OAI22_X1 U6753 ( .A1(n10161), .A2(n11244), .B1(n10160), .B2(n11241), .ZN(
        n3779) );
  OAI222_X1 U6754 ( .A1(n13928), .A2(n11220), .B1(n13864), .B2(n11217), .C1(
        n13896), .C2(n11214), .ZN(n3776) );
  OAI222_X1 U6755 ( .A1(n10155), .A2(n11229), .B1(n10154), .B2(n11226), .C1(
        n10156), .C2(n11223), .ZN(n3777) );
  NOR4_X1 U6756 ( .A1(n3785), .A2(n3786), .A3(n3787), .A4(n3788), .ZN(n3784)
         );
  OAI22_X1 U6757 ( .A1(n13960), .A2(n11178), .B1(n13992), .B2(n11175), .ZN(
        n3788) );
  OAI222_X1 U6758 ( .A1(n948), .A2(n11154), .B1(n14245), .B2(n11151), .C1(
        n14213), .C2(n11148), .ZN(n3785) );
  OAI222_X1 U6759 ( .A1(n14150), .A2(n11163), .B1(n14182), .B2(n11160), .C1(
        n14118), .C2(n11157), .ZN(n3786) );
  NOR4_X1 U6760 ( .A1(n5168), .A2(n5169), .A3(n5170), .A4(n5171), .ZN(n5167)
         );
  OAI22_X1 U6761 ( .A1(n10129), .A2(n10981), .B1(n10128), .B2(n10978), .ZN(
        n5171) );
  OAI222_X1 U6762 ( .A1(n13927), .A2(n10957), .B1(n13863), .B2(n10954), .C1(
        n13895), .C2(n10951), .ZN(n5168) );
  OAI222_X1 U6763 ( .A1(n10123), .A2(n10966), .B1(n10122), .B2(n10963), .C1(
        n10124), .C2(n10960), .ZN(n5169) );
  NOR4_X1 U6764 ( .A1(n5177), .A2(n5178), .A3(n5179), .A4(n5180), .ZN(n5176)
         );
  OAI22_X1 U6765 ( .A1(n13959), .A2(n10915), .B1(n13991), .B2(n10912), .ZN(
        n5180) );
  OAI222_X1 U6766 ( .A1(n944), .A2(n10891), .B1(n14244), .B2(n10888), .C1(
        n14212), .C2(n10885), .ZN(n5177) );
  OAI222_X1 U6767 ( .A1(n14149), .A2(n10900), .B1(n14181), .B2(n10897), .C1(
        n14117), .C2(n10894), .ZN(n5178) );
  NOR4_X1 U6768 ( .A1(n3735), .A2(n3736), .A3(n3737), .A4(n3738), .ZN(n3734)
         );
  OAI22_X1 U6769 ( .A1(n10129), .A2(n11245), .B1(n10128), .B2(n11242), .ZN(
        n3738) );
  OAI222_X1 U6770 ( .A1(n13927), .A2(n11221), .B1(n13863), .B2(n11218), .C1(
        n13895), .C2(n11215), .ZN(n3735) );
  OAI222_X1 U6771 ( .A1(n10123), .A2(n11230), .B1(n10122), .B2(n11227), .C1(
        n10124), .C2(n11224), .ZN(n3736) );
  NOR4_X1 U6772 ( .A1(n3744), .A2(n3745), .A3(n3746), .A4(n3747), .ZN(n3743)
         );
  OAI22_X1 U6773 ( .A1(n13959), .A2(n11179), .B1(n13991), .B2(n11176), .ZN(
        n3747) );
  OAI222_X1 U6774 ( .A1(n944), .A2(n11155), .B1(n14244), .B2(n11152), .C1(
        n14212), .C2(n11149), .ZN(n3744) );
  OAI222_X1 U6775 ( .A1(n14149), .A2(n11164), .B1(n14181), .B2(n11161), .C1(
        n14117), .C2(n11158), .ZN(n3745) );
  NOR4_X1 U6776 ( .A1(n5127), .A2(n5128), .A3(n5129), .A4(n5130), .ZN(n5126)
         );
  OAI22_X1 U6777 ( .A1(n10097), .A2(n10981), .B1(n10096), .B2(n10978), .ZN(
        n5130) );
  OAI222_X1 U6778 ( .A1(n13926), .A2(n10957), .B1(n13862), .B2(n10954), .C1(
        n13894), .C2(n10951), .ZN(n5127) );
  OAI222_X1 U6779 ( .A1(n10091), .A2(n10966), .B1(n10090), .B2(n10963), .C1(
        n10092), .C2(n10960), .ZN(n5128) );
  NOR4_X1 U6780 ( .A1(n5136), .A2(n5137), .A3(n5138), .A4(n5139), .ZN(n5135)
         );
  OAI22_X1 U6781 ( .A1(n13958), .A2(n10915), .B1(n13990), .B2(n10912), .ZN(
        n5139) );
  OAI222_X1 U6782 ( .A1(n940), .A2(n10891), .B1(n14243), .B2(n10888), .C1(
        n14211), .C2(n10885), .ZN(n5136) );
  OAI222_X1 U6783 ( .A1(n14148), .A2(n10900), .B1(n14180), .B2(n10897), .C1(
        n14116), .C2(n10894), .ZN(n5137) );
  NOR4_X1 U6784 ( .A1(n3694), .A2(n3695), .A3(n3696), .A4(n3697), .ZN(n3693)
         );
  OAI22_X1 U6785 ( .A1(n10097), .A2(n11245), .B1(n10096), .B2(n11242), .ZN(
        n3697) );
  OAI222_X1 U6786 ( .A1(n13926), .A2(n11221), .B1(n13862), .B2(n11218), .C1(
        n13894), .C2(n11215), .ZN(n3694) );
  OAI222_X1 U6787 ( .A1(n10091), .A2(n11230), .B1(n10090), .B2(n11227), .C1(
        n10092), .C2(n11224), .ZN(n3695) );
  NOR4_X1 U6788 ( .A1(n3703), .A2(n3704), .A3(n3705), .A4(n3706), .ZN(n3702)
         );
  OAI22_X1 U6789 ( .A1(n13958), .A2(n11179), .B1(n13990), .B2(n11176), .ZN(
        n3706) );
  OAI222_X1 U6790 ( .A1(n940), .A2(n11155), .B1(n14243), .B2(n11152), .C1(
        n14211), .C2(n11149), .ZN(n3703) );
  OAI222_X1 U6791 ( .A1(n14148), .A2(n11164), .B1(n14180), .B2(n11161), .C1(
        n14116), .C2(n11158), .ZN(n3704) );
  NOR4_X1 U6792 ( .A1(n5086), .A2(n5087), .A3(n5088), .A4(n5089), .ZN(n5085)
         );
  OAI22_X1 U6793 ( .A1(n10065), .A2(n10981), .B1(n10064), .B2(n10978), .ZN(
        n5089) );
  OAI222_X1 U6794 ( .A1(n13925), .A2(n10957), .B1(n13861), .B2(n10954), .C1(
        n13893), .C2(n10951), .ZN(n5086) );
  OAI222_X1 U6795 ( .A1(n10059), .A2(n10966), .B1(n10058), .B2(n10963), .C1(
        n10060), .C2(n10960), .ZN(n5087) );
  NOR4_X1 U6796 ( .A1(n5095), .A2(n5096), .A3(n5097), .A4(n5098), .ZN(n5094)
         );
  OAI22_X1 U6797 ( .A1(n13957), .A2(n10915), .B1(n13989), .B2(n10912), .ZN(
        n5098) );
  OAI222_X1 U6798 ( .A1(n936), .A2(n10891), .B1(n14242), .B2(n10888), .C1(
        n14210), .C2(n10885), .ZN(n5095) );
  OAI222_X1 U6799 ( .A1(n14147), .A2(n10900), .B1(n14179), .B2(n10897), .C1(
        n14115), .C2(n10894), .ZN(n5096) );
  NOR4_X1 U6800 ( .A1(n3653), .A2(n3654), .A3(n3655), .A4(n3656), .ZN(n3652)
         );
  OAI22_X1 U6801 ( .A1(n10065), .A2(n11245), .B1(n10064), .B2(n11242), .ZN(
        n3656) );
  OAI222_X1 U6802 ( .A1(n13925), .A2(n11221), .B1(n13861), .B2(n11218), .C1(
        n13893), .C2(n11215), .ZN(n3653) );
  OAI222_X1 U6803 ( .A1(n10059), .A2(n11230), .B1(n10058), .B2(n11227), .C1(
        n10060), .C2(n11224), .ZN(n3654) );
  NOR4_X1 U6804 ( .A1(n3662), .A2(n3663), .A3(n3664), .A4(n3665), .ZN(n3661)
         );
  OAI22_X1 U6805 ( .A1(n13957), .A2(n11179), .B1(n13989), .B2(n11176), .ZN(
        n3665) );
  OAI222_X1 U6806 ( .A1(n936), .A2(n11155), .B1(n14242), .B2(n11152), .C1(
        n14210), .C2(n11149), .ZN(n3662) );
  OAI222_X1 U6807 ( .A1(n14147), .A2(n11164), .B1(n14179), .B2(n11161), .C1(
        n14115), .C2(n11158), .ZN(n3663) );
  NOR4_X1 U6808 ( .A1(n5045), .A2(n5046), .A3(n5047), .A4(n5048), .ZN(n5044)
         );
  OAI22_X1 U6809 ( .A1(n10033), .A2(n10981), .B1(n10032), .B2(n10978), .ZN(
        n5048) );
  OAI222_X1 U6810 ( .A1(n13924), .A2(n10957), .B1(n13860), .B2(n10954), .C1(
        n13892), .C2(n10951), .ZN(n5045) );
  OAI222_X1 U6811 ( .A1(n10027), .A2(n10966), .B1(n10026), .B2(n10963), .C1(
        n10028), .C2(n10960), .ZN(n5046) );
  NOR4_X1 U6812 ( .A1(n5054), .A2(n5055), .A3(n5056), .A4(n5057), .ZN(n5053)
         );
  OAI22_X1 U6813 ( .A1(n13956), .A2(n10915), .B1(n13988), .B2(n10912), .ZN(
        n5057) );
  OAI222_X1 U6814 ( .A1(n932), .A2(n10891), .B1(n14241), .B2(n10888), .C1(
        n14209), .C2(n10885), .ZN(n5054) );
  OAI222_X1 U6815 ( .A1(n14146), .A2(n10900), .B1(n14178), .B2(n10897), .C1(
        n14114), .C2(n10894), .ZN(n5055) );
  NOR4_X1 U6816 ( .A1(n3612), .A2(n3613), .A3(n3614), .A4(n3615), .ZN(n3611)
         );
  OAI22_X1 U6817 ( .A1(n10033), .A2(n11245), .B1(n10032), .B2(n11242), .ZN(
        n3615) );
  OAI222_X1 U6818 ( .A1(n13924), .A2(n11221), .B1(n13860), .B2(n11218), .C1(
        n13892), .C2(n11215), .ZN(n3612) );
  OAI222_X1 U6819 ( .A1(n10027), .A2(n11230), .B1(n10026), .B2(n11227), .C1(
        n10028), .C2(n11224), .ZN(n3613) );
  NOR4_X1 U6820 ( .A1(n3621), .A2(n3622), .A3(n3623), .A4(n3624), .ZN(n3620)
         );
  OAI22_X1 U6821 ( .A1(n13956), .A2(n11179), .B1(n13988), .B2(n11176), .ZN(
        n3624) );
  OAI222_X1 U6822 ( .A1(n932), .A2(n11155), .B1(n14241), .B2(n11152), .C1(
        n14209), .C2(n11149), .ZN(n3621) );
  OAI222_X1 U6823 ( .A1(n14146), .A2(n11164), .B1(n14178), .B2(n11161), .C1(
        n14114), .C2(n11158), .ZN(n3622) );
  NOR4_X1 U6824 ( .A1(n5004), .A2(n5005), .A3(n5006), .A4(n5007), .ZN(n5003)
         );
  OAI22_X1 U6825 ( .A1(n10001), .A2(n10981), .B1(n10000), .B2(n10978), .ZN(
        n5007) );
  OAI222_X1 U6826 ( .A1(n13923), .A2(n10957), .B1(n13859), .B2(n10954), .C1(
        n13891), .C2(n10951), .ZN(n5004) );
  OAI222_X1 U6827 ( .A1(n9697), .A2(n10966), .B1(n9696), .B2(n10963), .C1(
        n9698), .C2(n10960), .ZN(n5005) );
  NOR4_X1 U6828 ( .A1(n5013), .A2(n5014), .A3(n5015), .A4(n5016), .ZN(n5012)
         );
  OAI22_X1 U6829 ( .A1(n13955), .A2(n10915), .B1(n13987), .B2(n10912), .ZN(
        n5016) );
  OAI222_X1 U6830 ( .A1(n928), .A2(n10891), .B1(n14240), .B2(n10888), .C1(
        n14208), .C2(n10885), .ZN(n5013) );
  OAI222_X1 U6831 ( .A1(n14145), .A2(n10900), .B1(n14177), .B2(n10897), .C1(
        n14113), .C2(n10894), .ZN(n5014) );
  NOR4_X1 U6832 ( .A1(n3571), .A2(n3572), .A3(n3573), .A4(n3574), .ZN(n3570)
         );
  OAI22_X1 U6833 ( .A1(n10001), .A2(n11245), .B1(n10000), .B2(n11242), .ZN(
        n3574) );
  OAI222_X1 U6834 ( .A1(n13923), .A2(n11221), .B1(n13859), .B2(n11218), .C1(
        n13891), .C2(n11215), .ZN(n3571) );
  OAI222_X1 U6835 ( .A1(n9697), .A2(n11230), .B1(n9696), .B2(n11227), .C1(
        n9698), .C2(n11224), .ZN(n3572) );
  NOR4_X1 U6836 ( .A1(n3580), .A2(n3581), .A3(n3582), .A4(n3583), .ZN(n3579)
         );
  OAI22_X1 U6837 ( .A1(n13955), .A2(n11179), .B1(n13987), .B2(n11176), .ZN(
        n3583) );
  OAI222_X1 U6838 ( .A1(n928), .A2(n11155), .B1(n14240), .B2(n11152), .C1(
        n14208), .C2(n11149), .ZN(n3580) );
  OAI222_X1 U6839 ( .A1(n14145), .A2(n11164), .B1(n14177), .B2(n11161), .C1(
        n14113), .C2(n11158), .ZN(n3581) );
  NOR4_X1 U6840 ( .A1(n4963), .A2(n4964), .A3(n4965), .A4(n4966), .ZN(n4962)
         );
  OAI22_X1 U6841 ( .A1(n9639), .A2(n10981), .B1(n9638), .B2(n10978), .ZN(n4966) );
  OAI222_X1 U6842 ( .A1(n13922), .A2(n10957), .B1(n13858), .B2(n10954), .C1(
        n13890), .C2(n10951), .ZN(n4963) );
  OAI222_X1 U6843 ( .A1(n9633), .A2(n10966), .B1(n9632), .B2(n10963), .C1(
        n9634), .C2(n10960), .ZN(n4964) );
  NOR4_X1 U6844 ( .A1(n4972), .A2(n4973), .A3(n4974), .A4(n4975), .ZN(n4971)
         );
  OAI22_X1 U6845 ( .A1(n13954), .A2(n10915), .B1(n13986), .B2(n10912), .ZN(
        n4975) );
  OAI222_X1 U6846 ( .A1(n924), .A2(n10891), .B1(n14239), .B2(n10888), .C1(
        n14207), .C2(n10885), .ZN(n4972) );
  OAI222_X1 U6847 ( .A1(n14144), .A2(n10900), .B1(n14176), .B2(n10897), .C1(
        n14112), .C2(n10894), .ZN(n4973) );
  NOR4_X1 U6848 ( .A1(n3530), .A2(n3531), .A3(n3532), .A4(n3533), .ZN(n3529)
         );
  OAI22_X1 U6849 ( .A1(n9639), .A2(n11245), .B1(n9638), .B2(n11242), .ZN(n3533) );
  OAI222_X1 U6850 ( .A1(n13922), .A2(n11221), .B1(n13858), .B2(n11218), .C1(
        n13890), .C2(n11215), .ZN(n3530) );
  OAI222_X1 U6851 ( .A1(n9633), .A2(n11230), .B1(n9632), .B2(n11227), .C1(
        n9634), .C2(n11224), .ZN(n3531) );
  NOR4_X1 U6852 ( .A1(n3539), .A2(n3540), .A3(n3541), .A4(n3542), .ZN(n3538)
         );
  OAI22_X1 U6853 ( .A1(n13954), .A2(n11179), .B1(n13986), .B2(n11176), .ZN(
        n3542) );
  OAI222_X1 U6854 ( .A1(n924), .A2(n11155), .B1(n14239), .B2(n11152), .C1(
        n14207), .C2(n11149), .ZN(n3539) );
  OAI222_X1 U6855 ( .A1(n14144), .A2(n11164), .B1(n14176), .B2(n11161), .C1(
        n14112), .C2(n11158), .ZN(n3540) );
  NOR4_X1 U6856 ( .A1(n4922), .A2(n4923), .A3(n4924), .A4(n4925), .ZN(n4921)
         );
  OAI22_X1 U6857 ( .A1(n9607), .A2(n10981), .B1(n9606), .B2(n10978), .ZN(n4925) );
  OAI222_X1 U6858 ( .A1(n13921), .A2(n10957), .B1(n13857), .B2(n10954), .C1(
        n13889), .C2(n10951), .ZN(n4922) );
  OAI222_X1 U6859 ( .A1(n9601), .A2(n10966), .B1(n9600), .B2(n10963), .C1(
        n9602), .C2(n10960), .ZN(n4923) );
  NOR4_X1 U6860 ( .A1(n4931), .A2(n4932), .A3(n4933), .A4(n4934), .ZN(n4930)
         );
  OAI22_X1 U6861 ( .A1(n13953), .A2(n10915), .B1(n13985), .B2(n10912), .ZN(
        n4934) );
  OAI222_X1 U6862 ( .A1(n920), .A2(n10891), .B1(n14238), .B2(n10888), .C1(
        n14206), .C2(n10885), .ZN(n4931) );
  OAI222_X1 U6863 ( .A1(n14143), .A2(n10900), .B1(n14175), .B2(n10897), .C1(
        n14111), .C2(n10894), .ZN(n4932) );
  NOR4_X1 U6864 ( .A1(n3489), .A2(n3490), .A3(n3491), .A4(n3492), .ZN(n3488)
         );
  OAI22_X1 U6865 ( .A1(n9607), .A2(n11245), .B1(n9606), .B2(n11242), .ZN(n3492) );
  OAI222_X1 U6866 ( .A1(n13921), .A2(n11221), .B1(n13857), .B2(n11218), .C1(
        n13889), .C2(n11215), .ZN(n3489) );
  OAI222_X1 U6867 ( .A1(n9601), .A2(n11230), .B1(n9600), .B2(n11227), .C1(
        n9602), .C2(n11224), .ZN(n3490) );
  NOR4_X1 U6868 ( .A1(n3498), .A2(n3499), .A3(n3500), .A4(n3501), .ZN(n3497)
         );
  OAI22_X1 U6869 ( .A1(n13953), .A2(n11179), .B1(n13985), .B2(n11176), .ZN(
        n3501) );
  OAI222_X1 U6870 ( .A1(n920), .A2(n11155), .B1(n14238), .B2(n11152), .C1(
        n14206), .C2(n11149), .ZN(n3498) );
  OAI222_X1 U6871 ( .A1(n14143), .A2(n11164), .B1(n14175), .B2(n11161), .C1(
        n14111), .C2(n11158), .ZN(n3499) );
  NOR4_X1 U6872 ( .A1(n4881), .A2(n4882), .A3(n4883), .A4(n4884), .ZN(n4880)
         );
  OAI22_X1 U6873 ( .A1(n9575), .A2(n10981), .B1(n9574), .B2(n10978), .ZN(n4884) );
  OAI222_X1 U6874 ( .A1(n13920), .A2(n10957), .B1(n13856), .B2(n10954), .C1(
        n13888), .C2(n10951), .ZN(n4881) );
  OAI222_X1 U6875 ( .A1(n9569), .A2(n10966), .B1(n9568), .B2(n10963), .C1(
        n9570), .C2(n10960), .ZN(n4882) );
  NOR4_X1 U6876 ( .A1(n4890), .A2(n4891), .A3(n4892), .A4(n4893), .ZN(n4889)
         );
  OAI22_X1 U6877 ( .A1(n13952), .A2(n10915), .B1(n13984), .B2(n10912), .ZN(
        n4893) );
  OAI222_X1 U6878 ( .A1(n916), .A2(n10891), .B1(n14237), .B2(n10888), .C1(
        n14205), .C2(n10885), .ZN(n4890) );
  OAI222_X1 U6879 ( .A1(n14142), .A2(n10900), .B1(n14174), .B2(n10897), .C1(
        n14110), .C2(n10894), .ZN(n4891) );
  NOR4_X1 U6880 ( .A1(n3448), .A2(n3449), .A3(n3450), .A4(n3451), .ZN(n3447)
         );
  OAI22_X1 U6881 ( .A1(n9575), .A2(n11245), .B1(n9574), .B2(n11242), .ZN(n3451) );
  OAI222_X1 U6882 ( .A1(n13920), .A2(n11221), .B1(n13856), .B2(n11218), .C1(
        n13888), .C2(n11215), .ZN(n3448) );
  OAI222_X1 U6883 ( .A1(n9569), .A2(n11230), .B1(n9568), .B2(n11227), .C1(
        n9570), .C2(n11224), .ZN(n3449) );
  NOR4_X1 U6884 ( .A1(n3457), .A2(n3458), .A3(n3459), .A4(n3460), .ZN(n3456)
         );
  OAI22_X1 U6885 ( .A1(n13952), .A2(n11179), .B1(n13984), .B2(n11176), .ZN(
        n3460) );
  OAI222_X1 U6886 ( .A1(n916), .A2(n11155), .B1(n14237), .B2(n11152), .C1(
        n14205), .C2(n11149), .ZN(n3457) );
  OAI222_X1 U6887 ( .A1(n14142), .A2(n11164), .B1(n14174), .B2(n11161), .C1(
        n14110), .C2(n11158), .ZN(n3458) );
  NOR4_X1 U6888 ( .A1(n4840), .A2(n4841), .A3(n4842), .A4(n4843), .ZN(n4839)
         );
  OAI22_X1 U6889 ( .A1(n9209), .A2(n10981), .B1(n9208), .B2(n10978), .ZN(n4843) );
  OAI222_X1 U6890 ( .A1(n13919), .A2(n10957), .B1(n13855), .B2(n10954), .C1(
        n13887), .C2(n10951), .ZN(n4840) );
  OAI222_X1 U6891 ( .A1(n9203), .A2(n10966), .B1(n9202), .B2(n10963), .C1(
        n9204), .C2(n10960), .ZN(n4841) );
  NOR4_X1 U6892 ( .A1(n4849), .A2(n4850), .A3(n4851), .A4(n4852), .ZN(n4848)
         );
  OAI22_X1 U6893 ( .A1(n13951), .A2(n10915), .B1(n13983), .B2(n10912), .ZN(
        n4852) );
  OAI222_X1 U6894 ( .A1(n912), .A2(n10891), .B1(n14236), .B2(n10888), .C1(
        n14204), .C2(n10885), .ZN(n4849) );
  OAI222_X1 U6895 ( .A1(n14141), .A2(n10900), .B1(n14173), .B2(n10897), .C1(
        n14109), .C2(n10894), .ZN(n4850) );
  NOR4_X1 U6896 ( .A1(n3407), .A2(n3408), .A3(n3409), .A4(n3410), .ZN(n3406)
         );
  OAI22_X1 U6897 ( .A1(n9209), .A2(n11245), .B1(n9208), .B2(n11242), .ZN(n3410) );
  OAI222_X1 U6898 ( .A1(n13919), .A2(n11221), .B1(n13855), .B2(n11218), .C1(
        n13887), .C2(n11215), .ZN(n3407) );
  OAI222_X1 U6899 ( .A1(n9203), .A2(n11230), .B1(n9202), .B2(n11227), .C1(
        n9204), .C2(n11224), .ZN(n3408) );
  NOR4_X1 U6900 ( .A1(n3416), .A2(n3417), .A3(n3418), .A4(n3419), .ZN(n3415)
         );
  OAI22_X1 U6901 ( .A1(n13951), .A2(n11179), .B1(n13983), .B2(n11176), .ZN(
        n3419) );
  OAI222_X1 U6902 ( .A1(n912), .A2(n11155), .B1(n14236), .B2(n11152), .C1(
        n14204), .C2(n11149), .ZN(n3416) );
  OAI222_X1 U6903 ( .A1(n14141), .A2(n11164), .B1(n14173), .B2(n11161), .C1(
        n14109), .C2(n11158), .ZN(n3417) );
  NOR4_X1 U6904 ( .A1(n4799), .A2(n4800), .A3(n4801), .A4(n4802), .ZN(n4798)
         );
  OAI22_X1 U6905 ( .A1(n9177), .A2(n10981), .B1(n9176), .B2(n10978), .ZN(n4802) );
  OAI222_X1 U6906 ( .A1(n13918), .A2(n10957), .B1(n13854), .B2(n10954), .C1(
        n13886), .C2(n10951), .ZN(n4799) );
  OAI222_X1 U6907 ( .A1(n9171), .A2(n10966), .B1(n9170), .B2(n10963), .C1(
        n9172), .C2(n10960), .ZN(n4800) );
  NOR4_X1 U6908 ( .A1(n4808), .A2(n4809), .A3(n4810), .A4(n4811), .ZN(n4807)
         );
  OAI22_X1 U6909 ( .A1(n13950), .A2(n10915), .B1(n13982), .B2(n10912), .ZN(
        n4811) );
  OAI222_X1 U6910 ( .A1(n908), .A2(n10891), .B1(n14235), .B2(n10888), .C1(
        n14203), .C2(n10885), .ZN(n4808) );
  OAI222_X1 U6911 ( .A1(n14140), .A2(n10900), .B1(n14172), .B2(n10897), .C1(
        n14108), .C2(n10894), .ZN(n4809) );
  NOR4_X1 U6912 ( .A1(n3366), .A2(n3367), .A3(n3368), .A4(n3369), .ZN(n3365)
         );
  OAI22_X1 U6913 ( .A1(n9177), .A2(n11245), .B1(n9176), .B2(n11242), .ZN(n3369) );
  OAI222_X1 U6914 ( .A1(n13918), .A2(n11221), .B1(n13854), .B2(n11218), .C1(
        n13886), .C2(n11215), .ZN(n3366) );
  OAI222_X1 U6915 ( .A1(n9171), .A2(n11230), .B1(n9170), .B2(n11227), .C1(
        n9172), .C2(n11224), .ZN(n3367) );
  NOR4_X1 U6916 ( .A1(n3375), .A2(n3376), .A3(n3377), .A4(n3378), .ZN(n3374)
         );
  OAI22_X1 U6917 ( .A1(n13950), .A2(n11179), .B1(n13982), .B2(n11176), .ZN(
        n3378) );
  OAI222_X1 U6918 ( .A1(n908), .A2(n11155), .B1(n14235), .B2(n11152), .C1(
        n14203), .C2(n11149), .ZN(n3375) );
  OAI222_X1 U6919 ( .A1(n14140), .A2(n11164), .B1(n14172), .B2(n11161), .C1(
        n14108), .C2(n11158), .ZN(n3376) );
  NOR4_X1 U6920 ( .A1(n4758), .A2(n4759), .A3(n4760), .A4(n4761), .ZN(n4757)
         );
  OAI22_X1 U6921 ( .A1(n9145), .A2(n10981), .B1(n9144), .B2(n10978), .ZN(n4761) );
  OAI222_X1 U6922 ( .A1(n13917), .A2(n10957), .B1(n13853), .B2(n10954), .C1(
        n13885), .C2(n10951), .ZN(n4758) );
  OAI222_X1 U6923 ( .A1(n9139), .A2(n10966), .B1(n9138), .B2(n10963), .C1(
        n9140), .C2(n10960), .ZN(n4759) );
  NOR4_X1 U6924 ( .A1(n4767), .A2(n4768), .A3(n4769), .A4(n4770), .ZN(n4766)
         );
  OAI22_X1 U6925 ( .A1(n13949), .A2(n10915), .B1(n13981), .B2(n10912), .ZN(
        n4770) );
  OAI222_X1 U6926 ( .A1(n904), .A2(n10891), .B1(n14234), .B2(n10888), .C1(
        n14202), .C2(n10885), .ZN(n4767) );
  OAI222_X1 U6927 ( .A1(n14139), .A2(n10900), .B1(n14171), .B2(n10897), .C1(
        n14107), .C2(n10894), .ZN(n4768) );
  NOR4_X1 U6928 ( .A1(n3325), .A2(n3326), .A3(n3327), .A4(n3328), .ZN(n3324)
         );
  OAI22_X1 U6929 ( .A1(n9145), .A2(n11245), .B1(n9144), .B2(n11242), .ZN(n3328) );
  OAI222_X1 U6930 ( .A1(n13917), .A2(n11221), .B1(n13853), .B2(n11218), .C1(
        n13885), .C2(n11215), .ZN(n3325) );
  OAI222_X1 U6931 ( .A1(n9139), .A2(n11230), .B1(n9138), .B2(n11227), .C1(
        n9140), .C2(n11224), .ZN(n3326) );
  NOR4_X1 U6932 ( .A1(n3334), .A2(n3335), .A3(n3336), .A4(n3337), .ZN(n3333)
         );
  OAI22_X1 U6933 ( .A1(n13949), .A2(n11179), .B1(n13981), .B2(n11176), .ZN(
        n3337) );
  OAI222_X1 U6934 ( .A1(n904), .A2(n11155), .B1(n14234), .B2(n11152), .C1(
        n14202), .C2(n11149), .ZN(n3334) );
  OAI222_X1 U6935 ( .A1(n14139), .A2(n11164), .B1(n14171), .B2(n11161), .C1(
        n14107), .C2(n11158), .ZN(n3335) );
  NOR4_X1 U6936 ( .A1(n4717), .A2(n4718), .A3(n4719), .A4(n4720), .ZN(n4716)
         );
  OAI22_X1 U6937 ( .A1(n6010), .A2(n10981), .B1(n6009), .B2(n10978), .ZN(n4720) );
  OAI222_X1 U6938 ( .A1(n13916), .A2(n10957), .B1(n13852), .B2(n10954), .C1(
        n13884), .C2(n10951), .ZN(n4717) );
  OAI222_X1 U6939 ( .A1(n6004), .A2(n10966), .B1(n6003), .B2(n10963), .C1(
        n6005), .C2(n10960), .ZN(n4718) );
  NOR4_X1 U6940 ( .A1(n4726), .A2(n4727), .A3(n4728), .A4(n4729), .ZN(n4725)
         );
  OAI22_X1 U6941 ( .A1(n13948), .A2(n10915), .B1(n13980), .B2(n10912), .ZN(
        n4729) );
  OAI222_X1 U6942 ( .A1(n900), .A2(n10891), .B1(n14233), .B2(n10888), .C1(
        n14201), .C2(n10885), .ZN(n4726) );
  OAI222_X1 U6943 ( .A1(n14138), .A2(n10900), .B1(n14170), .B2(n10897), .C1(
        n14106), .C2(n10894), .ZN(n4727) );
  NOR4_X1 U6944 ( .A1(n3284), .A2(n3285), .A3(n3286), .A4(n3287), .ZN(n3283)
         );
  OAI22_X1 U6945 ( .A1(n6010), .A2(n11245), .B1(n6009), .B2(n11242), .ZN(n3287) );
  OAI222_X1 U6946 ( .A1(n13916), .A2(n11221), .B1(n13852), .B2(n11218), .C1(
        n13884), .C2(n11215), .ZN(n3284) );
  OAI222_X1 U6947 ( .A1(n6004), .A2(n11230), .B1(n6003), .B2(n11227), .C1(
        n6005), .C2(n11224), .ZN(n3285) );
  NOR4_X1 U6948 ( .A1(n3293), .A2(n3294), .A3(n3295), .A4(n3296), .ZN(n3292)
         );
  OAI22_X1 U6949 ( .A1(n13948), .A2(n11179), .B1(n13980), .B2(n11176), .ZN(
        n3296) );
  OAI222_X1 U6950 ( .A1(n900), .A2(n11155), .B1(n14233), .B2(n11152), .C1(
        n14201), .C2(n11149), .ZN(n3293) );
  OAI222_X1 U6951 ( .A1(n14138), .A2(n11164), .B1(n14170), .B2(n11161), .C1(
        n14106), .C2(n11158), .ZN(n3294) );
  NOR4_X1 U6952 ( .A1(n4676), .A2(n4677), .A3(n4678), .A4(n4679), .ZN(n4675)
         );
  OAI22_X1 U6953 ( .A1(n5946), .A2(n10982), .B1(n5945), .B2(n10979), .ZN(n4679) );
  OAI222_X1 U6954 ( .A1(n13915), .A2(n10958), .B1(n13851), .B2(n10955), .C1(
        n13883), .C2(n10952), .ZN(n4676) );
  OAI222_X1 U6955 ( .A1(n5940), .A2(n10967), .B1(n5939), .B2(n10964), .C1(
        n5941), .C2(n10961), .ZN(n4677) );
  NOR4_X1 U6956 ( .A1(n4685), .A2(n4686), .A3(n4687), .A4(n4688), .ZN(n4684)
         );
  OAI22_X1 U6957 ( .A1(n13947), .A2(n10916), .B1(n13979), .B2(n10913), .ZN(
        n4688) );
  OAI222_X1 U6958 ( .A1(n896), .A2(n10892), .B1(n14232), .B2(n10889), .C1(
        n14200), .C2(n10886), .ZN(n4685) );
  OAI222_X1 U6959 ( .A1(n14137), .A2(n10901), .B1(n14169), .B2(n10898), .C1(
        n14105), .C2(n10895), .ZN(n4686) );
  NOR4_X1 U6960 ( .A1(n3243), .A2(n3244), .A3(n3245), .A4(n3246), .ZN(n3242)
         );
  OAI22_X1 U6961 ( .A1(n5946), .A2(n11246), .B1(n5945), .B2(n11243), .ZN(n3246) );
  OAI222_X1 U6962 ( .A1(n13915), .A2(n11222), .B1(n13851), .B2(n11219), .C1(
        n13883), .C2(n11216), .ZN(n3243) );
  OAI222_X1 U6963 ( .A1(n5940), .A2(n11231), .B1(n5939), .B2(n11228), .C1(
        n5941), .C2(n11225), .ZN(n3244) );
  NOR4_X1 U6964 ( .A1(n3252), .A2(n3253), .A3(n3254), .A4(n3255), .ZN(n3251)
         );
  OAI22_X1 U6965 ( .A1(n13947), .A2(n11180), .B1(n13979), .B2(n11177), .ZN(
        n3255) );
  OAI222_X1 U6966 ( .A1(n896), .A2(n11156), .B1(n14232), .B2(n11153), .C1(
        n14200), .C2(n11150), .ZN(n3252) );
  OAI222_X1 U6967 ( .A1(n14137), .A2(n11165), .B1(n14169), .B2(n11162), .C1(
        n14105), .C2(n11159), .ZN(n3253) );
  NOR4_X1 U6968 ( .A1(n4635), .A2(n4636), .A3(n4637), .A4(n4638), .ZN(n4634)
         );
  OAI22_X1 U6969 ( .A1(n5914), .A2(n10982), .B1(n5913), .B2(n10979), .ZN(n4638) );
  OAI222_X1 U6970 ( .A1(n13914), .A2(n10958), .B1(n13850), .B2(n10955), .C1(
        n13882), .C2(n10952), .ZN(n4635) );
  OAI222_X1 U6971 ( .A1(n5908), .A2(n10967), .B1(n5907), .B2(n10964), .C1(
        n5909), .C2(n10961), .ZN(n4636) );
  NOR4_X1 U6972 ( .A1(n4644), .A2(n4645), .A3(n4646), .A4(n4647), .ZN(n4643)
         );
  OAI22_X1 U6973 ( .A1(n13946), .A2(n10916), .B1(n13978), .B2(n10913), .ZN(
        n4647) );
  OAI222_X1 U6974 ( .A1(n892), .A2(n10892), .B1(n14231), .B2(n10889), .C1(
        n14199), .C2(n10886), .ZN(n4644) );
  OAI222_X1 U6975 ( .A1(n14136), .A2(n10901), .B1(n14168), .B2(n10898), .C1(
        n14104), .C2(n10895), .ZN(n4645) );
  NOR4_X1 U6976 ( .A1(n3202), .A2(n3203), .A3(n3204), .A4(n3205), .ZN(n3201)
         );
  OAI22_X1 U6977 ( .A1(n5914), .A2(n11246), .B1(n5913), .B2(n11243), .ZN(n3205) );
  OAI222_X1 U6978 ( .A1(n13914), .A2(n11222), .B1(n13850), .B2(n11219), .C1(
        n13882), .C2(n11216), .ZN(n3202) );
  OAI222_X1 U6979 ( .A1(n5908), .A2(n11231), .B1(n5907), .B2(n11228), .C1(
        n5909), .C2(n11225), .ZN(n3203) );
  NOR4_X1 U6980 ( .A1(n3211), .A2(n3212), .A3(n3213), .A4(n3214), .ZN(n3210)
         );
  OAI22_X1 U6981 ( .A1(n13946), .A2(n11180), .B1(n13978), .B2(n11177), .ZN(
        n3214) );
  OAI222_X1 U6982 ( .A1(n892), .A2(n11156), .B1(n14231), .B2(n11153), .C1(
        n14199), .C2(n11150), .ZN(n3211) );
  OAI222_X1 U6983 ( .A1(n14136), .A2(n11165), .B1(n14168), .B2(n11162), .C1(
        n14104), .C2(n11159), .ZN(n3212) );
  NOR4_X1 U6984 ( .A1(n4594), .A2(n4595), .A3(n4596), .A4(n4597), .ZN(n4593)
         );
  OAI22_X1 U6985 ( .A1(n5882), .A2(n10982), .B1(n5881), .B2(n10979), .ZN(n4597) );
  OAI222_X1 U6986 ( .A1(n13913), .A2(n10958), .B1(n13849), .B2(n10955), .C1(
        n13881), .C2(n10952), .ZN(n4594) );
  OAI222_X1 U6987 ( .A1(n5876), .A2(n10967), .B1(n5875), .B2(n10964), .C1(
        n5877), .C2(n10961), .ZN(n4595) );
  NOR4_X1 U6988 ( .A1(n4603), .A2(n4604), .A3(n4605), .A4(n4606), .ZN(n4602)
         );
  OAI22_X1 U6989 ( .A1(n13945), .A2(n10916), .B1(n13977), .B2(n10913), .ZN(
        n4606) );
  OAI222_X1 U6990 ( .A1(n888), .A2(n10892), .B1(n14230), .B2(n10889), .C1(
        n14198), .C2(n10886), .ZN(n4603) );
  OAI222_X1 U6991 ( .A1(n14135), .A2(n10901), .B1(n14167), .B2(n10898), .C1(
        n14103), .C2(n10895), .ZN(n4604) );
  NOR4_X1 U6992 ( .A1(n3161), .A2(n3162), .A3(n3163), .A4(n3164), .ZN(n3160)
         );
  OAI22_X1 U6993 ( .A1(n5882), .A2(n11246), .B1(n5881), .B2(n11243), .ZN(n3164) );
  OAI222_X1 U6994 ( .A1(n13913), .A2(n11222), .B1(n13849), .B2(n11219), .C1(
        n13881), .C2(n11216), .ZN(n3161) );
  OAI222_X1 U6995 ( .A1(n5876), .A2(n11231), .B1(n5875), .B2(n11228), .C1(
        n5877), .C2(n11225), .ZN(n3162) );
  NOR4_X1 U6996 ( .A1(n3170), .A2(n3171), .A3(n3172), .A4(n3173), .ZN(n3169)
         );
  OAI22_X1 U6997 ( .A1(n13945), .A2(n11180), .B1(n13977), .B2(n11177), .ZN(
        n3173) );
  OAI222_X1 U6998 ( .A1(n888), .A2(n11156), .B1(n14230), .B2(n11153), .C1(
        n14198), .C2(n11150), .ZN(n3170) );
  OAI222_X1 U6999 ( .A1(n14135), .A2(n11165), .B1(n14167), .B2(n11162), .C1(
        n14103), .C2(n11159), .ZN(n3171) );
  NOR4_X1 U7000 ( .A1(n4553), .A2(n4554), .A3(n4555), .A4(n4556), .ZN(n4552)
         );
  OAI22_X1 U7001 ( .A1(n5850), .A2(n10982), .B1(n5849), .B2(n10979), .ZN(n4556) );
  OAI222_X1 U7002 ( .A1(n13912), .A2(n10958), .B1(n13848), .B2(n10955), .C1(
        n13880), .C2(n10952), .ZN(n4553) );
  OAI222_X1 U7003 ( .A1(n5844), .A2(n10967), .B1(n5843), .B2(n10964), .C1(
        n5845), .C2(n10961), .ZN(n4554) );
  NOR4_X1 U7004 ( .A1(n4562), .A2(n4563), .A3(n4564), .A4(n4565), .ZN(n4561)
         );
  OAI22_X1 U7005 ( .A1(n13944), .A2(n10916), .B1(n13976), .B2(n10913), .ZN(
        n4565) );
  OAI222_X1 U7006 ( .A1(n884), .A2(n10892), .B1(n14229), .B2(n10889), .C1(
        n14197), .C2(n10886), .ZN(n4562) );
  OAI222_X1 U7007 ( .A1(n14134), .A2(n10901), .B1(n14166), .B2(n10898), .C1(
        n14102), .C2(n10895), .ZN(n4563) );
  NOR4_X1 U7008 ( .A1(n3120), .A2(n3121), .A3(n3122), .A4(n3123), .ZN(n3119)
         );
  OAI22_X1 U7009 ( .A1(n5850), .A2(n11246), .B1(n5849), .B2(n11243), .ZN(n3123) );
  OAI222_X1 U7010 ( .A1(n13912), .A2(n11222), .B1(n13848), .B2(n11219), .C1(
        n13880), .C2(n11216), .ZN(n3120) );
  OAI222_X1 U7011 ( .A1(n5844), .A2(n11231), .B1(n5843), .B2(n11228), .C1(
        n5845), .C2(n11225), .ZN(n3121) );
  NOR4_X1 U7012 ( .A1(n3129), .A2(n3130), .A3(n3131), .A4(n3132), .ZN(n3128)
         );
  OAI22_X1 U7013 ( .A1(n13944), .A2(n11180), .B1(n13976), .B2(n11177), .ZN(
        n3132) );
  OAI222_X1 U7014 ( .A1(n884), .A2(n11156), .B1(n14229), .B2(n11153), .C1(
        n14197), .C2(n11150), .ZN(n3129) );
  OAI222_X1 U7015 ( .A1(n14134), .A2(n11165), .B1(n14166), .B2(n11162), .C1(
        n14102), .C2(n11159), .ZN(n3130) );
  NOR4_X1 U7016 ( .A1(n4512), .A2(n4513), .A3(n4514), .A4(n4515), .ZN(n4511)
         );
  OAI22_X1 U7017 ( .A1(n5818), .A2(n10982), .B1(n5817), .B2(n10979), .ZN(n4515) );
  OAI222_X1 U7018 ( .A1(n13911), .A2(n10958), .B1(n13847), .B2(n10955), .C1(
        n13879), .C2(n10952), .ZN(n4512) );
  OAI222_X1 U7019 ( .A1(n5812), .A2(n10967), .B1(n5811), .B2(n10964), .C1(
        n5813), .C2(n10961), .ZN(n4513) );
  NOR4_X1 U7020 ( .A1(n4521), .A2(n4522), .A3(n4523), .A4(n4524), .ZN(n4520)
         );
  OAI22_X1 U7021 ( .A1(n13943), .A2(n10916), .B1(n13975), .B2(n10913), .ZN(
        n4524) );
  OAI222_X1 U7022 ( .A1(n880), .A2(n10892), .B1(n14228), .B2(n10889), .C1(
        n14196), .C2(n10886), .ZN(n4521) );
  OAI222_X1 U7023 ( .A1(n14133), .A2(n10901), .B1(n14165), .B2(n10898), .C1(
        n14101), .C2(n10895), .ZN(n4522) );
  NOR4_X1 U7024 ( .A1(n3079), .A2(n3080), .A3(n3081), .A4(n3082), .ZN(n3078)
         );
  OAI22_X1 U7025 ( .A1(n5818), .A2(n11246), .B1(n5817), .B2(n11243), .ZN(n3082) );
  OAI222_X1 U7026 ( .A1(n13911), .A2(n11222), .B1(n13847), .B2(n11219), .C1(
        n13879), .C2(n11216), .ZN(n3079) );
  OAI222_X1 U7027 ( .A1(n5812), .A2(n11231), .B1(n5811), .B2(n11228), .C1(
        n5813), .C2(n11225), .ZN(n3080) );
  NOR4_X1 U7028 ( .A1(n3088), .A2(n3089), .A3(n3090), .A4(n3091), .ZN(n3087)
         );
  OAI22_X1 U7029 ( .A1(n13943), .A2(n11180), .B1(n13975), .B2(n11177), .ZN(
        n3091) );
  OAI222_X1 U7030 ( .A1(n880), .A2(n11156), .B1(n14228), .B2(n11153), .C1(
        n14196), .C2(n11150), .ZN(n3088) );
  OAI222_X1 U7031 ( .A1(n14133), .A2(n11165), .B1(n14165), .B2(n11162), .C1(
        n14101), .C2(n11159), .ZN(n3089) );
  NOR4_X1 U7032 ( .A1(n4471), .A2(n4472), .A3(n4473), .A4(n4474), .ZN(n4470)
         );
  OAI22_X1 U7033 ( .A1(n5786), .A2(n10982), .B1(n5785), .B2(n10979), .ZN(n4474) );
  OAI222_X1 U7034 ( .A1(n13910), .A2(n10958), .B1(n13846), .B2(n10955), .C1(
        n13878), .C2(n10952), .ZN(n4471) );
  OAI222_X1 U7035 ( .A1(n5780), .A2(n10967), .B1(n5779), .B2(n10964), .C1(
        n5781), .C2(n10961), .ZN(n4472) );
  NOR4_X1 U7036 ( .A1(n4480), .A2(n4481), .A3(n4482), .A4(n4483), .ZN(n4479)
         );
  OAI22_X1 U7037 ( .A1(n13942), .A2(n10916), .B1(n13974), .B2(n10913), .ZN(
        n4483) );
  OAI222_X1 U7038 ( .A1(n876), .A2(n10892), .B1(n14227), .B2(n10889), .C1(
        n14195), .C2(n10886), .ZN(n4480) );
  OAI222_X1 U7039 ( .A1(n14132), .A2(n10901), .B1(n14164), .B2(n10898), .C1(
        n14100), .C2(n10895), .ZN(n4481) );
  NOR4_X1 U7040 ( .A1(n3038), .A2(n3039), .A3(n3040), .A4(n3041), .ZN(n3037)
         );
  OAI22_X1 U7041 ( .A1(n5786), .A2(n11246), .B1(n5785), .B2(n11243), .ZN(n3041) );
  OAI222_X1 U7042 ( .A1(n13910), .A2(n11222), .B1(n13846), .B2(n11219), .C1(
        n13878), .C2(n11216), .ZN(n3038) );
  OAI222_X1 U7043 ( .A1(n5780), .A2(n11231), .B1(n5779), .B2(n11228), .C1(
        n5781), .C2(n11225), .ZN(n3039) );
  NOR4_X1 U7044 ( .A1(n3047), .A2(n3048), .A3(n3049), .A4(n3050), .ZN(n3046)
         );
  OAI22_X1 U7045 ( .A1(n13942), .A2(n11180), .B1(n13974), .B2(n11177), .ZN(
        n3050) );
  OAI222_X1 U7046 ( .A1(n876), .A2(n11156), .B1(n14227), .B2(n11153), .C1(
        n14195), .C2(n11150), .ZN(n3047) );
  OAI222_X1 U7047 ( .A1(n14132), .A2(n11165), .B1(n14164), .B2(n11162), .C1(
        n14100), .C2(n11159), .ZN(n3048) );
  NOR4_X1 U7048 ( .A1(n4430), .A2(n4431), .A3(n4432), .A4(n4433), .ZN(n4429)
         );
  OAI22_X1 U7049 ( .A1(n5754), .A2(n10982), .B1(n5753), .B2(n10979), .ZN(n4433) );
  OAI222_X1 U7050 ( .A1(n13909), .A2(n10958), .B1(n13845), .B2(n10955), .C1(
        n13877), .C2(n10952), .ZN(n4430) );
  OAI222_X1 U7051 ( .A1(n5748), .A2(n10967), .B1(n5747), .B2(n10964), .C1(
        n5749), .C2(n10961), .ZN(n4431) );
  NOR4_X1 U7052 ( .A1(n4439), .A2(n4440), .A3(n4441), .A4(n4442), .ZN(n4438)
         );
  OAI22_X1 U7053 ( .A1(n13941), .A2(n10916), .B1(n13973), .B2(n10913), .ZN(
        n4442) );
  OAI222_X1 U7054 ( .A1(n872), .A2(n10892), .B1(n14226), .B2(n10889), .C1(
        n14194), .C2(n10886), .ZN(n4439) );
  OAI222_X1 U7055 ( .A1(n14131), .A2(n10901), .B1(n14163), .B2(n10898), .C1(
        n14099), .C2(n10895), .ZN(n4440) );
  NOR4_X1 U7056 ( .A1(n2997), .A2(n2998), .A3(n2999), .A4(n3000), .ZN(n2996)
         );
  OAI22_X1 U7057 ( .A1(n5754), .A2(n11246), .B1(n5753), .B2(n11243), .ZN(n3000) );
  OAI222_X1 U7058 ( .A1(n13909), .A2(n11222), .B1(n13845), .B2(n11219), .C1(
        n13877), .C2(n11216), .ZN(n2997) );
  OAI222_X1 U7059 ( .A1(n5748), .A2(n11231), .B1(n5747), .B2(n11228), .C1(
        n5749), .C2(n11225), .ZN(n2998) );
  NOR4_X1 U7060 ( .A1(n3006), .A2(n3007), .A3(n3008), .A4(n3009), .ZN(n3005)
         );
  OAI22_X1 U7061 ( .A1(n13941), .A2(n11180), .B1(n13973), .B2(n11177), .ZN(
        n3009) );
  OAI222_X1 U7062 ( .A1(n872), .A2(n11156), .B1(n14226), .B2(n11153), .C1(
        n14194), .C2(n11150), .ZN(n3006) );
  OAI222_X1 U7063 ( .A1(n14131), .A2(n11165), .B1(n14163), .B2(n11162), .C1(
        n14099), .C2(n11159), .ZN(n3007) );
  NOR4_X1 U7064 ( .A1(n4345), .A2(n4346), .A3(n4347), .A4(n4348), .ZN(n4344)
         );
  OAI22_X1 U7065 ( .A1(n5722), .A2(n10982), .B1(n5721), .B2(n10979), .ZN(n4348) );
  OAI222_X1 U7066 ( .A1(n13908), .A2(n10958), .B1(n13844), .B2(n10955), .C1(
        n13876), .C2(n10952), .ZN(n4345) );
  OAI222_X1 U7067 ( .A1(n5716), .A2(n10967), .B1(n5715), .B2(n10964), .C1(
        n5717), .C2(n10961), .ZN(n4346) );
  NOR4_X1 U7068 ( .A1(n4376), .A2(n4377), .A3(n4378), .A4(n4379), .ZN(n4375)
         );
  OAI22_X1 U7069 ( .A1(n13940), .A2(n10916), .B1(n13972), .B2(n10913), .ZN(
        n4379) );
  OAI222_X1 U7070 ( .A1(n868), .A2(n10892), .B1(n14225), .B2(n10889), .C1(n996), .C2(n10886), .ZN(n4376) );
  OAI222_X1 U7071 ( .A1(n14130), .A2(n10901), .B1(n14162), .B2(n10898), .C1(
        n997), .C2(n10895), .ZN(n4377) );
  NOR4_X1 U7072 ( .A1(n2877), .A2(n2878), .A3(n2879), .A4(n2880), .ZN(n2876)
         );
  OAI22_X1 U7073 ( .A1(n5722), .A2(n11246), .B1(n5721), .B2(n11243), .ZN(n2880) );
  OAI222_X1 U7074 ( .A1(n13908), .A2(n11222), .B1(n13844), .B2(n11219), .C1(
        n13876), .C2(n11216), .ZN(n2877) );
  OAI222_X1 U7075 ( .A1(n5716), .A2(n11231), .B1(n5715), .B2(n11228), .C1(
        n5717), .C2(n11225), .ZN(n2878) );
  NOR4_X1 U7076 ( .A1(n2943), .A2(n2944), .A3(n2945), .A4(n2946), .ZN(n2942)
         );
  OAI22_X1 U7077 ( .A1(n13940), .A2(n11180), .B1(n13972), .B2(n11177), .ZN(
        n2946) );
  OAI222_X1 U7078 ( .A1(n868), .A2(n11156), .B1(n14225), .B2(n11153), .C1(n996), .C2(n11150), .ZN(n2943) );
  OAI222_X1 U7079 ( .A1(n14130), .A2(n11165), .B1(n14162), .B2(n11162), .C1(
        n997), .C2(n11159), .ZN(n2944) );
  AOI221_X1 U7080 ( .B1(n10947), .B2(n9504), .C1(n10944), .C2(n9536), .A(n5691), .ZN(n5681) );
  OAI222_X1 U7081 ( .A1(n13619), .A2(n10941), .B1(n13651), .B2(n10938), .C1(
        n13587), .C2(n10935), .ZN(n5691) );
  AOI221_X1 U7082 ( .B1(n10881), .B2(n14288), .C1(n10878), .C2(n14480), .A(
        n5704), .ZN(n5695) );
  OAI222_X1 U7083 ( .A1(n10510), .A2(n10875), .B1(n10509), .B2(n10872), .C1(
        n10511), .C2(n10869), .ZN(n5704) );
  AOI221_X1 U7084 ( .B1(n11211), .B2(n9504), .C1(n11208), .C2(n9536), .A(n4258), .ZN(n4248) );
  OAI222_X1 U7085 ( .A1(n13619), .A2(n11205), .B1(n13651), .B2(n11202), .C1(
        n13587), .C2(n11199), .ZN(n4258) );
  AOI221_X1 U7086 ( .B1(n11145), .B2(n14288), .C1(n11142), .C2(n14480), .A(
        n4271), .ZN(n4262) );
  OAI222_X1 U7087 ( .A1(n10510), .A2(n11139), .B1(n10509), .B2(n11136), .C1(
        n10511), .C2(n11133), .ZN(n4271) );
  AOI221_X1 U7088 ( .B1(n10947), .B2(n9505), .C1(n10944), .C2(n9537), .A(n5623), .ZN(n5617) );
  OAI222_X1 U7089 ( .A1(n13618), .A2(n10941), .B1(n13650), .B2(n10938), .C1(
        n13586), .C2(n10935), .ZN(n5623) );
  AOI221_X1 U7090 ( .B1(n10881), .B2(n14287), .C1(n10878), .C2(n14479), .A(
        n5632), .ZN(n5626) );
  OAI222_X1 U7091 ( .A1(n10478), .A2(n10875), .B1(n10477), .B2(n10872), .C1(
        n10479), .C2(n10869), .ZN(n5632) );
  AOI221_X1 U7092 ( .B1(n11211), .B2(n9505), .C1(n11208), .C2(n9537), .A(n4190), .ZN(n4184) );
  OAI222_X1 U7093 ( .A1(n13618), .A2(n11205), .B1(n13650), .B2(n11202), .C1(
        n13586), .C2(n11199), .ZN(n4190) );
  AOI221_X1 U7094 ( .B1(n11145), .B2(n14287), .C1(n11142), .C2(n14479), .A(
        n4199), .ZN(n4193) );
  OAI222_X1 U7095 ( .A1(n10478), .A2(n11139), .B1(n10477), .B2(n11136), .C1(
        n10479), .C2(n11133), .ZN(n4199) );
  AOI221_X1 U7096 ( .B1(n10947), .B2(n9506), .C1(n10944), .C2(n9538), .A(n5582), .ZN(n5576) );
  OAI222_X1 U7097 ( .A1(n13617), .A2(n10941), .B1(n13649), .B2(n10938), .C1(
        n13585), .C2(n10935), .ZN(n5582) );
  AOI221_X1 U7098 ( .B1(n10881), .B2(n14286), .C1(n10878), .C2(n14478), .A(
        n5591), .ZN(n5585) );
  OAI222_X1 U7099 ( .A1(n10446), .A2(n10875), .B1(n10445), .B2(n10872), .C1(
        n10447), .C2(n10869), .ZN(n5591) );
  AOI221_X1 U7100 ( .B1(n11211), .B2(n9506), .C1(n11208), .C2(n9538), .A(n4149), .ZN(n4143) );
  OAI222_X1 U7101 ( .A1(n13617), .A2(n11205), .B1(n13649), .B2(n11202), .C1(
        n13585), .C2(n11199), .ZN(n4149) );
  AOI221_X1 U7102 ( .B1(n11145), .B2(n14286), .C1(n11142), .C2(n14478), .A(
        n4158), .ZN(n4152) );
  OAI222_X1 U7103 ( .A1(n10446), .A2(n11139), .B1(n10445), .B2(n11136), .C1(
        n10447), .C2(n11133), .ZN(n4158) );
  AOI221_X1 U7104 ( .B1(n10947), .B2(n9507), .C1(n10944), .C2(n9539), .A(n5541), .ZN(n5535) );
  OAI222_X1 U7105 ( .A1(n13616), .A2(n10941), .B1(n13648), .B2(n10938), .C1(
        n13584), .C2(n10935), .ZN(n5541) );
  AOI221_X1 U7106 ( .B1(n10881), .B2(n14285), .C1(n10878), .C2(n14477), .A(
        n5550), .ZN(n5544) );
  OAI222_X1 U7107 ( .A1(n10414), .A2(n10875), .B1(n10413), .B2(n10872), .C1(
        n10415), .C2(n10869), .ZN(n5550) );
  AOI221_X1 U7108 ( .B1(n11211), .B2(n9507), .C1(n11208), .C2(n9539), .A(n4108), .ZN(n4102) );
  OAI222_X1 U7109 ( .A1(n13616), .A2(n11205), .B1(n13648), .B2(n11202), .C1(
        n13584), .C2(n11199), .ZN(n4108) );
  AOI221_X1 U7110 ( .B1(n11145), .B2(n14285), .C1(n11142), .C2(n14477), .A(
        n4117), .ZN(n4111) );
  OAI222_X1 U7111 ( .A1(n10414), .A2(n11139), .B1(n10413), .B2(n11136), .C1(
        n10415), .C2(n11133), .ZN(n4117) );
  AOI221_X1 U7112 ( .B1(n10947), .B2(n9508), .C1(n10944), .C2(n9540), .A(n5500), .ZN(n5494) );
  OAI222_X1 U7113 ( .A1(n13615), .A2(n10941), .B1(n13647), .B2(n10938), .C1(
        n13583), .C2(n10935), .ZN(n5500) );
  AOI221_X1 U7114 ( .B1(n10881), .B2(n14284), .C1(n10878), .C2(n14476), .A(
        n5509), .ZN(n5503) );
  OAI222_X1 U7115 ( .A1(n10379), .A2(n10875), .B1(n10378), .B2(n10872), .C1(
        n10380), .C2(n10869), .ZN(n5509) );
  AOI221_X1 U7116 ( .B1(n11211), .B2(n9508), .C1(n11208), .C2(n9540), .A(n4067), .ZN(n4061) );
  OAI222_X1 U7117 ( .A1(n13615), .A2(n11205), .B1(n13647), .B2(n11202), .C1(
        n13583), .C2(n11199), .ZN(n4067) );
  AOI221_X1 U7118 ( .B1(n11145), .B2(n14284), .C1(n11142), .C2(n14476), .A(
        n4076), .ZN(n4070) );
  OAI222_X1 U7119 ( .A1(n10379), .A2(n11139), .B1(n10378), .B2(n11136), .C1(
        n10380), .C2(n11133), .ZN(n4076) );
  AOI221_X1 U7120 ( .B1(n10947), .B2(n9509), .C1(n10944), .C2(n9541), .A(n5459), .ZN(n5453) );
  OAI222_X1 U7121 ( .A1(n13614), .A2(n10941), .B1(n13646), .B2(n10938), .C1(
        n13582), .C2(n10935), .ZN(n5459) );
  AOI221_X1 U7122 ( .B1(n10881), .B2(n14283), .C1(n10878), .C2(n14475), .A(
        n5468), .ZN(n5462) );
  OAI222_X1 U7123 ( .A1(n10347), .A2(n10875), .B1(n10346), .B2(n10872), .C1(
        n10348), .C2(n10869), .ZN(n5468) );
  AOI221_X1 U7124 ( .B1(n11211), .B2(n9509), .C1(n11208), .C2(n9541), .A(n4026), .ZN(n4020) );
  OAI222_X1 U7125 ( .A1(n13614), .A2(n11205), .B1(n13646), .B2(n11202), .C1(
        n13582), .C2(n11199), .ZN(n4026) );
  AOI221_X1 U7126 ( .B1(n11145), .B2(n14283), .C1(n11142), .C2(n14475), .A(
        n4035), .ZN(n4029) );
  OAI222_X1 U7127 ( .A1(n10347), .A2(n11139), .B1(n10346), .B2(n11136), .C1(
        n10348), .C2(n11133), .ZN(n4035) );
  AOI221_X1 U7128 ( .B1(n10947), .B2(n9510), .C1(n10944), .C2(n9542), .A(n5418), .ZN(n5412) );
  OAI222_X1 U7129 ( .A1(n13613), .A2(n10941), .B1(n13645), .B2(n10938), .C1(
        n13581), .C2(n10935), .ZN(n5418) );
  AOI221_X1 U7130 ( .B1(n10881), .B2(n14282), .C1(n10878), .C2(n14474), .A(
        n5427), .ZN(n5421) );
  OAI222_X1 U7131 ( .A1(n10315), .A2(n10875), .B1(n10314), .B2(n10872), .C1(
        n10316), .C2(n10869), .ZN(n5427) );
  AOI221_X1 U7132 ( .B1(n11211), .B2(n9510), .C1(n11208), .C2(n9542), .A(n3985), .ZN(n3979) );
  OAI222_X1 U7133 ( .A1(n13613), .A2(n11205), .B1(n13645), .B2(n11202), .C1(
        n13581), .C2(n11199), .ZN(n3985) );
  AOI221_X1 U7134 ( .B1(n11145), .B2(n14282), .C1(n11142), .C2(n14474), .A(
        n3994), .ZN(n3988) );
  OAI222_X1 U7135 ( .A1(n10315), .A2(n11139), .B1(n10314), .B2(n11136), .C1(
        n10316), .C2(n11133), .ZN(n3994) );
  AOI221_X1 U7136 ( .B1(n10947), .B2(n9511), .C1(n10944), .C2(n9543), .A(n5377), .ZN(n5371) );
  OAI222_X1 U7137 ( .A1(n13612), .A2(n10941), .B1(n13644), .B2(n10938), .C1(
        n13580), .C2(n10935), .ZN(n5377) );
  AOI221_X1 U7138 ( .B1(n10881), .B2(n14281), .C1(n10878), .C2(n14473), .A(
        n5386), .ZN(n5380) );
  OAI222_X1 U7139 ( .A1(n10280), .A2(n10875), .B1(n10279), .B2(n10872), .C1(
        n10281), .C2(n10869), .ZN(n5386) );
  AOI221_X1 U7140 ( .B1(n11211), .B2(n9511), .C1(n11208), .C2(n9543), .A(n3944), .ZN(n3938) );
  OAI222_X1 U7141 ( .A1(n13612), .A2(n11205), .B1(n13644), .B2(n11202), .C1(
        n13580), .C2(n11199), .ZN(n3944) );
  AOI221_X1 U7142 ( .B1(n11145), .B2(n14281), .C1(n11142), .C2(n14473), .A(
        n3953), .ZN(n3947) );
  OAI222_X1 U7143 ( .A1(n10280), .A2(n11139), .B1(n10279), .B2(n11136), .C1(
        n10281), .C2(n11133), .ZN(n3953) );
  AOI221_X1 U7144 ( .B1(n10947), .B2(n9512), .C1(n10944), .C2(n9544), .A(n5336), .ZN(n5330) );
  OAI222_X1 U7145 ( .A1(n13611), .A2(n10941), .B1(n13643), .B2(n10938), .C1(
        n13579), .C2(n10935), .ZN(n5336) );
  AOI221_X1 U7146 ( .B1(n10881), .B2(n14280), .C1(n10878), .C2(n14472), .A(
        n5345), .ZN(n5339) );
  OAI222_X1 U7147 ( .A1(n10248), .A2(n10875), .B1(n10247), .B2(n10872), .C1(
        n10249), .C2(n10869), .ZN(n5345) );
  AOI221_X1 U7148 ( .B1(n11211), .B2(n9512), .C1(n11208), .C2(n9544), .A(n3903), .ZN(n3897) );
  OAI222_X1 U7149 ( .A1(n13611), .A2(n11205), .B1(n13643), .B2(n11202), .C1(
        n13579), .C2(n11199), .ZN(n3903) );
  AOI221_X1 U7150 ( .B1(n11145), .B2(n14280), .C1(n11142), .C2(n14472), .A(
        n3912), .ZN(n3906) );
  OAI222_X1 U7151 ( .A1(n10248), .A2(n11139), .B1(n10247), .B2(n11136), .C1(
        n10249), .C2(n11133), .ZN(n3912) );
  AOI221_X1 U7152 ( .B1(n10947), .B2(n9513), .C1(n10944), .C2(n9545), .A(n5295), .ZN(n5289) );
  OAI222_X1 U7153 ( .A1(n13610), .A2(n10941), .B1(n13642), .B2(n10938), .C1(
        n13578), .C2(n10935), .ZN(n5295) );
  AOI221_X1 U7154 ( .B1(n10881), .B2(n14279), .C1(n10878), .C2(n14471), .A(
        n5304), .ZN(n5298) );
  OAI222_X1 U7155 ( .A1(n10216), .A2(n10875), .B1(n10215), .B2(n10872), .C1(
        n10217), .C2(n10869), .ZN(n5304) );
  AOI221_X1 U7156 ( .B1(n11211), .B2(n9513), .C1(n11208), .C2(n9545), .A(n3862), .ZN(n3856) );
  OAI222_X1 U7157 ( .A1(n13610), .A2(n11205), .B1(n13642), .B2(n11202), .C1(
        n13578), .C2(n11199), .ZN(n3862) );
  AOI221_X1 U7158 ( .B1(n11145), .B2(n14279), .C1(n11142), .C2(n14471), .A(
        n3871), .ZN(n3865) );
  OAI222_X1 U7159 ( .A1(n10216), .A2(n11139), .B1(n10215), .B2(n11136), .C1(
        n10217), .C2(n11133), .ZN(n3871) );
  AOI221_X1 U7160 ( .B1(n10947), .B2(n9514), .C1(n10944), .C2(n9546), .A(n5254), .ZN(n5248) );
  OAI222_X1 U7161 ( .A1(n13609), .A2(n10941), .B1(n13641), .B2(n10938), .C1(
        n13577), .C2(n10935), .ZN(n5254) );
  AOI221_X1 U7162 ( .B1(n10881), .B2(n14278), .C1(n10878), .C2(n14470), .A(
        n5263), .ZN(n5257) );
  OAI222_X1 U7163 ( .A1(n10182), .A2(n10875), .B1(n10181), .B2(n10872), .C1(
        n10183), .C2(n10869), .ZN(n5263) );
  AOI221_X1 U7164 ( .B1(n11211), .B2(n9514), .C1(n11208), .C2(n9546), .A(n3821), .ZN(n3815) );
  OAI222_X1 U7165 ( .A1(n13609), .A2(n11205), .B1(n13641), .B2(n11202), .C1(
        n13577), .C2(n11199), .ZN(n3821) );
  AOI221_X1 U7166 ( .B1(n11145), .B2(n14278), .C1(n11142), .C2(n14470), .A(
        n3830), .ZN(n3824) );
  OAI222_X1 U7167 ( .A1(n10182), .A2(n11139), .B1(n10181), .B2(n11136), .C1(
        n10183), .C2(n11133), .ZN(n3830) );
  AOI221_X1 U7168 ( .B1(n10947), .B2(n9515), .C1(n10944), .C2(n9547), .A(n5213), .ZN(n5207) );
  OAI222_X1 U7169 ( .A1(n13608), .A2(n10941), .B1(n13640), .B2(n10938), .C1(
        n13576), .C2(n10935), .ZN(n5213) );
  AOI221_X1 U7170 ( .B1(n10881), .B2(n14277), .C1(n10878), .C2(n14469), .A(
        n5222), .ZN(n5216) );
  OAI222_X1 U7171 ( .A1(n10150), .A2(n10875), .B1(n10149), .B2(n10872), .C1(
        n10151), .C2(n10869), .ZN(n5222) );
  AOI221_X1 U7172 ( .B1(n11211), .B2(n9515), .C1(n11208), .C2(n9547), .A(n3780), .ZN(n3774) );
  OAI222_X1 U7173 ( .A1(n13608), .A2(n11205), .B1(n13640), .B2(n11202), .C1(
        n13576), .C2(n11199), .ZN(n3780) );
  AOI221_X1 U7174 ( .B1(n11145), .B2(n14277), .C1(n11142), .C2(n14469), .A(
        n3789), .ZN(n3783) );
  OAI222_X1 U7175 ( .A1(n10150), .A2(n11139), .B1(n10149), .B2(n11136), .C1(
        n10151), .C2(n11133), .ZN(n3789) );
  AOI221_X1 U7176 ( .B1(n10948), .B2(n9516), .C1(n10945), .C2(n9548), .A(n5172), .ZN(n5166) );
  OAI222_X1 U7177 ( .A1(n13607), .A2(n10942), .B1(n13639), .B2(n10939), .C1(
        n13575), .C2(n10936), .ZN(n5172) );
  AOI221_X1 U7178 ( .B1(n10882), .B2(n14276), .C1(n10879), .C2(n14468), .A(
        n5181), .ZN(n5175) );
  OAI222_X1 U7179 ( .A1(n10118), .A2(n10876), .B1(n10117), .B2(n10873), .C1(
        n10119), .C2(n10870), .ZN(n5181) );
  AOI221_X1 U7180 ( .B1(n11212), .B2(n9516), .C1(n11209), .C2(n9548), .A(n3739), .ZN(n3733) );
  OAI222_X1 U7181 ( .A1(n13607), .A2(n11206), .B1(n13639), .B2(n11203), .C1(
        n13575), .C2(n11200), .ZN(n3739) );
  AOI221_X1 U7182 ( .B1(n11146), .B2(n14276), .C1(n11143), .C2(n14468), .A(
        n3748), .ZN(n3742) );
  OAI222_X1 U7183 ( .A1(n10118), .A2(n11140), .B1(n10117), .B2(n11137), .C1(
        n10119), .C2(n11134), .ZN(n3748) );
  AOI221_X1 U7184 ( .B1(n10948), .B2(n9517), .C1(n10945), .C2(n9549), .A(n5131), .ZN(n5125) );
  OAI222_X1 U7185 ( .A1(n13606), .A2(n10942), .B1(n13638), .B2(n10939), .C1(
        n13574), .C2(n10936), .ZN(n5131) );
  AOI221_X1 U7186 ( .B1(n10882), .B2(n14275), .C1(n10879), .C2(n14467), .A(
        n5140), .ZN(n5134) );
  OAI222_X1 U7187 ( .A1(n10086), .A2(n10876), .B1(n10085), .B2(n10873), .C1(
        n10087), .C2(n10870), .ZN(n5140) );
  AOI221_X1 U7188 ( .B1(n11212), .B2(n9517), .C1(n11209), .C2(n9549), .A(n3698), .ZN(n3692) );
  OAI222_X1 U7189 ( .A1(n13606), .A2(n11206), .B1(n13638), .B2(n11203), .C1(
        n13574), .C2(n11200), .ZN(n3698) );
  AOI221_X1 U7190 ( .B1(n11146), .B2(n14275), .C1(n11143), .C2(n14467), .A(
        n3707), .ZN(n3701) );
  OAI222_X1 U7191 ( .A1(n10086), .A2(n11140), .B1(n10085), .B2(n11137), .C1(
        n10087), .C2(n11134), .ZN(n3707) );
  AOI221_X1 U7192 ( .B1(n10948), .B2(n9518), .C1(n10945), .C2(n9550), .A(n5090), .ZN(n5084) );
  OAI222_X1 U7193 ( .A1(n13605), .A2(n10942), .B1(n13637), .B2(n10939), .C1(
        n13573), .C2(n10936), .ZN(n5090) );
  AOI221_X1 U7194 ( .B1(n10882), .B2(n14274), .C1(n10879), .C2(n14466), .A(
        n5099), .ZN(n5093) );
  OAI222_X1 U7195 ( .A1(n10054), .A2(n10876), .B1(n10053), .B2(n10873), .C1(
        n10055), .C2(n10870), .ZN(n5099) );
  AOI221_X1 U7196 ( .B1(n11212), .B2(n9518), .C1(n11209), .C2(n9550), .A(n3657), .ZN(n3651) );
  OAI222_X1 U7197 ( .A1(n13605), .A2(n11206), .B1(n13637), .B2(n11203), .C1(
        n13573), .C2(n11200), .ZN(n3657) );
  AOI221_X1 U7198 ( .B1(n11146), .B2(n14274), .C1(n11143), .C2(n14466), .A(
        n3666), .ZN(n3660) );
  OAI222_X1 U7199 ( .A1(n10054), .A2(n11140), .B1(n10053), .B2(n11137), .C1(
        n10055), .C2(n11134), .ZN(n3666) );
  AOI221_X1 U7200 ( .B1(n10948), .B2(n9519), .C1(n10945), .C2(n9551), .A(n5049), .ZN(n5043) );
  OAI222_X1 U7201 ( .A1(n13604), .A2(n10942), .B1(n13636), .B2(n10939), .C1(
        n13572), .C2(n10936), .ZN(n5049) );
  AOI221_X1 U7202 ( .B1(n10882), .B2(n14273), .C1(n10879), .C2(n14465), .A(
        n5058), .ZN(n5052) );
  OAI222_X1 U7203 ( .A1(n10022), .A2(n10876), .B1(n10021), .B2(n10873), .C1(
        n10023), .C2(n10870), .ZN(n5058) );
  AOI221_X1 U7204 ( .B1(n11212), .B2(n9519), .C1(n11209), .C2(n9551), .A(n3616), .ZN(n3610) );
  OAI222_X1 U7205 ( .A1(n13604), .A2(n11206), .B1(n13636), .B2(n11203), .C1(
        n13572), .C2(n11200), .ZN(n3616) );
  AOI221_X1 U7206 ( .B1(n11146), .B2(n14273), .C1(n11143), .C2(n14465), .A(
        n3625), .ZN(n3619) );
  OAI222_X1 U7207 ( .A1(n10022), .A2(n11140), .B1(n10021), .B2(n11137), .C1(
        n10023), .C2(n11134), .ZN(n3625) );
  AOI221_X1 U7208 ( .B1(n10948), .B2(n9520), .C1(n10945), .C2(n9552), .A(n5008), .ZN(n5002) );
  OAI222_X1 U7209 ( .A1(n13603), .A2(n10942), .B1(n13635), .B2(n10939), .C1(
        n13571), .C2(n10936), .ZN(n5008) );
  AOI221_X1 U7210 ( .B1(n10882), .B2(n14272), .C1(n10879), .C2(n14464), .A(
        n5017), .ZN(n5011) );
  OAI222_X1 U7211 ( .A1(n9660), .A2(n10876), .B1(n9659), .B2(n10873), .C1(
        n9661), .C2(n10870), .ZN(n5017) );
  AOI221_X1 U7212 ( .B1(n11212), .B2(n9520), .C1(n11209), .C2(n9552), .A(n3575), .ZN(n3569) );
  OAI222_X1 U7213 ( .A1(n13603), .A2(n11206), .B1(n13635), .B2(n11203), .C1(
        n13571), .C2(n11200), .ZN(n3575) );
  AOI221_X1 U7214 ( .B1(n11146), .B2(n14272), .C1(n11143), .C2(n14464), .A(
        n3584), .ZN(n3578) );
  OAI222_X1 U7215 ( .A1(n9660), .A2(n11140), .B1(n9659), .B2(n11137), .C1(
        n9661), .C2(n11134), .ZN(n3584) );
  AOI221_X1 U7216 ( .B1(n10948), .B2(n9521), .C1(n10945), .C2(n9553), .A(n4967), .ZN(n4961) );
  OAI222_X1 U7217 ( .A1(n13602), .A2(n10942), .B1(n13634), .B2(n10939), .C1(
        n13570), .C2(n10936), .ZN(n4967) );
  AOI221_X1 U7218 ( .B1(n10882), .B2(n14271), .C1(n10879), .C2(n14463), .A(
        n4976), .ZN(n4970) );
  OAI222_X1 U7219 ( .A1(n9628), .A2(n10876), .B1(n9627), .B2(n10873), .C1(
        n9629), .C2(n10870), .ZN(n4976) );
  AOI221_X1 U7220 ( .B1(n11212), .B2(n9521), .C1(n11209), .C2(n9553), .A(n3534), .ZN(n3528) );
  OAI222_X1 U7221 ( .A1(n13602), .A2(n11206), .B1(n13634), .B2(n11203), .C1(
        n13570), .C2(n11200), .ZN(n3534) );
  AOI221_X1 U7222 ( .B1(n11146), .B2(n14271), .C1(n11143), .C2(n14463), .A(
        n3543), .ZN(n3537) );
  OAI222_X1 U7223 ( .A1(n9628), .A2(n11140), .B1(n9627), .B2(n11137), .C1(
        n9629), .C2(n11134), .ZN(n3543) );
  AOI221_X1 U7224 ( .B1(n10948), .B2(n9522), .C1(n10945), .C2(n9554), .A(n4926), .ZN(n4920) );
  OAI222_X1 U7225 ( .A1(n13601), .A2(n10942), .B1(n13633), .B2(n10939), .C1(
        n13569), .C2(n10936), .ZN(n4926) );
  AOI221_X1 U7226 ( .B1(n10882), .B2(n14270), .C1(n10879), .C2(n14462), .A(
        n4935), .ZN(n4929) );
  OAI222_X1 U7227 ( .A1(n9596), .A2(n10876), .B1(n9595), .B2(n10873), .C1(
        n9597), .C2(n10870), .ZN(n4935) );
  AOI221_X1 U7228 ( .B1(n11212), .B2(n9522), .C1(n11209), .C2(n9554), .A(n3493), .ZN(n3487) );
  OAI222_X1 U7229 ( .A1(n13601), .A2(n11206), .B1(n13633), .B2(n11203), .C1(
        n13569), .C2(n11200), .ZN(n3493) );
  AOI221_X1 U7230 ( .B1(n11146), .B2(n14270), .C1(n11143), .C2(n14462), .A(
        n3502), .ZN(n3496) );
  OAI222_X1 U7231 ( .A1(n9596), .A2(n11140), .B1(n9595), .B2(n11137), .C1(
        n9597), .C2(n11134), .ZN(n3502) );
  AOI221_X1 U7232 ( .B1(n10948), .B2(n9523), .C1(n10945), .C2(n9555), .A(n4885), .ZN(n4879) );
  OAI222_X1 U7233 ( .A1(n13600), .A2(n10942), .B1(n13632), .B2(n10939), .C1(
        n13568), .C2(n10936), .ZN(n4885) );
  AOI221_X1 U7234 ( .B1(n10882), .B2(n14269), .C1(n10879), .C2(n14461), .A(
        n4894), .ZN(n4888) );
  OAI222_X1 U7235 ( .A1(n9262), .A2(n10876), .B1(n9261), .B2(n10873), .C1(
        n9263), .C2(n10870), .ZN(n4894) );
  AOI221_X1 U7236 ( .B1(n11212), .B2(n9523), .C1(n11209), .C2(n9555), .A(n3452), .ZN(n3446) );
  OAI222_X1 U7237 ( .A1(n13600), .A2(n11206), .B1(n13632), .B2(n11203), .C1(
        n13568), .C2(n11200), .ZN(n3452) );
  AOI221_X1 U7238 ( .B1(n11146), .B2(n14269), .C1(n11143), .C2(n14461), .A(
        n3461), .ZN(n3455) );
  OAI222_X1 U7239 ( .A1(n9262), .A2(n11140), .B1(n9261), .B2(n11137), .C1(
        n9263), .C2(n11134), .ZN(n3461) );
  AOI221_X1 U7240 ( .B1(n10948), .B2(n9524), .C1(n10945), .C2(n9556), .A(n4844), .ZN(n4838) );
  OAI222_X1 U7241 ( .A1(n13599), .A2(n10942), .B1(n13631), .B2(n10939), .C1(
        n13567), .C2(n10936), .ZN(n4844) );
  AOI221_X1 U7242 ( .B1(n10882), .B2(n14268), .C1(n10879), .C2(n14460), .A(
        n4853), .ZN(n4847) );
  OAI222_X1 U7243 ( .A1(n9198), .A2(n10876), .B1(n9197), .B2(n10873), .C1(
        n9199), .C2(n10870), .ZN(n4853) );
  AOI221_X1 U7244 ( .B1(n11212), .B2(n9524), .C1(n11209), .C2(n9556), .A(n3411), .ZN(n3405) );
  OAI222_X1 U7245 ( .A1(n13599), .A2(n11206), .B1(n13631), .B2(n11203), .C1(
        n13567), .C2(n11200), .ZN(n3411) );
  AOI221_X1 U7246 ( .B1(n11146), .B2(n14268), .C1(n11143), .C2(n14460), .A(
        n3420), .ZN(n3414) );
  OAI222_X1 U7247 ( .A1(n9198), .A2(n11140), .B1(n9197), .B2(n11137), .C1(
        n9199), .C2(n11134), .ZN(n3420) );
  AOI221_X1 U7248 ( .B1(n10948), .B2(n9525), .C1(n10945), .C2(n9557), .A(n4803), .ZN(n4797) );
  OAI222_X1 U7249 ( .A1(n13598), .A2(n10942), .B1(n13630), .B2(n10939), .C1(
        n13566), .C2(n10936), .ZN(n4803) );
  AOI221_X1 U7250 ( .B1(n10882), .B2(n14267), .C1(n10879), .C2(n14459), .A(
        n4812), .ZN(n4806) );
  OAI222_X1 U7251 ( .A1(n9166), .A2(n10876), .B1(n9165), .B2(n10873), .C1(
        n9167), .C2(n10870), .ZN(n4812) );
  AOI221_X1 U7252 ( .B1(n11212), .B2(n9525), .C1(n11209), .C2(n9557), .A(n3370), .ZN(n3364) );
  OAI222_X1 U7253 ( .A1(n13598), .A2(n11206), .B1(n13630), .B2(n11203), .C1(
        n13566), .C2(n11200), .ZN(n3370) );
  AOI221_X1 U7254 ( .B1(n11146), .B2(n14267), .C1(n11143), .C2(n14459), .A(
        n3379), .ZN(n3373) );
  OAI222_X1 U7255 ( .A1(n9166), .A2(n11140), .B1(n9165), .B2(n11137), .C1(
        n9167), .C2(n11134), .ZN(n3379) );
  AOI221_X1 U7256 ( .B1(n10948), .B2(n9526), .C1(n10945), .C2(n9558), .A(n4762), .ZN(n4756) );
  OAI222_X1 U7257 ( .A1(n13597), .A2(n10942), .B1(n13629), .B2(n10939), .C1(
        n13565), .C2(n10936), .ZN(n4762) );
  AOI221_X1 U7258 ( .B1(n10882), .B2(n14266), .C1(n10879), .C2(n14458), .A(
        n4771), .ZN(n4765) );
  OAI222_X1 U7259 ( .A1(n9134), .A2(n10876), .B1(n6315), .B2(n10873), .C1(
        n9135), .C2(n10870), .ZN(n4771) );
  AOI221_X1 U7260 ( .B1(n11212), .B2(n9526), .C1(n11209), .C2(n9558), .A(n3329), .ZN(n3323) );
  OAI222_X1 U7261 ( .A1(n13597), .A2(n11206), .B1(n13629), .B2(n11203), .C1(
        n13565), .C2(n11200), .ZN(n3329) );
  AOI221_X1 U7262 ( .B1(n11146), .B2(n14266), .C1(n11143), .C2(n14458), .A(
        n3338), .ZN(n3332) );
  OAI222_X1 U7263 ( .A1(n9134), .A2(n11140), .B1(n6315), .B2(n11137), .C1(
        n9135), .C2(n11134), .ZN(n3338) );
  AOI221_X1 U7264 ( .B1(n10948), .B2(n9527), .C1(n10945), .C2(n9559), .A(n4721), .ZN(n4715) );
  OAI222_X1 U7265 ( .A1(n13596), .A2(n10942), .B1(n13628), .B2(n10939), .C1(
        n13564), .C2(n10936), .ZN(n4721) );
  AOI221_X1 U7266 ( .B1(n10882), .B2(n14265), .C1(n10879), .C2(n14457), .A(
        n4730), .ZN(n4724) );
  OAI222_X1 U7267 ( .A1(n5999), .A2(n10876), .B1(n5998), .B2(n10873), .C1(
        n6000), .C2(n10870), .ZN(n4730) );
  AOI221_X1 U7268 ( .B1(n11212), .B2(n9527), .C1(n11209), .C2(n9559), .A(n3288), .ZN(n3282) );
  OAI222_X1 U7269 ( .A1(n13596), .A2(n11206), .B1(n13628), .B2(n11203), .C1(
        n13564), .C2(n11200), .ZN(n3288) );
  AOI221_X1 U7270 ( .B1(n11146), .B2(n14265), .C1(n11143), .C2(n14457), .A(
        n3297), .ZN(n3291) );
  OAI222_X1 U7271 ( .A1(n5999), .A2(n11140), .B1(n5998), .B2(n11137), .C1(
        n6000), .C2(n11134), .ZN(n3297) );
  AOI221_X1 U7272 ( .B1(n10949), .B2(n9528), .C1(n10946), .C2(n9560), .A(n4680), .ZN(n4674) );
  OAI222_X1 U7273 ( .A1(n13595), .A2(n10943), .B1(n13627), .B2(n10940), .C1(
        n13563), .C2(n10937), .ZN(n4680) );
  AOI221_X1 U7274 ( .B1(n10883), .B2(n14264), .C1(n10880), .C2(n14456), .A(
        n4689), .ZN(n4683) );
  OAI222_X1 U7275 ( .A1(n5935), .A2(n10877), .B1(n5934), .B2(n10874), .C1(
        n5936), .C2(n10871), .ZN(n4689) );
  AOI221_X1 U7276 ( .B1(n11213), .B2(n9528), .C1(n11210), .C2(n9560), .A(n3247), .ZN(n3241) );
  OAI222_X1 U7277 ( .A1(n13595), .A2(n11207), .B1(n13627), .B2(n11204), .C1(
        n13563), .C2(n11201), .ZN(n3247) );
  AOI221_X1 U7278 ( .B1(n11147), .B2(n14264), .C1(n11144), .C2(n14456), .A(
        n3256), .ZN(n3250) );
  OAI222_X1 U7279 ( .A1(n5935), .A2(n11141), .B1(n5934), .B2(n11138), .C1(
        n5936), .C2(n11135), .ZN(n3256) );
  AOI221_X1 U7280 ( .B1(n10949), .B2(n9529), .C1(n10946), .C2(n9561), .A(n4639), .ZN(n4633) );
  OAI222_X1 U7281 ( .A1(n13594), .A2(n10943), .B1(n13626), .B2(n10940), .C1(
        n13562), .C2(n10937), .ZN(n4639) );
  AOI221_X1 U7282 ( .B1(n10883), .B2(n14263), .C1(n10880), .C2(n14455), .A(
        n4648), .ZN(n4642) );
  OAI222_X1 U7283 ( .A1(n5903), .A2(n10877), .B1(n5902), .B2(n10874), .C1(
        n5904), .C2(n10871), .ZN(n4648) );
  AOI221_X1 U7284 ( .B1(n11213), .B2(n9529), .C1(n11210), .C2(n9561), .A(n3206), .ZN(n3200) );
  OAI222_X1 U7285 ( .A1(n13594), .A2(n11207), .B1(n13626), .B2(n11204), .C1(
        n13562), .C2(n11201), .ZN(n3206) );
  AOI221_X1 U7286 ( .B1(n11147), .B2(n14263), .C1(n11144), .C2(n14455), .A(
        n3215), .ZN(n3209) );
  OAI222_X1 U7287 ( .A1(n5903), .A2(n11141), .B1(n5902), .B2(n11138), .C1(
        n5904), .C2(n11135), .ZN(n3215) );
  AOI221_X1 U7288 ( .B1(n10949), .B2(n9530), .C1(n10946), .C2(n9562), .A(n4598), .ZN(n4592) );
  OAI222_X1 U7289 ( .A1(n13593), .A2(n10943), .B1(n13625), .B2(n10940), .C1(
        n13561), .C2(n10937), .ZN(n4598) );
  AOI221_X1 U7290 ( .B1(n10883), .B2(n14262), .C1(n10880), .C2(n14454), .A(
        n4607), .ZN(n4601) );
  OAI222_X1 U7291 ( .A1(n5871), .A2(n10877), .B1(n5870), .B2(n10874), .C1(
        n5872), .C2(n10871), .ZN(n4607) );
  AOI221_X1 U7292 ( .B1(n11213), .B2(n9530), .C1(n11210), .C2(n9562), .A(n3165), .ZN(n3159) );
  OAI222_X1 U7293 ( .A1(n13593), .A2(n11207), .B1(n13625), .B2(n11204), .C1(
        n13561), .C2(n11201), .ZN(n3165) );
  AOI221_X1 U7294 ( .B1(n11147), .B2(n14262), .C1(n11144), .C2(n14454), .A(
        n3174), .ZN(n3168) );
  OAI222_X1 U7295 ( .A1(n5871), .A2(n11141), .B1(n5870), .B2(n11138), .C1(
        n5872), .C2(n11135), .ZN(n3174) );
  AOI221_X1 U7296 ( .B1(n10949), .B2(n9531), .C1(n10946), .C2(n9563), .A(n4557), .ZN(n4551) );
  OAI222_X1 U7297 ( .A1(n13592), .A2(n10943), .B1(n13624), .B2(n10940), .C1(
        n13560), .C2(n10937), .ZN(n4557) );
  AOI221_X1 U7298 ( .B1(n10883), .B2(n14261), .C1(n10880), .C2(n14453), .A(
        n4566), .ZN(n4560) );
  OAI222_X1 U7299 ( .A1(n5839), .A2(n10877), .B1(n5838), .B2(n10874), .C1(
        n5840), .C2(n10871), .ZN(n4566) );
  AOI221_X1 U7300 ( .B1(n11213), .B2(n9531), .C1(n11210), .C2(n9563), .A(n3124), .ZN(n3118) );
  OAI222_X1 U7301 ( .A1(n13592), .A2(n11207), .B1(n13624), .B2(n11204), .C1(
        n13560), .C2(n11201), .ZN(n3124) );
  AOI221_X1 U7302 ( .B1(n11147), .B2(n14261), .C1(n11144), .C2(n14453), .A(
        n3133), .ZN(n3127) );
  OAI222_X1 U7303 ( .A1(n5839), .A2(n11141), .B1(n5838), .B2(n11138), .C1(
        n5840), .C2(n11135), .ZN(n3133) );
  AOI221_X1 U7304 ( .B1(n10949), .B2(n9532), .C1(n10946), .C2(n9564), .A(n4516), .ZN(n4510) );
  OAI222_X1 U7305 ( .A1(n13591), .A2(n10943), .B1(n13623), .B2(n10940), .C1(
        n13559), .C2(n10937), .ZN(n4516) );
  AOI221_X1 U7306 ( .B1(n10883), .B2(n14260), .C1(n10880), .C2(n14452), .A(
        n4525), .ZN(n4519) );
  OAI222_X1 U7307 ( .A1(n5807), .A2(n10877), .B1(n5806), .B2(n10874), .C1(
        n5808), .C2(n10871), .ZN(n4525) );
  AOI221_X1 U7308 ( .B1(n11213), .B2(n9532), .C1(n11210), .C2(n9564), .A(n3083), .ZN(n3077) );
  OAI222_X1 U7309 ( .A1(n13591), .A2(n11207), .B1(n13623), .B2(n11204), .C1(
        n13559), .C2(n11201), .ZN(n3083) );
  AOI221_X1 U7310 ( .B1(n11147), .B2(n14260), .C1(n11144), .C2(n14452), .A(
        n3092), .ZN(n3086) );
  OAI222_X1 U7311 ( .A1(n5807), .A2(n11141), .B1(n5806), .B2(n11138), .C1(
        n5808), .C2(n11135), .ZN(n3092) );
  AOI221_X1 U7312 ( .B1(n10949), .B2(n9533), .C1(n10946), .C2(n9565), .A(n4475), .ZN(n4469) );
  OAI222_X1 U7313 ( .A1(n13590), .A2(n10943), .B1(n13622), .B2(n10940), .C1(
        n13558), .C2(n10937), .ZN(n4475) );
  AOI221_X1 U7314 ( .B1(n10883), .B2(n14259), .C1(n10880), .C2(n14451), .A(
        n4484), .ZN(n4478) );
  OAI222_X1 U7315 ( .A1(n5775), .A2(n10877), .B1(n5774), .B2(n10874), .C1(
        n5776), .C2(n10871), .ZN(n4484) );
  AOI221_X1 U7316 ( .B1(n11213), .B2(n9533), .C1(n11210), .C2(n9565), .A(n3042), .ZN(n3036) );
  OAI222_X1 U7317 ( .A1(n13590), .A2(n11207), .B1(n13622), .B2(n11204), .C1(
        n13558), .C2(n11201), .ZN(n3042) );
  AOI221_X1 U7318 ( .B1(n11147), .B2(n14259), .C1(n11144), .C2(n14451), .A(
        n3051), .ZN(n3045) );
  OAI222_X1 U7319 ( .A1(n5775), .A2(n11141), .B1(n5774), .B2(n11138), .C1(
        n5776), .C2(n11135), .ZN(n3051) );
  AOI221_X1 U7320 ( .B1(n10949), .B2(n9534), .C1(n10946), .C2(n9566), .A(n4434), .ZN(n4428) );
  OAI222_X1 U7321 ( .A1(n13589), .A2(n10943), .B1(n13621), .B2(n10940), .C1(
        n13557), .C2(n10937), .ZN(n4434) );
  AOI221_X1 U7322 ( .B1(n10883), .B2(n14258), .C1(n10880), .C2(n14450), .A(
        n4443), .ZN(n4437) );
  OAI222_X1 U7323 ( .A1(n5743), .A2(n10877), .B1(n5742), .B2(n10874), .C1(
        n5744), .C2(n10871), .ZN(n4443) );
  AOI221_X1 U7324 ( .B1(n11213), .B2(n9534), .C1(n11210), .C2(n9566), .A(n3001), .ZN(n2995) );
  OAI222_X1 U7325 ( .A1(n13589), .A2(n11207), .B1(n13621), .B2(n11204), .C1(
        n13557), .C2(n11201), .ZN(n3001) );
  AOI221_X1 U7326 ( .B1(n11147), .B2(n14258), .C1(n11144), .C2(n14450), .A(
        n3010), .ZN(n3004) );
  OAI222_X1 U7327 ( .A1(n5743), .A2(n11141), .B1(n5742), .B2(n11138), .C1(
        n5744), .C2(n11135), .ZN(n3010) );
  AOI221_X1 U7328 ( .B1(n10949), .B2(n9535), .C1(n10946), .C2(n9567), .A(n4362), .ZN(n4343) );
  OAI222_X1 U7329 ( .A1(n13588), .A2(n10943), .B1(n13620), .B2(n10940), .C1(
        n13556), .C2(n10937), .ZN(n4362) );
  AOI221_X1 U7330 ( .B1(n10883), .B2(n14257), .C1(n10880), .C2(n14449), .A(
        n4393), .ZN(n4374) );
  OAI222_X1 U7331 ( .A1(n5711), .A2(n10877), .B1(n5710), .B2(n10874), .C1(
        n5712), .C2(n10871), .ZN(n4393) );
  AOI221_X1 U7332 ( .B1(n11213), .B2(n9535), .C1(n11210), .C2(n9567), .A(n2926), .ZN(n2875) );
  OAI222_X1 U7333 ( .A1(n13588), .A2(n11207), .B1(n13620), .B2(n11204), .C1(
        n13556), .C2(n11201), .ZN(n2926) );
  AOI221_X1 U7334 ( .B1(n11147), .B2(n14257), .C1(n11144), .C2(n14449), .A(
        n2960), .ZN(n2941) );
  OAI222_X1 U7335 ( .A1(n5711), .A2(n11141), .B1(n5710), .B2(n11138), .C1(
        n5712), .C2(n11135), .ZN(n2960) );
  NOR2_X1 U7336 ( .A1(N8431), .A2(N8434), .ZN(n5654) );
  NOR2_X1 U7337 ( .A1(N8575), .A2(N8578), .ZN(n4221) );
  OAI22_X1 U7338 ( .A1(n1955), .A2(n11114), .B1(n227), .B2(n11111), .ZN(n4661)
         );
  OAI22_X1 U7339 ( .A1(n5986), .A2(n11048), .B1(n5985), .B2(n11045), .ZN(n4670) );
  OAI22_X1 U7340 ( .A1(n1955), .A2(n11378), .B1(n227), .B2(n11375), .ZN(n3228)
         );
  OAI22_X1 U7341 ( .A1(n5986), .A2(n11312), .B1(n5985), .B2(n11309), .ZN(n3237) );
  OAI22_X1 U7342 ( .A1(n1943), .A2(n11114), .B1(n215), .B2(n11111), .ZN(n4620)
         );
  OAI22_X1 U7343 ( .A1(n5922), .A2(n11048), .B1(n5921), .B2(n11045), .ZN(n4629) );
  OAI22_X1 U7344 ( .A1(n1943), .A2(n11378), .B1(n215), .B2(n11375), .ZN(n3187)
         );
  OAI22_X1 U7345 ( .A1(n5922), .A2(n11312), .B1(n5921), .B2(n11309), .ZN(n3196) );
  OAI22_X1 U7346 ( .A1(n1931), .A2(n11114), .B1(n203), .B2(n11111), .ZN(n4579)
         );
  OAI22_X1 U7347 ( .A1(n5890), .A2(n11048), .B1(n5889), .B2(n11045), .ZN(n4588) );
  OAI22_X1 U7348 ( .A1(n1931), .A2(n11378), .B1(n203), .B2(n11375), .ZN(n3146)
         );
  OAI22_X1 U7349 ( .A1(n5890), .A2(n11312), .B1(n5889), .B2(n11309), .ZN(n3155) );
  OAI22_X1 U7350 ( .A1(n1919), .A2(n11114), .B1(n191), .B2(n11111), .ZN(n4538)
         );
  OAI22_X1 U7351 ( .A1(n5858), .A2(n11048), .B1(n5857), .B2(n11045), .ZN(n4547) );
  OAI22_X1 U7352 ( .A1(n1919), .A2(n11378), .B1(n191), .B2(n11375), .ZN(n3105)
         );
  OAI22_X1 U7353 ( .A1(n5858), .A2(n11312), .B1(n5857), .B2(n11309), .ZN(n3114) );
  OAI22_X1 U7354 ( .A1(n1907), .A2(n11114), .B1(n179), .B2(n11111), .ZN(n4497)
         );
  OAI22_X1 U7355 ( .A1(n5826), .A2(n11048), .B1(n5825), .B2(n11045), .ZN(n4506) );
  OAI22_X1 U7356 ( .A1(n1907), .A2(n11378), .B1(n179), .B2(n11375), .ZN(n3064)
         );
  OAI22_X1 U7357 ( .A1(n5826), .A2(n11312), .B1(n5825), .B2(n11309), .ZN(n3073) );
  OAI22_X1 U7358 ( .A1(n1895), .A2(n11114), .B1(n167), .B2(n11111), .ZN(n4456)
         );
  OAI22_X1 U7359 ( .A1(n5794), .A2(n11048), .B1(n5793), .B2(n11045), .ZN(n4465) );
  OAI22_X1 U7360 ( .A1(n1895), .A2(n11378), .B1(n167), .B2(n11375), .ZN(n3023)
         );
  OAI22_X1 U7361 ( .A1(n5794), .A2(n11312), .B1(n5793), .B2(n11309), .ZN(n3032) );
  OAI22_X1 U7362 ( .A1(n1883), .A2(n11114), .B1(n155), .B2(n11111), .ZN(n4415)
         );
  OAI22_X1 U7363 ( .A1(n5762), .A2(n11048), .B1(n5761), .B2(n11045), .ZN(n4424) );
  OAI22_X1 U7364 ( .A1(n1883), .A2(n11378), .B1(n155), .B2(n11375), .ZN(n2982)
         );
  OAI22_X1 U7365 ( .A1(n5762), .A2(n11312), .B1(n5761), .B2(n11309), .ZN(n2991) );
  OAI22_X1 U7366 ( .A1(n1871), .A2(n11114), .B1(n143), .B2(n11111), .ZN(n4286)
         );
  OAI22_X1 U7367 ( .A1(n5730), .A2(n11048), .B1(n5729), .B2(n11045), .ZN(n4317) );
  OAI22_X1 U7368 ( .A1(n1871), .A2(n11378), .B1(n143), .B2(n11375), .ZN(n2786)
         );
  OAI22_X1 U7369 ( .A1(n5730), .A2(n11312), .B1(n5729), .B2(n11309), .ZN(n2817) );
  OAI22_X1 U7370 ( .A1(n2339), .A2(n11112), .B1(n515), .B2(n11109), .ZN(n5645)
         );
  OAI22_X1 U7371 ( .A1(n10529), .A2(n11046), .B1(n10528), .B2(n11043), .ZN(
        n5673) );
  OAI22_X1 U7372 ( .A1(n2339), .A2(n11376), .B1(n515), .B2(n11373), .ZN(n4212)
         );
  OAI22_X1 U7373 ( .A1(n10529), .A2(n11310), .B1(n10528), .B2(n11307), .ZN(
        n4240) );
  OAI22_X1 U7374 ( .A1(n2327), .A2(n11112), .B1(n503), .B2(n11109), .ZN(n5604)
         );
  OAI22_X1 U7375 ( .A1(n10497), .A2(n11046), .B1(n10496), .B2(n11043), .ZN(
        n5613) );
  OAI22_X1 U7376 ( .A1(n2327), .A2(n11376), .B1(n503), .B2(n11373), .ZN(n4171)
         );
  OAI22_X1 U7377 ( .A1(n10497), .A2(n11310), .B1(n10496), .B2(n11307), .ZN(
        n4180) );
  OAI22_X1 U7378 ( .A1(n2315), .A2(n11112), .B1(n491), .B2(n11109), .ZN(n5563)
         );
  OAI22_X1 U7379 ( .A1(n10465), .A2(n11046), .B1(n10464), .B2(n11043), .ZN(
        n5572) );
  OAI22_X1 U7380 ( .A1(n2315), .A2(n11376), .B1(n491), .B2(n11373), .ZN(n4130)
         );
  OAI22_X1 U7381 ( .A1(n10465), .A2(n11310), .B1(n10464), .B2(n11307), .ZN(
        n4139) );
  OAI22_X1 U7382 ( .A1(n2303), .A2(n11112), .B1(n479), .B2(n11109), .ZN(n5522)
         );
  OAI22_X1 U7383 ( .A1(n10433), .A2(n11046), .B1(n10432), .B2(n11043), .ZN(
        n5531) );
  OAI22_X1 U7384 ( .A1(n2303), .A2(n11376), .B1(n479), .B2(n11373), .ZN(n4089)
         );
  OAI22_X1 U7385 ( .A1(n10433), .A2(n11310), .B1(n10432), .B2(n11307), .ZN(
        n4098) );
  OAI22_X1 U7386 ( .A1(n2291), .A2(n11112), .B1(n467), .B2(n11109), .ZN(n5481)
         );
  OAI22_X1 U7387 ( .A1(n10401), .A2(n11046), .B1(n10400), .B2(n11043), .ZN(
        n5490) );
  OAI22_X1 U7388 ( .A1(n2291), .A2(n11376), .B1(n467), .B2(n11373), .ZN(n4048)
         );
  OAI22_X1 U7389 ( .A1(n10401), .A2(n11310), .B1(n10400), .B2(n11307), .ZN(
        n4057) );
  OAI22_X1 U7390 ( .A1(n2279), .A2(n11112), .B1(n455), .B2(n11109), .ZN(n5440)
         );
  OAI22_X1 U7391 ( .A1(n10366), .A2(n11046), .B1(n10365), .B2(n11043), .ZN(
        n5449) );
  OAI22_X1 U7392 ( .A1(n2279), .A2(n11376), .B1(n455), .B2(n11373), .ZN(n4007)
         );
  OAI22_X1 U7393 ( .A1(n10366), .A2(n11310), .B1(n10365), .B2(n11307), .ZN(
        n4016) );
  OAI22_X1 U7394 ( .A1(n2267), .A2(n11112), .B1(n443), .B2(n11109), .ZN(n5399)
         );
  OAI22_X1 U7395 ( .A1(n10334), .A2(n11046), .B1(n10333), .B2(n11043), .ZN(
        n5408) );
  OAI22_X1 U7396 ( .A1(n2267), .A2(n11376), .B1(n443), .B2(n11373), .ZN(n3966)
         );
  OAI22_X1 U7397 ( .A1(n10334), .A2(n11310), .B1(n10333), .B2(n11307), .ZN(
        n3975) );
  OAI22_X1 U7398 ( .A1(n2255), .A2(n11112), .B1(n431), .B2(n11109), .ZN(n5358)
         );
  OAI22_X1 U7399 ( .A1(n10299), .A2(n11046), .B1(n10298), .B2(n11043), .ZN(
        n5367) );
  OAI22_X1 U7400 ( .A1(n2255), .A2(n11376), .B1(n431), .B2(n11373), .ZN(n3925)
         );
  OAI22_X1 U7401 ( .A1(n10299), .A2(n11310), .B1(n10298), .B2(n11307), .ZN(
        n3934) );
  OAI22_X1 U7402 ( .A1(n2243), .A2(n11112), .B1(n419), .B2(n11109), .ZN(n5317)
         );
  OAI22_X1 U7403 ( .A1(n10267), .A2(n11046), .B1(n10266), .B2(n11043), .ZN(
        n5326) );
  OAI22_X1 U7404 ( .A1(n2243), .A2(n11376), .B1(n419), .B2(n11373), .ZN(n3884)
         );
  OAI22_X1 U7405 ( .A1(n10267), .A2(n11310), .B1(n10266), .B2(n11307), .ZN(
        n3893) );
  OAI22_X1 U7406 ( .A1(n2231), .A2(n11112), .B1(n407), .B2(n11109), .ZN(n5276)
         );
  OAI22_X1 U7407 ( .A1(n10235), .A2(n11046), .B1(n10234), .B2(n11043), .ZN(
        n5285) );
  OAI22_X1 U7408 ( .A1(n2231), .A2(n11376), .B1(n407), .B2(n11373), .ZN(n3843)
         );
  OAI22_X1 U7409 ( .A1(n10235), .A2(n11310), .B1(n10234), .B2(n11307), .ZN(
        n3852) );
  OAI22_X1 U7410 ( .A1(n2219), .A2(n11112), .B1(n395), .B2(n11109), .ZN(n5235)
         );
  OAI22_X1 U7411 ( .A1(n10201), .A2(n11046), .B1(n10200), .B2(n11043), .ZN(
        n5244) );
  OAI22_X1 U7412 ( .A1(n2219), .A2(n11376), .B1(n395), .B2(n11373), .ZN(n3802)
         );
  OAI22_X1 U7413 ( .A1(n10201), .A2(n11310), .B1(n10200), .B2(n11307), .ZN(
        n3811) );
  OAI22_X1 U7414 ( .A1(n2175), .A2(n11112), .B1(n383), .B2(n11109), .ZN(n5194)
         );
  OAI22_X1 U7415 ( .A1(n10169), .A2(n11046), .B1(n10168), .B2(n11043), .ZN(
        n5203) );
  OAI22_X1 U7416 ( .A1(n2175), .A2(n11376), .B1(n383), .B2(n11373), .ZN(n3761)
         );
  OAI22_X1 U7417 ( .A1(n10169), .A2(n11310), .B1(n10168), .B2(n11307), .ZN(
        n3770) );
  OAI22_X1 U7418 ( .A1(n2163), .A2(n11113), .B1(n371), .B2(n11110), .ZN(n5153)
         );
  OAI22_X1 U7419 ( .A1(n10137), .A2(n11047), .B1(n10136), .B2(n11044), .ZN(
        n5162) );
  OAI22_X1 U7420 ( .A1(n2163), .A2(n11377), .B1(n371), .B2(n11374), .ZN(n3720)
         );
  OAI22_X1 U7421 ( .A1(n10137), .A2(n11311), .B1(n10136), .B2(n11308), .ZN(
        n3729) );
  OAI22_X1 U7422 ( .A1(n2151), .A2(n11113), .B1(n359), .B2(n11110), .ZN(n5112)
         );
  OAI22_X1 U7423 ( .A1(n10105), .A2(n11047), .B1(n10104), .B2(n11044), .ZN(
        n5121) );
  OAI22_X1 U7424 ( .A1(n2151), .A2(n11377), .B1(n359), .B2(n11374), .ZN(n3679)
         );
  OAI22_X1 U7425 ( .A1(n10105), .A2(n11311), .B1(n10104), .B2(n11308), .ZN(
        n3688) );
  OAI22_X1 U7426 ( .A1(n2107), .A2(n11113), .B1(n347), .B2(n11110), .ZN(n5071)
         );
  OAI22_X1 U7427 ( .A1(n10073), .A2(n11047), .B1(n10072), .B2(n11044), .ZN(
        n5080) );
  OAI22_X1 U7428 ( .A1(n2107), .A2(n11377), .B1(n347), .B2(n11374), .ZN(n3638)
         );
  OAI22_X1 U7429 ( .A1(n10073), .A2(n11311), .B1(n10072), .B2(n11308), .ZN(
        n3647) );
  OAI22_X1 U7430 ( .A1(n2095), .A2(n11113), .B1(n335), .B2(n11110), .ZN(n5030)
         );
  OAI22_X1 U7431 ( .A1(n10041), .A2(n11047), .B1(n10040), .B2(n11044), .ZN(
        n5039) );
  OAI22_X1 U7432 ( .A1(n2095), .A2(n11377), .B1(n335), .B2(n11374), .ZN(n3597)
         );
  OAI22_X1 U7433 ( .A1(n10041), .A2(n11311), .B1(n10040), .B2(n11308), .ZN(
        n3606) );
  OAI22_X1 U7434 ( .A1(n2083), .A2(n11113), .B1(n323), .B2(n11110), .ZN(n4989)
         );
  OAI22_X1 U7435 ( .A1(n10009), .A2(n11047), .B1(n10008), .B2(n11044), .ZN(
        n4998) );
  OAI22_X1 U7436 ( .A1(n2083), .A2(n11377), .B1(n323), .B2(n11374), .ZN(n3556)
         );
  OAI22_X1 U7437 ( .A1(n10009), .A2(n11311), .B1(n10008), .B2(n11308), .ZN(
        n3565) );
  OAI22_X1 U7438 ( .A1(n2039), .A2(n11113), .B1(n311), .B2(n11110), .ZN(n4948)
         );
  OAI22_X1 U7439 ( .A1(n9647), .A2(n11047), .B1(n9646), .B2(n11044), .ZN(n4957) );
  OAI22_X1 U7440 ( .A1(n2039), .A2(n11377), .B1(n311), .B2(n11374), .ZN(n3515)
         );
  OAI22_X1 U7441 ( .A1(n9647), .A2(n11311), .B1(n9646), .B2(n11308), .ZN(n3524) );
  OAI22_X1 U7442 ( .A1(n2027), .A2(n11113), .B1(n299), .B2(n11110), .ZN(n4907)
         );
  OAI22_X1 U7443 ( .A1(n9615), .A2(n11047), .B1(n9614), .B2(n11044), .ZN(n4916) );
  OAI22_X1 U7444 ( .A1(n2027), .A2(n11377), .B1(n299), .B2(n11374), .ZN(n3474)
         );
  OAI22_X1 U7445 ( .A1(n9615), .A2(n11311), .B1(n9614), .B2(n11308), .ZN(n3483) );
  OAI22_X1 U7446 ( .A1(n2015), .A2(n11113), .B1(n287), .B2(n11110), .ZN(n4866)
         );
  OAI22_X1 U7447 ( .A1(n9583), .A2(n11047), .B1(n9582), .B2(n11044), .ZN(n4875) );
  OAI22_X1 U7448 ( .A1(n2015), .A2(n11377), .B1(n287), .B2(n11374), .ZN(n3433)
         );
  OAI22_X1 U7449 ( .A1(n9583), .A2(n11311), .B1(n9582), .B2(n11308), .ZN(n3442) );
  OAI22_X1 U7450 ( .A1(n2003), .A2(n11113), .B1(n275), .B2(n11110), .ZN(n4825)
         );
  OAI22_X1 U7451 ( .A1(n9249), .A2(n11047), .B1(n9248), .B2(n11044), .ZN(n4834) );
  OAI22_X1 U7452 ( .A1(n2003), .A2(n11377), .B1(n275), .B2(n11374), .ZN(n3392)
         );
  OAI22_X1 U7453 ( .A1(n9249), .A2(n11311), .B1(n9248), .B2(n11308), .ZN(n3401) );
  OAI22_X1 U7454 ( .A1(n1991), .A2(n11113), .B1(n263), .B2(n11110), .ZN(n4784)
         );
  OAI22_X1 U7455 ( .A1(n9185), .A2(n11047), .B1(n9184), .B2(n11044), .ZN(n4793) );
  OAI22_X1 U7456 ( .A1(n1991), .A2(n11377), .B1(n263), .B2(n11374), .ZN(n3351)
         );
  OAI22_X1 U7457 ( .A1(n9185), .A2(n11311), .B1(n9184), .B2(n11308), .ZN(n3360) );
  OAI22_X1 U7458 ( .A1(n1979), .A2(n11113), .B1(n251), .B2(n11110), .ZN(n4743)
         );
  OAI22_X1 U7459 ( .A1(n9153), .A2(n11047), .B1(n9152), .B2(n11044), .ZN(n4752) );
  OAI22_X1 U7460 ( .A1(n1979), .A2(n11377), .B1(n251), .B2(n11374), .ZN(n3310)
         );
  OAI22_X1 U7461 ( .A1(n9153), .A2(n11311), .B1(n9152), .B2(n11308), .ZN(n3319) );
  OAI22_X1 U7462 ( .A1(n1967), .A2(n11113), .B1(n239), .B2(n11110), .ZN(n4702)
         );
  OAI22_X1 U7463 ( .A1(n6303), .A2(n11047), .B1(n6302), .B2(n11044), .ZN(n4711) );
  OAI22_X1 U7464 ( .A1(n1967), .A2(n11377), .B1(n239), .B2(n11374), .ZN(n3269)
         );
  OAI22_X1 U7465 ( .A1(n6303), .A2(n11311), .B1(n6302), .B2(n11308), .ZN(n3278) );
  AND2_X1 U7466 ( .A1(N8432), .A2(N8433), .ZN(n5651) );
  AND2_X1 U7467 ( .A1(N8576), .A2(N8577), .ZN(n4218) );
  AND2_X1 U7468 ( .A1(N8433), .A2(n14513), .ZN(n5650) );
  AND2_X1 U7469 ( .A1(N8577), .A2(n14515), .ZN(n4217) );
  NOR2_X1 U7470 ( .A1(n12772), .A2(N8431), .ZN(n5703) );
  NOR2_X1 U7471 ( .A1(n12776), .A2(N8575), .ZN(n4270) );
  XNOR2_X1 U7472 ( .A(\U3/U97/Z_6 ), .B(\r472/n4 ), .ZN(N2173) );
  NAND2_X1 U7473 ( .A1(\U3/U97/Z_5 ), .A2(\r472/carry[5] ), .ZN(\r472/n4 ) );
  NOR2_X1 U7474 ( .A1(n2935), .A2(\r472/B[3] ), .ZN(\U3/U97/Z_6 ) );
  NOR2_X1 U7475 ( .A1(n12735), .A2(N2167), .ZN(n2719) );
  NOR2_X1 U7476 ( .A1(n12736), .A2(N2168), .ZN(n2721) );
  NOR2_X1 U7477 ( .A1(N2167), .A2(N2168), .ZN(n2723) );
  NOR2_X1 U7478 ( .A1(N2169), .A2(N2170), .ZN(n2735) );
  NAND4_X1 U7479 ( .A1(n5666), .A2(n5667), .A3(n5668), .A4(n5669), .ZN(n5636)
         );
  AOI221_X1 U7480 ( .B1(n11013), .B2(n9952), .C1(n11010), .C2(n9984), .A(n5677), .ZN(n5668) );
  NOR4_X1 U7481 ( .A1(n5670), .A2(n5671), .A3(n5672), .A4(n5673), .ZN(n5669)
         );
  AOI222_X1 U7482 ( .A1(n10989), .A2(n9824), .B1(n10986), .B2(n9760), .C1(
        n10983), .C2(n9792), .ZN(n5666) );
  NAND4_X1 U7483 ( .A1(n4233), .A2(n4234), .A3(n4235), .A4(n4236), .ZN(n4203)
         );
  AOI221_X1 U7484 ( .B1(n11277), .B2(n9952), .C1(n11274), .C2(n9984), .A(n4244), .ZN(n4235) );
  NOR4_X1 U7485 ( .A1(n4237), .A2(n4238), .A3(n4239), .A4(n4240), .ZN(n4236)
         );
  AOI222_X1 U7486 ( .A1(n11253), .A2(n9824), .B1(n11250), .B2(n9760), .C1(
        n11247), .C2(n9792), .ZN(n4233) );
  NAND4_X1 U7487 ( .A1(n5606), .A2(n5607), .A3(n5608), .A4(n5609), .ZN(n5595)
         );
  AOI221_X1 U7488 ( .B1(n11013), .B2(n9953), .C1(n11010), .C2(n9985), .A(n5614), .ZN(n5608) );
  NOR4_X1 U7489 ( .A1(n5610), .A2(n5611), .A3(n5612), .A4(n5613), .ZN(n5609)
         );
  AOI222_X1 U7490 ( .A1(n10989), .A2(n9825), .B1(n10986), .B2(n9761), .C1(
        n10983), .C2(n9793), .ZN(n5606) );
  NAND4_X1 U7491 ( .A1(n4173), .A2(n4174), .A3(n4175), .A4(n4176), .ZN(n4162)
         );
  AOI221_X1 U7492 ( .B1(n11277), .B2(n9953), .C1(n11274), .C2(n9985), .A(n4181), .ZN(n4175) );
  NOR4_X1 U7493 ( .A1(n4177), .A2(n4178), .A3(n4179), .A4(n4180), .ZN(n4176)
         );
  AOI222_X1 U7494 ( .A1(n11253), .A2(n9825), .B1(n11250), .B2(n9761), .C1(
        n11247), .C2(n9793), .ZN(n4173) );
  NAND4_X1 U7495 ( .A1(n5565), .A2(n5566), .A3(n5567), .A4(n5568), .ZN(n5554)
         );
  AOI221_X1 U7496 ( .B1(n11013), .B2(n9954), .C1(n11010), .C2(n9986), .A(n5573), .ZN(n5567) );
  NOR4_X1 U7497 ( .A1(n5569), .A2(n5570), .A3(n5571), .A4(n5572), .ZN(n5568)
         );
  AOI222_X1 U7498 ( .A1(n10989), .A2(n9826), .B1(n10986), .B2(n9762), .C1(
        n10983), .C2(n9794), .ZN(n5565) );
  NAND4_X1 U7499 ( .A1(n4132), .A2(n4133), .A3(n4134), .A4(n4135), .ZN(n4121)
         );
  AOI221_X1 U7500 ( .B1(n11277), .B2(n9954), .C1(n11274), .C2(n9986), .A(n4140), .ZN(n4134) );
  NOR4_X1 U7501 ( .A1(n4136), .A2(n4137), .A3(n4138), .A4(n4139), .ZN(n4135)
         );
  AOI222_X1 U7502 ( .A1(n11253), .A2(n9826), .B1(n11250), .B2(n9762), .C1(
        n11247), .C2(n9794), .ZN(n4132) );
  NAND4_X1 U7503 ( .A1(n5524), .A2(n5525), .A3(n5526), .A4(n5527), .ZN(n5513)
         );
  AOI221_X1 U7504 ( .B1(n11013), .B2(n9955), .C1(n11010), .C2(n9987), .A(n5532), .ZN(n5526) );
  NOR4_X1 U7505 ( .A1(n5528), .A2(n5529), .A3(n5530), .A4(n5531), .ZN(n5527)
         );
  AOI222_X1 U7506 ( .A1(n10989), .A2(n9827), .B1(n10986), .B2(n9763), .C1(
        n10983), .C2(n9795), .ZN(n5524) );
  NAND4_X1 U7507 ( .A1(n4091), .A2(n4092), .A3(n4093), .A4(n4094), .ZN(n4080)
         );
  AOI221_X1 U7508 ( .B1(n11277), .B2(n9955), .C1(n11274), .C2(n9987), .A(n4099), .ZN(n4093) );
  NOR4_X1 U7509 ( .A1(n4095), .A2(n4096), .A3(n4097), .A4(n4098), .ZN(n4094)
         );
  AOI222_X1 U7510 ( .A1(n11253), .A2(n9827), .B1(n11250), .B2(n9763), .C1(
        n11247), .C2(n9795), .ZN(n4091) );
  NAND4_X1 U7511 ( .A1(n5483), .A2(n5484), .A3(n5485), .A4(n5486), .ZN(n5472)
         );
  AOI221_X1 U7512 ( .B1(n11013), .B2(n9956), .C1(n11010), .C2(n9988), .A(n5491), .ZN(n5485) );
  NOR4_X1 U7513 ( .A1(n5487), .A2(n5488), .A3(n5489), .A4(n5490), .ZN(n5486)
         );
  AOI222_X1 U7514 ( .A1(n10989), .A2(n9828), .B1(n10986), .B2(n9764), .C1(
        n10983), .C2(n9796), .ZN(n5483) );
  NAND4_X1 U7515 ( .A1(n4050), .A2(n4051), .A3(n4052), .A4(n4053), .ZN(n4039)
         );
  AOI221_X1 U7516 ( .B1(n11277), .B2(n9956), .C1(n11274), .C2(n9988), .A(n4058), .ZN(n4052) );
  NOR4_X1 U7517 ( .A1(n4054), .A2(n4055), .A3(n4056), .A4(n4057), .ZN(n4053)
         );
  AOI222_X1 U7518 ( .A1(n11253), .A2(n9828), .B1(n11250), .B2(n9764), .C1(
        n11247), .C2(n9796), .ZN(n4050) );
  NAND4_X1 U7519 ( .A1(n5442), .A2(n5443), .A3(n5444), .A4(n5445), .ZN(n5431)
         );
  AOI221_X1 U7520 ( .B1(n11013), .B2(n9957), .C1(n11010), .C2(n9989), .A(n5450), .ZN(n5444) );
  NOR4_X1 U7521 ( .A1(n5446), .A2(n5447), .A3(n5448), .A4(n5449), .ZN(n5445)
         );
  AOI222_X1 U7522 ( .A1(n10989), .A2(n9829), .B1(n10986), .B2(n9765), .C1(
        n10983), .C2(n9797), .ZN(n5442) );
  NAND4_X1 U7523 ( .A1(n4009), .A2(n4010), .A3(n4011), .A4(n4012), .ZN(n3998)
         );
  AOI221_X1 U7524 ( .B1(n11277), .B2(n9957), .C1(n11274), .C2(n9989), .A(n4017), .ZN(n4011) );
  NOR4_X1 U7525 ( .A1(n4013), .A2(n4014), .A3(n4015), .A4(n4016), .ZN(n4012)
         );
  AOI222_X1 U7526 ( .A1(n11253), .A2(n9829), .B1(n11250), .B2(n9765), .C1(
        n11247), .C2(n9797), .ZN(n4009) );
  NAND4_X1 U7527 ( .A1(n5401), .A2(n5402), .A3(n5403), .A4(n5404), .ZN(n5390)
         );
  AOI221_X1 U7528 ( .B1(n11013), .B2(n9958), .C1(n11010), .C2(n9990), .A(n5409), .ZN(n5403) );
  NOR4_X1 U7529 ( .A1(n5405), .A2(n5406), .A3(n5407), .A4(n5408), .ZN(n5404)
         );
  AOI222_X1 U7530 ( .A1(n10989), .A2(n9830), .B1(n10986), .B2(n9766), .C1(
        n10983), .C2(n9798), .ZN(n5401) );
  NAND4_X1 U7531 ( .A1(n3968), .A2(n3969), .A3(n3970), .A4(n3971), .ZN(n3957)
         );
  AOI221_X1 U7532 ( .B1(n11277), .B2(n9958), .C1(n11274), .C2(n9990), .A(n3976), .ZN(n3970) );
  NOR4_X1 U7533 ( .A1(n3972), .A2(n3973), .A3(n3974), .A4(n3975), .ZN(n3971)
         );
  AOI222_X1 U7534 ( .A1(n11253), .A2(n9830), .B1(n11250), .B2(n9766), .C1(
        n11247), .C2(n9798), .ZN(n3968) );
  NAND4_X1 U7535 ( .A1(n5360), .A2(n5361), .A3(n5362), .A4(n5363), .ZN(n5349)
         );
  AOI221_X1 U7536 ( .B1(n11013), .B2(n9959), .C1(n11010), .C2(n9991), .A(n5368), .ZN(n5362) );
  NOR4_X1 U7537 ( .A1(n5364), .A2(n5365), .A3(n5366), .A4(n5367), .ZN(n5363)
         );
  AOI222_X1 U7538 ( .A1(n10989), .A2(n9831), .B1(n10986), .B2(n9767), .C1(
        n10983), .C2(n9799), .ZN(n5360) );
  NAND4_X1 U7539 ( .A1(n3927), .A2(n3928), .A3(n3929), .A4(n3930), .ZN(n3916)
         );
  AOI221_X1 U7540 ( .B1(n11277), .B2(n9959), .C1(n11274), .C2(n9991), .A(n3935), .ZN(n3929) );
  NOR4_X1 U7541 ( .A1(n3931), .A2(n3932), .A3(n3933), .A4(n3934), .ZN(n3930)
         );
  AOI222_X1 U7542 ( .A1(n11253), .A2(n9831), .B1(n11250), .B2(n9767), .C1(
        n11247), .C2(n9799), .ZN(n3927) );
  NAND4_X1 U7543 ( .A1(n5319), .A2(n5320), .A3(n5321), .A4(n5322), .ZN(n5308)
         );
  AOI221_X1 U7544 ( .B1(n11013), .B2(n9960), .C1(n11010), .C2(n9992), .A(n5327), .ZN(n5321) );
  NOR4_X1 U7545 ( .A1(n5323), .A2(n5324), .A3(n5325), .A4(n5326), .ZN(n5322)
         );
  AOI222_X1 U7546 ( .A1(n10989), .A2(n9832), .B1(n10986), .B2(n9768), .C1(
        n10983), .C2(n9800), .ZN(n5319) );
  NAND4_X1 U7547 ( .A1(n3886), .A2(n3887), .A3(n3888), .A4(n3889), .ZN(n3875)
         );
  AOI221_X1 U7548 ( .B1(n11277), .B2(n9960), .C1(n11274), .C2(n9992), .A(n3894), .ZN(n3888) );
  NOR4_X1 U7549 ( .A1(n3890), .A2(n3891), .A3(n3892), .A4(n3893), .ZN(n3889)
         );
  AOI222_X1 U7550 ( .A1(n11253), .A2(n9832), .B1(n11250), .B2(n9768), .C1(
        n11247), .C2(n9800), .ZN(n3886) );
  NAND4_X1 U7551 ( .A1(n5278), .A2(n5279), .A3(n5280), .A4(n5281), .ZN(n5267)
         );
  AOI221_X1 U7552 ( .B1(n11013), .B2(n9961), .C1(n11010), .C2(n9993), .A(n5286), .ZN(n5280) );
  NOR4_X1 U7553 ( .A1(n5282), .A2(n5283), .A3(n5284), .A4(n5285), .ZN(n5281)
         );
  AOI222_X1 U7554 ( .A1(n10989), .A2(n9833), .B1(n10986), .B2(n9769), .C1(
        n10983), .C2(n9801), .ZN(n5278) );
  NAND4_X1 U7555 ( .A1(n3845), .A2(n3846), .A3(n3847), .A4(n3848), .ZN(n3834)
         );
  AOI221_X1 U7556 ( .B1(n11277), .B2(n9961), .C1(n11274), .C2(n9993), .A(n3853), .ZN(n3847) );
  NOR4_X1 U7557 ( .A1(n3849), .A2(n3850), .A3(n3851), .A4(n3852), .ZN(n3848)
         );
  AOI222_X1 U7558 ( .A1(n11253), .A2(n9833), .B1(n11250), .B2(n9769), .C1(
        n11247), .C2(n9801), .ZN(n3845) );
  NAND4_X1 U7559 ( .A1(n5237), .A2(n5238), .A3(n5239), .A4(n5240), .ZN(n5226)
         );
  AOI221_X1 U7560 ( .B1(n11013), .B2(n9962), .C1(n11010), .C2(n9994), .A(n5245), .ZN(n5239) );
  NOR4_X1 U7561 ( .A1(n5241), .A2(n5242), .A3(n5243), .A4(n5244), .ZN(n5240)
         );
  AOI222_X1 U7562 ( .A1(n10989), .A2(n9834), .B1(n10986), .B2(n9770), .C1(
        n10983), .C2(n9802), .ZN(n5237) );
  NAND4_X1 U7563 ( .A1(n3804), .A2(n3805), .A3(n3806), .A4(n3807), .ZN(n3793)
         );
  AOI221_X1 U7564 ( .B1(n11277), .B2(n9962), .C1(n11274), .C2(n9994), .A(n3812), .ZN(n3806) );
  NOR4_X1 U7565 ( .A1(n3808), .A2(n3809), .A3(n3810), .A4(n3811), .ZN(n3807)
         );
  AOI222_X1 U7566 ( .A1(n11253), .A2(n9834), .B1(n11250), .B2(n9770), .C1(
        n11247), .C2(n9802), .ZN(n3804) );
  NAND4_X1 U7567 ( .A1(n5196), .A2(n5197), .A3(n5198), .A4(n5199), .ZN(n5185)
         );
  AOI221_X1 U7568 ( .B1(n11013), .B2(n9963), .C1(n11010), .C2(n9995), .A(n5204), .ZN(n5198) );
  NOR4_X1 U7569 ( .A1(n5200), .A2(n5201), .A3(n5202), .A4(n5203), .ZN(n5199)
         );
  AOI222_X1 U7570 ( .A1(n10989), .A2(n9835), .B1(n10986), .B2(n9771), .C1(
        n10983), .C2(n9803), .ZN(n5196) );
  NAND4_X1 U7571 ( .A1(n3763), .A2(n3764), .A3(n3765), .A4(n3766), .ZN(n3752)
         );
  AOI221_X1 U7572 ( .B1(n11277), .B2(n9963), .C1(n11274), .C2(n9995), .A(n3771), .ZN(n3765) );
  NOR4_X1 U7573 ( .A1(n3767), .A2(n3768), .A3(n3769), .A4(n3770), .ZN(n3766)
         );
  AOI222_X1 U7574 ( .A1(n11253), .A2(n9835), .B1(n11250), .B2(n9771), .C1(
        n11247), .C2(n9803), .ZN(n3763) );
  NAND4_X1 U7575 ( .A1(n5155), .A2(n5156), .A3(n5157), .A4(n5158), .ZN(n5144)
         );
  AOI221_X1 U7576 ( .B1(n11014), .B2(n9964), .C1(n11011), .C2(n9996), .A(n5163), .ZN(n5157) );
  NOR4_X1 U7577 ( .A1(n5159), .A2(n5160), .A3(n5161), .A4(n5162), .ZN(n5158)
         );
  AOI222_X1 U7578 ( .A1(n10990), .A2(n9836), .B1(n10987), .B2(n9772), .C1(
        n10984), .C2(n9804), .ZN(n5155) );
  NAND4_X1 U7579 ( .A1(n3722), .A2(n3723), .A3(n3724), .A4(n3725), .ZN(n3711)
         );
  AOI221_X1 U7580 ( .B1(n11278), .B2(n9964), .C1(n11275), .C2(n9996), .A(n3730), .ZN(n3724) );
  NOR4_X1 U7581 ( .A1(n3726), .A2(n3727), .A3(n3728), .A4(n3729), .ZN(n3725)
         );
  AOI222_X1 U7582 ( .A1(n11254), .A2(n9836), .B1(n11251), .B2(n9772), .C1(
        n11248), .C2(n9804), .ZN(n3722) );
  NAND4_X1 U7583 ( .A1(n5114), .A2(n5115), .A3(n5116), .A4(n5117), .ZN(n5103)
         );
  AOI221_X1 U7584 ( .B1(n11014), .B2(n9965), .C1(n11011), .C2(n9997), .A(n5122), .ZN(n5116) );
  NOR4_X1 U7585 ( .A1(n5118), .A2(n5119), .A3(n5120), .A4(n5121), .ZN(n5117)
         );
  AOI222_X1 U7586 ( .A1(n10990), .A2(n9837), .B1(n10987), .B2(n9773), .C1(
        n10984), .C2(n9805), .ZN(n5114) );
  NAND4_X1 U7587 ( .A1(n3681), .A2(n3682), .A3(n3683), .A4(n3684), .ZN(n3670)
         );
  AOI221_X1 U7588 ( .B1(n11278), .B2(n9965), .C1(n11275), .C2(n9997), .A(n3689), .ZN(n3683) );
  NOR4_X1 U7589 ( .A1(n3685), .A2(n3686), .A3(n3687), .A4(n3688), .ZN(n3684)
         );
  AOI222_X1 U7590 ( .A1(n11254), .A2(n9837), .B1(n11251), .B2(n9773), .C1(
        n11248), .C2(n9805), .ZN(n3681) );
  NAND4_X1 U7591 ( .A1(n5073), .A2(n5074), .A3(n5075), .A4(n5076), .ZN(n5062)
         );
  AOI221_X1 U7592 ( .B1(n11014), .B2(n9966), .C1(n11011), .C2(n9998), .A(n5081), .ZN(n5075) );
  NOR4_X1 U7593 ( .A1(n5077), .A2(n5078), .A3(n5079), .A4(n5080), .ZN(n5076)
         );
  AOI222_X1 U7594 ( .A1(n10990), .A2(n9838), .B1(n10987), .B2(n9774), .C1(
        n10984), .C2(n9806), .ZN(n5073) );
  NAND4_X1 U7595 ( .A1(n3640), .A2(n3641), .A3(n3642), .A4(n3643), .ZN(n3629)
         );
  AOI221_X1 U7596 ( .B1(n11278), .B2(n9966), .C1(n11275), .C2(n9998), .A(n3648), .ZN(n3642) );
  NOR4_X1 U7597 ( .A1(n3644), .A2(n3645), .A3(n3646), .A4(n3647), .ZN(n3643)
         );
  AOI222_X1 U7598 ( .A1(n11254), .A2(n9838), .B1(n11251), .B2(n9774), .C1(
        n11248), .C2(n9806), .ZN(n3640) );
  NAND4_X1 U7599 ( .A1(n5032), .A2(n5033), .A3(n5034), .A4(n5035), .ZN(n5021)
         );
  AOI221_X1 U7600 ( .B1(n11014), .B2(n9967), .C1(n11011), .C2(n9999), .A(n5040), .ZN(n5034) );
  NOR4_X1 U7601 ( .A1(n5036), .A2(n5037), .A3(n5038), .A4(n5039), .ZN(n5035)
         );
  AOI222_X1 U7602 ( .A1(n10990), .A2(n9839), .B1(n10987), .B2(n9775), .C1(
        n10984), .C2(n9807), .ZN(n5032) );
  NAND4_X1 U7603 ( .A1(n3599), .A2(n3600), .A3(n3601), .A4(n3602), .ZN(n3588)
         );
  AOI221_X1 U7604 ( .B1(n11278), .B2(n9967), .C1(n11275), .C2(n9999), .A(n3607), .ZN(n3601) );
  NOR4_X1 U7605 ( .A1(n3603), .A2(n3604), .A3(n3605), .A4(n3606), .ZN(n3602)
         );
  AOI222_X1 U7606 ( .A1(n11254), .A2(n9839), .B1(n11251), .B2(n9775), .C1(
        n11248), .C2(n9807), .ZN(n3599) );
  NAND4_X1 U7607 ( .A1(n4991), .A2(n4992), .A3(n4993), .A4(n4994), .ZN(n4980)
         );
  AOI221_X1 U7608 ( .B1(n11014), .B2(n9968), .C1(n11011), .C2(n13059), .A(
        n4999), .ZN(n4993) );
  NOR4_X1 U7609 ( .A1(n4995), .A2(n4996), .A3(n4997), .A4(n4998), .ZN(n4994)
         );
  AOI222_X1 U7610 ( .A1(n10990), .A2(n9840), .B1(n10987), .B2(n9776), .C1(
        n10984), .C2(n9808), .ZN(n4991) );
  NAND4_X1 U7611 ( .A1(n3558), .A2(n3559), .A3(n3560), .A4(n3561), .ZN(n3547)
         );
  AOI221_X1 U7612 ( .B1(n11278), .B2(n9968), .C1(n11275), .C2(n13059), .A(
        n3566), .ZN(n3560) );
  NOR4_X1 U7613 ( .A1(n3562), .A2(n3563), .A3(n3564), .A4(n3565), .ZN(n3561)
         );
  AOI222_X1 U7614 ( .A1(n11254), .A2(n9840), .B1(n11251), .B2(n9776), .C1(
        n11248), .C2(n9808), .ZN(n3558) );
  NAND4_X1 U7615 ( .A1(n4950), .A2(n4951), .A3(n4952), .A4(n4953), .ZN(n4939)
         );
  AOI221_X1 U7616 ( .B1(n11014), .B2(n9969), .C1(n11011), .C2(n13058), .A(
        n4958), .ZN(n4952) );
  NOR4_X1 U7617 ( .A1(n4954), .A2(n4955), .A3(n4956), .A4(n4957), .ZN(n4953)
         );
  AOI222_X1 U7618 ( .A1(n10990), .A2(n9841), .B1(n10987), .B2(n9777), .C1(
        n10984), .C2(n9809), .ZN(n4950) );
  NAND4_X1 U7619 ( .A1(n3517), .A2(n3518), .A3(n3519), .A4(n3520), .ZN(n3506)
         );
  AOI221_X1 U7620 ( .B1(n11278), .B2(n9969), .C1(n11275), .C2(n13058), .A(
        n3525), .ZN(n3519) );
  NOR4_X1 U7621 ( .A1(n3521), .A2(n3522), .A3(n3523), .A4(n3524), .ZN(n3520)
         );
  AOI222_X1 U7622 ( .A1(n11254), .A2(n9841), .B1(n11251), .B2(n9777), .C1(
        n11248), .C2(n9809), .ZN(n3517) );
  NAND4_X1 U7623 ( .A1(n4909), .A2(n4910), .A3(n4911), .A4(n4912), .ZN(n4898)
         );
  AOI221_X1 U7624 ( .B1(n11014), .B2(n9970), .C1(n11011), .C2(n13057), .A(
        n4917), .ZN(n4911) );
  NOR4_X1 U7625 ( .A1(n4913), .A2(n4914), .A3(n4915), .A4(n4916), .ZN(n4912)
         );
  AOI222_X1 U7626 ( .A1(n10990), .A2(n9842), .B1(n10987), .B2(n9778), .C1(
        n10984), .C2(n9810), .ZN(n4909) );
  NAND4_X1 U7627 ( .A1(n3476), .A2(n3477), .A3(n3478), .A4(n3479), .ZN(n3465)
         );
  AOI221_X1 U7628 ( .B1(n11278), .B2(n9970), .C1(n11275), .C2(n13057), .A(
        n3484), .ZN(n3478) );
  NOR4_X1 U7629 ( .A1(n3480), .A2(n3481), .A3(n3482), .A4(n3483), .ZN(n3479)
         );
  AOI222_X1 U7630 ( .A1(n11254), .A2(n9842), .B1(n11251), .B2(n9778), .C1(
        n11248), .C2(n9810), .ZN(n3476) );
  NAND4_X1 U7631 ( .A1(n4868), .A2(n4869), .A3(n4870), .A4(n4871), .ZN(n4857)
         );
  AOI221_X1 U7632 ( .B1(n11014), .B2(n9971), .C1(n11011), .C2(n13056), .A(
        n4876), .ZN(n4870) );
  NOR4_X1 U7633 ( .A1(n4872), .A2(n4873), .A3(n4874), .A4(n4875), .ZN(n4871)
         );
  AOI222_X1 U7634 ( .A1(n10990), .A2(n9843), .B1(n10987), .B2(n9779), .C1(
        n10984), .C2(n9811), .ZN(n4868) );
  NAND4_X1 U7635 ( .A1(n3435), .A2(n3436), .A3(n3437), .A4(n3438), .ZN(n3424)
         );
  AOI221_X1 U7636 ( .B1(n11278), .B2(n9971), .C1(n11275), .C2(n13056), .A(
        n3443), .ZN(n3437) );
  NOR4_X1 U7637 ( .A1(n3439), .A2(n3440), .A3(n3441), .A4(n3442), .ZN(n3438)
         );
  AOI222_X1 U7638 ( .A1(n11254), .A2(n9843), .B1(n11251), .B2(n9779), .C1(
        n11248), .C2(n9811), .ZN(n3435) );
  NAND4_X1 U7639 ( .A1(n4827), .A2(n4828), .A3(n4829), .A4(n4830), .ZN(n4816)
         );
  AOI221_X1 U7640 ( .B1(n11014), .B2(n9972), .C1(n11011), .C2(n13055), .A(
        n4835), .ZN(n4829) );
  NOR4_X1 U7641 ( .A1(n4831), .A2(n4832), .A3(n4833), .A4(n4834), .ZN(n4830)
         );
  AOI222_X1 U7642 ( .A1(n10990), .A2(n9844), .B1(n10987), .B2(n9780), .C1(
        n10984), .C2(n9812), .ZN(n4827) );
  NAND4_X1 U7643 ( .A1(n3394), .A2(n3395), .A3(n3396), .A4(n3397), .ZN(n3383)
         );
  AOI221_X1 U7644 ( .B1(n11278), .B2(n9972), .C1(n11275), .C2(n13055), .A(
        n3402), .ZN(n3396) );
  NOR4_X1 U7645 ( .A1(n3398), .A2(n3399), .A3(n3400), .A4(n3401), .ZN(n3397)
         );
  AOI222_X1 U7646 ( .A1(n11254), .A2(n9844), .B1(n11251), .B2(n9780), .C1(
        n11248), .C2(n9812), .ZN(n3394) );
  NAND4_X1 U7647 ( .A1(n4786), .A2(n4787), .A3(n4788), .A4(n4789), .ZN(n4775)
         );
  AOI221_X1 U7648 ( .B1(n11014), .B2(n9973), .C1(n11011), .C2(n13054), .A(
        n4794), .ZN(n4788) );
  NOR4_X1 U7649 ( .A1(n4790), .A2(n4791), .A3(n4792), .A4(n4793), .ZN(n4789)
         );
  AOI222_X1 U7650 ( .A1(n10990), .A2(n9845), .B1(n10987), .B2(n9781), .C1(
        n10984), .C2(n9813), .ZN(n4786) );
  NAND4_X1 U7651 ( .A1(n3353), .A2(n3354), .A3(n3355), .A4(n3356), .ZN(n3342)
         );
  AOI221_X1 U7652 ( .B1(n11278), .B2(n9973), .C1(n11275), .C2(n13054), .A(
        n3361), .ZN(n3355) );
  NOR4_X1 U7653 ( .A1(n3357), .A2(n3358), .A3(n3359), .A4(n3360), .ZN(n3356)
         );
  AOI222_X1 U7654 ( .A1(n11254), .A2(n9845), .B1(n11251), .B2(n9781), .C1(
        n11248), .C2(n9813), .ZN(n3353) );
  NAND4_X1 U7655 ( .A1(n4745), .A2(n4746), .A3(n4747), .A4(n4748), .ZN(n4734)
         );
  AOI221_X1 U7656 ( .B1(n11014), .B2(n9974), .C1(n11011), .C2(n13053), .A(
        n4753), .ZN(n4747) );
  NOR4_X1 U7657 ( .A1(n4749), .A2(n4750), .A3(n4751), .A4(n4752), .ZN(n4748)
         );
  AOI222_X1 U7658 ( .A1(n10990), .A2(n9846), .B1(n10987), .B2(n9782), .C1(
        n10984), .C2(n9814), .ZN(n4745) );
  NAND4_X1 U7659 ( .A1(n3312), .A2(n3313), .A3(n3314), .A4(n3315), .ZN(n3301)
         );
  AOI221_X1 U7660 ( .B1(n11278), .B2(n9974), .C1(n11275), .C2(n13053), .A(
        n3320), .ZN(n3314) );
  NOR4_X1 U7661 ( .A1(n3316), .A2(n3317), .A3(n3318), .A4(n3319), .ZN(n3315)
         );
  AOI222_X1 U7662 ( .A1(n11254), .A2(n9846), .B1(n11251), .B2(n9782), .C1(
        n11248), .C2(n9814), .ZN(n3312) );
  NAND4_X1 U7663 ( .A1(n4704), .A2(n4705), .A3(n4706), .A4(n4707), .ZN(n4693)
         );
  AOI221_X1 U7664 ( .B1(n11014), .B2(n9975), .C1(n11011), .C2(n13052), .A(
        n4712), .ZN(n4706) );
  NOR4_X1 U7665 ( .A1(n4708), .A2(n4709), .A3(n4710), .A4(n4711), .ZN(n4707)
         );
  AOI222_X1 U7666 ( .A1(n10990), .A2(n9847), .B1(n10987), .B2(n9783), .C1(
        n10984), .C2(n9815), .ZN(n4704) );
  NAND4_X1 U7667 ( .A1(n3271), .A2(n3272), .A3(n3273), .A4(n3274), .ZN(n3260)
         );
  AOI221_X1 U7668 ( .B1(n11278), .B2(n9975), .C1(n11275), .C2(n13052), .A(
        n3279), .ZN(n3273) );
  NOR4_X1 U7669 ( .A1(n3275), .A2(n3276), .A3(n3277), .A4(n3278), .ZN(n3274)
         );
  AOI222_X1 U7670 ( .A1(n11254), .A2(n9847), .B1(n11251), .B2(n9783), .C1(
        n11248), .C2(n9815), .ZN(n3271) );
  NAND4_X1 U7671 ( .A1(n4663), .A2(n4664), .A3(n4665), .A4(n4666), .ZN(n4652)
         );
  AOI221_X1 U7672 ( .B1(n11015), .B2(n9976), .C1(n11012), .C2(n13051), .A(
        n4671), .ZN(n4665) );
  NOR4_X1 U7673 ( .A1(n4667), .A2(n4668), .A3(n4669), .A4(n4670), .ZN(n4666)
         );
  AOI222_X1 U7674 ( .A1(n10991), .A2(n9848), .B1(n10988), .B2(n9784), .C1(
        n10985), .C2(n9816), .ZN(n4663) );
  NAND4_X1 U7675 ( .A1(n3230), .A2(n3231), .A3(n3232), .A4(n3233), .ZN(n3219)
         );
  AOI221_X1 U7676 ( .B1(n11279), .B2(n9976), .C1(n11276), .C2(n13051), .A(
        n3238), .ZN(n3232) );
  NOR4_X1 U7677 ( .A1(n3234), .A2(n3235), .A3(n3236), .A4(n3237), .ZN(n3233)
         );
  AOI222_X1 U7678 ( .A1(n11255), .A2(n9848), .B1(n11252), .B2(n9784), .C1(
        n11249), .C2(n9816), .ZN(n3230) );
  NAND4_X1 U7679 ( .A1(n4622), .A2(n4623), .A3(n4624), .A4(n4625), .ZN(n4611)
         );
  AOI221_X1 U7680 ( .B1(n11015), .B2(n9977), .C1(n11012), .C2(n13050), .A(
        n4630), .ZN(n4624) );
  NOR4_X1 U7681 ( .A1(n4626), .A2(n4627), .A3(n4628), .A4(n4629), .ZN(n4625)
         );
  AOI222_X1 U7682 ( .A1(n10991), .A2(n9849), .B1(n10988), .B2(n9785), .C1(
        n10985), .C2(n9817), .ZN(n4622) );
  NAND4_X1 U7683 ( .A1(n3189), .A2(n3190), .A3(n3191), .A4(n3192), .ZN(n3178)
         );
  AOI221_X1 U7684 ( .B1(n11279), .B2(n9977), .C1(n11276), .C2(n13050), .A(
        n3197), .ZN(n3191) );
  NOR4_X1 U7685 ( .A1(n3193), .A2(n3194), .A3(n3195), .A4(n3196), .ZN(n3192)
         );
  AOI222_X1 U7686 ( .A1(n11255), .A2(n9849), .B1(n11252), .B2(n9785), .C1(
        n11249), .C2(n9817), .ZN(n3189) );
  NAND4_X1 U7687 ( .A1(n4581), .A2(n4582), .A3(n4583), .A4(n4584), .ZN(n4570)
         );
  AOI221_X1 U7688 ( .B1(n11015), .B2(n9978), .C1(n11012), .C2(n13049), .A(
        n4589), .ZN(n4583) );
  NOR4_X1 U7689 ( .A1(n4585), .A2(n4586), .A3(n4587), .A4(n4588), .ZN(n4584)
         );
  AOI222_X1 U7690 ( .A1(n10991), .A2(n9850), .B1(n10988), .B2(n9786), .C1(
        n10985), .C2(n9818), .ZN(n4581) );
  NAND4_X1 U7691 ( .A1(n3148), .A2(n3149), .A3(n3150), .A4(n3151), .ZN(n3137)
         );
  AOI221_X1 U7692 ( .B1(n11279), .B2(n9978), .C1(n11276), .C2(n13049), .A(
        n3156), .ZN(n3150) );
  NOR4_X1 U7693 ( .A1(n3152), .A2(n3153), .A3(n3154), .A4(n3155), .ZN(n3151)
         );
  AOI222_X1 U7694 ( .A1(n11255), .A2(n9850), .B1(n11252), .B2(n9786), .C1(
        n11249), .C2(n9818), .ZN(n3148) );
  NAND4_X1 U7695 ( .A1(n4540), .A2(n4541), .A3(n4542), .A4(n4543), .ZN(n4529)
         );
  AOI221_X1 U7696 ( .B1(n11015), .B2(n9979), .C1(n11012), .C2(n13048), .A(
        n4548), .ZN(n4542) );
  NOR4_X1 U7697 ( .A1(n4544), .A2(n4545), .A3(n4546), .A4(n4547), .ZN(n4543)
         );
  AOI222_X1 U7698 ( .A1(n10991), .A2(n9851), .B1(n10988), .B2(n9787), .C1(
        n10985), .C2(n9819), .ZN(n4540) );
  NAND4_X1 U7699 ( .A1(n3107), .A2(n3108), .A3(n3109), .A4(n3110), .ZN(n3096)
         );
  AOI221_X1 U7700 ( .B1(n11279), .B2(n9979), .C1(n11276), .C2(n13048), .A(
        n3115), .ZN(n3109) );
  NOR4_X1 U7701 ( .A1(n3111), .A2(n3112), .A3(n3113), .A4(n3114), .ZN(n3110)
         );
  AOI222_X1 U7702 ( .A1(n11255), .A2(n9851), .B1(n11252), .B2(n9787), .C1(
        n11249), .C2(n9819), .ZN(n3107) );
  NAND4_X1 U7703 ( .A1(n4499), .A2(n4500), .A3(n4501), .A4(n4502), .ZN(n4488)
         );
  AOI221_X1 U7704 ( .B1(n11015), .B2(n9980), .C1(n11012), .C2(n13047), .A(
        n4507), .ZN(n4501) );
  NOR4_X1 U7705 ( .A1(n4503), .A2(n4504), .A3(n4505), .A4(n4506), .ZN(n4502)
         );
  AOI222_X1 U7706 ( .A1(n10991), .A2(n9852), .B1(n10988), .B2(n9788), .C1(
        n10985), .C2(n9820), .ZN(n4499) );
  NAND4_X1 U7707 ( .A1(n3066), .A2(n3067), .A3(n3068), .A4(n3069), .ZN(n3055)
         );
  AOI221_X1 U7708 ( .B1(n11279), .B2(n9980), .C1(n11276), .C2(n13047), .A(
        n3074), .ZN(n3068) );
  NOR4_X1 U7709 ( .A1(n3070), .A2(n3071), .A3(n3072), .A4(n3073), .ZN(n3069)
         );
  AOI222_X1 U7710 ( .A1(n11255), .A2(n9852), .B1(n11252), .B2(n9788), .C1(
        n11249), .C2(n9820), .ZN(n3066) );
  NAND4_X1 U7711 ( .A1(n4458), .A2(n4459), .A3(n4460), .A4(n4461), .ZN(n4447)
         );
  AOI221_X1 U7712 ( .B1(n11015), .B2(n9981), .C1(n11012), .C2(n13046), .A(
        n4466), .ZN(n4460) );
  NOR4_X1 U7713 ( .A1(n4462), .A2(n4463), .A3(n4464), .A4(n4465), .ZN(n4461)
         );
  AOI222_X1 U7714 ( .A1(n10991), .A2(n9853), .B1(n10988), .B2(n9789), .C1(
        n10985), .C2(n9821), .ZN(n4458) );
  NAND4_X1 U7715 ( .A1(n3025), .A2(n3026), .A3(n3027), .A4(n3028), .ZN(n3014)
         );
  AOI221_X1 U7716 ( .B1(n11279), .B2(n9981), .C1(n11276), .C2(n13046), .A(
        n3033), .ZN(n3027) );
  NOR4_X1 U7717 ( .A1(n3029), .A2(n3030), .A3(n3031), .A4(n3032), .ZN(n3028)
         );
  AOI222_X1 U7718 ( .A1(n11255), .A2(n9853), .B1(n11252), .B2(n9789), .C1(
        n11249), .C2(n9821), .ZN(n3025) );
  NAND4_X1 U7719 ( .A1(n4417), .A2(n4418), .A3(n4419), .A4(n4420), .ZN(n4406)
         );
  AOI221_X1 U7720 ( .B1(n11015), .B2(n9982), .C1(n11012), .C2(n13045), .A(
        n4425), .ZN(n4419) );
  NOR4_X1 U7721 ( .A1(n4421), .A2(n4422), .A3(n4423), .A4(n4424), .ZN(n4420)
         );
  AOI222_X1 U7722 ( .A1(n10991), .A2(n9854), .B1(n10988), .B2(n9790), .C1(
        n10985), .C2(n9822), .ZN(n4417) );
  NAND4_X1 U7723 ( .A1(n2984), .A2(n2985), .A3(n2986), .A4(n2987), .ZN(n2973)
         );
  AOI221_X1 U7724 ( .B1(n11279), .B2(n9982), .C1(n11276), .C2(n13045), .A(
        n2992), .ZN(n2986) );
  NOR4_X1 U7725 ( .A1(n2988), .A2(n2989), .A3(n2990), .A4(n2991), .ZN(n2987)
         );
  AOI222_X1 U7726 ( .A1(n11255), .A2(n9854), .B1(n11252), .B2(n9790), .C1(
        n11249), .C2(n9822), .ZN(n2984) );
  NAND4_X1 U7727 ( .A1(n4310), .A2(n4311), .A3(n4312), .A4(n4313), .ZN(n4277)
         );
  AOI221_X1 U7728 ( .B1(n11015), .B2(n9983), .C1(n11012), .C2(n13044), .A(
        n4331), .ZN(n4312) );
  NOR4_X1 U7729 ( .A1(n4314), .A2(n4315), .A3(n4316), .A4(n4317), .ZN(n4313)
         );
  AOI222_X1 U7730 ( .A1(n10991), .A2(n9855), .B1(n10988), .B2(n9791), .C1(
        n10985), .C2(n9823), .ZN(n4310) );
  NAND4_X1 U7731 ( .A1(n2810), .A2(n2811), .A3(n2812), .A4(n2813), .ZN(n2745)
         );
  AOI221_X1 U7732 ( .B1(n11279), .B2(n9983), .C1(n11276), .C2(n13044), .A(
        n2863), .ZN(n2812) );
  NOR4_X1 U7733 ( .A1(n2814), .A2(n2815), .A3(n2816), .A4(n2817), .ZN(n2813)
         );
  AOI222_X1 U7734 ( .A1(n11255), .A2(n9855), .B1(n11252), .B2(n9791), .C1(
        n11249), .C2(n9823), .ZN(n2810) );
  NAND2_X1 U7735 ( .A1(n2937), .A2(n2740), .ZN(\U3/U98/Z_4 ) );
  NAND2_X1 U7736 ( .A1(n2937), .A2(n2739), .ZN(\U3/U99/Z_4 ) );
  NAND2_X1 U7737 ( .A1(n2937), .A2(n2741), .ZN(\U3/U97/Z_4 ) );
  NAND2_X1 U7738 ( .A1(n2936), .A2(n2740), .ZN(\U3/U98/Z_5 ) );
  NAND2_X1 U7739 ( .A1(n2936), .A2(n2739), .ZN(\U3/U99/Z_5 ) );
  NAND2_X1 U7740 ( .A1(n2936), .A2(n2741), .ZN(\U3/U97/Z_5 ) );
  INV_X1 U7741 ( .A(DATAIN[0]), .ZN(n12768) );
  INV_X1 U7742 ( .A(DATAIN[1]), .ZN(n12767) );
  INV_X1 U7743 ( .A(DATAIN[2]), .ZN(n12766) );
  INV_X1 U7744 ( .A(DATAIN[3]), .ZN(n12765) );
  INV_X1 U7745 ( .A(DATAIN[4]), .ZN(n12764) );
  INV_X1 U7746 ( .A(DATAIN[5]), .ZN(n12763) );
  INV_X1 U7747 ( .A(DATAIN[6]), .ZN(n12762) );
  INV_X1 U7748 ( .A(DATAIN[7]), .ZN(n12761) );
  INV_X1 U7749 ( .A(DATAIN[8]), .ZN(n12760) );
  INV_X1 U7750 ( .A(DATAIN[9]), .ZN(n12759) );
  INV_X1 U7751 ( .A(DATAIN[10]), .ZN(n12758) );
  INV_X1 U7752 ( .A(DATAIN[11]), .ZN(n12757) );
  INV_X1 U7753 ( .A(DATAIN[12]), .ZN(n12756) );
  INV_X1 U7754 ( .A(DATAIN[13]), .ZN(n12755) );
  INV_X1 U7755 ( .A(DATAIN[14]), .ZN(n12754) );
  INV_X1 U7756 ( .A(DATAIN[15]), .ZN(n12753) );
  INV_X1 U7757 ( .A(DATAIN[16]), .ZN(n12752) );
  INV_X1 U7758 ( .A(DATAIN[17]), .ZN(n12751) );
  INV_X1 U7759 ( .A(DATAIN[18]), .ZN(n12750) );
  INV_X1 U7760 ( .A(DATAIN[19]), .ZN(n12749) );
  INV_X1 U7761 ( .A(DATAIN[20]), .ZN(n12748) );
  INV_X1 U7762 ( .A(DATAIN[21]), .ZN(n12747) );
  INV_X1 U7763 ( .A(DATAIN[22]), .ZN(n12746) );
  INV_X1 U7764 ( .A(DATAIN[23]), .ZN(n12745) );
  INV_X1 U7765 ( .A(DATAIN[24]), .ZN(n12744) );
  INV_X1 U7766 ( .A(DATAIN[25]), .ZN(n12743) );
  INV_X1 U7767 ( .A(DATAIN[26]), .ZN(n12742) );
  INV_X1 U7768 ( .A(DATAIN[27]), .ZN(n12741) );
  INV_X1 U7769 ( .A(DATAIN[28]), .ZN(n12740) );
  INV_X1 U7770 ( .A(DATAIN[29]), .ZN(n12739) );
  INV_X1 U7771 ( .A(DATAIN[30]), .ZN(n12738) );
  INV_X1 U7772 ( .A(DATAIN[31]), .ZN(n12737) );
  NAND2_X1 U7773 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n2740) );
  NAND2_X1 U7774 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n2739) );
  NAND2_X1 U7775 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .ZN(n2741) );
  INV_X1 U7776 ( .A(N8431), .ZN(n14514) );
  INV_X1 U7777 ( .A(N8575), .ZN(n14516) );
  INV_X1 U7778 ( .A(N8432), .ZN(n14513) );
  INV_X1 U7779 ( .A(N8576), .ZN(n14515) );
  AND2_X1 U7780 ( .A1(N2170), .A2(N2169), .ZN(n2716) );
  INV_X1 U7781 ( .A(N2167), .ZN(n12736) );
  INV_X1 U7782 ( .A(N2168), .ZN(n12735) );
  INV_X1 U7783 ( .A(N2169), .ZN(n12734) );
  OR2_X1 U7784 ( .A1(RD1), .A2(n12712), .ZN(N8702) );
  OR2_X1 U7785 ( .A1(RD2), .A2(n12712), .ZN(N8735) );
  INV_X1 U7786 ( .A(n11390), .ZN(n11381) );
  INV_X1 U7787 ( .A(n11402), .ZN(n11393) );
  INV_X1 U7788 ( .A(n11414), .ZN(n11405) );
  INV_X1 U7789 ( .A(n11426), .ZN(n11417) );
  INV_X1 U7790 ( .A(n11438), .ZN(n11429) );
  INV_X1 U7791 ( .A(n11450), .ZN(n11441) );
  INV_X1 U7792 ( .A(n11462), .ZN(n11453) );
  INV_X1 U7793 ( .A(n11474), .ZN(n11465) );
  INV_X1 U7794 ( .A(n11486), .ZN(n11477) );
  INV_X1 U7795 ( .A(n11498), .ZN(n11489) );
  INV_X1 U7796 ( .A(n11510), .ZN(n11501) );
  INV_X1 U7797 ( .A(n11522), .ZN(n11513) );
  INV_X1 U7798 ( .A(n11534), .ZN(n11525) );
  INV_X1 U7799 ( .A(n11546), .ZN(n11537) );
  INV_X1 U7800 ( .A(n11558), .ZN(n11549) );
  INV_X1 U7801 ( .A(n11570), .ZN(n11561) );
  INV_X1 U7802 ( .A(n11582), .ZN(n11573) );
  INV_X1 U7803 ( .A(n11594), .ZN(n11585) );
  INV_X1 U7804 ( .A(n11606), .ZN(n11597) );
  INV_X1 U7805 ( .A(n11618), .ZN(n11609) );
  INV_X1 U7806 ( .A(n11630), .ZN(n11621) );
  INV_X1 U7807 ( .A(n11642), .ZN(n11633) );
  INV_X1 U7808 ( .A(n11654), .ZN(n11645) );
  INV_X1 U7809 ( .A(n11666), .ZN(n11657) );
  INV_X1 U7810 ( .A(n11678), .ZN(n11669) );
  INV_X1 U7811 ( .A(n11690), .ZN(n11681) );
  INV_X1 U7812 ( .A(n11702), .ZN(n11693) );
  INV_X1 U7813 ( .A(n11714), .ZN(n11705) );
  INV_X1 U7814 ( .A(n11726), .ZN(n11717) );
  INV_X1 U7815 ( .A(n11738), .ZN(n11729) );
  INV_X1 U7816 ( .A(n11750), .ZN(n11741) );
  INV_X1 U7817 ( .A(n11762), .ZN(n11753) );
  INV_X1 U7818 ( .A(n11774), .ZN(n11765) );
  INV_X1 U7819 ( .A(n11786), .ZN(n11777) );
  INV_X1 U7820 ( .A(n11798), .ZN(n11789) );
  INV_X1 U7821 ( .A(n11810), .ZN(n11801) );
  INV_X1 U7822 ( .A(n11822), .ZN(n11813) );
  INV_X1 U7823 ( .A(n11834), .ZN(n11825) );
  INV_X1 U7824 ( .A(n11846), .ZN(n11837) );
  INV_X1 U7825 ( .A(n11858), .ZN(n11849) );
  INV_X1 U7826 ( .A(n11870), .ZN(n11861) );
  INV_X1 U7827 ( .A(n11882), .ZN(n11873) );
  INV_X1 U7828 ( .A(n11894), .ZN(n11885) );
  INV_X1 U7829 ( .A(n11906), .ZN(n11897) );
  INV_X1 U7830 ( .A(n11918), .ZN(n11909) );
  INV_X1 U7831 ( .A(n11930), .ZN(n11921) );
  INV_X1 U7832 ( .A(n11942), .ZN(n11933) );
  INV_X1 U7833 ( .A(n11954), .ZN(n11945) );
  INV_X1 U7834 ( .A(n11966), .ZN(n11957) );
  INV_X1 U7839 ( .A(n11978), .ZN(n11969) );
  INV_X1 U7840 ( .A(n11990), .ZN(n11981) );
  INV_X1 U7841 ( .A(n12002), .ZN(n11993) );
  INV_X1 U7842 ( .A(n12014), .ZN(n12005) );
  INV_X1 U7843 ( .A(n12026), .ZN(n12017) );
  INV_X1 U7844 ( .A(n12038), .ZN(n12029) );
  INV_X1 U7845 ( .A(n12050), .ZN(n12041) );
  INV_X1 U7846 ( .A(n12062), .ZN(n12053) );
  INV_X1 U7847 ( .A(n12074), .ZN(n12065) );
  INV_X1 U7848 ( .A(n12086), .ZN(n12077) );
  INV_X1 U7849 ( .A(n12098), .ZN(n12089) );
  INV_X1 U7850 ( .A(n12110), .ZN(n12101) );
  INV_X1 U7851 ( .A(n12122), .ZN(n12113) );
  INV_X1 U7852 ( .A(n12134), .ZN(n12125) );
  INV_X1 U7853 ( .A(n12146), .ZN(n12137) );
  INV_X1 U7854 ( .A(n12158), .ZN(n12149) );
  INV_X1 U7855 ( .A(n12170), .ZN(n12161) );
  INV_X1 U7856 ( .A(n12182), .ZN(n12173) );
  INV_X1 U7857 ( .A(n12194), .ZN(n12185) );
  INV_X1 U7858 ( .A(n12206), .ZN(n12197) );
  INV_X1 U7859 ( .A(n12218), .ZN(n12209) );
  INV_X1 U7860 ( .A(n12230), .ZN(n12221) );
  INV_X1 U7861 ( .A(n12242), .ZN(n12233) );
  INV_X1 U7862 ( .A(n12254), .ZN(n12245) );
  INV_X1 U7863 ( .A(n12266), .ZN(n12257) );
  INV_X1 U7864 ( .A(n12278), .ZN(n12269) );
  INV_X1 U7865 ( .A(n12290), .ZN(n12281) );
  INV_X1 U7866 ( .A(n12302), .ZN(n12293) );
  INV_X1 U7867 ( .A(n12314), .ZN(n12305) );
  INV_X1 U7868 ( .A(n12326), .ZN(n12317) );
  INV_X1 U7869 ( .A(n12338), .ZN(n12329) );
  INV_X1 U7870 ( .A(n12425), .ZN(n12418) );
  INV_X1 U7871 ( .A(n12691), .ZN(n12433) );
  INV_X1 U7872 ( .A(n12691), .ZN(n12434) );
  INV_X1 U7873 ( .A(n12690), .ZN(n12435) );
  INV_X1 U7874 ( .A(n12690), .ZN(n12436) );
  INV_X1 U7875 ( .A(n12690), .ZN(n12437) );
  INV_X1 U7876 ( .A(n12690), .ZN(n12438) );
  INV_X1 U7877 ( .A(n12690), .ZN(n12439) );
  INV_X1 U7878 ( .A(n12690), .ZN(n12440) );
  INV_X1 U7879 ( .A(n12690), .ZN(n12441) );
  INV_X1 U7880 ( .A(n12689), .ZN(n12442) );
  INV_X1 U7881 ( .A(n12689), .ZN(n12443) );
  INV_X1 U7882 ( .A(n12689), .ZN(n12444) );
  INV_X1 U7883 ( .A(n12689), .ZN(n12445) );
  INV_X1 U7884 ( .A(n12689), .ZN(n12446) );
  INV_X1 U7885 ( .A(n12689), .ZN(n12447) );
  INV_X1 U7886 ( .A(n12689), .ZN(n12448) );
  INV_X1 U7887 ( .A(n12688), .ZN(n12449) );
  INV_X1 U7888 ( .A(n12688), .ZN(n12450) );
  INV_X1 U7889 ( .A(n12688), .ZN(n12451) );
  INV_X1 U7890 ( .A(n12688), .ZN(n12452) );
  INV_X1 U7891 ( .A(n12688), .ZN(n12453) );
  INV_X1 U7892 ( .A(n12688), .ZN(n12454) );
  INV_X1 U7893 ( .A(n12687), .ZN(n12455) );
  INV_X1 U7894 ( .A(n12687), .ZN(n12456) );
  INV_X1 U7895 ( .A(n12687), .ZN(n12457) );
  INV_X1 U7896 ( .A(n12687), .ZN(n12458) );
  INV_X1 U7897 ( .A(n12687), .ZN(n12459) );
  INV_X1 U7898 ( .A(n12687), .ZN(n12460) );
  INV_X1 U7899 ( .A(n12687), .ZN(n12461) );
  INV_X1 U7900 ( .A(n12686), .ZN(n12462) );
  INV_X1 U7901 ( .A(n12686), .ZN(n12463) );
  INV_X1 U7902 ( .A(n12686), .ZN(n12464) );
  INV_X1 U7903 ( .A(n12686), .ZN(n12465) );
  INV_X1 U7904 ( .A(n12686), .ZN(n12466) );
  INV_X1 U7905 ( .A(n12686), .ZN(n12467) );
  INV_X1 U7906 ( .A(n12686), .ZN(n12468) );
  INV_X1 U7907 ( .A(n12685), .ZN(n12469) );
  INV_X1 U7908 ( .A(n12685), .ZN(n12470) );
  INV_X1 U7909 ( .A(n12685), .ZN(n12471) );
  INV_X1 U7910 ( .A(n12685), .ZN(n12472) );
  INV_X1 U7911 ( .A(n12685), .ZN(n12473) );
  INV_X1 U7912 ( .A(n12685), .ZN(n12474) );
  INV_X1 U7913 ( .A(n12684), .ZN(n12475) );
  INV_X1 U7914 ( .A(n12684), .ZN(n12476) );
  INV_X1 U7915 ( .A(n12684), .ZN(n12477) );
  INV_X1 U7916 ( .A(n12684), .ZN(n12478) );
  INV_X1 U7917 ( .A(n12684), .ZN(n12479) );
  INV_X1 U7918 ( .A(n12684), .ZN(n12480) );
  INV_X1 U7919 ( .A(n12684), .ZN(n12481) );
  INV_X1 U7920 ( .A(n12683), .ZN(n12482) );
  INV_X1 U7921 ( .A(n12683), .ZN(n12483) );
  INV_X1 U7922 ( .A(n12683), .ZN(n12484) );
  INV_X1 U7923 ( .A(n12683), .ZN(n12485) );
  INV_X1 U7924 ( .A(n12683), .ZN(n12486) );
  INV_X1 U7925 ( .A(n12683), .ZN(n12487) );
  INV_X1 U7926 ( .A(n12683), .ZN(n12488) );
  INV_X1 U7927 ( .A(n12682), .ZN(n12489) );
  INV_X1 U7928 ( .A(n12682), .ZN(n12490) );
  INV_X1 U7929 ( .A(n12682), .ZN(n12491) );
  INV_X1 U7930 ( .A(n12682), .ZN(n12492) );
  INV_X1 U7931 ( .A(n12682), .ZN(n12493) );
  INV_X1 U7932 ( .A(n12682), .ZN(n12494) );
  INV_X1 U7933 ( .A(n12682), .ZN(n12495) );
  INV_X1 U7934 ( .A(n12681), .ZN(n12496) );
  INV_X1 U7935 ( .A(n12681), .ZN(n12497) );
  INV_X1 U7936 ( .A(n12681), .ZN(n12498) );
  INV_X1 U7937 ( .A(n12681), .ZN(n12499) );
  INV_X1 U7938 ( .A(n12681), .ZN(n12500) );
  INV_X1 U7939 ( .A(n12681), .ZN(n12501) );
  INV_X1 U7940 ( .A(n12681), .ZN(n12502) );
  INV_X1 U7941 ( .A(n12680), .ZN(n12503) );
  INV_X1 U7942 ( .A(n12680), .ZN(n12504) );
  INV_X1 U7943 ( .A(n12680), .ZN(n12505) );
  INV_X1 U7944 ( .A(n12680), .ZN(n12506) );
  INV_X1 U7945 ( .A(n12680), .ZN(n12507) );
  INV_X1 U7946 ( .A(n12680), .ZN(n12508) );
  INV_X1 U7947 ( .A(n12680), .ZN(n12509) );
  INV_X1 U7948 ( .A(n12679), .ZN(n12510) );
  INV_X1 U7949 ( .A(n12679), .ZN(n12511) );
  INV_X1 U7950 ( .A(n12679), .ZN(n12512) );
  INV_X1 U7951 ( .A(n12679), .ZN(n12513) );
  INV_X1 U7952 ( .A(n12679), .ZN(n12514) );
  INV_X1 U7953 ( .A(n12679), .ZN(n12515) );
  INV_X1 U7954 ( .A(n12685), .ZN(n12516) );
  INV_X1 U7955 ( .A(n12711), .ZN(n12517) );
  INV_X1 U7956 ( .A(n12711), .ZN(n12518) );
  INV_X1 U7957 ( .A(n12711), .ZN(n12519) );
  INV_X1 U7958 ( .A(n12711), .ZN(n12520) );
  INV_X1 U7959 ( .A(n12711), .ZN(n12521) );
  INV_X1 U7960 ( .A(n12711), .ZN(n12522) );
  INV_X1 U7961 ( .A(n12710), .ZN(n12523) );
  INV_X1 U7962 ( .A(n12711), .ZN(n12524) );
  INV_X1 U7963 ( .A(n12710), .ZN(n12525) );
  INV_X1 U7964 ( .A(n12710), .ZN(n12526) );
  INV_X1 U7965 ( .A(n12710), .ZN(n12527) );
  INV_X1 U7966 ( .A(n12710), .ZN(n12528) );
  INV_X1 U7967 ( .A(n12710), .ZN(n12529) );
  INV_X1 U7968 ( .A(n12710), .ZN(n12530) );
  INV_X1 U7969 ( .A(n12709), .ZN(n12531) );
  INV_X1 U7970 ( .A(n12709), .ZN(n12532) );
  INV_X1 U7971 ( .A(n12709), .ZN(n12533) );
  INV_X1 U7972 ( .A(n12709), .ZN(n12534) );
  INV_X1 U7973 ( .A(n12709), .ZN(n12535) );
  INV_X1 U7974 ( .A(n12709), .ZN(n12536) );
  INV_X1 U7975 ( .A(n12708), .ZN(n12537) );
  INV_X1 U7976 ( .A(n12709), .ZN(n12538) );
  INV_X1 U7977 ( .A(n12708), .ZN(n12539) );
  INV_X1 U7978 ( .A(n12708), .ZN(n12540) );
  INV_X1 U7979 ( .A(n12708), .ZN(n12541) );
  INV_X1 U7980 ( .A(n12708), .ZN(n12542) );
  INV_X1 U7981 ( .A(n12708), .ZN(n12543) );
  INV_X1 U7982 ( .A(n12708), .ZN(n12544) );
  INV_X1 U7983 ( .A(n12707), .ZN(n12545) );
  INV_X1 U7984 ( .A(n12707), .ZN(n12546) );
  INV_X1 U7985 ( .A(n12707), .ZN(n12547) );
  INV_X1 U7986 ( .A(n12707), .ZN(n12548) );
  INV_X1 U7987 ( .A(n12707), .ZN(n12549) );
  INV_X1 U7988 ( .A(n12707), .ZN(n12550) );
  INV_X1 U7989 ( .A(n12707), .ZN(n12551) );
  INV_X1 U7990 ( .A(n12706), .ZN(n12552) );
  INV_X1 U7991 ( .A(n12706), .ZN(n12553) );
  INV_X1 U7992 ( .A(n12706), .ZN(n12554) );
  INV_X1 U7993 ( .A(n12706), .ZN(n12555) );
  INV_X1 U7994 ( .A(n12706), .ZN(n12556) );
  INV_X1 U7995 ( .A(n12706), .ZN(n12557) );
  INV_X1 U7996 ( .A(n12706), .ZN(n12558) );
  INV_X1 U7997 ( .A(n12705), .ZN(n12559) );
  INV_X1 U7998 ( .A(n12705), .ZN(n12560) );
  INV_X1 U7999 ( .A(n12705), .ZN(n12561) );
  INV_X1 U8000 ( .A(n12705), .ZN(n12562) );
  INV_X1 U8001 ( .A(n12705), .ZN(n12563) );
  INV_X1 U8002 ( .A(n12705), .ZN(n12564) );
  INV_X1 U8003 ( .A(n12705), .ZN(n12565) );
  INV_X1 U8004 ( .A(n12704), .ZN(n12566) );
  INV_X1 U8005 ( .A(n12704), .ZN(n12567) );
  INV_X1 U8006 ( .A(n12704), .ZN(n12568) );
  INV_X1 U8007 ( .A(n12704), .ZN(n12569) );
  INV_X1 U8008 ( .A(n12704), .ZN(n12570) );
  INV_X1 U8009 ( .A(n12704), .ZN(n12571) );
  INV_X1 U8010 ( .A(n12704), .ZN(n12572) );
  INV_X1 U8011 ( .A(n12703), .ZN(n12573) );
  INV_X1 U8012 ( .A(n12703), .ZN(n12574) );
  INV_X1 U8013 ( .A(n12703), .ZN(n12575) );
  INV_X1 U8014 ( .A(n12703), .ZN(n12576) );
  INV_X1 U8015 ( .A(n12703), .ZN(n12577) );
  INV_X1 U8016 ( .A(n12703), .ZN(n12578) );
  INV_X1 U8017 ( .A(n12703), .ZN(n12579) );
  INV_X1 U8018 ( .A(n12702), .ZN(n12580) );
  INV_X1 U8019 ( .A(n12702), .ZN(n12581) );
  INV_X1 U8020 ( .A(n12702), .ZN(n12582) );
  INV_X1 U8021 ( .A(n12702), .ZN(n12583) );
  INV_X1 U8022 ( .A(n12702), .ZN(n12584) );
  INV_X1 U8023 ( .A(n12702), .ZN(n12585) );
  INV_X1 U8024 ( .A(n12702), .ZN(n12586) );
  INV_X1 U8025 ( .A(n12701), .ZN(n12587) );
  INV_X1 U8026 ( .A(n12701), .ZN(n12588) );
  INV_X1 U8027 ( .A(n12701), .ZN(n12589) );
  INV_X1 U8028 ( .A(n12701), .ZN(n12590) );
  INV_X1 U8029 ( .A(n12701), .ZN(n12591) );
  INV_X1 U8030 ( .A(n12701), .ZN(n12592) );
  INV_X1 U8031 ( .A(n12700), .ZN(n12593) );
  INV_X1 U8032 ( .A(n12700), .ZN(n12594) );
  INV_X1 U8033 ( .A(n12700), .ZN(n12595) );
  INV_X1 U8034 ( .A(n12700), .ZN(n12596) );
  INV_X1 U8035 ( .A(n12700), .ZN(n12597) );
  INV_X1 U8036 ( .A(n12700), .ZN(n12598) );
  INV_X1 U8037 ( .A(n12700), .ZN(n12599) );
  INV_X1 U8038 ( .A(n12699), .ZN(n12600) );
  INV_X1 U8039 ( .A(n12699), .ZN(n12601) );
  INV_X1 U8040 ( .A(n12699), .ZN(n12602) );
  INV_X1 U8041 ( .A(n12699), .ZN(n12603) );
  INV_X1 U8042 ( .A(n12699), .ZN(n12604) );
  INV_X1 U8043 ( .A(n12699), .ZN(n12605) );
  INV_X1 U8044 ( .A(n12699), .ZN(n12606) );
  INV_X1 U8045 ( .A(n12698), .ZN(n12607) );
  INV_X1 U8046 ( .A(n12698), .ZN(n12608) );
  INV_X1 U8047 ( .A(n12698), .ZN(n12609) );
  INV_X1 U8048 ( .A(n12698), .ZN(n12610) );
  INV_X1 U8049 ( .A(n12698), .ZN(n12611) );
  INV_X1 U8050 ( .A(n12698), .ZN(n12612) );
  INV_X1 U8051 ( .A(n12698), .ZN(n12613) );
  INV_X1 U8052 ( .A(n12697), .ZN(n12614) );
  INV_X1 U8053 ( .A(n12697), .ZN(n12615) );
  INV_X1 U8054 ( .A(n12697), .ZN(n12616) );
  INV_X1 U8055 ( .A(n12697), .ZN(n12617) );
  INV_X1 U8056 ( .A(n12697), .ZN(n12618) );
  INV_X1 U8057 ( .A(n12697), .ZN(n12619) );
  INV_X1 U8058 ( .A(n12697), .ZN(n12620) );
  INV_X1 U8059 ( .A(n12696), .ZN(n12621) );
  INV_X1 U8060 ( .A(n12696), .ZN(n12622) );
  INV_X1 U8061 ( .A(n12696), .ZN(n12623) );
  INV_X1 U8062 ( .A(n12696), .ZN(n12624) );
  INV_X1 U8063 ( .A(n12696), .ZN(n12625) );
  INV_X1 U8064 ( .A(n12696), .ZN(n12626) );
  INV_X1 U8065 ( .A(n12696), .ZN(n12627) );
  INV_X1 U8066 ( .A(n12695), .ZN(n12628) );
  INV_X1 U8067 ( .A(n12695), .ZN(n12629) );
  INV_X1 U8068 ( .A(n12695), .ZN(n12630) );
  INV_X1 U8069 ( .A(n12695), .ZN(n12631) );
  INV_X1 U8070 ( .A(n12695), .ZN(n12632) );
  INV_X1 U8071 ( .A(n12695), .ZN(n12633) );
  INV_X1 U8072 ( .A(n12695), .ZN(n12634) );
  INV_X1 U8073 ( .A(n12694), .ZN(n12635) );
  INV_X1 U8074 ( .A(n12694), .ZN(n12636) );
  INV_X1 U8075 ( .A(n12694), .ZN(n12637) );
  INV_X1 U8076 ( .A(n12694), .ZN(n12638) );
  INV_X1 U8077 ( .A(n12694), .ZN(n12639) );
  INV_X1 U8078 ( .A(n12694), .ZN(n12640) );
  INV_X1 U8079 ( .A(n12694), .ZN(n12641) );
  INV_X1 U8080 ( .A(n12693), .ZN(n12642) );
  INV_X1 U8081 ( .A(n12693), .ZN(n12643) );
  INV_X1 U8082 ( .A(n12693), .ZN(n12644) );
  INV_X1 U8083 ( .A(n12693), .ZN(n12645) );
  INV_X1 U8084 ( .A(n12693), .ZN(n12646) );
  INV_X1 U8085 ( .A(n12693), .ZN(n12647) );
  INV_X1 U8086 ( .A(n12693), .ZN(n12648) );
  INV_X1 U8087 ( .A(n12692), .ZN(n12649) );
  INV_X1 U8088 ( .A(n12692), .ZN(n12650) );
  INV_X1 U8089 ( .A(n12692), .ZN(n12651) );
  INV_X1 U8090 ( .A(n12692), .ZN(n12652) );
  INV_X1 U8091 ( .A(n12692), .ZN(n12653) );
  INV_X1 U8092 ( .A(n12692), .ZN(n12654) );
  INV_X1 U8093 ( .A(n12692), .ZN(n12655) );
  INV_X1 U8094 ( .A(n12691), .ZN(n12656) );
  INV_X1 U8095 ( .A(n12691), .ZN(n12657) );
  INV_X1 U8096 ( .A(n12691), .ZN(n12658) );
  INV_X1 U8097 ( .A(n12691), .ZN(n12659) );
  INV_X1 U8098 ( .A(n12701), .ZN(n12660) );
  INV_X1 U8099 ( .A(n12679), .ZN(n12661) );
  INV_X1 U8100 ( .A(n12691), .ZN(n12662) );
  AND2_X1 U8101 ( .A1(\r480/A[3] ), .A2(ADD_RD1[3]), .ZN(\r480/carry[4] ) );
  XOR2_X1 U8102 ( .A(ADD_RD1[3]), .B(\r480/A[3] ), .Z(N8434) );
  AND2_X1 U8103 ( .A1(\r486/A[3] ), .A2(ADD_RD2[3]), .ZN(\r486/carry[4] ) );
  XOR2_X1 U8104 ( .A(ADD_RD2[3]), .B(\r486/A[3] ), .Z(N8578) );
  AND2_X1 U8105 ( .A1(ADD_WR[3]), .A2(\r472/B[3] ), .ZN(\r472/carry[4] ) );
  XOR2_X1 U8106 ( .A(\r472/B[3] ), .B(ADD_WR[3]), .Z(N2170) );
endmodule


module FF_0 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n2, n4, n3, n5;

  DFF_X1 Q_reg ( .D(n2), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n4), .A2(n3), .ZN(n2) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n5), .B2(Q), .ZN(n4) );
  INV_X1 U5 ( .A(EN), .ZN(n5) );
  INV_X1 U6 ( .A(RESET), .ZN(n3) );
endmodule


module regFFD_NBIT32_11 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U7 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U8 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U9 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U10 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U11 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U12 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U13 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U14 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U15 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U16 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U17 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U18 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U19 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U20 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U21 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U22 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U23 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U24 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U25 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U26 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U27 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U28 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U29 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U30 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U31 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U32 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U33 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U34 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U35 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U36 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U37 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U38 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U39 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U40 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U41 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U42 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U43 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U44 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U45 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U46 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U47 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U48 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U49 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U50 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U51 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U52 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module regFFD_NBIT32_10 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n65) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n66) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n67) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n68) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n98), .Q(Q[27]), .QN(n69) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n98), .Q(Q[26]), .QN(n70) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n98), .Q(Q[25]), .QN(n71) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n98), .Q(Q[24]), .QN(n72) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n99), .Q(Q[23]), .QN(n73) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n74) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n75) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n97), .Q(Q[20]), .QN(n76) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n99), .Q(Q[19]), .QN(n77) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n97), .Q(Q[18]), .QN(n78) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n97), .Q(Q[17]), .QN(n79) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n97), .Q(Q[16]), .QN(n80) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n99), .Q(Q[15]), .QN(n81) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n97), .Q(Q[14]), .QN(n82) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n97), .Q(Q[13]), .QN(n83) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n97), .Q(Q[12]), .QN(n84) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n85) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n86) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n98), .Q(Q[9]), .QN(n87) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n98), .Q(Q[8]), .QN(n88) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n89) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n90) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n91) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n92) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n98), .Q(Q[3]), .QN(n93) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n94) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n95) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n96) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n96), .B2(ENABLE), .A(n39), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n39) );
  OAI21_X1 U7 ( .B1(n95), .B2(ENABLE), .A(n40), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n40) );
  OAI21_X1 U9 ( .B1(n94), .B2(ENABLE), .A(n41), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n41) );
  OAI21_X1 U11 ( .B1(n93), .B2(ENABLE), .A(n43), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n43) );
  OAI21_X1 U13 ( .B1(n92), .B2(ENABLE), .A(n44), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n91), .B2(ENABLE), .A(n45), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n45) );
  OAI21_X1 U17 ( .B1(n90), .B2(ENABLE), .A(n46), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n46) );
  OAI21_X1 U19 ( .B1(n89), .B2(ENABLE), .A(n47), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n47) );
  OAI21_X1 U21 ( .B1(n88), .B2(ENABLE), .A(n48), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n48) );
  OAI21_X1 U23 ( .B1(n87), .B2(ENABLE), .A(n49), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n49) );
  OAI21_X1 U25 ( .B1(n86), .B2(ENABLE), .A(n50), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n50) );
  OAI21_X1 U27 ( .B1(n85), .B2(ENABLE), .A(n51), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n51) );
  OAI21_X1 U29 ( .B1(n84), .B2(ENABLE), .A(n52), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n52) );
  OAI21_X1 U31 ( .B1(n83), .B2(ENABLE), .A(n54), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n82), .B2(ENABLE), .A(n55), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n55) );
  OAI21_X1 U35 ( .B1(n81), .B2(ENABLE), .A(n56), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n56) );
  OAI21_X1 U37 ( .B1(n80), .B2(ENABLE), .A(n57), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n57) );
  OAI21_X1 U39 ( .B1(n79), .B2(ENABLE), .A(n58), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n58) );
  OAI21_X1 U41 ( .B1(n78), .B2(ENABLE), .A(n59), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n59) );
  OAI21_X1 U43 ( .B1(n77), .B2(ENABLE), .A(n60), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n60) );
  OAI21_X1 U45 ( .B1(n76), .B2(ENABLE), .A(n61), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n61) );
  OAI21_X1 U47 ( .B1(n75), .B2(ENABLE), .A(n62), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n62) );
  OAI21_X1 U49 ( .B1(n74), .B2(ENABLE), .A(n63), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n63) );
  OAI21_X1 U51 ( .B1(n73), .B2(ENABLE), .A(n33), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U53 ( .B1(n72), .B2(ENABLE), .A(n34), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n34) );
  OAI21_X1 U55 ( .B1(n71), .B2(ENABLE), .A(n35), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n35) );
  OAI21_X1 U57 ( .B1(n70), .B2(ENABLE), .A(n36), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n36) );
  OAI21_X1 U59 ( .B1(n69), .B2(ENABLE), .A(n37), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n37) );
  OAI21_X1 U61 ( .B1(n68), .B2(ENABLE), .A(n38), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n38) );
  OAI21_X1 U63 ( .B1(n67), .B2(ENABLE), .A(n42), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n42) );
  OAI21_X1 U65 ( .B1(n66), .B2(ENABLE), .A(n53), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n65), .B2(ENABLE), .A(n64), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n64) );
endmodule


module regFFD_NBIT32_9 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n65) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n66) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n67) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n68) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n69) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n70) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n71) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n72) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n99), .Q(Q[23]), .QN(n73) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n74) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n75) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n97), .Q(Q[20]), .QN(n76) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n99), .Q(Q[19]), .QN(n77) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n78) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n79) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n80) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n99), .Q(Q[15]), .QN(n81) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n82) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n83) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n84) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n97), .Q(Q[11]), .QN(n85) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n97), .Q(Q[10]), .QN(n86) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n87) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n97), .Q(Q[8]), .QN(n88) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n89) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n90) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n98), .Q(Q[5]), .QN(n91) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n98), .Q(Q[4]), .QN(n92) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n93) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n98), .Q(Q[2]), .QN(n94) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n98), .Q(Q[1]), .QN(n95) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n96) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n96), .B2(ENABLE), .A(n39), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n39) );
  OAI21_X1 U7 ( .B1(n95), .B2(ENABLE), .A(n40), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n40) );
  OAI21_X1 U9 ( .B1(n94), .B2(ENABLE), .A(n41), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n41) );
  OAI21_X1 U11 ( .B1(n93), .B2(ENABLE), .A(n43), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n43) );
  OAI21_X1 U13 ( .B1(n92), .B2(ENABLE), .A(n44), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n91), .B2(ENABLE), .A(n45), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n45) );
  OAI21_X1 U17 ( .B1(n90), .B2(ENABLE), .A(n46), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n46) );
  OAI21_X1 U19 ( .B1(n89), .B2(ENABLE), .A(n47), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n47) );
  OAI21_X1 U21 ( .B1(n88), .B2(ENABLE), .A(n48), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n48) );
  OAI21_X1 U23 ( .B1(n87), .B2(ENABLE), .A(n49), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n49) );
  OAI21_X1 U25 ( .B1(n86), .B2(ENABLE), .A(n50), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n50) );
  OAI21_X1 U27 ( .B1(n85), .B2(ENABLE), .A(n51), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n51) );
  OAI21_X1 U29 ( .B1(n84), .B2(ENABLE), .A(n52), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n52) );
  OAI21_X1 U31 ( .B1(n83), .B2(ENABLE), .A(n54), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n82), .B2(ENABLE), .A(n55), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n55) );
  OAI21_X1 U35 ( .B1(n81), .B2(ENABLE), .A(n56), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n56) );
  OAI21_X1 U37 ( .B1(n80), .B2(ENABLE), .A(n57), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n57) );
  OAI21_X1 U39 ( .B1(n79), .B2(ENABLE), .A(n58), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n58) );
  OAI21_X1 U41 ( .B1(n78), .B2(ENABLE), .A(n59), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n59) );
  OAI21_X1 U43 ( .B1(n77), .B2(ENABLE), .A(n60), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n60) );
  OAI21_X1 U45 ( .B1(n76), .B2(ENABLE), .A(n61), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n61) );
  OAI21_X1 U47 ( .B1(n75), .B2(ENABLE), .A(n62), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n62) );
  OAI21_X1 U49 ( .B1(n74), .B2(ENABLE), .A(n63), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n63) );
  OAI21_X1 U51 ( .B1(n73), .B2(ENABLE), .A(n33), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U53 ( .B1(n72), .B2(ENABLE), .A(n34), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n34) );
  OAI21_X1 U55 ( .B1(n71), .B2(ENABLE), .A(n35), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n35) );
  OAI21_X1 U57 ( .B1(n70), .B2(ENABLE), .A(n36), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n36) );
  OAI21_X1 U59 ( .B1(n69), .B2(ENABLE), .A(n37), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n37) );
  OAI21_X1 U61 ( .B1(n68), .B2(ENABLE), .A(n38), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n38) );
  OAI21_X1 U63 ( .B1(n67), .B2(ENABLE), .A(n42), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n42) );
  OAI21_X1 U65 ( .B1(n66), .B2(ENABLE), .A(n53), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n65), .B2(ENABLE), .A(n64), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n64) );
endmodule


module regFFD_NBIT32_8 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n65) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n66) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n67) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n68) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n69) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n70) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n71) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n98), .Q(Q[24]), .QN(n72) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n73) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n74) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n75) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n76) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n97), .Q(Q[19]), .QN(n77) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n78) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n97), .Q(Q[17]), .QN(n79) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n80) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n81) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n82) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n83) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n84) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n85) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n86) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n87) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n88) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n89) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n90) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n91) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n92) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n93) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n94) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n95) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n96) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n96), .B2(ENABLE), .A(n39), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n39) );
  OAI21_X1 U7 ( .B1(n95), .B2(ENABLE), .A(n40), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n40) );
  OAI21_X1 U9 ( .B1(n94), .B2(ENABLE), .A(n41), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n41) );
  OAI21_X1 U11 ( .B1(n93), .B2(ENABLE), .A(n43), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n43) );
  OAI21_X1 U13 ( .B1(n92), .B2(ENABLE), .A(n44), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n91), .B2(ENABLE), .A(n45), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n45) );
  OAI21_X1 U17 ( .B1(n90), .B2(ENABLE), .A(n46), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n46) );
  OAI21_X1 U19 ( .B1(n89), .B2(ENABLE), .A(n47), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n47) );
  OAI21_X1 U21 ( .B1(n88), .B2(ENABLE), .A(n48), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n48) );
  OAI21_X1 U23 ( .B1(n87), .B2(ENABLE), .A(n49), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n49) );
  OAI21_X1 U25 ( .B1(n86), .B2(ENABLE), .A(n50), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n50) );
  OAI21_X1 U27 ( .B1(n85), .B2(ENABLE), .A(n51), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n51) );
  OAI21_X1 U29 ( .B1(n84), .B2(ENABLE), .A(n52), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n52) );
  OAI21_X1 U31 ( .B1(n83), .B2(ENABLE), .A(n54), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n82), .B2(ENABLE), .A(n55), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n55) );
  OAI21_X1 U35 ( .B1(n81), .B2(ENABLE), .A(n56), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n56) );
  OAI21_X1 U37 ( .B1(n80), .B2(ENABLE), .A(n57), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n57) );
  OAI21_X1 U39 ( .B1(n79), .B2(ENABLE), .A(n58), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n58) );
  OAI21_X1 U41 ( .B1(n78), .B2(ENABLE), .A(n59), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n59) );
  OAI21_X1 U43 ( .B1(n77), .B2(ENABLE), .A(n60), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n60) );
  OAI21_X1 U45 ( .B1(n76), .B2(ENABLE), .A(n61), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n61) );
  OAI21_X1 U47 ( .B1(n75), .B2(ENABLE), .A(n62), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n62) );
  OAI21_X1 U49 ( .B1(n74), .B2(ENABLE), .A(n63), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n63) );
  OAI21_X1 U51 ( .B1(n73), .B2(ENABLE), .A(n33), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U53 ( .B1(n72), .B2(ENABLE), .A(n34), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n34) );
  OAI21_X1 U55 ( .B1(n71), .B2(ENABLE), .A(n35), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n35) );
  OAI21_X1 U57 ( .B1(n70), .B2(ENABLE), .A(n36), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n36) );
  OAI21_X1 U59 ( .B1(n69), .B2(ENABLE), .A(n37), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n37) );
  OAI21_X1 U61 ( .B1(n68), .B2(ENABLE), .A(n38), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n38) );
  OAI21_X1 U63 ( .B1(n67), .B2(ENABLE), .A(n42), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n42) );
  OAI21_X1 U65 ( .B1(n66), .B2(ENABLE), .A(n53), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n53) );
  OAI21_X1 U67 ( .B1(n65), .B2(ENABLE), .A(n64), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n64) );
endmodule


module regFFD_NBIT5_0 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n11) );
  DFFR_X1 \Q_reg[3]  ( .D(n2), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n12) );
  DFFR_X1 \Q_reg[2]  ( .D(n3), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n13) );
  DFFR_X1 \Q_reg[1]  ( .D(n4), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n14) );
  DFFR_X1 \Q_reg[0]  ( .D(n5), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n15) );
  OAI21_X1 U2 ( .B1(n14), .B2(ENABLE), .A(n7), .ZN(n4) );
  NAND2_X1 U3 ( .A1(D[1]), .A2(ENABLE), .ZN(n7) );
  OAI21_X1 U4 ( .B1(n13), .B2(ENABLE), .A(n8), .ZN(n3) );
  NAND2_X1 U5 ( .A1(D[2]), .A2(ENABLE), .ZN(n8) );
  OAI21_X1 U6 ( .B1(n12), .B2(ENABLE), .A(n9), .ZN(n2) );
  NAND2_X1 U7 ( .A1(D[3]), .A2(ENABLE), .ZN(n9) );
  OAI21_X1 U8 ( .B1(n11), .B2(ENABLE), .A(n10), .ZN(n1) );
  NAND2_X1 U9 ( .A1(D[4]), .A2(ENABLE), .ZN(n10) );
  OAI21_X1 U10 ( .B1(n15), .B2(ENABLE), .A(n6), .ZN(n5) );
  NAND2_X1 U11 ( .A1(ENABLE), .A2(D[0]), .ZN(n6) );
endmodule


module FF_7 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n2, n3, n5, n6;

  DFF_X1 Q_reg ( .D(n2), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n3), .ZN(n2) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n5), .B2(Q), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n5) );
  INV_X1 U6 ( .A(RESET), .ZN(n3) );
endmodule


module regFFD_NBIT6_0 ( CK, RESET, ENABLE, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  DFFR_X1 \Q_reg[5]  ( .D(n1), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n13) );
  DFFR_X1 \Q_reg[4]  ( .D(n2), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n14) );
  DFFR_X1 \Q_reg[3]  ( .D(n3), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n15) );
  DFFR_X1 \Q_reg[2]  ( .D(n4), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n16) );
  DFFR_X1 \Q_reg[1]  ( .D(n5), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n17) );
  DFFR_X1 \Q_reg[0]  ( .D(n6), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n18) );
  OAI21_X1 U2 ( .B1(n13), .B2(ENABLE), .A(n12), .ZN(n1) );
  NAND2_X1 U3 ( .A1(D[5]), .A2(ENABLE), .ZN(n12) );
  OAI21_X1 U4 ( .B1(n16), .B2(ENABLE), .A(n9), .ZN(n4) );
  NAND2_X1 U5 ( .A1(D[2]), .A2(ENABLE), .ZN(n9) );
  OAI21_X1 U6 ( .B1(n14), .B2(ENABLE), .A(n11), .ZN(n2) );
  NAND2_X1 U7 ( .A1(D[4]), .A2(ENABLE), .ZN(n11) );
  OAI21_X1 U8 ( .B1(n15), .B2(ENABLE), .A(n10), .ZN(n3) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n10) );
  OAI21_X1 U10 ( .B1(n17), .B2(ENABLE), .A(n8), .ZN(n5) );
  NAND2_X1 U11 ( .A1(D[1]), .A2(ENABLE), .ZN(n8) );
  OAI21_X1 U12 ( .B1(n18), .B2(ENABLE), .A(n7), .ZN(n6) );
  NAND2_X1 U13 ( .A1(ENABLE), .A2(D[0]), .ZN(n7) );
endmodule


module regFFD_NBIT32_7 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U7 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U8 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U9 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U10 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U11 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U12 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U13 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U14 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U15 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U16 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U17 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U18 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U19 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U20 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U21 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U22 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U23 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U24 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U25 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U26 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U27 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U28 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U29 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U30 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U31 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U32 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U33 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U34 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U35 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U36 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
  OAI21_X1 U37 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U38 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U39 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U40 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U41 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U42 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U43 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U44 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U45 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U46 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U47 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U48 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U49 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U50 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U51 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U52 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U53 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U54 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U55 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U56 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U57 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U58 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U59 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U60 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U61 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U62 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U63 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U64 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U65 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U66 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U67 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U68 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
endmodule


module regFFD_NBIT32_6 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U7 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U8 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U9 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U10 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U11 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U12 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U13 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U14 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U15 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U16 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U17 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U18 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U19 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U20 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U21 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U22 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U23 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U24 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U25 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U26 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U27 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U28 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U29 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U30 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U31 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U32 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U33 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U34 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U35 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U36 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U37 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U38 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U39 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U40 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U41 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U42 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U43 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U44 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U45 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U46 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U47 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U48 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U49 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U50 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U51 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U52 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module IV_224 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_672 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_671 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_670 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_224 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_224 UIV ( .A(S), .Y(SB) );
  ND2_672 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_671 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_670 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_223 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_669 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_668 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_667 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_223 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_223 UIV ( .A(S), .Y(SB) );
  ND2_669 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_668 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_667 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_222 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_666 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_665 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_664 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_222 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_222 UIV ( .A(S), .Y(SB) );
  ND2_666 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_665 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_664 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_221 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_663 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_662 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_661 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_221 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_221 UIV ( .A(S), .Y(SB) );
  ND2_663 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_662 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_661 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_220 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_660 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_659 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_658 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_220 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_220 UIV ( .A(S), .Y(SB) );
  ND2_660 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_659 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_658 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_219 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_657 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_656 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_655 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_219 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_219 UIV ( .A(S), .Y(SB) );
  ND2_657 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_656 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_655 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_218 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_654 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_653 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_652 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_218 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_218 UIV ( .A(S), .Y(SB) );
  ND2_654 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_653 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_652 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_217 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_651 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_650 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_649 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_217 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_217 UIV ( .A(S), .Y(SB) );
  ND2_651 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_650 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_649 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_216 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_648 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_647 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_646 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_216 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_216 UIV ( .A(S), .Y(SB) );
  ND2_648 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_647 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_646 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_215 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_645 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_644 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_643 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_215 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_215 UIV ( .A(S), .Y(SB) );
  ND2_645 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_644 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_643 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_214 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_642 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_641 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_640 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_214 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_214 UIV ( .A(S), .Y(SB) );
  ND2_642 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_641 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_640 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_213 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_639 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_638 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_637 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_213 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_213 UIV ( .A(S), .Y(SB) );
  ND2_639 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_638 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_637 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_212 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_636 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_635 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_634 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_212 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_212 UIV ( .A(S), .Y(SB) );
  ND2_636 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_635 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_634 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_211 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_633 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_632 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_631 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_211 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_211 UIV ( .A(S), .Y(SB) );
  ND2_633 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_632 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_631 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_210 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_630 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_629 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_628 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_210 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_210 UIV ( .A(S), .Y(SB) );
  ND2_630 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_629 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_628 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_209 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_627 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_626 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_625 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_209 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_209 UIV ( .A(S), .Y(SB) );
  ND2_627 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_626 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_625 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_208 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_624 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_623 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_622 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_208 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_208 UIV ( .A(S), .Y(SB) );
  ND2_624 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_623 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_622 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_207 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_621 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_620 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_619 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_207 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_207 UIV ( .A(S), .Y(SB) );
  ND2_621 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_620 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_619 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_206 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_618 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_617 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_616 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_206 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_206 UIV ( .A(S), .Y(SB) );
  ND2_618 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_617 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_616 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_205 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_615 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_614 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_205 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_205 UIV ( .A(S), .Y(SB) );
  ND2_615 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_614 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_613 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_204 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_204 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_204 UIV ( .A(S), .Y(SB) );
  ND2_612 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_611 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_610 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_203 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_203 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_203 UIV ( .A(S), .Y(SB) );
  ND2_609 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_608 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_607 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_202 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_202 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_202 UIV ( .A(S), .Y(SB) );
  ND2_606 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_605 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_604 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_201 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_201 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_201 UIV ( .A(S), .Y(SB) );
  ND2_603 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_602 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_601 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_200 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_200 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_200 UIV ( .A(S), .Y(SB) );
  ND2_600 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_599 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_598 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_199 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_199 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_199 UIV ( .A(S), .Y(SB) );
  ND2_597 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_596 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_595 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_198 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_198 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_198 UIV ( .A(S), .Y(SB) );
  ND2_594 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_593 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_592 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_197 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_197 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_197 UIV ( .A(S), .Y(SB) );
  ND2_591 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_590 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_589 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_196 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_196 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_196 UIV ( .A(S), .Y(SB) );
  ND2_588 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_587 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_586 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_195 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_195 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_195 UIV ( .A(S), .Y(SB) );
  ND2_585 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_584 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_583 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_194 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_194 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_194 UIV ( .A(S), .Y(SB) );
  ND2_582 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_581 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_580 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_193 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_193 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_193 UIV ( .A(S), .Y(SB) );
  ND2_579 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_578 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_577 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_6 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_224 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_223 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_222 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_221 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_220 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_219 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_218 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_217 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_216 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_215 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_214 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_213 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_212 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_211 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_210 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_209 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_208 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_207 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_206 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_205 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_204 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_203 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_202 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_201 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_200 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_199 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_198 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_197 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_196 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_195 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_194 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_193 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_192 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_192 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_192 UIV ( .A(S), .Y(SB) );
  ND2_576 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_575 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_574 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_191 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_191 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_191 UIV ( .A(S), .Y(SB) );
  ND2_573 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_572 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_571 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_190 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_190 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_190 UIV ( .A(S), .Y(SB) );
  ND2_570 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_569 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_568 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_189 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_189 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_189 UIV ( .A(S), .Y(SB) );
  ND2_567 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_566 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_565 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_188 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_188 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_188 UIV ( .A(S), .Y(SB) );
  ND2_564 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_563 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_562 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_187 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_187 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_187 UIV ( .A(S), .Y(SB) );
  ND2_561 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_560 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_559 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_186 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_186 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_186 UIV ( .A(S), .Y(SB) );
  ND2_558 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_557 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_556 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_185 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_185 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_185 UIV ( .A(S), .Y(SB) );
  ND2_555 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_554 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_553 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_184 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_184 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_184 UIV ( .A(S), .Y(SB) );
  ND2_552 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_551 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_550 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_183 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_183 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_183 UIV ( .A(S), .Y(SB) );
  ND2_549 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_548 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_547 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_182 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_182 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_182 UIV ( .A(S), .Y(SB) );
  ND2_546 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_545 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_544 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_181 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_181 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_181 UIV ( .A(S), .Y(SB) );
  ND2_543 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_542 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_541 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_180 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_180 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_180 UIV ( .A(S), .Y(SB) );
  ND2_540 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_539 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_538 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_179 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_179 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_179 UIV ( .A(S), .Y(SB) );
  ND2_537 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_536 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_535 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_178 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_178 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_178 UIV ( .A(S), .Y(SB) );
  ND2_534 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_533 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_532 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_177 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_177 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_177 UIV ( .A(S), .Y(SB) );
  ND2_531 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_530 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_529 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_176 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_176 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_176 UIV ( .A(S), .Y(SB) );
  ND2_528 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_527 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_526 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_175 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_175 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_175 UIV ( .A(S), .Y(SB) );
  ND2_525 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_524 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_523 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_174 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_174 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_174 UIV ( .A(S), .Y(SB) );
  ND2_522 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_521 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_520 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_173 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_173 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_173 UIV ( .A(S), .Y(SB) );
  ND2_519 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_518 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_517 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_172 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_172 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_172 UIV ( .A(S), .Y(SB) );
  ND2_516 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_515 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_514 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_171 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_171 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_171 UIV ( .A(S), .Y(SB) );
  ND2_513 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_512 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_511 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_170 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_170 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_170 UIV ( .A(S), .Y(SB) );
  ND2_510 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_509 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_508 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_169 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_169 UIV ( .A(S), .Y(SB) );
  ND2_507 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_506 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_505 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_168 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_168 UIV ( .A(S), .Y(SB) );
  ND2_504 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_503 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_502 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_167 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_167 UIV ( .A(S), .Y(SB) );
  ND2_501 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_500 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_499 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_166 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_166 UIV ( .A(S), .Y(SB) );
  ND2_498 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_497 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_496 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_165 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_165 UIV ( .A(S), .Y(SB) );
  ND2_495 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_494 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_493 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_164 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_164 UIV ( .A(S), .Y(SB) );
  ND2_492 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_491 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_490 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_163 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_163 UIV ( .A(S), .Y(SB) );
  ND2_489 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_488 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_487 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_162 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_162 UIV ( .A(S), .Y(SB) );
  ND2_486 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_485 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_484 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_161 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_161 UIV ( .A(S), .Y(SB) );
  ND2_483 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_482 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_481 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_5 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_192 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_191 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_190 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_189 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_188 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_187 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_186 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_185 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_184 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_183 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_182 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_181 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_180 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_179 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_178 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_177 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_176 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_175 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_174 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_173 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_172 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_171 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_170 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_169 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_168 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_167 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_166 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_165 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_164 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_163 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_162 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_161 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module logic_N32 ( .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , 
        \FUNC[1] , \FUNC[0] }), DATA1, DATA2, OUT_ALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUT_ALU;
  input \FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258;
  wire   [5:0] FUNC;

  NAND3_X1 U172 ( .A1(n258), .A2(n257), .A3(FUNC[3]), .ZN(n139) );
  BUF_X1 U2 ( .A(n177), .Z(n180) );
  BUF_X1 U3 ( .A(n177), .Z(n179) );
  BUF_X1 U4 ( .A(n178), .Z(n182) );
  BUF_X1 U5 ( .A(n178), .Z(n183) );
  BUF_X1 U6 ( .A(n177), .Z(n181) );
  AOI21_X1 U7 ( .B1(n191), .B2(n245), .A(n183), .ZN(n122) );
  AOI21_X1 U8 ( .B1(n191), .B2(n246), .A(n183), .ZN(n124) );
  AOI21_X1 U9 ( .B1(n191), .B2(n247), .A(n183), .ZN(n126) );
  AOI21_X1 U10 ( .B1(n191), .B2(n248), .A(n183), .ZN(n128) );
  AOI21_X1 U11 ( .B1(n191), .B2(n249), .A(n184), .ZN(n130) );
  AOI21_X1 U12 ( .B1(n191), .B2(n250), .A(n184), .ZN(n132) );
  AOI21_X1 U13 ( .B1(n190), .B2(n193), .A(n183), .ZN(n112) );
  AOI21_X1 U14 ( .B1(n189), .B2(n194), .A(n182), .ZN(n90) );
  AOI21_X1 U15 ( .B1(n189), .B2(n229), .A(n182), .ZN(n86) );
  AOI21_X1 U16 ( .B1(n189), .B2(n230), .A(n182), .ZN(n88) );
  AOI21_X1 U17 ( .B1(n189), .B2(n231), .A(n182), .ZN(n92) );
  AOI21_X1 U18 ( .B1(n189), .B2(n232), .A(n182), .ZN(n94) );
  AOI21_X1 U19 ( .B1(n189), .B2(n233), .A(n182), .ZN(n96) );
  AOI21_X1 U20 ( .B1(n190), .B2(n234), .A(n182), .ZN(n98) );
  AOI21_X1 U21 ( .B1(n190), .B2(n235), .A(n182), .ZN(n100) );
  AOI21_X1 U22 ( .B1(n190), .B2(n236), .A(n182), .ZN(n102) );
  AOI21_X1 U23 ( .B1(n190), .B2(n237), .A(n183), .ZN(n104) );
  AOI21_X1 U24 ( .B1(n190), .B2(n238), .A(n183), .ZN(n106) );
  AOI21_X1 U25 ( .B1(n190), .B2(n239), .A(n183), .ZN(n108) );
  AOI21_X1 U26 ( .B1(n190), .B2(n240), .A(n183), .ZN(n110) );
  AOI21_X1 U27 ( .B1(n190), .B2(n241), .A(n183), .ZN(n114) );
  AOI21_X1 U28 ( .B1(n190), .B2(n242), .A(n183), .ZN(n116) );
  AOI21_X1 U29 ( .B1(n190), .B2(n243), .A(n183), .ZN(n118) );
  AOI21_X1 U30 ( .B1(n190), .B2(n244), .A(n183), .ZN(n120) );
  AOI21_X1 U31 ( .B1(n189), .B2(n251), .A(n182), .ZN(n69) );
  AOI21_X1 U32 ( .B1(n188), .B2(n252), .A(n181), .ZN(n74) );
  AOI21_X1 U33 ( .B1(n189), .B2(n253), .A(n182), .ZN(n76) );
  AOI21_X1 U34 ( .B1(n189), .B2(n254), .A(n181), .ZN(n78) );
  AOI21_X1 U35 ( .B1(n189), .B2(n255), .A(n181), .ZN(n80) );
  AOI21_X1 U36 ( .B1(n189), .B2(n196), .A(n182), .ZN(n82) );
  AOI21_X1 U37 ( .B1(n189), .B2(n195), .A(n182), .ZN(n84) );
  OAI22_X1 U38 ( .A1(n85), .A2(n229), .B1(n86), .B2(n197), .ZN(OUT_ALU[31]) );
  OAI22_X1 U39 ( .A1(n87), .A2(n230), .B1(n88), .B2(n198), .ZN(OUT_ALU[30]) );
  OAI22_X1 U40 ( .A1(n91), .A2(n231), .B1(n92), .B2(n199), .ZN(OUT_ALU[29]) );
  OAI22_X1 U41 ( .A1(n93), .A2(n232), .B1(n94), .B2(n200), .ZN(OUT_ALU[28]) );
  OAI22_X1 U42 ( .A1(n95), .A2(n233), .B1(n96), .B2(n201), .ZN(OUT_ALU[27]) );
  OAI22_X1 U43 ( .A1(n97), .A2(n234), .B1(n98), .B2(n202), .ZN(OUT_ALU[26]) );
  OAI22_X1 U44 ( .A1(n99), .A2(n235), .B1(n100), .B2(n203), .ZN(OUT_ALU[25])
         );
  OAI22_X1 U45 ( .A1(n101), .A2(n236), .B1(n102), .B2(n204), .ZN(OUT_ALU[24])
         );
  OAI22_X1 U46 ( .A1(n103), .A2(n237), .B1(n104), .B2(n205), .ZN(OUT_ALU[23])
         );
  OAI22_X1 U47 ( .A1(n105), .A2(n238), .B1(n106), .B2(n206), .ZN(OUT_ALU[22])
         );
  OAI22_X1 U48 ( .A1(n107), .A2(n239), .B1(n108), .B2(n207), .ZN(OUT_ALU[21])
         );
  OAI22_X1 U49 ( .A1(n109), .A2(n240), .B1(n110), .B2(n208), .ZN(OUT_ALU[20])
         );
  OAI22_X1 U50 ( .A1(n113), .A2(n241), .B1(n114), .B2(n209), .ZN(OUT_ALU[19])
         );
  OAI22_X1 U51 ( .A1(n115), .A2(n242), .B1(n116), .B2(n210), .ZN(OUT_ALU[18])
         );
  OAI22_X1 U52 ( .A1(n117), .A2(n243), .B1(n118), .B2(n211), .ZN(OUT_ALU[17])
         );
  OAI22_X1 U53 ( .A1(n119), .A2(n244), .B1(n120), .B2(n212), .ZN(OUT_ALU[16])
         );
  OAI22_X1 U54 ( .A1(n121), .A2(n245), .B1(n122), .B2(n213), .ZN(OUT_ALU[15])
         );
  OAI22_X1 U55 ( .A1(n123), .A2(n246), .B1(n124), .B2(n214), .ZN(OUT_ALU[14])
         );
  OAI22_X1 U56 ( .A1(n125), .A2(n247), .B1(n126), .B2(n215), .ZN(OUT_ALU[13])
         );
  OAI22_X1 U57 ( .A1(n127), .A2(n248), .B1(n128), .B2(n216), .ZN(OUT_ALU[12])
         );
  OAI22_X1 U58 ( .A1(n129), .A2(n249), .B1(n130), .B2(n217), .ZN(OUT_ALU[11])
         );
  OAI22_X1 U59 ( .A1(n131), .A2(n250), .B1(n132), .B2(n218), .ZN(OUT_ALU[10])
         );
  OAI22_X1 U60 ( .A1(n68), .A2(n251), .B1(n69), .B2(n219), .ZN(OUT_ALU[9]) );
  OAI22_X1 U61 ( .A1(n73), .A2(n252), .B1(n74), .B2(n220), .ZN(OUT_ALU[8]) );
  OAI22_X1 U62 ( .A1(n75), .A2(n253), .B1(n76), .B2(n221), .ZN(OUT_ALU[7]) );
  OAI22_X1 U63 ( .A1(n77), .A2(n254), .B1(n78), .B2(n222), .ZN(OUT_ALU[6]) );
  OAI22_X1 U64 ( .A1(n79), .A2(n255), .B1(n80), .B2(n223), .ZN(OUT_ALU[5]) );
  OAI22_X1 U65 ( .A1(n81), .A2(n196), .B1(n82), .B2(n224), .ZN(OUT_ALU[4]) );
  BUF_X1 U66 ( .A(n178), .Z(n184) );
  AOI221_X1 U67 ( .B1(n186), .B2(n219), .C1(n176), .C2(DATA1[9]), .A(n179), 
        .ZN(n68) );
  AOI221_X1 U68 ( .B1(n188), .B2(n200), .C1(DATA1[28]), .C2(n175), .A(n181), 
        .ZN(n93) );
  AOI221_X1 U69 ( .B1(n188), .B2(n202), .C1(DATA1[26]), .C2(n175), .A(n180), 
        .ZN(n97) );
  AOI221_X1 U70 ( .B1(n188), .B2(n203), .C1(DATA1[25]), .C2(n175), .A(n181), 
        .ZN(n99) );
  AOI221_X1 U71 ( .B1(n188), .B2(n204), .C1(DATA1[24]), .C2(n175), .A(n181), 
        .ZN(n101) );
  AOI221_X1 U72 ( .B1(n187), .B2(n205), .C1(DATA1[23]), .C2(n175), .A(n180), 
        .ZN(n103) );
  AOI221_X1 U73 ( .B1(n188), .B2(n206), .C1(DATA1[22]), .C2(n175), .A(n180), 
        .ZN(n105) );
  AOI221_X1 U74 ( .B1(n187), .B2(n211), .C1(DATA1[17]), .C2(n174), .A(n180), 
        .ZN(n117) );
  AOI221_X1 U75 ( .B1(n187), .B2(n212), .C1(DATA1[16]), .C2(n174), .A(n179), 
        .ZN(n119) );
  AOI221_X1 U76 ( .B1(n186), .B2(n213), .C1(DATA1[15]), .C2(n174), .A(n179), 
        .ZN(n121) );
  AOI221_X1 U77 ( .B1(n186), .B2(n214), .C1(DATA1[14]), .C2(n174), .A(n179), 
        .ZN(n123) );
  AOI221_X1 U78 ( .B1(n186), .B2(n215), .C1(DATA1[13]), .C2(n174), .A(n179), 
        .ZN(n125) );
  AOI221_X1 U79 ( .B1(n186), .B2(n216), .C1(DATA1[12]), .C2(n174), .A(n179), 
        .ZN(n127) );
  AOI221_X1 U80 ( .B1(n188), .B2(n197), .C1(DATA1[31]), .C2(n176), .A(n181), 
        .ZN(n85) );
  AOI221_X1 U81 ( .B1(n188), .B2(n199), .C1(DATA1[29]), .C2(n175), .A(n181), 
        .ZN(n91) );
  AOI221_X1 U82 ( .B1(n188), .B2(n201), .C1(DATA1[27]), .C2(n175), .A(n181), 
        .ZN(n95) );
  AOI221_X1 U83 ( .B1(n187), .B2(n207), .C1(DATA1[21]), .C2(n175), .A(n180), 
        .ZN(n107) );
  AOI221_X1 U84 ( .B1(n187), .B2(n208), .C1(DATA1[20]), .C2(n175), .A(n180), 
        .ZN(n109) );
  AOI221_X1 U85 ( .B1(n187), .B2(n209), .C1(DATA1[19]), .C2(n174), .A(n180), 
        .ZN(n113) );
  AOI221_X1 U86 ( .B1(n186), .B2(n217), .C1(DATA1[11]), .C2(n174), .A(n179), 
        .ZN(n129) );
  AOI221_X1 U87 ( .B1(n186), .B2(n218), .C1(DATA1[10]), .C2(n174), .A(n179), 
        .ZN(n131) );
  AOI221_X1 U88 ( .B1(n186), .B2(n220), .C1(DATA1[8]), .C2(n176), .A(n179), 
        .ZN(n73) );
  AOI221_X1 U89 ( .B1(n186), .B2(n221), .C1(DATA1[7]), .C2(n176), .A(n179), 
        .ZN(n75) );
  AOI221_X1 U90 ( .B1(n186), .B2(n222), .C1(DATA1[6]), .C2(n176), .A(n179), 
        .ZN(n77) );
  AOI221_X1 U91 ( .B1(n187), .B2(n223), .C1(DATA1[5]), .C2(n176), .A(n180), 
        .ZN(n79) );
  AOI221_X1 U92 ( .B1(n187), .B2(n224), .C1(DATA1[4]), .C2(n176), .A(n180), 
        .ZN(n81) );
  AOI221_X1 U93 ( .B1(n187), .B2(n225), .C1(DATA1[3]), .C2(n176), .A(n180), 
        .ZN(n83) );
  AOI221_X1 U94 ( .B1(n188), .B2(n226), .C1(DATA1[2]), .C2(n175), .A(n181), 
        .ZN(n89) );
  AOI221_X1 U95 ( .B1(n188), .B2(n198), .C1(DATA1[30]), .C2(n175), .A(n181), 
        .ZN(n87) );
  AOI221_X1 U96 ( .B1(n187), .B2(n210), .C1(DATA1[18]), .C2(n174), .A(n180), 
        .ZN(n115) );
  AOI221_X1 U97 ( .B1(n187), .B2(n227), .C1(DATA1[1]), .C2(n174), .A(n180), 
        .ZN(n111) );
  BUF_X1 U98 ( .A(n72), .Z(n175) );
  BUF_X1 U99 ( .A(n72), .Z(n174) );
  OAI22_X1 U100 ( .A1(n133), .A2(n192), .B1(n134), .B2(n228), .ZN(OUT_ALU[0])
         );
  AOI21_X1 U101 ( .B1(n188), .B2(n192), .A(n181), .ZN(n134) );
  AOI221_X1 U102 ( .B1(n186), .B2(n228), .C1(DATA1[0]), .C2(n174), .A(n179), 
        .ZN(n133) );
  BUF_X1 U103 ( .A(n185), .Z(n188) );
  BUF_X1 U104 ( .A(n185), .Z(n189) );
  BUF_X1 U105 ( .A(n185), .Z(n190) );
  BUF_X1 U106 ( .A(n72), .Z(n176) );
  BUF_X1 U107 ( .A(n185), .Z(n187) );
  BUF_X1 U108 ( .A(n185), .Z(n186) );
  INV_X1 U109 ( .A(DATA1[12]), .ZN(n216) );
  INV_X1 U110 ( .A(DATA1[13]), .ZN(n215) );
  INV_X1 U111 ( .A(DATA1[14]), .ZN(n214) );
  INV_X1 U112 ( .A(DATA1[23]), .ZN(n205) );
  INV_X1 U113 ( .A(DATA1[22]), .ZN(n206) );
  INV_X1 U114 ( .A(DATA1[17]), .ZN(n211) );
  INV_X1 U115 ( .A(DATA1[16]), .ZN(n212) );
  INV_X1 U116 ( .A(DATA1[15]), .ZN(n213) );
  INV_X1 U117 ( .A(DATA1[21]), .ZN(n207) );
  INV_X1 U118 ( .A(DATA1[9]), .ZN(n219) );
  INV_X1 U119 ( .A(DATA1[11]), .ZN(n217) );
  INV_X1 U120 ( .A(DATA1[10]), .ZN(n218) );
  INV_X1 U121 ( .A(DATA1[8]), .ZN(n220) );
  INV_X1 U122 ( .A(DATA1[7]), .ZN(n221) );
  INV_X1 U123 ( .A(DATA1[2]), .ZN(n226) );
  INV_X1 U124 ( .A(DATA1[3]), .ZN(n225) );
  INV_X1 U125 ( .A(DATA1[28]), .ZN(n200) );
  INV_X1 U126 ( .A(DATA1[27]), .ZN(n201) );
  INV_X1 U127 ( .A(DATA1[26]), .ZN(n202) );
  INV_X1 U128 ( .A(DATA1[25]), .ZN(n203) );
  INV_X1 U129 ( .A(DATA1[24]), .ZN(n204) );
  INV_X1 U130 ( .A(DATA1[18]), .ZN(n210) );
  INV_X1 U131 ( .A(DATA1[0]), .ZN(n228) );
  INV_X1 U132 ( .A(DATA1[6]), .ZN(n222) );
  INV_X1 U133 ( .A(DATA1[29]), .ZN(n199) );
  INV_X1 U134 ( .A(DATA1[4]), .ZN(n224) );
  INV_X1 U135 ( .A(DATA1[1]), .ZN(n227) );
  INV_X1 U136 ( .A(DATA1[19]), .ZN(n209) );
  INV_X1 U137 ( .A(DATA1[20]), .ZN(n208) );
  INV_X1 U138 ( .A(DATA1[31]), .ZN(n197) );
  INV_X1 U139 ( .A(DATA1[5]), .ZN(n223) );
  INV_X1 U140 ( .A(DATA1[30]), .ZN(n198) );
  BUF_X1 U141 ( .A(n71), .Z(n177) );
  BUF_X1 U142 ( .A(n71), .Z(n178) );
  INV_X1 U143 ( .A(DATA2[31]), .ZN(n229) );
  INV_X1 U144 ( .A(DATA2[30]), .ZN(n230) );
  INV_X1 U145 ( .A(DATA2[29]), .ZN(n231) );
  INV_X1 U146 ( .A(DATA2[28]), .ZN(n232) );
  INV_X1 U147 ( .A(DATA2[27]), .ZN(n233) );
  INV_X1 U148 ( .A(DATA2[26]), .ZN(n234) );
  INV_X1 U149 ( .A(DATA2[25]), .ZN(n235) );
  INV_X1 U150 ( .A(DATA2[24]), .ZN(n236) );
  INV_X1 U151 ( .A(DATA2[23]), .ZN(n237) );
  INV_X1 U152 ( .A(DATA2[22]), .ZN(n238) );
  INV_X1 U153 ( .A(DATA2[21]), .ZN(n239) );
  INV_X1 U154 ( .A(DATA2[20]), .ZN(n240) );
  INV_X1 U155 ( .A(DATA2[19]), .ZN(n241) );
  INV_X1 U156 ( .A(DATA2[18]), .ZN(n242) );
  INV_X1 U157 ( .A(DATA2[17]), .ZN(n243) );
  INV_X1 U158 ( .A(DATA2[16]), .ZN(n244) );
  INV_X1 U159 ( .A(DATA2[15]), .ZN(n245) );
  INV_X1 U160 ( .A(DATA2[14]), .ZN(n246) );
  INV_X1 U161 ( .A(DATA2[13]), .ZN(n247) );
  INV_X1 U162 ( .A(DATA2[12]), .ZN(n248) );
  INV_X1 U163 ( .A(DATA2[11]), .ZN(n249) );
  INV_X1 U164 ( .A(DATA2[10]), .ZN(n250) );
  INV_X1 U165 ( .A(DATA2[9]), .ZN(n251) );
  INV_X1 U166 ( .A(DATA2[8]), .ZN(n252) );
  INV_X1 U167 ( .A(DATA2[7]), .ZN(n253) );
  INV_X1 U168 ( .A(DATA2[6]), .ZN(n254) );
  INV_X1 U169 ( .A(DATA2[5]), .ZN(n255) );
  OAI22_X1 U170 ( .A1(n83), .A2(n195), .B1(n84), .B2(n225), .ZN(OUT_ALU[3]) );
  OAI22_X1 U171 ( .A1(n89), .A2(n194), .B1(n90), .B2(n226), .ZN(OUT_ALU[2]) );
  OAI22_X1 U173 ( .A1(n111), .A2(n193), .B1(n112), .B2(n227), .ZN(OUT_ALU[1])
         );
  AOI211_X1 U174 ( .C1(n135), .C2(n136), .A(FUNC[3]), .B(FUNC[5]), .ZN(n71) );
  OR4_X1 U175 ( .A1(FUNC[2]), .A2(FUNC[1]), .A3(FUNC[0]), .A4(n257), .ZN(n135)
         );
  NAND4_X1 U176 ( .A1(n257), .A2(FUNC[0]), .A3(FUNC[1]), .A4(FUNC[2]), .ZN(
        n136) );
  INV_X1 U177 ( .A(FUNC[4]), .ZN(n257) );
  INV_X1 U178 ( .A(FUNC[0]), .ZN(n258) );
  AND3_X1 U179 ( .A1(FUNC[2]), .A2(FUNC[1]), .A3(n137), .ZN(n72) );
  AOI211_X1 U180 ( .C1(FUNC[3]), .C2(n258), .A(FUNC[5]), .B(FUNC[4]), .ZN(n137) );
  BUF_X1 U181 ( .A(n70), .Z(n185) );
  NOR4_X1 U182 ( .A1(n256), .A2(FUNC[1]), .A3(FUNC[2]), .A4(FUNC[5]), .ZN(n70)
         );
  INV_X1 U183 ( .A(n138), .ZN(n256) );
  OAI21_X1 U184 ( .B1(FUNC[3]), .B2(n257), .A(n139), .ZN(n138) );
  CLKBUF_X1 U185 ( .A(n185), .Z(n191) );
  INV_X1 U186 ( .A(DATA2[0]), .ZN(n192) );
  INV_X1 U187 ( .A(DATA2[1]), .ZN(n193) );
  INV_X1 U188 ( .A(DATA2[2]), .ZN(n194) );
  INV_X1 U189 ( .A(DATA2[3]), .ZN(n195) );
  INV_X1 U190 ( .A(DATA2[4]), .ZN(n196) );
endmodule


module comparator ( DATA1, DATA2i, .tipo({\tipo[5] , \tipo[4] , \tipo[3] , 
        \tipo[2] , \tipo[1] , \tipo[0] }), OUTALU );
  input [31:0] DATA1;
  output [31:0] OUTALU;
  input DATA2i, \tipo[5] , \tipo[4] , \tipo[3] , \tipo[2] , \tipo[1] ,
         \tipo[0] ;
  wire   N57, N58, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63;
  wire   [5:0] tipo;
  assign OUTALU[31] = 1'b0;
  assign OUTALU[30] = 1'b0;
  assign OUTALU[29] = 1'b0;
  assign OUTALU[28] = 1'b0;
  assign OUTALU[27] = 1'b0;
  assign OUTALU[26] = 1'b0;
  assign OUTALU[25] = 1'b0;
  assign OUTALU[24] = 1'b0;
  assign OUTALU[23] = 1'b0;
  assign OUTALU[22] = 1'b0;
  assign OUTALU[21] = 1'b0;
  assign OUTALU[20] = 1'b0;
  assign OUTALU[19] = 1'b0;
  assign OUTALU[18] = 1'b0;
  assign OUTALU[17] = 1'b0;
  assign OUTALU[16] = 1'b0;
  assign OUTALU[15] = 1'b0;
  assign OUTALU[14] = 1'b0;
  assign OUTALU[13] = 1'b0;
  assign OUTALU[12] = 1'b0;
  assign OUTALU[11] = 1'b0;
  assign OUTALU[10] = 1'b0;
  assign OUTALU[9] = 1'b0;
  assign OUTALU[8] = 1'b0;
  assign OUTALU[7] = 1'b0;
  assign OUTALU[6] = 1'b0;
  assign OUTALU[5] = 1'b0;
  assign OUTALU[4] = 1'b0;
  assign OUTALU[3] = 1'b0;
  assign OUTALU[2] = 1'b0;
  assign OUTALU[1] = 1'b0;

  DLH_X1 \OUTALU_reg[0]  ( .G(N57), .D(N58), .Q(OUTALU[0]) );
  NAND3_X1 U85 ( .A1(tipo[5]), .A2(n44), .A3(n45), .ZN(n43) );
  OR4_X1 U33 ( .A1(tipo[4]), .A2(n61), .A3(n62), .A4(n57), .ZN(n52) );
  INV_X1 U34 ( .A(n19), .ZN(n53) );
  NOR4_X1 U35 ( .A1(DATA1[23]), .A2(DATA1[22]), .A3(DATA1[21]), .A4(DATA1[20]), 
        .ZN(n27) );
  NOR4_X1 U36 ( .A1(DATA1[9]), .A2(DATA1[8]), .A3(DATA1[7]), .A4(DATA1[6]), 
        .ZN(n31) );
  NOR4_X1 U37 ( .A1(DATA1[16]), .A2(DATA1[15]), .A3(DATA1[14]), .A4(DATA1[13]), 
        .ZN(n25) );
  NOR2_X1 U38 ( .A1(n22), .A2(n23), .ZN(n19) );
  NAND4_X1 U39 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n22) );
  NAND4_X1 U40 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n23) );
  NOR4_X1 U41 ( .A1(DATA1[27]), .A2(DATA1[26]), .A3(DATA1[25]), .A4(DATA1[24]), 
        .ZN(n28) );
  INV_X1 U42 ( .A(DATA2i), .ZN(n54) );
  NOR4_X1 U43 ( .A1(DATA1[1]), .A2(DATA1[19]), .A3(DATA1[18]), .A4(DATA1[17]), 
        .ZN(n26) );
  NOR4_X1 U44 ( .A1(DATA1[5]), .A2(DATA1[4]), .A3(DATA1[3]), .A4(DATA1[31]), 
        .ZN(n30) );
  NOR4_X1 U45 ( .A1(DATA1[30]), .A2(DATA1[2]), .A3(DATA1[29]), .A4(DATA1[28]), 
        .ZN(n29) );
  NOR4_X1 U46 ( .A1(DATA1[12]), .A2(DATA1[11]), .A3(DATA1[10]), .A4(DATA1[0]), 
        .ZN(n24) );
  OAI221_X1 U47 ( .B1(n13), .B2(n54), .C1(n58), .C2(n53), .A(n14), .ZN(N58) );
  INV_X1 U48 ( .A(n20), .ZN(n58) );
  AOI21_X1 U49 ( .B1(n56), .B2(n53), .A(n21), .ZN(n13) );
  AOI22_X1 U50 ( .A1(n15), .A2(n55), .B1(n16), .B2(n54), .ZN(n14) );
  OAI21_X1 U51 ( .B1(n17), .B2(n63), .A(n18), .ZN(n16) );
  INV_X1 U52 ( .A(n34), .ZN(n55) );
  INV_X1 U53 ( .A(n32), .ZN(n56) );
  OR3_X1 U54 ( .A1(n20), .A2(n21), .A3(n33), .ZN(N57) );
  OAI211_X1 U55 ( .C1(n63), .C2(n17), .A(n34), .B(n32), .ZN(n33) );
  NOR4_X1 U56 ( .A1(n57), .A2(tipo[2]), .A3(tipo[3]), .A4(tipo[4]), .ZN(n35)
         );
  OAI221_X1 U57 ( .B1(tipo[5]), .B2(tipo[1]), .C1(tipo[4]), .C2(n62), .A(n51), 
        .ZN(n40) );
  AOI22_X1 U58 ( .A1(tipo[4]), .A2(n61), .B1(tipo[5]), .B2(tipo[2]), .ZN(n51)
         );
  OAI211_X1 U59 ( .C1(tipo[4]), .C2(tipo[3]), .A(n49), .B(n50), .ZN(n18) );
  AOI211_X1 U60 ( .C1(tipo[4]), .C2(n63), .A(tipo[5]), .B(n44), .ZN(n50) );
  AOI22_X1 U61 ( .A1(tipo[3]), .A2(n62), .B1(tipo[1]), .B2(tipo[2]), .ZN(n49)
         );
  INV_X1 U62 ( .A(tipo[1]), .ZN(n62) );
  INV_X1 U63 ( .A(tipo[2]), .ZN(n61) );
  NOR2_X1 U64 ( .A1(n63), .A2(tipo[2]), .ZN(n44) );
  INV_X1 U65 ( .A(tipo[5]), .ZN(n57) );
  INV_X1 U66 ( .A(tipo[4]), .ZN(n59) );
  INV_X1 U67 ( .A(tipo[0]), .ZN(n63) );
  AOI21_X1 U68 ( .B1(n62), .B2(n35), .A(n39), .ZN(n17) );
  AOI21_X1 U69 ( .B1(n52), .B2(n40), .A(n60), .ZN(n39) );
  INV_X1 U70 ( .A(tipo[3]), .ZN(n60) );
  OAI21_X1 U71 ( .B1(n40), .B2(n48), .A(n18), .ZN(n20) );
  NAND2_X1 U72 ( .A1(tipo[3]), .A2(n63), .ZN(n48) );
  NOR2_X1 U73 ( .A1(tipo[1]), .A2(n19), .ZN(n15) );
  OAI21_X1 U74 ( .B1(n35), .B2(n36), .A(n63), .ZN(n32) );
  AOI211_X1 U75 ( .C1(tipo[4]), .C2(n37), .A(n38), .B(tipo[2]), .ZN(n36) );
  OR2_X1 U76 ( .A1(tipo[3]), .A2(tipo[1]), .ZN(n37) );
  OAI21_X1 U77 ( .B1(tipo[4]), .B2(tipo[1]), .A(tipo[5]), .ZN(n38) );
  OAI21_X1 U78 ( .B1(n46), .B2(n47), .A(n57), .ZN(n34) );
  AND3_X1 U79 ( .A1(tipo[3]), .A2(n59), .A3(n44), .ZN(n47) );
  NOR4_X1 U80 ( .A1(tipo[3]), .A2(tipo[0]), .A3(n61), .A4(n59), .ZN(n46) );
  OAI21_X1 U81 ( .B1(n42), .B2(n62), .A(n43), .ZN(n21) );
  AOI21_X1 U82 ( .B1(n35), .B2(tipo[0]), .A(n55), .ZN(n42) );
  NOR3_X1 U83 ( .A1(n59), .A2(tipo[3]), .A3(tipo[1]), .ZN(n45) );
endmodule


module SHIFTER_GENERIC_N32_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[5][31] , \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] ,
         \ML_int[5][15] , \ML_int[5][14] , \ML_int[5][13] , \ML_int[5][12] ,
         \ML_int[5][11] , \ML_int[5][10] , \ML_int[5][9] , \ML_int[5][8] ,
         \ML_int[5][7] , \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] ,
         \ML_int[5][3] , \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;
  assign B[31] = \ML_int[5][31] ;
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[8] = \ML_int[5][8] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n34), .Z(
        \ML_int[5][31] ) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n34), .Z(
        \ML_int[5][30] ) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n34), .Z(
        \ML_int[5][29] ) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n34), .Z(
        \ML_int[5][28] ) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n34), .Z(
        \ML_int[5][27] ) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n34), .Z(
        \ML_int[5][26] ) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(SH[4]), .Z(
        \ML_int[5][25] ) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n34), .Z(
        \ML_int[5][24] ) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(n36), .S(SH[4]), .Z(
        \ML_int[5][23] ) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(n37), .S(n34), .Z(\ML_int[5][22] )
         );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(n38), .S(SH[4]), .Z(
        \ML_int[5][21] ) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(n39), .S(n34), .Z(\ML_int[5][20] )
         );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(n40), .S(SH[4]), .Z(
        \ML_int[5][19] ) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(n41), .S(SH[4]), .Z(
        \ML_int[5][18] ) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(n42), .S(SH[4]), .Z(
        \ML_int[5][17] ) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(n43), .S(SH[4]), .Z(
        \ML_int[5][16] ) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n32), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n32), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n32), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n32), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n32), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n32), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n32), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(SH[3]), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n32), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(SH[3]), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n32), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(SH[3]), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n32), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n32), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n32), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n32), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n32), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n32), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n32), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n32), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n32), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n32), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n32), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n32), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n30), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n29), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n30), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n29), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n30), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n29), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n30), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n30), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n30), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n30), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n30), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n30), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n30), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n30), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n30), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n30), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n30), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n29), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n29), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n29), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n29), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n29), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n29), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n29), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n29), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n29), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n29), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n29), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n27), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n26), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n27), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n26), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n27), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n26), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n27), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n26), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n27), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n27), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n27), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n27), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n27), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n27), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n27), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n27), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n27), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n27), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n27), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n26), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n26), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n26), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n26), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n26), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n26), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n26), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n26), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n26), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n26), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n26), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n24), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n23), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n24), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n23), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n24), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n23), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n24), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n23), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n24), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n24), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n24), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n24), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n24), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n24), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n24), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n24), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n24), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n24), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n24), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n24), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n23), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n23), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n23), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n23), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n23), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n23), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n23), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n23), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n23), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n23), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n23), .Z(\ML_int[1][1] ) );
  INV_X1 U3 ( .A(n15), .ZN(n36) );
  INV_X1 U4 ( .A(n16), .ZN(n37) );
  INV_X1 U5 ( .A(n17), .ZN(n38) );
  INV_X1 U6 ( .A(n18), .ZN(n39) );
  INV_X1 U7 ( .A(n19), .ZN(n40) );
  INV_X1 U8 ( .A(n20), .ZN(n41) );
  INV_X1 U9 ( .A(n21), .ZN(n42) );
  INV_X1 U10 ( .A(n22), .ZN(n43) );
  INV_X1 U11 ( .A(n33), .ZN(n32) );
  NAND2_X1 U12 ( .A1(\ML_int[3][7] ), .A2(n33), .ZN(n15) );
  NAND2_X1 U13 ( .A1(\ML_int[3][6] ), .A2(n33), .ZN(n16) );
  NAND2_X1 U14 ( .A1(\ML_int[3][5] ), .A2(n33), .ZN(n17) );
  NAND2_X1 U15 ( .A1(\ML_int[3][4] ), .A2(n33), .ZN(n18) );
  NAND2_X1 U16 ( .A1(\ML_int[3][3] ), .A2(n33), .ZN(n19) );
  NAND2_X1 U17 ( .A1(\ML_int[3][2] ), .A2(n33), .ZN(n20) );
  NAND2_X1 U18 ( .A1(\ML_int[3][1] ), .A2(n33), .ZN(n21) );
  NAND2_X1 U19 ( .A1(\ML_int[3][0] ), .A2(n33), .ZN(n22) );
  INV_X1 U20 ( .A(n25), .ZN(n24) );
  INV_X1 U21 ( .A(n25), .ZN(n23) );
  INV_X1 U22 ( .A(n28), .ZN(n27) );
  INV_X1 U23 ( .A(n28), .ZN(n26) );
  INV_X1 U24 ( .A(n31), .ZN(n30) );
  INV_X1 U25 ( .A(SH[4]), .ZN(n35) );
  AND2_X1 U26 ( .A1(\ML_int[2][3] ), .A2(n31), .ZN(\ML_int[3][3] ) );
  AND2_X1 U27 ( .A1(\ML_int[2][2] ), .A2(n31), .ZN(\ML_int[3][2] ) );
  AND2_X1 U28 ( .A1(\ML_int[2][1] ), .A2(n31), .ZN(\ML_int[3][1] ) );
  AND2_X1 U29 ( .A1(\ML_int[2][0] ), .A2(n31), .ZN(\ML_int[3][0] ) );
  AND2_X1 U30 ( .A1(\ML_int[4][15] ), .A2(n35), .ZN(\ML_int[5][15] ) );
  AND2_X1 U31 ( .A1(\ML_int[4][14] ), .A2(n35), .ZN(\ML_int[5][14] ) );
  AND2_X1 U32 ( .A1(\ML_int[4][13] ), .A2(n35), .ZN(\ML_int[5][13] ) );
  AND2_X1 U33 ( .A1(\ML_int[4][12] ), .A2(n35), .ZN(\ML_int[5][12] ) );
  AND2_X1 U34 ( .A1(\ML_int[4][11] ), .A2(n35), .ZN(\ML_int[5][11] ) );
  AND2_X1 U35 ( .A1(\ML_int[4][10] ), .A2(n35), .ZN(\ML_int[5][10] ) );
  NOR2_X1 U36 ( .A1(n34), .A2(n20), .ZN(\ML_int[5][2] ) );
  NOR2_X1 U37 ( .A1(n34), .A2(n21), .ZN(\ML_int[5][1] ) );
  NOR2_X1 U38 ( .A1(n34), .A2(n22), .ZN(\ML_int[5][0] ) );
  AND2_X1 U39 ( .A1(\ML_int[4][9] ), .A2(n35), .ZN(\ML_int[5][9] ) );
  AND2_X1 U40 ( .A1(\ML_int[4][8] ), .A2(n35), .ZN(\ML_int[5][8] ) );
  NOR2_X1 U41 ( .A1(n34), .A2(n15), .ZN(\ML_int[5][7] ) );
  NOR2_X1 U42 ( .A1(n34), .A2(n16), .ZN(\ML_int[5][6] ) );
  NOR2_X1 U43 ( .A1(n34), .A2(n17), .ZN(\ML_int[5][5] ) );
  NOR2_X1 U44 ( .A1(n34), .A2(n18), .ZN(\ML_int[5][4] ) );
  NOR2_X1 U45 ( .A1(n34), .A2(n19), .ZN(\ML_int[5][3] ) );
  INV_X1 U46 ( .A(SH[0]), .ZN(n25) );
  INV_X1 U47 ( .A(SH[1]), .ZN(n28) );
  INV_X1 U48 ( .A(SH[2]), .ZN(n31) );
  AND2_X1 U49 ( .A1(\ML_int[1][1] ), .A2(n28), .ZN(\ML_int[2][1] ) );
  AND2_X1 U50 ( .A1(\ML_int[1][0] ), .A2(n28), .ZN(\ML_int[2][0] ) );
  AND2_X1 U51 ( .A1(A[0]), .A2(n25), .ZN(\ML_int[1][0] ) );
  INV_X1 U52 ( .A(n31), .ZN(n29) );
  INV_X1 U53 ( .A(SH[3]), .ZN(n33) );
  INV_X1 U54 ( .A(n35), .ZN(n34) );
endmodule


module SHIFTER_GENERIC_N32_DW_sla_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[0] , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251;
  assign B[0] = \A[0] ;
  assign \A[0]  = A[0];

  NOR2_X2 U10 ( .A1(n189), .A2(SH[3]), .ZN(n114) );
  NOR2_X2 U12 ( .A1(SH[2]), .A2(SH[3]), .ZN(n116) );
  MUX2_X1 U181 ( .A(\A[0] ), .B(A[1]), .S(n178), .Z(n119) );
  NAND2_X1 U2 ( .A1(n196), .A2(\A[0] ), .ZN(n62) );
  INV_X1 U3 ( .A(n196), .ZN(n192) );
  INV_X1 U4 ( .A(n69), .ZN(n250) );
  NAND2_X1 U5 ( .A1(n114), .A2(n192), .ZN(n69) );
  INV_X1 U6 ( .A(n100), .ZN(n251) );
  BUF_X1 U7 ( .A(n190), .Z(n193) );
  BUF_X1 U8 ( .A(n191), .Z(n195) );
  BUF_X1 U9 ( .A(n190), .Z(n194) );
  BUF_X1 U11 ( .A(n191), .Z(n196) );
  NAND2_X1 U13 ( .A1(n116), .A2(n192), .ZN(n100) );
  AND2_X1 U14 ( .A1(n152), .A2(n189), .ZN(n75) );
  AND2_X1 U15 ( .A1(SH[3]), .A2(n189), .ZN(n118) );
  BUF_X1 U16 ( .A(n80), .Z(n180) );
  BUF_X1 U17 ( .A(n80), .Z(n179) );
  BUF_X1 U18 ( .A(n77), .Z(n186) );
  BUF_X1 U19 ( .A(n77), .Z(n185) );
  BUF_X1 U20 ( .A(n175), .Z(n177) );
  BUF_X1 U21 ( .A(n175), .Z(n176) );
  BUF_X1 U22 ( .A(n78), .Z(n182) );
  BUF_X1 U23 ( .A(n78), .Z(n183) );
  BUF_X1 U24 ( .A(n175), .Z(n178) );
  BUF_X1 U25 ( .A(n80), .Z(n181) );
  BUF_X1 U26 ( .A(n77), .Z(n187) );
  BUF_X1 U27 ( .A(n78), .Z(n184) );
  AND2_X1 U28 ( .A1(SH[3]), .A2(n192), .ZN(n152) );
  BUF_X1 U29 ( .A(SH[4]), .Z(n191) );
  BUF_X1 U30 ( .A(SH[4]), .Z(n190) );
  AND2_X1 U31 ( .A1(n152), .A2(SH[2]), .ZN(n72) );
  AOI221_X1 U32 ( .B1(n125), .B2(n114), .C1(n126), .C2(n116), .A(n249), .ZN(
        n63) );
  AOI221_X1 U33 ( .B1(n131), .B2(n114), .C1(n132), .C2(n116), .A(n249), .ZN(
        n64) );
  AOI221_X1 U34 ( .B1(n244), .B2(n114), .C1(n136), .C2(n116), .A(n249), .ZN(
        n65) );
  AOI221_X1 U35 ( .B1(n119), .B2(n114), .C1(n113), .C2(n116), .A(n249), .ZN(
        n66) );
  AOI221_X1 U36 ( .B1(n130), .B2(n114), .C1(n103), .C2(n116), .A(n234), .ZN(
        n70) );
  INV_X1 U37 ( .A(n154), .ZN(n234) );
  AOI22_X1 U38 ( .A1(n155), .A2(n131), .B1(n118), .B2(n132), .ZN(n154) );
  AOI221_X1 U39 ( .B1(n135), .B2(n114), .C1(n108), .C2(n116), .A(n236), .ZN(
        n81) );
  INV_X1 U40 ( .A(n157), .ZN(n236) );
  AOI22_X1 U41 ( .A1(n155), .A2(n244), .B1(n118), .B2(n136), .ZN(n157) );
  AOI221_X1 U42 ( .B1(n119), .B2(n155), .C1(n113), .C2(n118), .A(n226), .ZN(
        n88) );
  INV_X1 U43 ( .A(n159), .ZN(n226) );
  AOI22_X1 U44 ( .A1(n114), .A2(n115), .B1(n116), .B2(n112), .ZN(n159) );
  AOI221_X1 U45 ( .B1(n126), .B2(n114), .C1(n124), .C2(n116), .A(n239), .ZN(
        n94) );
  INV_X1 U46 ( .A(n163), .ZN(n239) );
  AOI21_X1 U47 ( .B1(n118), .B2(n125), .A(n120), .ZN(n163) );
  AOI221_X1 U48 ( .B1(n132), .B2(n114), .C1(n130), .C2(n116), .A(n241), .ZN(
        n101) );
  INV_X1 U49 ( .A(n167), .ZN(n241) );
  AOI21_X1 U50 ( .B1(n118), .B2(n131), .A(n120), .ZN(n167) );
  AOI221_X1 U51 ( .B1(n136), .B2(n114), .C1(n135), .C2(n116), .A(n243), .ZN(
        n106) );
  INV_X1 U52 ( .A(n171), .ZN(n243) );
  AOI21_X1 U53 ( .B1(n118), .B2(n244), .A(n120), .ZN(n171) );
  AOI221_X1 U54 ( .B1(n113), .B2(n114), .C1(n115), .C2(n116), .A(n246), .ZN(
        n61) );
  INV_X1 U55 ( .A(n117), .ZN(n246) );
  AOI21_X1 U56 ( .B1(n118), .B2(n119), .A(n120), .ZN(n117) );
  AOI222_X1 U57 ( .A1(n250), .A2(n76), .B1(n75), .B2(n73), .C1(n72), .C2(n103), 
        .ZN(n102) );
  AOI222_X1 U58 ( .A1(n250), .A2(n85), .B1(n75), .B2(n83), .C1(n72), .C2(n108), 
        .ZN(n107) );
  AOI222_X1 U59 ( .A1(n250), .A2(n92), .B1(n75), .B2(n90), .C1(n72), .C2(n112), 
        .ZN(n111) );
  AOI222_X1 U60 ( .A1(n250), .A2(n98), .B1(n75), .B2(n96), .C1(n72), .C2(n124), 
        .ZN(n123) );
  AOI222_X1 U61 ( .A1(n250), .A2(n73), .B1(n75), .B2(n103), .C1(n72), .C2(n130), .ZN(n129) );
  AOI222_X1 U62 ( .A1(n250), .A2(n83), .B1(n75), .B2(n108), .C1(n72), .C2(n135), .ZN(n134) );
  AOI222_X1 U63 ( .A1(n250), .A2(n90), .B1(n75), .B2(n112), .C1(n72), .C2(n115), .ZN(n138) );
  AOI222_X1 U64 ( .A1(n250), .A2(n96), .B1(n75), .B2(n124), .C1(n72), .C2(n126), .ZN(n141) );
  AOI222_X1 U65 ( .A1(n250), .A2(n103), .B1(n75), .B2(n130), .C1(n72), .C2(
        n132), .ZN(n145) );
  AOI222_X1 U66 ( .A1(n250), .A2(n108), .B1(n75), .B2(n135), .C1(n72), .C2(
        n136), .ZN(n147) );
  AOI222_X1 U67 ( .A1(n250), .A2(n112), .B1(n75), .B2(n115), .C1(n72), .C2(
        n113), .ZN(n149) );
  OAI221_X1 U68 ( .B1(n202), .B2(n69), .C1(n81), .C2(n192), .A(n82), .ZN(B[30]) );
  OAI221_X1 U69 ( .B1(n204), .B2(n69), .C1(n88), .C2(n192), .A(n89), .ZN(B[29]) );
  OAI221_X1 U70 ( .B1(n206), .B2(n69), .C1(n94), .C2(n192), .A(n95), .ZN(B[28]) );
  OAI221_X1 U71 ( .B1(n200), .B2(n100), .C1(n101), .C2(n192), .A(n102), .ZN(
        B[27]) );
  OAI221_X1 U72 ( .B1(n202), .B2(n100), .C1(n106), .C2(n192), .A(n107), .ZN(
        B[26]) );
  OAI221_X1 U73 ( .B1(n204), .B2(n100), .C1(n61), .C2(n192), .A(n111), .ZN(
        B[25]) );
  OAI221_X1 U74 ( .B1(n206), .B2(n100), .C1(n63), .C2(n192), .A(n123), .ZN(
        B[24]) );
  OAI221_X1 U75 ( .B1(n208), .B2(n100), .C1(n64), .C2(n192), .A(n129), .ZN(
        B[23]) );
  OAI221_X1 U76 ( .B1(n210), .B2(n100), .C1(n65), .C2(n192), .A(n134), .ZN(
        B[22]) );
  OAI221_X1 U77 ( .B1(n212), .B2(n100), .C1(n66), .C2(n192), .A(n138), .ZN(
        B[21]) );
  OAI221_X1 U78 ( .B1(n214), .B2(n100), .C1(n67), .C2(n192), .A(n141), .ZN(
        B[20]) );
  OAI221_X1 U79 ( .B1(n216), .B2(n100), .C1(n68), .C2(n192), .A(n145), .ZN(
        B[19]) );
  OAI221_X1 U80 ( .B1(n218), .B2(n100), .C1(n87), .C2(n192), .A(n147), .ZN(
        B[18]) );
  OAI221_X1 U81 ( .B1(n220), .B2(n100), .C1(n144), .C2(n192), .A(n149), .ZN(
        B[17]) );
  OAI221_X1 U82 ( .B1(n228), .B2(n69), .C1(n222), .C2(n100), .A(n151), .ZN(
        B[16]) );
  OAI21_X1 U83 ( .B1(n193), .B2(n70), .A(n62), .ZN(B[15]) );
  OAI21_X1 U84 ( .B1(n193), .B2(n81), .A(n62), .ZN(B[14]) );
  OAI21_X1 U85 ( .B1(n194), .B2(n88), .A(n62), .ZN(B[13]) );
  OAI21_X1 U86 ( .B1(n193), .B2(n94), .A(n62), .ZN(B[12]) );
  OAI21_X1 U87 ( .B1(n193), .B2(n101), .A(n62), .ZN(B[11]) );
  OAI21_X1 U88 ( .B1(n193), .B2(n106), .A(n62), .ZN(B[10]) );
  OAI21_X1 U89 ( .B1(n194), .B2(n87), .A(n62), .ZN(B[2]) );
  OAI21_X1 U90 ( .B1(n194), .B2(n144), .A(n62), .ZN(B[1]) );
  OAI21_X1 U91 ( .B1(n195), .B2(n61), .A(n62), .ZN(B[9]) );
  OAI21_X1 U92 ( .B1(n195), .B2(n63), .A(n62), .ZN(B[8]) );
  OAI21_X1 U93 ( .B1(n195), .B2(n64), .A(n62), .ZN(B[7]) );
  OAI21_X1 U94 ( .B1(n195), .B2(n65), .A(n62), .ZN(B[6]) );
  OAI21_X1 U95 ( .B1(n195), .B2(n66), .A(n62), .ZN(B[5]) );
  OAI21_X1 U96 ( .B1(n194), .B2(n67), .A(n62), .ZN(B[4]) );
  OAI21_X1 U97 ( .B1(n194), .B2(n68), .A(n62), .ZN(B[3]) );
  OAI21_X1 U98 ( .B1(n247), .B2(n189), .A(n139), .ZN(n142) );
  AOI221_X1 U99 ( .B1(n72), .B2(n125), .C1(n75), .C2(n126), .A(n248), .ZN(n151) );
  INV_X1 U100 ( .A(n62), .ZN(n248) );
  NOR2_X1 U101 ( .A1(n189), .A2(n139), .ZN(n120) );
  AOI21_X1 U102 ( .B1(n125), .B2(n116), .A(n142), .ZN(n67) );
  AOI21_X1 U103 ( .B1(n131), .B2(n116), .A(n142), .ZN(n68) );
  AOI21_X1 U104 ( .B1(n244), .B2(n116), .A(n142), .ZN(n87) );
  AOI21_X1 U105 ( .B1(n119), .B2(n116), .A(n142), .ZN(n144) );
  NAND2_X1 U106 ( .A1(SH[0]), .A2(SH[1]), .ZN(n78) );
  NAND2_X1 U107 ( .A1(SH[1]), .A2(n188), .ZN(n77) );
  INV_X1 U108 ( .A(n139), .ZN(n249) );
  NOR2_X1 U109 ( .A1(n188), .A2(SH[1]), .ZN(n80) );
  AND2_X1 U110 ( .A1(SH[2]), .A2(SH[3]), .ZN(n155) );
  INV_X1 U111 ( .A(n124), .ZN(n228) );
  INV_X1 U112 ( .A(n73), .ZN(n216) );
  INV_X1 U113 ( .A(n83), .ZN(n218) );
  INV_X1 U114 ( .A(n90), .ZN(n220) );
  INV_X1 U115 ( .A(n96), .ZN(n222) );
  NOR2_X1 U116 ( .A1(SH[0]), .A2(SH[1]), .ZN(n175) );
  INV_X1 U117 ( .A(n76), .ZN(n208) );
  INV_X1 U118 ( .A(n85), .ZN(n210) );
  INV_X1 U119 ( .A(n92), .ZN(n212) );
  INV_X1 U120 ( .A(n98), .ZN(n214) );
  OAI221_X1 U121 ( .B1(n185), .B2(n229), .C1(n182), .C2(n230), .A(n160), .ZN(
        n112) );
  AOI22_X1 U122 ( .A1(A[12]), .A2(n179), .B1(A[13]), .B2(n176), .ZN(n160) );
  OAI221_X1 U123 ( .B1(n185), .B2(n233), .C1(n182), .C2(n235), .A(n161), .ZN(
        n115) );
  AOI22_X1 U124 ( .A1(A[8]), .A2(n179), .B1(A[9]), .B2(n176), .ZN(n161) );
  OAI221_X1 U125 ( .B1(n245), .B2(n187), .C1(n247), .C2(n182), .A(n168), .ZN(
        n131) );
  AOI22_X1 U126 ( .A1(n181), .A2(A[2]), .B1(A[3]), .B2(n176), .ZN(n168) );
  OAI221_X1 U127 ( .B1(n187), .B2(n235), .C1(n184), .C2(n237), .A(n166), .ZN(
        n126) );
  AOI22_X1 U128 ( .A1(A[7]), .A2(n179), .B1(A[8]), .B2(n176), .ZN(n166) );
  OAI221_X1 U129 ( .B1(n187), .B2(n237), .C1(n184), .C2(n238), .A(n170), .ZN(
        n132) );
  AOI22_X1 U130 ( .A1(A[6]), .A2(n179), .B1(A[7]), .B2(n176), .ZN(n170) );
  OAI221_X1 U131 ( .B1(n186), .B2(n238), .C1(n240), .C2(n182), .A(n174), .ZN(
        n136) );
  AOI22_X1 U132 ( .A1(A[5]), .A2(n180), .B1(A[6]), .B2(n176), .ZN(n174) );
  OAI221_X1 U133 ( .B1(n185), .B2(n230), .C1(n184), .C2(n231), .A(n165), .ZN(
        n124) );
  AOI22_X1 U134 ( .A1(A[11]), .A2(n179), .B1(A[12]), .B2(n176), .ZN(n165) );
  OAI221_X1 U135 ( .B1(n187), .B2(n231), .C1(n184), .C2(n232), .A(n169), .ZN(
        n130) );
  AOI22_X1 U136 ( .A1(A[10]), .A2(n179), .B1(A[11]), .B2(n176), .ZN(n169) );
  OAI221_X1 U137 ( .B1(n187), .B2(n232), .C1(n184), .C2(n233), .A(n173), .ZN(
        n135) );
  AOI22_X1 U138 ( .A1(A[9]), .A2(n179), .B1(A[10]), .B2(n176), .ZN(n173) );
  OAI221_X1 U139 ( .B1(n185), .B2(n219), .C1(n182), .C2(n221), .A(n146), .ZN(
        n73) );
  AOI22_X1 U140 ( .A1(A[18]), .A2(n180), .B1(A[19]), .B2(n177), .ZN(n146) );
  OAI221_X1 U141 ( .B1(n185), .B2(n221), .C1(n182), .C2(n223), .A(n148), .ZN(
        n83) );
  AOI22_X1 U142 ( .A1(A[17]), .A2(n180), .B1(A[18]), .B2(n177), .ZN(n148) );
  OAI221_X1 U143 ( .B1(n185), .B2(n223), .C1(n182), .C2(n224), .A(n150), .ZN(
        n90) );
  AOI22_X1 U144 ( .A1(A[16]), .A2(n180), .B1(A[17]), .B2(n177), .ZN(n150) );
  OAI221_X1 U145 ( .B1(n185), .B2(n224), .C1(n182), .C2(n225), .A(n153), .ZN(
        n96) );
  AOI22_X1 U146 ( .A1(A[15]), .A2(n179), .B1(A[16]), .B2(n177), .ZN(n153) );
  OAI221_X1 U147 ( .B1(n185), .B2(n225), .C1(n182), .C2(n227), .A(n156), .ZN(
        n103) );
  AOI22_X1 U148 ( .A1(A[14]), .A2(n179), .B1(A[15]), .B2(n177), .ZN(n156) );
  OAI221_X1 U149 ( .B1(n185), .B2(n227), .C1(n182), .C2(n229), .A(n158), .ZN(
        n108) );
  AOI22_X1 U150 ( .A1(A[13]), .A2(n179), .B1(A[14]), .B2(n176), .ZN(n158) );
  OAI221_X1 U151 ( .B1(n185), .B2(n242), .C1(n245), .C2(n182), .A(n164), .ZN(
        n125) );
  AOI22_X1 U152 ( .A1(n181), .A2(A[3]), .B1(A[4]), .B2(n176), .ZN(n164) );
  OAI221_X1 U153 ( .B1(n185), .B2(n240), .C1(n182), .C2(n242), .A(n162), .ZN(
        n113) );
  AOI22_X1 U154 ( .A1(A[4]), .A2(n179), .B1(A[5]), .B2(n176), .ZN(n162) );
  OAI221_X1 U155 ( .B1(n186), .B2(n211), .C1(n183), .C2(n213), .A(n133), .ZN(
        n76) );
  AOI22_X1 U156 ( .A1(A[22]), .A2(n180), .B1(A[23]), .B2(n177), .ZN(n133) );
  OAI221_X1 U157 ( .B1(n186), .B2(n213), .C1(n183), .C2(n215), .A(n137), .ZN(
        n85) );
  AOI22_X1 U158 ( .A1(A[21]), .A2(n180), .B1(A[22]), .B2(n177), .ZN(n137) );
  OAI221_X1 U159 ( .B1(n186), .B2(n215), .C1(n183), .C2(n217), .A(n140), .ZN(
        n92) );
  AOI22_X1 U160 ( .A1(A[20]), .A2(n180), .B1(A[21]), .B2(n177), .ZN(n140) );
  OAI221_X1 U161 ( .B1(n185), .B2(n217), .C1(n183), .C2(n219), .A(n143), .ZN(
        n98) );
  AOI22_X1 U162 ( .A1(A[19]), .A2(n180), .B1(A[20]), .B2(n177), .ZN(n143) );
  AOI222_X1 U163 ( .A1(n72), .A2(n83), .B1(n251), .B2(n84), .C1(n75), .C2(n85), 
        .ZN(n82) );
  OAI221_X1 U164 ( .B1(n186), .B2(n198), .C1(n183), .C2(n199), .A(n86), .ZN(
        n84) );
  AOI22_X1 U165 ( .A1(A[29]), .A2(n181), .B1(A[30]), .B2(n178), .ZN(n86) );
  AOI222_X1 U166 ( .A1(n72), .A2(n90), .B1(n251), .B2(n91), .C1(n75), .C2(n92), 
        .ZN(n89) );
  OAI221_X1 U167 ( .B1(n186), .B2(n199), .C1(n183), .C2(n201), .A(n93), .ZN(
        n91) );
  AOI22_X1 U168 ( .A1(A[28]), .A2(n181), .B1(A[29]), .B2(n178), .ZN(n93) );
  AOI222_X1 U169 ( .A1(n72), .A2(n96), .B1(n251), .B2(n97), .C1(n75), .C2(n98), 
        .ZN(n95) );
  OAI221_X1 U170 ( .B1(n186), .B2(n201), .C1(n183), .C2(n203), .A(n99), .ZN(
        n97) );
  AOI22_X1 U171 ( .A1(A[27]), .A2(n181), .B1(A[28]), .B2(n178), .ZN(n99) );
  OAI221_X1 U172 ( .B1(n200), .B2(n69), .C1(n70), .C2(n192), .A(n71), .ZN(
        B[31]) );
  AOI222_X1 U173 ( .A1(n72), .A2(n73), .B1(n251), .B2(n74), .C1(n75), .C2(n76), 
        .ZN(n71) );
  OAI221_X1 U174 ( .B1(n186), .B2(n197), .C1(n183), .C2(n198), .A(n79), .ZN(
        n74) );
  INV_X1 U175 ( .A(A[29]), .ZN(n197) );
  AOI22_X1 U176 ( .A1(A[30]), .A2(n179), .B1(A[31]), .B2(n177), .ZN(n79) );
  NAND2_X1 U177 ( .A1(SH[3]), .A2(\A[0] ), .ZN(n139) );
  INV_X1 U178 ( .A(n172), .ZN(n244) );
  AOI222_X1 U179 ( .A1(n178), .A2(A[2]), .B1(A[1]), .B2(n181), .C1(\A[0] ), 
        .C2(SH[1]), .ZN(n172) );
  INV_X1 U180 ( .A(A[12]), .ZN(n227) );
  INV_X1 U182 ( .A(A[13]), .ZN(n225) );
  INV_X1 U183 ( .A(A[14]), .ZN(n224) );
  INV_X1 U184 ( .A(A[23]), .ZN(n207) );
  INV_X1 U185 ( .A(A[22]), .ZN(n209) );
  INV_X1 U186 ( .A(A[17]), .ZN(n219) );
  INV_X1 U187 ( .A(A[16]), .ZN(n221) );
  INV_X1 U188 ( .A(A[15]), .ZN(n223) );
  INV_X1 U189 ( .A(A[21]), .ZN(n211) );
  INV_X1 U190 ( .A(A[9]), .ZN(n231) );
  INV_X1 U191 ( .A(A[11]), .ZN(n229) );
  INV_X1 U192 ( .A(A[10]), .ZN(n230) );
  INV_X1 U193 ( .A(A[8]), .ZN(n232) );
  INV_X1 U194 ( .A(A[7]), .ZN(n233) );
  INV_X1 U195 ( .A(A[2]), .ZN(n242) );
  INV_X1 U196 ( .A(A[28]), .ZN(n198) );
  INV_X1 U197 ( .A(A[27]), .ZN(n199) );
  INV_X1 U198 ( .A(A[26]), .ZN(n201) );
  INV_X1 U199 ( .A(A[25]), .ZN(n203) );
  INV_X1 U200 ( .A(A[24]), .ZN(n205) );
  INV_X1 U201 ( .A(A[3]), .ZN(n240) );
  INV_X1 U202 ( .A(A[18]), .ZN(n217) );
  INV_X1 U203 ( .A(\A[0] ), .ZN(n247) );
  INV_X1 U204 ( .A(A[6]), .ZN(n235) );
  INV_X1 U205 ( .A(A[4]), .ZN(n238) );
  INV_X1 U206 ( .A(A[1]), .ZN(n245) );
  INV_X1 U207 ( .A(A[19]), .ZN(n215) );
  INV_X1 U208 ( .A(A[20]), .ZN(n213) );
  INV_X1 U209 ( .A(A[5]), .ZN(n237) );
  INV_X1 U210 ( .A(n127), .ZN(n206) );
  OAI221_X1 U211 ( .B1(n186), .B2(n209), .C1(n183), .C2(n211), .A(n128), .ZN(
        n127) );
  AOI22_X1 U212 ( .A1(A[23]), .A2(n180), .B1(A[24]), .B2(n177), .ZN(n128) );
  INV_X1 U213 ( .A(n104), .ZN(n200) );
  OAI221_X1 U214 ( .B1(n186), .B2(n203), .C1(n183), .C2(n205), .A(n105), .ZN(
        n104) );
  AOI22_X1 U215 ( .A1(A[26]), .A2(n180), .B1(A[27]), .B2(n178), .ZN(n105) );
  INV_X1 U216 ( .A(n109), .ZN(n202) );
  OAI221_X1 U217 ( .B1(n186), .B2(n205), .C1(n183), .C2(n207), .A(n110), .ZN(
        n109) );
  AOI22_X1 U218 ( .A1(A[25]), .A2(n180), .B1(A[26]), .B2(n178), .ZN(n110) );
  INV_X1 U219 ( .A(n121), .ZN(n204) );
  OAI221_X1 U220 ( .B1(n186), .B2(n207), .C1(n183), .C2(n209), .A(n122), .ZN(
        n121) );
  AOI22_X1 U221 ( .A1(A[24]), .A2(n180), .B1(A[25]), .B2(n177), .ZN(n122) );
  INV_X1 U222 ( .A(SH[0]), .ZN(n188) );
  INV_X1 U223 ( .A(SH[2]), .ZN(n189) );
endmodule


module SHIFTER_GENERIC_N32_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228;

  NOR2_X2 U3 ( .A1(SH[0]), .A2(SH[1]), .ZN(n96) );
  NOR2_X2 U5 ( .A1(n167), .A2(SH[1]), .ZN(n95) );
  MUX2_X1 U141 ( .A(n112), .B(n98), .S(SH[2]), .Z(n123) );
  INV_X1 U4 ( .A(n57), .ZN(n223) );
  NAND2_X1 U6 ( .A1(n224), .A2(n177), .ZN(n57) );
  INV_X1 U7 ( .A(n174), .ZN(n177) );
  INV_X1 U8 ( .A(n87), .ZN(n222) );
  NAND2_X1 U9 ( .A1(n110), .A2(n177), .ZN(n87) );
  NOR2_X1 U10 ( .A1(n177), .A2(n138), .ZN(n129) );
  INV_X1 U11 ( .A(n138), .ZN(n224) );
  NOR2_X1 U12 ( .A1(n170), .A2(n171), .ZN(n155) );
  BUF_X1 U13 ( .A(n176), .Z(n171) );
  BUF_X1 U14 ( .A(n175), .Z(n173) );
  BUF_X1 U15 ( .A(n176), .Z(n172) );
  BUF_X1 U16 ( .A(n175), .Z(n174) );
  INV_X1 U17 ( .A(n96), .ZN(n227) );
  INV_X1 U18 ( .A(n95), .ZN(n228) );
  NOR2_X2 U19 ( .A1(n168), .A2(n169), .ZN(n110) );
  INV_X1 U20 ( .A(n92), .ZN(n226) );
  INV_X1 U21 ( .A(n93), .ZN(n225) );
  AND2_X1 U22 ( .A1(n155), .A2(n168), .ZN(n61) );
  NOR2_X1 U23 ( .A1(n168), .A2(n170), .ZN(n125) );
  INV_X1 U24 ( .A(SH[3]), .ZN(n170) );
  NAND2_X1 U25 ( .A1(n168), .A2(n170), .ZN(n138) );
  BUF_X1 U26 ( .A(n93), .Z(n164) );
  BUF_X1 U27 ( .A(n93), .Z(n165) );
  BUF_X1 U28 ( .A(n93), .Z(n166) );
  INV_X1 U29 ( .A(n123), .ZN(n182) );
  BUF_X1 U30 ( .A(SH[4]), .Z(n175) );
  BUF_X1 U31 ( .A(SH[4]), .Z(n176) );
  NAND2_X1 U32 ( .A1(SH[1]), .A2(SH[0]), .ZN(n92) );
  OAI222_X1 U33 ( .A1(n228), .A2(n185), .B1(n164), .B2(n184), .C1(n227), .C2(
        n186), .ZN(n106) );
  AND2_X1 U34 ( .A1(SH[2]), .A2(n155), .ZN(n63) );
  NOR2_X1 U35 ( .A1(n170), .A2(SH[2]), .ZN(n113) );
  OAI22_X1 U36 ( .A1(n227), .A2(n185), .B1(n228), .B2(n184), .ZN(n99) );
  AOI222_X1 U37 ( .A1(n112), .A2(n110), .B1(n98), .B2(n113), .C1(n114), .C2(
        n224), .ZN(n72) );
  AOI222_X1 U38 ( .A1(n115), .A2(n110), .B1(n99), .B2(n113), .C1(n116), .C2(
        n224), .ZN(n77) );
  AOI222_X1 U39 ( .A1(n109), .A2(n110), .B1(n106), .B2(n113), .C1(n64), .C2(
        n224), .ZN(n82) );
  AOI222_X1 U40 ( .A1(n111), .A2(n110), .B1(n107), .B2(n113), .C1(n70), .C2(
        n224), .ZN(n85) );
  AOI222_X1 U41 ( .A1(n75), .A2(n224), .B1(n114), .B2(n110), .C1(n123), .C2(
        n169), .ZN(n88) );
  AOI221_X1 U42 ( .B1(n116), .B2(n110), .C1(n80), .C2(n224), .A(n181), .ZN(
        n100) );
  INV_X1 U43 ( .A(n124), .ZN(n181) );
  AOI22_X1 U44 ( .A1(n125), .A2(n99), .B1(n113), .B2(n115), .ZN(n124) );
  AOI221_X1 U45 ( .B1(n64), .B2(n110), .C1(n62), .C2(n224), .A(n183), .ZN(n117) );
  INV_X1 U46 ( .A(n126), .ZN(n183) );
  AOI22_X1 U47 ( .A1(n125), .A2(n106), .B1(n113), .B2(n109), .ZN(n126) );
  AOI221_X1 U48 ( .B1(n70), .B2(n110), .C1(n69), .C2(n224), .A(n180), .ZN(n127) );
  INV_X1 U49 ( .A(n158), .ZN(n180) );
  AOI22_X1 U50 ( .A1(n125), .A2(n107), .B1(n113), .B2(n111), .ZN(n158) );
  AOI222_X1 U51 ( .A1(n63), .A2(n109), .B1(n129), .B2(n106), .C1(n61), .C2(n64), .ZN(n131) );
  AOI222_X1 U52 ( .A1(n222), .A2(n79), .B1(n61), .B2(n80), .C1(n63), .C2(n116), 
        .ZN(n146) );
  AOI222_X1 U53 ( .A1(n222), .A2(n60), .B1(n61), .B2(n62), .C1(n63), .C2(n64), 
        .ZN(n59) );
  AOI222_X1 U54 ( .A1(n222), .A2(n68), .B1(n61), .B2(n69), .C1(n63), .C2(n70), 
        .ZN(n67) );
  AOI222_X1 U55 ( .A1(n222), .A2(n208), .B1(n61), .B2(n79), .C1(n63), .C2(n80), 
        .ZN(n78) );
  AOI222_X1 U56 ( .A1(n222), .A2(n210), .B1(n61), .B2(n60), .C1(n63), .C2(n62), 
        .ZN(n83) );
  AOI222_X1 U57 ( .A1(n222), .A2(n212), .B1(n61), .B2(n68), .C1(n63), .C2(n69), 
        .ZN(n86) );
  AOI222_X1 U58 ( .A1(n63), .A2(n115), .B1(n129), .B2(n99), .C1(n61), .C2(n116), .ZN(n130) );
  AOI222_X1 U59 ( .A1(n222), .A2(n207), .B1(n61), .B2(n74), .C1(n63), .C2(n75), 
        .ZN(n73) );
  AOI222_X1 U60 ( .A1(n63), .A2(n112), .B1(n129), .B2(n98), .C1(n61), .C2(n114), .ZN(n128) );
  AND2_X1 U61 ( .A1(n99), .A2(n223), .ZN(B[30]) );
  AND2_X1 U62 ( .A1(n106), .A2(n223), .ZN(B[29]) );
  AND2_X1 U63 ( .A1(n107), .A2(n223), .ZN(B[28]) );
  NOR3_X1 U64 ( .A1(n182), .A2(n171), .A3(n169), .ZN(B[27]) );
  NOR2_X1 U65 ( .A1(n171), .A2(n108), .ZN(B[26]) );
  NOR2_X1 U66 ( .A1(n172), .A2(n58), .ZN(B[25]) );
  NOR2_X1 U67 ( .A1(n172), .A2(n66), .ZN(B[24]) );
  NOR2_X1 U68 ( .A1(n172), .A2(n72), .ZN(B[23]) );
  NOR2_X1 U69 ( .A1(n173), .A2(n77), .ZN(B[22]) );
  NOR2_X1 U70 ( .A1(n173), .A2(n82), .ZN(B[21]) );
  NOR2_X1 U71 ( .A1(n173), .A2(n85), .ZN(B[20]) );
  NOR2_X1 U72 ( .A1(n173), .A2(n88), .ZN(B[19]) );
  NOR2_X1 U73 ( .A1(n174), .A2(n100), .ZN(B[18]) );
  NOR2_X1 U74 ( .A1(n172), .A2(n117), .ZN(B[17]) );
  NOR2_X1 U75 ( .A1(n171), .A2(n127), .ZN(B[16]) );
  OAI221_X1 U76 ( .B1(n193), .B2(n87), .C1(n199), .C2(n57), .A(n128), .ZN(
        B[15]) );
  OAI221_X1 U77 ( .B1(n194), .B2(n87), .C1(n201), .C2(n57), .A(n130), .ZN(
        B[14]) );
  OAI221_X1 U78 ( .B1(n196), .B2(n87), .C1(n203), .C2(n57), .A(n131), .ZN(
        B[13]) );
  INV_X1 U79 ( .A(n136), .ZN(B[12]) );
  OAI221_X1 U80 ( .B1(n199), .B2(n87), .C1(n91), .C2(n57), .A(n139), .ZN(B[11]) );
  OAI221_X1 U81 ( .B1(n103), .B2(n57), .C1(n108), .C2(n177), .A(n146), .ZN(
        B[10]) );
  OAI221_X1 U82 ( .B1(n76), .B2(n87), .C1(n100), .C2(n177), .A(n101), .ZN(B[2]) );
  OAI221_X1 U83 ( .B1(n81), .B2(n87), .C1(n117), .C2(n177), .A(n118), .ZN(B[1]) );
  OAI221_X1 U84 ( .B1(n56), .B2(n57), .C1(n58), .C2(n177), .A(n59), .ZN(B[9])
         );
  OAI221_X1 U85 ( .B1(n65), .B2(n57), .C1(n66), .C2(n177), .A(n67), .ZN(B[8])
         );
  OAI221_X1 U86 ( .B1(n71), .B2(n57), .C1(n72), .C2(n177), .A(n73), .ZN(B[7])
         );
  OAI221_X1 U87 ( .B1(n76), .B2(n57), .C1(n77), .C2(n177), .A(n78), .ZN(B[6])
         );
  OAI221_X1 U88 ( .B1(n81), .B2(n57), .C1(n82), .C2(n177), .A(n83), .ZN(B[5])
         );
  OAI221_X1 U89 ( .B1(n84), .B2(n57), .C1(n85), .C2(n177), .A(n86), .ZN(B[4])
         );
  OAI221_X1 U90 ( .B1(n71), .B2(n87), .C1(n88), .C2(n177), .A(n89), .ZN(B[3])
         );
  AOI221_X1 U91 ( .B1(n63), .B2(n114), .C1(n61), .C2(n75), .A(n140), .ZN(n139)
         );
  NOR3_X1 U92 ( .A1(n177), .A2(n169), .A3(n182), .ZN(n140) );
  AOI221_X1 U93 ( .B1(n69), .B2(n222), .C1(n68), .C2(n223), .A(n179), .ZN(n136) );
  INV_X1 U94 ( .A(n137), .ZN(n179) );
  AOI222_X1 U95 ( .A1(n63), .A2(n111), .B1(n129), .B2(n107), .C1(n61), .C2(n70), .ZN(n137) );
  NOR2_X1 U96 ( .A1(n184), .A2(n227), .ZN(n98) );
  AOI22_X1 U97 ( .A1(n115), .A2(n224), .B1(n99), .B2(n110), .ZN(n108) );
  AOI22_X1 U98 ( .A1(n109), .A2(n224), .B1(n106), .B2(n110), .ZN(n58) );
  AOI22_X1 U99 ( .A1(n111), .A2(n224), .B1(n107), .B2(n110), .ZN(n66) );
  NAND2_X1 U100 ( .A1(SH[1]), .A2(n167), .ZN(n93) );
  INV_X1 U101 ( .A(n74), .ZN(n199) );
  INV_X1 U102 ( .A(n103), .ZN(n208) );
  INV_X1 U103 ( .A(n56), .ZN(n210) );
  INV_X1 U104 ( .A(n65), .ZN(n212) );
  INV_X1 U105 ( .A(n91), .ZN(n207) );
  INV_X1 U106 ( .A(n80), .ZN(n194) );
  INV_X1 U107 ( .A(n62), .ZN(n196) );
  INV_X1 U108 ( .A(n75), .ZN(n193) );
  INV_X1 U109 ( .A(n79), .ZN(n201) );
  INV_X1 U110 ( .A(n60), .ZN(n203) );
  OAI221_X1 U111 ( .B1(n92), .B2(n184), .C1(n165), .C2(n185), .A(n160), .ZN(
        n107) );
  AOI22_X1 U112 ( .A1(A[29]), .A2(n95), .B1(A[28]), .B2(n96), .ZN(n160) );
  OAI221_X1 U113 ( .B1(n92), .B2(n195), .C1(n197), .C2(n165), .A(n148), .ZN(
        n80) );
  AOI22_X1 U114 ( .A1(n95), .A2(A[19]), .B1(n96), .B2(A[18]), .ZN(n148) );
  OAI221_X1 U115 ( .B1(n92), .B2(n197), .C1(n165), .C2(n198), .A(n135), .ZN(
        n62) );
  AOI22_X1 U116 ( .A1(A[18]), .A2(n95), .B1(A[17]), .B2(n96), .ZN(n135) );
  OAI221_X1 U117 ( .B1(n92), .B2(n198), .C1(n165), .C2(n200), .A(n161), .ZN(
        n69) );
  AOI22_X1 U118 ( .A1(A[17]), .A2(n95), .B1(A[16]), .B2(n96), .ZN(n161) );
  OAI221_X1 U119 ( .B1(n92), .B2(n202), .C1(n166), .C2(n204), .A(n149), .ZN(
        n79) );
  AOI22_X1 U120 ( .A1(A[15]), .A2(n95), .B1(A[14]), .B2(n96), .ZN(n149) );
  OAI221_X1 U121 ( .B1(n92), .B2(n204), .C1(n164), .C2(n205), .A(n134), .ZN(
        n60) );
  AOI22_X1 U122 ( .A1(A[14]), .A2(n95), .B1(A[13]), .B2(n96), .ZN(n134) );
  OAI221_X1 U123 ( .B1(n92), .B2(n205), .C1(n164), .C2(n206), .A(n157), .ZN(
        n68) );
  INV_X1 U124 ( .A(A[14]), .ZN(n206) );
  AOI22_X1 U125 ( .A1(A[13]), .A2(n95), .B1(A[12]), .B2(n96), .ZN(n157) );
  OAI221_X1 U126 ( .B1(n92), .B2(n186), .C1(n164), .C2(n187), .A(n150), .ZN(
        n115) );
  AOI22_X1 U127 ( .A1(A[27]), .A2(n95), .B1(A[26]), .B2(n96), .ZN(n150) );
  OAI221_X1 U128 ( .B1(n92), .B2(n187), .C1(n164), .C2(n188), .A(n133), .ZN(
        n109) );
  AOI22_X1 U129 ( .A1(A[26]), .A2(n95), .B1(A[25]), .B2(n96), .ZN(n133) );
  OAI221_X1 U130 ( .B1(n92), .B2(n188), .C1(n165), .C2(n189), .A(n159), .ZN(
        n111) );
  AOI22_X1 U131 ( .A1(A[25]), .A2(n95), .B1(A[24]), .B2(n96), .ZN(n159) );
  OAI221_X1 U132 ( .B1(n92), .B2(n190), .C1(n166), .C2(n191), .A(n147), .ZN(
        n116) );
  AOI22_X1 U133 ( .A1(A[23]), .A2(n95), .B1(A[22]), .B2(n96), .ZN(n147) );
  OAI221_X1 U134 ( .B1(n92), .B2(n191), .C1(n164), .C2(n192), .A(n132), .ZN(
        n64) );
  INV_X1 U135 ( .A(A[23]), .ZN(n192) );
  AOI22_X1 U136 ( .A1(A[22]), .A2(n95), .B1(A[21]), .B2(n96), .ZN(n132) );
  OAI221_X1 U137 ( .B1(n92), .B2(n189), .C1(n165), .C2(n190), .A(n143), .ZN(
        n114) );
  AOI22_X1 U138 ( .A1(A[24]), .A2(n95), .B1(A[23]), .B2(n96), .ZN(n143) );
  OAI221_X1 U139 ( .B1(n197), .B2(n228), .C1(n198), .C2(n227), .A(n142), .ZN(
        n75) );
  AOI22_X1 U140 ( .A1(A[22]), .A2(n226), .B1(A[21]), .B2(n225), .ZN(n142) );
  OAI221_X1 U142 ( .B1(n228), .B2(n195), .C1(n197), .C2(n227), .A(n162), .ZN(
        n70) );
  AOI22_X1 U143 ( .A1(A[23]), .A2(n226), .B1(A[22]), .B2(n225), .ZN(n162) );
  OAI221_X1 U144 ( .B1(n92), .B2(n200), .C1(n166), .C2(n202), .A(n145), .ZN(
        n74) );
  AOI22_X1 U145 ( .A1(A[16]), .A2(n95), .B1(A[15]), .B2(n96), .ZN(n145) );
  AOI221_X1 U146 ( .B1(n226), .B2(A[10]), .C1(n225), .C2(A[9]), .A(n97), .ZN(
        n71) );
  OAI22_X1 U147 ( .A1(n215), .A2(n228), .B1(n216), .B2(n227), .ZN(n97) );
  AOI221_X1 U148 ( .B1(n226), .B2(A[9]), .C1(n225), .C2(A[8]), .A(n105), .ZN(
        n76) );
  OAI22_X1 U149 ( .A1(n216), .A2(n228), .B1(n217), .B2(n227), .ZN(n105) );
  AOI221_X1 U150 ( .B1(n226), .B2(A[8]), .C1(n225), .C2(A[7]), .A(n122), .ZN(
        n81) );
  OAI22_X1 U151 ( .A1(n217), .A2(n228), .B1(n218), .B2(n227), .ZN(n122) );
  AOI221_X1 U152 ( .B1(n226), .B2(A[7]), .C1(n225), .C2(A[6]), .A(n163), .ZN(
        n84) );
  OAI22_X1 U153 ( .A1(n218), .A2(n228), .B1(n219), .B2(n227), .ZN(n163) );
  AOI221_X1 U154 ( .B1(n226), .B2(A[13]), .C1(n225), .C2(A[12]), .A(n151), 
        .ZN(n103) );
  OAI22_X1 U155 ( .A1(n211), .A2(n228), .B1(n213), .B2(n227), .ZN(n151) );
  AOI221_X1 U156 ( .B1(n226), .B2(A[12]), .C1(n225), .C2(A[11]), .A(n120), 
        .ZN(n56) );
  OAI22_X1 U157 ( .A1(n213), .A2(n228), .B1(n214), .B2(n227), .ZN(n120) );
  AOI221_X1 U158 ( .B1(n226), .B2(A[11]), .C1(n225), .C2(A[10]), .A(n154), 
        .ZN(n65) );
  OAI22_X1 U159 ( .A1(n214), .A2(n228), .B1(n215), .B2(n227), .ZN(n154) );
  AOI221_X1 U160 ( .B1(n226), .B2(A[14]), .C1(n225), .C2(A[13]), .A(n144), 
        .ZN(n91) );
  OAI22_X1 U161 ( .A1(n209), .A2(n228), .B1(n211), .B2(n227), .ZN(n144) );
  INV_X1 U162 ( .A(A[12]), .ZN(n209) );
  OAI221_X1 U163 ( .B1(n92), .B2(n185), .C1(n165), .C2(n186), .A(n141), .ZN(
        n112) );
  AOI22_X1 U164 ( .A1(A[28]), .A2(n95), .B1(A[27]), .B2(n96), .ZN(n141) );
  AOI222_X1 U165 ( .A1(n63), .A2(n74), .B1(n223), .B2(n90), .C1(n61), .C2(n207), .ZN(n89) );
  OAI221_X1 U166 ( .B1(n92), .B2(n217), .C1(n166), .C2(n218), .A(n94), .ZN(n90) );
  AOI22_X1 U167 ( .A1(A[4]), .A2(n95), .B1(A[3]), .B2(n96), .ZN(n94) );
  AOI222_X1 U168 ( .A1(n63), .A2(n79), .B1(n223), .B2(n102), .C1(n61), .C2(
        n208), .ZN(n101) );
  OAI221_X1 U169 ( .B1(n92), .B2(n218), .C1(n166), .C2(n219), .A(n104), .ZN(
        n102) );
  AOI22_X1 U170 ( .A1(A[3]), .A2(n95), .B1(A[2]), .B2(n96), .ZN(n104) );
  AOI222_X1 U171 ( .A1(n63), .A2(n60), .B1(n223), .B2(n119), .C1(n61), .C2(
        n210), .ZN(n118) );
  OAI221_X1 U172 ( .B1(n92), .B2(n219), .C1(n166), .C2(n220), .A(n121), .ZN(
        n119) );
  AOI22_X1 U173 ( .A1(A[2]), .A2(n95), .B1(A[1]), .B2(n96), .ZN(n121) );
  OAI221_X1 U174 ( .B1(n84), .B2(n87), .C1(n127), .C2(n177), .A(n152), .ZN(
        B[0]) );
  AOI222_X1 U175 ( .A1(n63), .A2(n68), .B1(n223), .B2(n153), .C1(n61), .C2(
        n212), .ZN(n152) );
  AND2_X1 U176 ( .A1(n223), .A2(n98), .ZN(B[31]) );
  OAI221_X1 U177 ( .B1(n92), .B2(n220), .C1(n164), .C2(n221), .A(n156), .ZN(
        n153) );
  INV_X1 U178 ( .A(A[2]), .ZN(n221) );
  AOI22_X1 U179 ( .A1(A[1]), .A2(n95), .B1(A[0]), .B2(n96), .ZN(n156) );
  INV_X1 U180 ( .A(A[31]), .ZN(n184) );
  INV_X1 U181 ( .A(A[20]), .ZN(n197) );
  INV_X1 U182 ( .A(A[5]), .ZN(n218) );
  INV_X1 U183 ( .A(A[30]), .ZN(n185) );
  INV_X1 U184 ( .A(A[4]), .ZN(n219) );
  INV_X1 U185 ( .A(A[6]), .ZN(n217) );
  INV_X1 U186 ( .A(A[29]), .ZN(n186) );
  INV_X1 U187 ( .A(A[19]), .ZN(n198) );
  INV_X1 U188 ( .A(A[17]), .ZN(n202) );
  INV_X1 U189 ( .A(A[16]), .ZN(n204) );
  INV_X1 U190 ( .A(A[15]), .ZN(n205) );
  INV_X1 U191 ( .A(A[21]), .ZN(n195) );
  INV_X1 U192 ( .A(A[9]), .ZN(n214) );
  INV_X1 U193 ( .A(A[11]), .ZN(n211) );
  INV_X1 U194 ( .A(A[10]), .ZN(n213) );
  INV_X1 U195 ( .A(A[8]), .ZN(n215) );
  INV_X1 U196 ( .A(A[7]), .ZN(n216) );
  INV_X1 U197 ( .A(A[3]), .ZN(n220) );
  INV_X1 U198 ( .A(A[28]), .ZN(n187) );
  INV_X1 U199 ( .A(A[27]), .ZN(n188) );
  INV_X1 U200 ( .A(A[26]), .ZN(n189) );
  INV_X1 U201 ( .A(A[25]), .ZN(n190) );
  INV_X1 U202 ( .A(A[24]), .ZN(n191) );
  INV_X1 U203 ( .A(A[18]), .ZN(n200) );
  INV_X1 U204 ( .A(SH[0]), .ZN(n167) );
  INV_X1 U205 ( .A(SH[2]), .ZN(n168) );
  INV_X1 U206 ( .A(n170), .ZN(n169) );
endmodule


module SHIFTER_GENERIC_N32_DW_sra_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  NOR2_X2 U4 ( .A1(n174), .A2(SH[3]), .ZN(n109) );
  NOR2_X2 U7 ( .A1(SH[2]), .A2(SH[3]), .ZN(n111) );
  MUX2_X1 U174 ( .A(A[30]), .B(\A[31] ), .S(n95), .Z(n120) );
  NAND2_X1 U2 ( .A1(n181), .A2(\A[31] ), .ZN(n97) );
  INV_X1 U3 ( .A(n181), .ZN(n177) );
  INV_X1 U5 ( .A(n85), .ZN(n228) );
  INV_X1 U6 ( .A(n94), .ZN(n232) );
  INV_X1 U8 ( .A(n95), .ZN(n233) );
  INV_X1 U9 ( .A(n91), .ZN(n230) );
  INV_X1 U10 ( .A(n92), .ZN(n231) );
  NAND2_X1 U11 ( .A1(n109), .A2(n177), .ZN(n85) );
  INV_X1 U12 ( .A(n58), .ZN(n229) );
  BUF_X1 U13 ( .A(n176), .Z(n180) );
  BUF_X1 U14 ( .A(n175), .Z(n179) );
  BUF_X1 U15 ( .A(n175), .Z(n178) );
  BUF_X1 U16 ( .A(n176), .Z(n181) );
  NOR2_X2 U17 ( .A1(n173), .A2(SH[0]), .ZN(n91) );
  NOR2_X2 U18 ( .A1(n172), .A2(n173), .ZN(n92) );
  NAND2_X1 U19 ( .A1(n111), .A2(n177), .ZN(n58) );
  NAND2_X1 U20 ( .A1(n172), .A2(n173), .ZN(n95) );
  NAND2_X1 U21 ( .A1(SH[0]), .A2(n173), .ZN(n94) );
  AND2_X1 U22 ( .A1(n163), .A2(n174), .ZN(n61) );
  AND2_X1 U23 ( .A1(SH[3]), .A2(n174), .ZN(n119) );
  AOI21_X1 U24 ( .B1(n108), .B2(n111), .A(n140), .ZN(n104) );
  AND2_X1 U25 ( .A1(SH[3]), .A2(n177), .ZN(n163) );
  BUF_X1 U26 ( .A(SH[4]), .Z(n176) );
  BUF_X1 U27 ( .A(SH[4]), .Z(n175) );
  OAI222_X1 U28 ( .A1(n95), .A2(n192), .B1(n94), .B2(n191), .C1(n173), .C2(
        n186), .ZN(n108) );
  AND2_X1 U29 ( .A1(SH[2]), .A2(n163), .ZN(n63) );
  AOI221_X1 U30 ( .B1(n120), .B2(n109), .C1(n116), .C2(n111), .A(n188), .ZN(
        n107) );
  AOI221_X1 U31 ( .B1(n108), .B2(n109), .C1(n110), .C2(n111), .A(n188), .ZN(
        n59) );
  AOI221_X1 U32 ( .B1(n112), .B2(n109), .C1(n113), .C2(n111), .A(n188), .ZN(
        n66) );
  AOI221_X1 U33 ( .B1(n114), .B2(n109), .C1(n115), .C2(n111), .A(n188), .ZN(
        n71) );
  AOI221_X1 U34 ( .B1(n116), .B2(n109), .C1(n117), .C2(n111), .A(n189), .ZN(
        n76) );
  INV_X1 U35 ( .A(n118), .ZN(n189) );
  AOI21_X1 U36 ( .B1(n119), .B2(n120), .A(n121), .ZN(n118) );
  AOI221_X1 U37 ( .B1(n110), .B2(n109), .C1(n64), .C2(n111), .A(n184), .ZN(n80) );
  INV_X1 U38 ( .A(n122), .ZN(n184) );
  AOI21_X1 U39 ( .B1(n119), .B2(n108), .A(n121), .ZN(n122) );
  AOI221_X1 U40 ( .B1(n113), .B2(n109), .C1(n69), .C2(n111), .A(n182), .ZN(n83) );
  INV_X1 U41 ( .A(n123), .ZN(n182) );
  AOI21_X1 U42 ( .B1(n119), .B2(n112), .A(n121), .ZN(n123) );
  AOI221_X1 U43 ( .B1(n115), .B2(n109), .C1(n74), .C2(n111), .A(n190), .ZN(n86) );
  INV_X1 U44 ( .A(n131), .ZN(n190) );
  AOI21_X1 U45 ( .B1(n119), .B2(n114), .A(n121), .ZN(n131) );
  AOI221_X1 U46 ( .B1(n120), .B2(n133), .C1(n116), .C2(n119), .A(n196), .ZN(
        n98) );
  INV_X1 U47 ( .A(n134), .ZN(n196) );
  AOI22_X1 U48 ( .A1(n109), .A2(n117), .B1(n111), .B2(n78), .ZN(n134) );
  AOI221_X1 U49 ( .B1(n64), .B2(n109), .C1(n62), .C2(n111), .A(n185), .ZN(n124) );
  INV_X1 U50 ( .A(n135), .ZN(n185) );
  AOI22_X1 U51 ( .A1(n133), .A2(n108), .B1(n119), .B2(n110), .ZN(n135) );
  AOI221_X1 U52 ( .B1(n69), .B2(n109), .C1(n68), .C2(n111), .A(n183), .ZN(n136) );
  INV_X1 U53 ( .A(n166), .ZN(n183) );
  AOI22_X1 U54 ( .A1(n133), .A2(n112), .B1(n119), .B2(n113), .ZN(n166) );
  AOI222_X1 U55 ( .A1(n228), .A2(n68), .B1(n61), .B2(n69), .C1(n63), .C2(n113), 
        .ZN(n147) );
  AOI222_X1 U56 ( .A1(n228), .A2(n73), .B1(n61), .B2(n74), .C1(n63), .C2(n115), 
        .ZN(n148) );
  AOI222_X1 U57 ( .A1(n228), .A2(n207), .B1(n61), .B2(n78), .C1(n63), .C2(n117), .ZN(n154) );
  AOI222_X1 U58 ( .A1(n228), .A2(n78), .B1(n61), .B2(n117), .C1(n63), .C2(n116), .ZN(n139) );
  AOI222_X1 U59 ( .A1(n228), .A2(n209), .B1(n61), .B2(n68), .C1(n63), .C2(n69), 
        .ZN(n67) );
  AOI222_X1 U60 ( .A1(n228), .A2(n62), .B1(n61), .B2(n64), .C1(n63), .C2(n110), 
        .ZN(n141) );
  AOI222_X1 U61 ( .A1(n228), .A2(n208), .B1(n61), .B2(n62), .C1(n63), .C2(n64), 
        .ZN(n60) );
  AOI222_X1 U62 ( .A1(n228), .A2(n212), .B1(n61), .B2(n73), .C1(n63), .C2(n74), 
        .ZN(n72) );
  AOI222_X1 U63 ( .A1(n228), .A2(n213), .B1(n61), .B2(n207), .C1(n63), .C2(n78), .ZN(n77) );
  AOI222_X1 U64 ( .A1(n228), .A2(n216), .B1(n61), .B2(n208), .C1(n63), .C2(n62), .ZN(n81) );
  AOI222_X1 U65 ( .A1(n228), .A2(n218), .B1(n61), .B2(n209), .C1(n63), .C2(n68), .ZN(n84) );
  OAI21_X1 U66 ( .B1(n180), .B2(n96), .A(n97), .ZN(B[30]) );
  OAI21_X1 U67 ( .B1(n180), .B2(n104), .A(n97), .ZN(B[29]) );
  OAI21_X1 U68 ( .B1(n180), .B2(n105), .A(n97), .ZN(B[28]) );
  OAI21_X1 U69 ( .B1(n180), .B2(n106), .A(n97), .ZN(B[27]) );
  OAI21_X1 U70 ( .B1(n180), .B2(n107), .A(n97), .ZN(B[26]) );
  OAI21_X1 U71 ( .B1(n179), .B2(n59), .A(n97), .ZN(B[25]) );
  OAI21_X1 U72 ( .B1(n179), .B2(n66), .A(n97), .ZN(B[24]) );
  OAI21_X1 U73 ( .B1(n179), .B2(n71), .A(n97), .ZN(B[23]) );
  OAI21_X1 U74 ( .B1(n179), .B2(n76), .A(n97), .ZN(B[22]) );
  OAI21_X1 U75 ( .B1(n178), .B2(n80), .A(n97), .ZN(B[21]) );
  OAI21_X1 U76 ( .B1(n178), .B2(n83), .A(n97), .ZN(B[20]) );
  OAI21_X1 U77 ( .B1(n179), .B2(n86), .A(n97), .ZN(B[19]) );
  OAI21_X1 U78 ( .B1(n178), .B2(n98), .A(n97), .ZN(B[18]) );
  OAI21_X1 U79 ( .B1(n178), .B2(n124), .A(n97), .ZN(B[17]) );
  OAI21_X1 U80 ( .B1(n178), .B2(n136), .A(n97), .ZN(B[16]) );
  OAI221_X1 U81 ( .B1(n200), .B2(n85), .C1(n204), .C2(n58), .A(n137), .ZN(
        B[15]) );
  OAI221_X1 U82 ( .B1(n138), .B2(n58), .C1(n96), .C2(n177), .A(n139), .ZN(
        B[14]) );
  OAI221_X1 U83 ( .B1(n129), .B2(n58), .C1(n104), .C2(n177), .A(n141), .ZN(
        B[13]) );
  OAI221_X1 U84 ( .B1(n146), .B2(n58), .C1(n105), .C2(n177), .A(n147), .ZN(
        B[12]) );
  OAI221_X1 U85 ( .B1(n89), .B2(n58), .C1(n106), .C2(n177), .A(n148), .ZN(
        B[11]) );
  OAI221_X1 U86 ( .B1(n101), .B2(n58), .C1(n107), .C2(n177), .A(n154), .ZN(
        B[10]) );
  OAI221_X1 U87 ( .B1(n75), .B2(n85), .C1(n98), .C2(n177), .A(n99), .ZN(B[2])
         );
  OAI221_X1 U88 ( .B1(n79), .B2(n85), .C1(n124), .C2(n177), .A(n125), .ZN(B[1]) );
  OAI221_X1 U89 ( .B1(n57), .B2(n58), .C1(n59), .C2(n177), .A(n60), .ZN(B[9])
         );
  OAI221_X1 U90 ( .B1(n65), .B2(n58), .C1(n66), .C2(n177), .A(n67), .ZN(B[8])
         );
  OAI221_X1 U91 ( .B1(n70), .B2(n58), .C1(n71), .C2(n177), .A(n72), .ZN(B[7])
         );
  OAI221_X1 U92 ( .B1(n75), .B2(n58), .C1(n76), .C2(n177), .A(n77), .ZN(B[6])
         );
  OAI221_X1 U93 ( .B1(n79), .B2(n58), .C1(n80), .C2(n177), .A(n81), .ZN(B[5])
         );
  OAI221_X1 U94 ( .B1(n82), .B2(n58), .C1(n83), .C2(n177), .A(n84), .ZN(B[4])
         );
  OAI221_X1 U95 ( .B1(n70), .B2(n85), .C1(n86), .C2(n177), .A(n87), .ZN(B[3])
         );
  OAI21_X1 U96 ( .B1(n174), .B2(n186), .A(n132), .ZN(n140) );
  AOI221_X1 U97 ( .B1(n63), .B2(n114), .C1(n61), .C2(n115), .A(n187), .ZN(n137) );
  INV_X1 U98 ( .A(n97), .ZN(n187) );
  NOR2_X1 U99 ( .A1(n132), .A2(n174), .ZN(n121) );
  AOI21_X1 U100 ( .B1(n120), .B2(n111), .A(n140), .ZN(n96) );
  AOI21_X1 U101 ( .B1(n112), .B2(n111), .A(n140), .ZN(n105) );
  AOI21_X1 U102 ( .B1(n114), .B2(n111), .A(n140), .ZN(n106) );
  INV_X1 U103 ( .A(SH[0]), .ZN(n172) );
  INV_X1 U104 ( .A(n132), .ZN(n188) );
  INV_X1 U105 ( .A(n138), .ZN(n207) );
  INV_X1 U106 ( .A(n129), .ZN(n208) );
  INV_X1 U107 ( .A(n146), .ZN(n209) );
  AND2_X1 U108 ( .A1(SH[2]), .A2(SH[3]), .ZN(n133) );
  INV_X1 U109 ( .A(n57), .ZN(n216) );
  INV_X1 U110 ( .A(n101), .ZN(n213) );
  INV_X1 U111 ( .A(n89), .ZN(n212) );
  INV_X1 U112 ( .A(n65), .ZN(n218) );
  INV_X1 U113 ( .A(n74), .ZN(n200) );
  INV_X1 U114 ( .A(n73), .ZN(n204) );
  OAI221_X1 U115 ( .B1(n203), .B2(n94), .C1(n205), .C2(n95), .A(n156), .ZN(n78) );
  AOI22_X1 U116 ( .A1(A[20]), .A2(n91), .B1(A[21]), .B2(n92), .ZN(n156) );
  OAI221_X1 U117 ( .B1(n230), .B2(n198), .C1(n231), .C2(n197), .A(n155), .ZN(
        n117) );
  AOI22_X1 U118 ( .A1(A[23]), .A2(n232), .B1(A[22]), .B2(n233), .ZN(n155) );
  OAI221_X1 U119 ( .B1(n230), .B2(n191), .C1(n231), .C2(n186), .A(n168), .ZN(
        n112) );
  AOI22_X1 U120 ( .A1(A[29]), .A2(n232), .B1(A[28]), .B2(n233), .ZN(n168) );
  OAI221_X1 U121 ( .B1(n94), .B2(n201), .C1(n202), .C2(n95), .A(n170), .ZN(n69) );
  INV_X1 U122 ( .A(A[21]), .ZN(n201) );
  AOI22_X1 U123 ( .A1(A[22]), .A2(n91), .B1(A[23]), .B2(n92), .ZN(n170) );
  OAI221_X1 U124 ( .B1(n202), .B2(n94), .C1(n203), .C2(n95), .A(n150), .ZN(n74) );
  AOI22_X1 U125 ( .A1(A[21]), .A2(n91), .B1(A[22]), .B2(n92), .ZN(n150) );
  OAI221_X1 U126 ( .B1(n230), .B2(n197), .C1(n231), .C2(n195), .A(n149), .ZN(
        n115) );
  AOI22_X1 U127 ( .A1(A[24]), .A2(n232), .B1(A[23]), .B2(n233), .ZN(n149) );
  OAI221_X1 U128 ( .B1(n230), .B2(n194), .C1(n231), .C2(n193), .A(n142), .ZN(
        n110) );
  AOI22_X1 U129 ( .A1(A[26]), .A2(n232), .B1(A[25]), .B2(n233), .ZN(n142) );
  OAI221_X1 U130 ( .B1(n230), .B2(n195), .C1(n231), .C2(n194), .A(n167), .ZN(
        n113) );
  AOI22_X1 U131 ( .A1(A[25]), .A2(n232), .B1(A[24]), .B2(n233), .ZN(n167) );
  OAI221_X1 U132 ( .B1(n230), .B2(n199), .C1(n231), .C2(n198), .A(n143), .ZN(
        n64) );
  INV_X1 U133 ( .A(A[23]), .ZN(n199) );
  AOI22_X1 U134 ( .A1(A[22]), .A2(n232), .B1(A[21]), .B2(n233), .ZN(n143) );
  OAI221_X1 U135 ( .B1(n230), .B2(n206), .C1(n231), .C2(n205), .A(n151), .ZN(
        n73) );
  INV_X1 U136 ( .A(A[17]), .ZN(n206) );
  AOI22_X1 U137 ( .A1(A[16]), .A2(n232), .B1(A[15]), .B2(n233), .ZN(n151) );
  OAI221_X1 U138 ( .B1(n230), .B2(n203), .C1(n231), .C2(n202), .A(n144), .ZN(
        n62) );
  AOI22_X1 U139 ( .A1(A[18]), .A2(n232), .B1(A[17]), .B2(n233), .ZN(n144) );
  OAI221_X1 U140 ( .B1(n230), .B2(n205), .C1(n203), .C2(n231), .A(n169), .ZN(
        n68) );
  AOI22_X1 U141 ( .A1(A[17]), .A2(n232), .B1(A[16]), .B2(n233), .ZN(n169) );
  OAI221_X1 U142 ( .B1(n230), .B2(n192), .C1(n231), .C2(n191), .A(n152), .ZN(
        n114) );
  AOI22_X1 U143 ( .A1(A[28]), .A2(n232), .B1(A[27]), .B2(n233), .ZN(n152) );
  OAI221_X1 U144 ( .B1(n230), .B2(n193), .C1(n231), .C2(n192), .A(n158), .ZN(
        n116) );
  AOI22_X1 U145 ( .A1(A[27]), .A2(n232), .B1(A[26]), .B2(n233), .ZN(n158) );
  AOI221_X1 U146 ( .B1(n91), .B2(A[8]), .C1(n92), .C2(A[9]), .A(n103), .ZN(n75) );
  OAI22_X1 U147 ( .A1(n222), .A2(n94), .B1(n223), .B2(n95), .ZN(n103) );
  AOI221_X1 U148 ( .B1(n91), .B2(A[9]), .C1(n92), .C2(A[10]), .A(n93), .ZN(n70) );
  OAI22_X1 U149 ( .A1(n221), .A2(n94), .B1(n222), .B2(n95), .ZN(n93) );
  AOI221_X1 U150 ( .B1(n91), .B2(A[7]), .C1(n92), .C2(A[8]), .A(n130), .ZN(n79) );
  OAI22_X1 U151 ( .A1(n223), .A2(n94), .B1(n224), .B2(n95), .ZN(n130) );
  AOI221_X1 U152 ( .B1(n91), .B2(A[6]), .C1(n92), .C2(A[7]), .A(n171), .ZN(n82) );
  OAI22_X1 U153 ( .A1(n224), .A2(n94), .B1(n225), .B2(n95), .ZN(n171) );
  AOI221_X1 U154 ( .B1(n91), .B2(A[11]), .C1(n92), .C2(A[12]), .A(n127), .ZN(
        n57) );
  OAI22_X1 U155 ( .A1(n219), .A2(n94), .B1(n220), .B2(n95), .ZN(n127) );
  AOI221_X1 U156 ( .B1(n91), .B2(A[12]), .C1(n92), .C2(A[13]), .A(n159), .ZN(
        n101) );
  OAI22_X1 U157 ( .A1(n217), .A2(n94), .B1(n219), .B2(n95), .ZN(n159) );
  AOI221_X1 U158 ( .B1(n91), .B2(A[13]), .C1(n92), .C2(A[14]), .A(n153), .ZN(
        n89) );
  OAI22_X1 U159 ( .A1(n215), .A2(n94), .B1(n217), .B2(n95), .ZN(n153) );
  INV_X1 U160 ( .A(A[12]), .ZN(n215) );
  AOI221_X1 U161 ( .B1(n91), .B2(A[16]), .C1(n92), .C2(A[17]), .A(n210), .ZN(
        n138) );
  INV_X1 U162 ( .A(n157), .ZN(n210) );
  AOI22_X1 U163 ( .A1(A[15]), .A2(n232), .B1(A[14]), .B2(n233), .ZN(n157) );
  AOI221_X1 U164 ( .B1(n91), .B2(A[15]), .C1(n92), .C2(A[16]), .A(n211), .ZN(
        n129) );
  INV_X1 U165 ( .A(n145), .ZN(n211) );
  AOI22_X1 U166 ( .A1(A[14]), .A2(n232), .B1(A[13]), .B2(n233), .ZN(n145) );
  AOI221_X1 U167 ( .B1(n91), .B2(A[14]), .C1(n92), .C2(A[15]), .A(n214), .ZN(
        n146) );
  INV_X1 U168 ( .A(n165), .ZN(n214) );
  AOI22_X1 U169 ( .A1(A[13]), .A2(n232), .B1(A[12]), .B2(n233), .ZN(n165) );
  AOI221_X1 U170 ( .B1(n91), .B2(A[10]), .C1(n92), .C2(A[11]), .A(n162), .ZN(
        n65) );
  OAI22_X1 U171 ( .A1(n220), .A2(n94), .B1(n221), .B2(n95), .ZN(n162) );
  AOI222_X1 U172 ( .A1(n63), .A2(n73), .B1(n229), .B2(n88), .C1(n61), .C2(n212), .ZN(n87) );
  OAI221_X1 U173 ( .B1(n230), .B2(n224), .C1(n231), .C2(n223), .A(n90), .ZN(
        n88) );
  AOI22_X1 U175 ( .A1(A[4]), .A2(n232), .B1(A[3]), .B2(n233), .ZN(n90) );
  AOI222_X1 U176 ( .A1(n63), .A2(n208), .B1(n229), .B2(n126), .C1(n61), .C2(
        n216), .ZN(n125) );
  OAI221_X1 U177 ( .B1(n230), .B2(n226), .C1(n231), .C2(n225), .A(n128), .ZN(
        n126) );
  AOI22_X1 U178 ( .A1(A[2]), .A2(n232), .B1(A[1]), .B2(n233), .ZN(n128) );
  AOI222_X1 U179 ( .A1(n63), .A2(n209), .B1(n229), .B2(n161), .C1(n61), .C2(
        n218), .ZN(n160) );
  OAI221_X1 U180 ( .B1(n230), .B2(n227), .C1(n231), .C2(n226), .A(n164), .ZN(
        n161) );
  INV_X1 U181 ( .A(A[2]), .ZN(n227) );
  AOI22_X1 U182 ( .A1(A[1]), .A2(n232), .B1(A[0]), .B2(n233), .ZN(n164) );
  AOI222_X1 U183 ( .A1(n63), .A2(n207), .B1(n229), .B2(n100), .C1(n61), .C2(
        n213), .ZN(n99) );
  OAI221_X1 U184 ( .B1(n230), .B2(n225), .C1(n231), .C2(n224), .A(n102), .ZN(
        n100) );
  AOI22_X1 U185 ( .A1(A[3]), .A2(n232), .B1(A[2]), .B2(n233), .ZN(n102) );
  OAI221_X1 U186 ( .B1(n82), .B2(n85), .C1(n136), .C2(n177), .A(n160), .ZN(
        B[0]) );
  NAND2_X1 U187 ( .A1(\A[31] ), .A2(SH[3]), .ZN(n132) );
  INV_X1 U188 ( .A(A[19]), .ZN(n203) );
  INV_X1 U189 ( .A(A[5]), .ZN(n224) );
  INV_X1 U190 ( .A(A[18]), .ZN(n205) );
  INV_X1 U191 ( .A(A[6]), .ZN(n223) );
  INV_X1 U192 ( .A(A[4]), .ZN(n225) );
  INV_X1 U193 ( .A(A[29]), .ZN(n192) );
  INV_X1 U194 ( .A(A[20]), .ZN(n202) );
  INV_X1 U195 ( .A(\A[31] ), .ZN(n186) );
  INV_X1 U196 ( .A(A[9]), .ZN(n220) );
  INV_X1 U197 ( .A(A[11]), .ZN(n217) );
  INV_X1 U198 ( .A(A[10]), .ZN(n219) );
  INV_X1 U199 ( .A(A[8]), .ZN(n221) );
  INV_X1 U200 ( .A(A[7]), .ZN(n222) );
  INV_X1 U201 ( .A(A[3]), .ZN(n226) );
  INV_X1 U202 ( .A(A[27]), .ZN(n194) );
  INV_X1 U203 ( .A(A[26]), .ZN(n195) );
  INV_X1 U204 ( .A(A[25]), .ZN(n197) );
  INV_X1 U205 ( .A(A[28]), .ZN(n193) );
  INV_X1 U206 ( .A(A[24]), .ZN(n198) );
  INV_X1 U207 ( .A(A[30]), .ZN(n191) );
  INV_X1 U208 ( .A(SH[1]), .ZN(n173) );
  INV_X1 U209 ( .A(SH[2]), .ZN(n174) );
endmodule


module SHIFTER_GENERIC_N32_DW_lbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] ,
         \ML_int[5][31] , \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] ,
         \ML_int[5][15] , \ML_int[5][14] , \ML_int[5][13] , \ML_int[5][12] ,
         \ML_int[5][11] , \ML_int[5][10] , \ML_int[5][9] , \ML_int[5][8] ,
         \ML_int[5][7] , \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] ,
         \ML_int[5][3] , \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[31] = \ML_int[5][31] ;
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[15] = \ML_int[5][15] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[8] = \ML_int[5][8] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n18), .Z(
        \ML_int[5][31] ) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n18), .Z(
        \ML_int[5][30] ) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n18), .Z(
        \ML_int[5][29] ) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n18), .Z(
        \ML_int[5][28] ) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n18), .Z(
        \ML_int[5][27] ) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n18), .Z(
        \ML_int[5][26] ) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n18), .Z(
        \ML_int[5][25] ) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n18), .Z(
        \ML_int[5][24] ) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n18), .Z(
        \ML_int[5][23] ) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n18), .Z(
        \ML_int[5][22] ) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n16), .Z(
        \ML_int[5][21] ) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n16), .Z(
        \ML_int[5][20] ) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n16), .Z(
        \ML_int[5][19] ) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n16), .Z(
        \ML_int[5][18] ) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n16), .Z(
        \ML_int[5][17] ) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n16), .Z(
        \ML_int[5][16] ) );
  MUX2_X1 M0_4_15 ( .A(\ML_int[4][15] ), .B(\ML_int[4][31] ), .S(n16), .Z(
        \ML_int[5][15] ) );
  MUX2_X1 M0_4_14 ( .A(\ML_int[4][14] ), .B(\ML_int[4][30] ), .S(n16), .Z(
        \ML_int[5][14] ) );
  MUX2_X1 M0_4_13 ( .A(\ML_int[4][13] ), .B(\ML_int[4][29] ), .S(n16), .Z(
        \ML_int[5][13] ) );
  MUX2_X1 M0_4_12 ( .A(\ML_int[4][12] ), .B(\ML_int[4][28] ), .S(n16), .Z(
        \ML_int[5][12] ) );
  MUX2_X1 M0_4_11 ( .A(\ML_int[4][11] ), .B(\ML_int[4][27] ), .S(n16), .Z(
        \ML_int[5][11] ) );
  MUX2_X1 M0_4_10 ( .A(\ML_int[4][10] ), .B(\ML_int[4][26] ), .S(n17), .Z(
        \ML_int[5][10] ) );
  MUX2_X1 M0_4_9 ( .A(\ML_int[4][9] ), .B(\ML_int[4][25] ), .S(n17), .Z(
        \ML_int[5][9] ) );
  MUX2_X1 M0_4_8 ( .A(\ML_int[4][8] ), .B(\ML_int[4][24] ), .S(n17), .Z(
        \ML_int[5][8] ) );
  MUX2_X1 M0_4_7 ( .A(\ML_int[4][7] ), .B(\ML_int[4][23] ), .S(n17), .Z(
        \ML_int[5][7] ) );
  MUX2_X1 M0_4_6 ( .A(\ML_int[4][6] ), .B(\ML_int[4][22] ), .S(n17), .Z(
        \ML_int[5][6] ) );
  MUX2_X1 M0_4_5 ( .A(\ML_int[4][5] ), .B(\ML_int[4][21] ), .S(n17), .Z(
        \ML_int[5][5] ) );
  MUX2_X1 M0_4_4 ( .A(\ML_int[4][4] ), .B(\ML_int[4][20] ), .S(n17), .Z(
        \ML_int[5][4] ) );
  MUX2_X1 M0_4_3 ( .A(\ML_int[4][3] ), .B(\ML_int[4][19] ), .S(n17), .Z(
        \ML_int[5][3] ) );
  MUX2_X1 M0_4_2 ( .A(\ML_int[4][2] ), .B(\ML_int[4][18] ), .S(n17), .Z(
        \ML_int[5][2] ) );
  MUX2_X1 M0_4_1 ( .A(\ML_int[4][1] ), .B(\ML_int[4][17] ), .S(n17), .Z(
        \ML_int[5][1] ) );
  MUX2_X1 M0_4_0 ( .A(\ML_int[4][0] ), .B(\ML_int[4][16] ), .S(n17), .Z(
        \ML_int[5][0] ) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n15), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n15), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n15), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n15), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n15), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n15), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n15), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n15), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n15), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n15), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n14), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n14), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n14), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n14), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n14), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n14), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n14), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n14), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n14), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n14), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n14), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n13), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n13), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n13), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M0_3_7 ( .A(\ML_int[3][7] ), .B(\ML_int[3][31] ), .S(n13), .Z(
        \ML_int[4][7] ) );
  MUX2_X1 M0_3_6 ( .A(\ML_int[3][6] ), .B(\ML_int[3][30] ), .S(n13), .Z(
        \ML_int[4][6] ) );
  MUX2_X1 M0_3_5 ( .A(\ML_int[3][5] ), .B(\ML_int[3][29] ), .S(n13), .Z(
        \ML_int[4][5] ) );
  MUX2_X1 M0_3_4 ( .A(\ML_int[3][4] ), .B(\ML_int[3][28] ), .S(n13), .Z(
        \ML_int[4][4] ) );
  MUX2_X1 M0_3_3 ( .A(\ML_int[3][3] ), .B(\ML_int[3][27] ), .S(n13), .Z(
        \ML_int[4][3] ) );
  MUX2_X1 M0_3_2 ( .A(\ML_int[3][2] ), .B(\ML_int[3][26] ), .S(n13), .Z(
        \ML_int[4][2] ) );
  MUX2_X1 M0_3_1 ( .A(\ML_int[3][1] ), .B(\ML_int[3][25] ), .S(n13), .Z(
        \ML_int[4][1] ) );
  MUX2_X1 M0_3_0 ( .A(\ML_int[3][0] ), .B(\ML_int[3][24] ), .S(n13), .Z(
        \ML_int[4][0] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n12), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n12), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n12), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n12), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n12), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n12), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n12), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n12), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n12), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n12), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n11), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n11), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n11), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n11), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n11), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n11), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n11), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n11), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n11), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n11), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n11), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n10), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n10), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n10), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n10), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n10), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n10), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n10), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M0_2_3 ( .A(\ML_int[2][3] ), .B(\ML_int[2][31] ), .S(n10), .Z(
        \ML_int[3][3] ) );
  MUX2_X1 M0_2_2 ( .A(\ML_int[2][2] ), .B(\ML_int[2][30] ), .S(n10), .Z(
        \ML_int[3][2] ) );
  MUX2_X1 M0_2_1 ( .A(\ML_int[2][1] ), .B(\ML_int[2][29] ), .S(n10), .Z(
        \ML_int[3][1] ) );
  MUX2_X1 M0_2_0 ( .A(\ML_int[2][0] ), .B(\ML_int[2][28] ), .S(n10), .Z(
        \ML_int[3][0] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n9), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n9), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n9), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n9), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n9), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n9), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n9), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n9), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n9), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n9), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n8), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n8), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n8), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n8), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n8), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n8), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n8), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n8), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n8), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n8), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n8), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n7), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n7), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n7), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n7), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n7), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n7), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n7), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n7), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n7), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M0_1_1 ( .A(\ML_int[1][1] ), .B(\ML_int[1][31] ), .S(n7), .Z(
        \ML_int[2][1] ) );
  MUX2_X1 M0_1_0 ( .A(\ML_int[1][0] ), .B(\ML_int[1][30] ), .S(n7), .Z(
        \ML_int[2][0] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n6), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n6), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n6), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n6), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n6), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n6), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n6), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n6), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n6), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n6), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n5), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n5), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n5), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n5), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n5), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n5), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n5), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n5), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n5), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n5), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n5), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n4), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n4), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n4), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n4), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n4), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n4), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n4), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n4), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n4), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n4), .Z(\ML_int[1][1] ) );
  MUX2_X1 M0_0_0 ( .A(A[0]), .B(A[31]), .S(n4), .Z(\ML_int[1][0] ) );
  BUF_X1 U2 ( .A(SH[3]), .Z(n14) );
  BUF_X1 U3 ( .A(SH[3]), .Z(n13) );
  BUF_X1 U4 ( .A(SH[4]), .Z(n16) );
  BUF_X1 U5 ( .A(SH[4]), .Z(n17) );
  BUF_X1 U6 ( .A(SH[3]), .Z(n15) );
  BUF_X1 U7 ( .A(SH[4]), .Z(n18) );
  BUF_X1 U8 ( .A(SH[0]), .Z(n4) );
  BUF_X1 U9 ( .A(SH[0]), .Z(n5) );
  BUF_X1 U10 ( .A(SH[1]), .Z(n7) );
  BUF_X1 U11 ( .A(SH[1]), .Z(n8) );
  BUF_X1 U12 ( .A(SH[2]), .Z(n11) );
  BUF_X1 U13 ( .A(SH[2]), .Z(n10) );
  BUF_X1 U14 ( .A(SH[0]), .Z(n6) );
  BUF_X1 U15 ( .A(SH[1]), .Z(n9) );
  BUF_X1 U16 ( .A(SH[2]), .Z(n12) );
endmodule


module SHIFTER_GENERIC_N32_DW_rbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \MR_int[1][31] , \MR_int[1][30] , \MR_int[1][29] , \MR_int[1][28] ,
         \MR_int[1][27] , \MR_int[1][26] , \MR_int[1][25] , \MR_int[1][24] ,
         \MR_int[1][23] , \MR_int[1][22] , \MR_int[1][21] , \MR_int[1][20] ,
         \MR_int[1][19] , \MR_int[1][18] , \MR_int[1][17] , \MR_int[1][16] ,
         \MR_int[1][15] , \MR_int[1][14] , \MR_int[1][13] , \MR_int[1][12] ,
         \MR_int[1][11] , \MR_int[1][10] , \MR_int[1][9] , \MR_int[1][8] ,
         \MR_int[1][7] , \MR_int[1][6] , \MR_int[1][5] , \MR_int[1][4] ,
         \MR_int[1][3] , \MR_int[1][2] , \MR_int[1][1] , \MR_int[1][0] ,
         \MR_int[2][31] , \MR_int[2][30] , \MR_int[2][29] , \MR_int[2][28] ,
         \MR_int[2][27] , \MR_int[2][26] , \MR_int[2][25] , \MR_int[2][24] ,
         \MR_int[2][23] , \MR_int[2][22] , \MR_int[2][21] , \MR_int[2][20] ,
         \MR_int[2][19] , \MR_int[2][18] , \MR_int[2][17] , \MR_int[2][16] ,
         \MR_int[2][15] , \MR_int[2][14] , \MR_int[2][13] , \MR_int[2][12] ,
         \MR_int[2][11] , \MR_int[2][10] , \MR_int[2][9] , \MR_int[2][8] ,
         \MR_int[2][7] , \MR_int[2][6] , \MR_int[2][5] , \MR_int[2][4] ,
         \MR_int[2][3] , \MR_int[2][2] , \MR_int[2][1] , \MR_int[2][0] ,
         \MR_int[3][31] , \MR_int[3][30] , \MR_int[3][29] , \MR_int[3][28] ,
         \MR_int[3][27] , \MR_int[3][26] , \MR_int[3][25] , \MR_int[3][24] ,
         \MR_int[3][23] , \MR_int[3][22] , \MR_int[3][21] , \MR_int[3][20] ,
         \MR_int[3][19] , \MR_int[3][18] , \MR_int[3][17] , \MR_int[3][16] ,
         \MR_int[3][15] , \MR_int[3][14] , \MR_int[3][13] , \MR_int[3][12] ,
         \MR_int[3][11] , \MR_int[3][10] , \MR_int[3][9] , \MR_int[3][8] ,
         \MR_int[3][7] , \MR_int[3][6] , \MR_int[3][5] , \MR_int[3][4] ,
         \MR_int[3][3] , \MR_int[3][2] , \MR_int[3][1] , \MR_int[3][0] ,
         \MR_int[4][31] , \MR_int[4][30] , \MR_int[4][29] , \MR_int[4][28] ,
         \MR_int[4][27] , \MR_int[4][26] , \MR_int[4][25] , \MR_int[4][24] ,
         \MR_int[4][23] , \MR_int[4][22] , \MR_int[4][21] , \MR_int[4][20] ,
         \MR_int[4][19] , \MR_int[4][18] , \MR_int[4][17] , \MR_int[4][16] ,
         \MR_int[4][15] , \MR_int[4][14] , \MR_int[4][13] , \MR_int[4][12] ,
         \MR_int[4][11] , \MR_int[4][10] , \MR_int[4][9] , \MR_int[4][8] ,
         \MR_int[4][7] , \MR_int[4][6] , \MR_int[4][5] , \MR_int[4][4] ,
         \MR_int[4][3] , \MR_int[4][2] , \MR_int[4][1] , \MR_int[4][0] ,
         \MR_int[5][31] , \MR_int[5][30] , \MR_int[5][29] , \MR_int[5][28] ,
         \MR_int[5][27] , \MR_int[5][26] , \MR_int[5][25] , \MR_int[5][24] ,
         \MR_int[5][23] , \MR_int[5][22] , \MR_int[5][21] , \MR_int[5][20] ,
         \MR_int[5][19] , \MR_int[5][18] , \MR_int[5][17] , \MR_int[5][16] ,
         \MR_int[5][15] , \MR_int[5][14] , \MR_int[5][13] , \MR_int[5][12] ,
         \MR_int[5][11] , \MR_int[5][10] , \MR_int[5][9] , \MR_int[5][8] ,
         \MR_int[5][7] , \MR_int[5][6] , \MR_int[5][5] , \MR_int[5][4] ,
         \MR_int[5][3] , \MR_int[5][2] , \MR_int[5][1] , \MR_int[5][0] , n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18;
  assign B[31] = \MR_int[5][31] ;
  assign B[30] = \MR_int[5][30] ;
  assign B[29] = \MR_int[5][29] ;
  assign B[28] = \MR_int[5][28] ;
  assign B[27] = \MR_int[5][27] ;
  assign B[26] = \MR_int[5][26] ;
  assign B[25] = \MR_int[5][25] ;
  assign B[24] = \MR_int[5][24] ;
  assign B[23] = \MR_int[5][23] ;
  assign B[22] = \MR_int[5][22] ;
  assign B[21] = \MR_int[5][21] ;
  assign B[20] = \MR_int[5][20] ;
  assign B[19] = \MR_int[5][19] ;
  assign B[18] = \MR_int[5][18] ;
  assign B[17] = \MR_int[5][17] ;
  assign B[16] = \MR_int[5][16] ;
  assign B[15] = \MR_int[5][15] ;
  assign B[14] = \MR_int[5][14] ;
  assign B[13] = \MR_int[5][13] ;
  assign B[12] = \MR_int[5][12] ;
  assign B[11] = \MR_int[5][11] ;
  assign B[10] = \MR_int[5][10] ;
  assign B[9] = \MR_int[5][9] ;
  assign B[8] = \MR_int[5][8] ;
  assign B[7] = \MR_int[5][7] ;
  assign B[6] = \MR_int[5][6] ;
  assign B[5] = \MR_int[5][5] ;
  assign B[4] = \MR_int[5][4] ;
  assign B[3] = \MR_int[5][3] ;
  assign B[2] = \MR_int[5][2] ;
  assign B[1] = \MR_int[5][1] ;
  assign B[0] = \MR_int[5][0] ;

  MUX2_X1 M1_4_31 ( .A(\MR_int[4][31] ), .B(\MR_int[4][15] ), .S(n18), .Z(
        \MR_int[5][31] ) );
  MUX2_X1 M1_4_30 ( .A(\MR_int[4][30] ), .B(\MR_int[4][14] ), .S(n18), .Z(
        \MR_int[5][30] ) );
  MUX2_X1 M1_4_29 ( .A(\MR_int[4][29] ), .B(\MR_int[4][13] ), .S(n18), .Z(
        \MR_int[5][29] ) );
  MUX2_X1 M1_4_28 ( .A(\MR_int[4][28] ), .B(\MR_int[4][12] ), .S(n18), .Z(
        \MR_int[5][28] ) );
  MUX2_X1 M1_4_27 ( .A(\MR_int[4][27] ), .B(\MR_int[4][11] ), .S(n18), .Z(
        \MR_int[5][27] ) );
  MUX2_X1 M1_4_26 ( .A(\MR_int[4][26] ), .B(\MR_int[4][10] ), .S(n18), .Z(
        \MR_int[5][26] ) );
  MUX2_X1 M1_4_25 ( .A(\MR_int[4][25] ), .B(\MR_int[4][9] ), .S(n18), .Z(
        \MR_int[5][25] ) );
  MUX2_X1 M1_4_24 ( .A(\MR_int[4][24] ), .B(\MR_int[4][8] ), .S(n18), .Z(
        \MR_int[5][24] ) );
  MUX2_X1 M1_4_23 ( .A(\MR_int[4][23] ), .B(\MR_int[4][7] ), .S(n18), .Z(
        \MR_int[5][23] ) );
  MUX2_X1 M1_4_22 ( .A(\MR_int[4][22] ), .B(\MR_int[4][6] ), .S(n18), .Z(
        \MR_int[5][22] ) );
  MUX2_X1 M1_4_21 ( .A(\MR_int[4][21] ), .B(\MR_int[4][5] ), .S(n16), .Z(
        \MR_int[5][21] ) );
  MUX2_X1 M1_4_20 ( .A(\MR_int[4][20] ), .B(\MR_int[4][4] ), .S(n16), .Z(
        \MR_int[5][20] ) );
  MUX2_X1 M1_4_19 ( .A(\MR_int[4][19] ), .B(\MR_int[4][3] ), .S(n16), .Z(
        \MR_int[5][19] ) );
  MUX2_X1 M1_4_18 ( .A(\MR_int[4][18] ), .B(\MR_int[4][2] ), .S(n16), .Z(
        \MR_int[5][18] ) );
  MUX2_X1 M1_4_17 ( .A(\MR_int[4][17] ), .B(\MR_int[4][1] ), .S(n16), .Z(
        \MR_int[5][17] ) );
  MUX2_X1 M1_4_16 ( .A(\MR_int[4][16] ), .B(\MR_int[4][0] ), .S(n16), .Z(
        \MR_int[5][16] ) );
  MUX2_X1 M1_4_15 ( .A(\MR_int[4][15] ), .B(\MR_int[4][31] ), .S(n16), .Z(
        \MR_int[5][15] ) );
  MUX2_X1 M1_4_14 ( .A(\MR_int[4][14] ), .B(\MR_int[4][30] ), .S(n16), .Z(
        \MR_int[5][14] ) );
  MUX2_X1 M1_4_13 ( .A(\MR_int[4][13] ), .B(\MR_int[4][29] ), .S(n16), .Z(
        \MR_int[5][13] ) );
  MUX2_X1 M1_4_12 ( .A(\MR_int[4][12] ), .B(\MR_int[4][28] ), .S(n16), .Z(
        \MR_int[5][12] ) );
  MUX2_X1 M1_4_11 ( .A(\MR_int[4][11] ), .B(\MR_int[4][27] ), .S(n16), .Z(
        \MR_int[5][11] ) );
  MUX2_X1 M1_4_10 ( .A(\MR_int[4][10] ), .B(\MR_int[4][26] ), .S(n17), .Z(
        \MR_int[5][10] ) );
  MUX2_X1 M1_4_9 ( .A(\MR_int[4][9] ), .B(\MR_int[4][25] ), .S(n17), .Z(
        \MR_int[5][9] ) );
  MUX2_X1 M1_4_8 ( .A(\MR_int[4][8] ), .B(\MR_int[4][24] ), .S(n17), .Z(
        \MR_int[5][8] ) );
  MUX2_X1 M1_4_7 ( .A(\MR_int[4][7] ), .B(\MR_int[4][23] ), .S(n17), .Z(
        \MR_int[5][7] ) );
  MUX2_X1 M1_4_6 ( .A(\MR_int[4][6] ), .B(\MR_int[4][22] ), .S(n17), .Z(
        \MR_int[5][6] ) );
  MUX2_X1 M1_4_5 ( .A(\MR_int[4][5] ), .B(\MR_int[4][21] ), .S(n17), .Z(
        \MR_int[5][5] ) );
  MUX2_X1 M1_4_4 ( .A(\MR_int[4][4] ), .B(\MR_int[4][20] ), .S(n17), .Z(
        \MR_int[5][4] ) );
  MUX2_X1 M1_4_3 ( .A(\MR_int[4][3] ), .B(\MR_int[4][19] ), .S(n17), .Z(
        \MR_int[5][3] ) );
  MUX2_X1 M1_4_2 ( .A(\MR_int[4][2] ), .B(\MR_int[4][18] ), .S(n17), .Z(
        \MR_int[5][2] ) );
  MUX2_X1 M1_4_1 ( .A(\MR_int[4][1] ), .B(\MR_int[4][17] ), .S(n17), .Z(
        \MR_int[5][1] ) );
  MUX2_X1 M1_4_0 ( .A(\MR_int[4][0] ), .B(\MR_int[4][16] ), .S(n17), .Z(
        \MR_int[5][0] ) );
  MUX2_X1 M1_3_31_0 ( .A(\MR_int[3][31] ), .B(\MR_int[3][7] ), .S(n15), .Z(
        \MR_int[4][31] ) );
  MUX2_X1 M1_3_30_0 ( .A(\MR_int[3][30] ), .B(\MR_int[3][6] ), .S(n15), .Z(
        \MR_int[4][30] ) );
  MUX2_X1 M1_3_29_0 ( .A(\MR_int[3][29] ), .B(\MR_int[3][5] ), .S(n15), .Z(
        \MR_int[4][29] ) );
  MUX2_X1 M1_3_28_0 ( .A(\MR_int[3][28] ), .B(\MR_int[3][4] ), .S(n15), .Z(
        \MR_int[4][28] ) );
  MUX2_X1 M1_3_27_0 ( .A(\MR_int[3][27] ), .B(\MR_int[3][3] ), .S(n15), .Z(
        \MR_int[4][27] ) );
  MUX2_X1 M1_3_26_0 ( .A(\MR_int[3][26] ), .B(\MR_int[3][2] ), .S(n15), .Z(
        \MR_int[4][26] ) );
  MUX2_X1 M1_3_25_0 ( .A(\MR_int[3][25] ), .B(\MR_int[3][1] ), .S(n15), .Z(
        \MR_int[4][25] ) );
  MUX2_X1 M1_3_24_0 ( .A(\MR_int[3][24] ), .B(\MR_int[3][0] ), .S(n15), .Z(
        \MR_int[4][24] ) );
  MUX2_X1 M1_3_23_0 ( .A(\MR_int[3][23] ), .B(\MR_int[3][31] ), .S(n15), .Z(
        \MR_int[4][23] ) );
  MUX2_X1 M1_3_22_0 ( .A(\MR_int[3][22] ), .B(\MR_int[3][30] ), .S(n15), .Z(
        \MR_int[4][22] ) );
  MUX2_X1 M1_3_21_0 ( .A(\MR_int[3][21] ), .B(\MR_int[3][29] ), .S(n14), .Z(
        \MR_int[4][21] ) );
  MUX2_X1 M1_3_20_0 ( .A(\MR_int[3][20] ), .B(\MR_int[3][28] ), .S(n14), .Z(
        \MR_int[4][20] ) );
  MUX2_X1 M1_3_19_0 ( .A(\MR_int[3][19] ), .B(\MR_int[3][27] ), .S(n14), .Z(
        \MR_int[4][19] ) );
  MUX2_X1 M1_3_18_0 ( .A(\MR_int[3][18] ), .B(\MR_int[3][26] ), .S(n14), .Z(
        \MR_int[4][18] ) );
  MUX2_X1 M1_3_17_0 ( .A(\MR_int[3][17] ), .B(\MR_int[3][25] ), .S(n14), .Z(
        \MR_int[4][17] ) );
  MUX2_X1 M1_3_16_0 ( .A(\MR_int[3][16] ), .B(\MR_int[3][24] ), .S(n14), .Z(
        \MR_int[4][16] ) );
  MUX2_X1 M1_3_15_0 ( .A(\MR_int[3][15] ), .B(\MR_int[3][23] ), .S(n14), .Z(
        \MR_int[4][15] ) );
  MUX2_X1 M1_3_14_0 ( .A(\MR_int[3][14] ), .B(\MR_int[3][22] ), .S(n14), .Z(
        \MR_int[4][14] ) );
  MUX2_X1 M1_3_13_0 ( .A(\MR_int[3][13] ), .B(\MR_int[3][21] ), .S(n14), .Z(
        \MR_int[4][13] ) );
  MUX2_X1 M1_3_12_0 ( .A(\MR_int[3][12] ), .B(\MR_int[3][20] ), .S(n14), .Z(
        \MR_int[4][12] ) );
  MUX2_X1 M1_3_11_0 ( .A(\MR_int[3][11] ), .B(\MR_int[3][19] ), .S(n14), .Z(
        \MR_int[4][11] ) );
  MUX2_X1 M1_3_10_0 ( .A(\MR_int[3][10] ), .B(\MR_int[3][18] ), .S(n13), .Z(
        \MR_int[4][10] ) );
  MUX2_X1 M1_3_9_0 ( .A(\MR_int[3][9] ), .B(\MR_int[3][17] ), .S(n13), .Z(
        \MR_int[4][9] ) );
  MUX2_X1 M1_3_8_0 ( .A(\MR_int[3][8] ), .B(\MR_int[3][16] ), .S(n13), .Z(
        \MR_int[4][8] ) );
  MUX2_X1 M1_3_7 ( .A(\MR_int[3][7] ), .B(\MR_int[3][15] ), .S(n13), .Z(
        \MR_int[4][7] ) );
  MUX2_X1 M1_3_6 ( .A(\MR_int[3][6] ), .B(\MR_int[3][14] ), .S(n13), .Z(
        \MR_int[4][6] ) );
  MUX2_X1 M1_3_5 ( .A(\MR_int[3][5] ), .B(\MR_int[3][13] ), .S(n13), .Z(
        \MR_int[4][5] ) );
  MUX2_X1 M1_3_4 ( .A(\MR_int[3][4] ), .B(\MR_int[3][12] ), .S(n13), .Z(
        \MR_int[4][4] ) );
  MUX2_X1 M1_3_3 ( .A(\MR_int[3][3] ), .B(\MR_int[3][11] ), .S(n13), .Z(
        \MR_int[4][3] ) );
  MUX2_X1 M1_3_2 ( .A(\MR_int[3][2] ), .B(\MR_int[3][10] ), .S(n13), .Z(
        \MR_int[4][2] ) );
  MUX2_X1 M1_3_1 ( .A(\MR_int[3][1] ), .B(\MR_int[3][9] ), .S(n13), .Z(
        \MR_int[4][1] ) );
  MUX2_X1 M1_3_0 ( .A(\MR_int[3][0] ), .B(\MR_int[3][8] ), .S(n13), .Z(
        \MR_int[4][0] ) );
  MUX2_X1 M1_2_31_0 ( .A(\MR_int[2][31] ), .B(\MR_int[2][3] ), .S(n12), .Z(
        \MR_int[3][31] ) );
  MUX2_X1 M1_2_30_0 ( .A(\MR_int[2][30] ), .B(\MR_int[2][2] ), .S(n12), .Z(
        \MR_int[3][30] ) );
  MUX2_X1 M1_2_29_0 ( .A(\MR_int[2][29] ), .B(\MR_int[2][1] ), .S(n12), .Z(
        \MR_int[3][29] ) );
  MUX2_X1 M1_2_28_0 ( .A(\MR_int[2][28] ), .B(\MR_int[2][0] ), .S(n12), .Z(
        \MR_int[3][28] ) );
  MUX2_X1 M1_2_27_0 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n12), .Z(
        \MR_int[3][27] ) );
  MUX2_X1 M1_2_26_0 ( .A(\MR_int[2][26] ), .B(\MR_int[2][30] ), .S(n12), .Z(
        \MR_int[3][26] ) );
  MUX2_X1 M1_2_25_0 ( .A(\MR_int[2][25] ), .B(\MR_int[2][29] ), .S(n12), .Z(
        \MR_int[3][25] ) );
  MUX2_X1 M1_2_24_0 ( .A(\MR_int[2][24] ), .B(\MR_int[2][28] ), .S(n12), .Z(
        \MR_int[3][24] ) );
  MUX2_X1 M1_2_23_0 ( .A(\MR_int[2][23] ), .B(\MR_int[2][27] ), .S(n12), .Z(
        \MR_int[3][23] ) );
  MUX2_X1 M1_2_22_0 ( .A(\MR_int[2][22] ), .B(\MR_int[2][26] ), .S(n12), .Z(
        \MR_int[3][22] ) );
  MUX2_X1 M1_2_21_0 ( .A(\MR_int[2][21] ), .B(\MR_int[2][25] ), .S(n11), .Z(
        \MR_int[3][21] ) );
  MUX2_X1 M1_2_20_0 ( .A(\MR_int[2][20] ), .B(\MR_int[2][24] ), .S(n11), .Z(
        \MR_int[3][20] ) );
  MUX2_X1 M1_2_19_0 ( .A(\MR_int[2][19] ), .B(\MR_int[2][23] ), .S(n11), .Z(
        \MR_int[3][19] ) );
  MUX2_X1 M1_2_18_0 ( .A(\MR_int[2][18] ), .B(\MR_int[2][22] ), .S(n11), .Z(
        \MR_int[3][18] ) );
  MUX2_X1 M1_2_17_0 ( .A(\MR_int[2][17] ), .B(\MR_int[2][21] ), .S(n11), .Z(
        \MR_int[3][17] ) );
  MUX2_X1 M1_2_16_0 ( .A(\MR_int[2][16] ), .B(\MR_int[2][20] ), .S(n11), .Z(
        \MR_int[3][16] ) );
  MUX2_X1 M1_2_15_0 ( .A(\MR_int[2][15] ), .B(\MR_int[2][19] ), .S(n11), .Z(
        \MR_int[3][15] ) );
  MUX2_X1 M1_2_14_0 ( .A(\MR_int[2][14] ), .B(\MR_int[2][18] ), .S(n11), .Z(
        \MR_int[3][14] ) );
  MUX2_X1 M1_2_13_0 ( .A(\MR_int[2][13] ), .B(\MR_int[2][17] ), .S(n11), .Z(
        \MR_int[3][13] ) );
  MUX2_X1 M1_2_12_0 ( .A(\MR_int[2][12] ), .B(\MR_int[2][16] ), .S(n11), .Z(
        \MR_int[3][12] ) );
  MUX2_X1 M1_2_11_0 ( .A(\MR_int[2][11] ), .B(\MR_int[2][15] ), .S(n11), .Z(
        \MR_int[3][11] ) );
  MUX2_X1 M1_2_10_0 ( .A(\MR_int[2][10] ), .B(\MR_int[2][14] ), .S(n10), .Z(
        \MR_int[3][10] ) );
  MUX2_X1 M1_2_9_0 ( .A(\MR_int[2][9] ), .B(\MR_int[2][13] ), .S(n10), .Z(
        \MR_int[3][9] ) );
  MUX2_X1 M1_2_8_0 ( .A(\MR_int[2][8] ), .B(\MR_int[2][12] ), .S(n10), .Z(
        \MR_int[3][8] ) );
  MUX2_X1 M1_2_7_0 ( .A(\MR_int[2][7] ), .B(\MR_int[2][11] ), .S(n10), .Z(
        \MR_int[3][7] ) );
  MUX2_X1 M1_2_6_0 ( .A(\MR_int[2][6] ), .B(\MR_int[2][10] ), .S(n10), .Z(
        \MR_int[3][6] ) );
  MUX2_X1 M1_2_5_0 ( .A(\MR_int[2][5] ), .B(\MR_int[2][9] ), .S(n10), .Z(
        \MR_int[3][5] ) );
  MUX2_X1 M1_2_4_0 ( .A(\MR_int[2][4] ), .B(\MR_int[2][8] ), .S(n10), .Z(
        \MR_int[3][4] ) );
  MUX2_X1 M1_2_3 ( .A(\MR_int[2][3] ), .B(\MR_int[2][7] ), .S(n10), .Z(
        \MR_int[3][3] ) );
  MUX2_X1 M1_2_2 ( .A(\MR_int[2][2] ), .B(\MR_int[2][6] ), .S(n10), .Z(
        \MR_int[3][2] ) );
  MUX2_X1 M1_2_1 ( .A(\MR_int[2][1] ), .B(\MR_int[2][5] ), .S(n10), .Z(
        \MR_int[3][1] ) );
  MUX2_X1 M1_2_0 ( .A(\MR_int[2][0] ), .B(\MR_int[2][4] ), .S(n10), .Z(
        \MR_int[3][0] ) );
  MUX2_X1 M1_1_31_0 ( .A(\MR_int[1][31] ), .B(\MR_int[1][1] ), .S(n9), .Z(
        \MR_int[2][31] ) );
  MUX2_X1 M1_1_30_0 ( .A(\MR_int[1][30] ), .B(\MR_int[1][0] ), .S(n9), .Z(
        \MR_int[2][30] ) );
  MUX2_X1 M1_1_29_0 ( .A(\MR_int[1][29] ), .B(\MR_int[1][31] ), .S(n9), .Z(
        \MR_int[2][29] ) );
  MUX2_X1 M1_1_28_0 ( .A(\MR_int[1][28] ), .B(\MR_int[1][30] ), .S(n9), .Z(
        \MR_int[2][28] ) );
  MUX2_X1 M1_1_27_0 ( .A(\MR_int[1][27] ), .B(\MR_int[1][29] ), .S(n9), .Z(
        \MR_int[2][27] ) );
  MUX2_X1 M1_1_26_0 ( .A(\MR_int[1][26] ), .B(\MR_int[1][28] ), .S(n9), .Z(
        \MR_int[2][26] ) );
  MUX2_X1 M1_1_25_0 ( .A(\MR_int[1][25] ), .B(\MR_int[1][27] ), .S(n9), .Z(
        \MR_int[2][25] ) );
  MUX2_X1 M1_1_24_0 ( .A(\MR_int[1][24] ), .B(\MR_int[1][26] ), .S(n9), .Z(
        \MR_int[2][24] ) );
  MUX2_X1 M1_1_23_0 ( .A(\MR_int[1][23] ), .B(\MR_int[1][25] ), .S(n9), .Z(
        \MR_int[2][23] ) );
  MUX2_X1 M1_1_22_0 ( .A(\MR_int[1][22] ), .B(\MR_int[1][24] ), .S(n9), .Z(
        \MR_int[2][22] ) );
  MUX2_X1 M1_1_21_0 ( .A(\MR_int[1][21] ), .B(\MR_int[1][23] ), .S(n8), .Z(
        \MR_int[2][21] ) );
  MUX2_X1 M1_1_20_0 ( .A(\MR_int[1][20] ), .B(\MR_int[1][22] ), .S(n8), .Z(
        \MR_int[2][20] ) );
  MUX2_X1 M1_1_19_0 ( .A(\MR_int[1][19] ), .B(\MR_int[1][21] ), .S(n8), .Z(
        \MR_int[2][19] ) );
  MUX2_X1 M1_1_18_0 ( .A(\MR_int[1][18] ), .B(\MR_int[1][20] ), .S(n8), .Z(
        \MR_int[2][18] ) );
  MUX2_X1 M1_1_17_0 ( .A(\MR_int[1][17] ), .B(\MR_int[1][19] ), .S(n8), .Z(
        \MR_int[2][17] ) );
  MUX2_X1 M1_1_16_0 ( .A(\MR_int[1][16] ), .B(\MR_int[1][18] ), .S(n8), .Z(
        \MR_int[2][16] ) );
  MUX2_X1 M1_1_15_0 ( .A(\MR_int[1][15] ), .B(\MR_int[1][17] ), .S(n8), .Z(
        \MR_int[2][15] ) );
  MUX2_X1 M1_1_14_0 ( .A(\MR_int[1][14] ), .B(\MR_int[1][16] ), .S(n8), .Z(
        \MR_int[2][14] ) );
  MUX2_X1 M1_1_13_0 ( .A(\MR_int[1][13] ), .B(\MR_int[1][15] ), .S(n8), .Z(
        \MR_int[2][13] ) );
  MUX2_X1 M1_1_12_0 ( .A(\MR_int[1][12] ), .B(\MR_int[1][14] ), .S(n8), .Z(
        \MR_int[2][12] ) );
  MUX2_X1 M1_1_11_0 ( .A(\MR_int[1][11] ), .B(\MR_int[1][13] ), .S(n8), .Z(
        \MR_int[2][11] ) );
  MUX2_X1 M1_1_10_0 ( .A(\MR_int[1][10] ), .B(\MR_int[1][12] ), .S(n7), .Z(
        \MR_int[2][10] ) );
  MUX2_X1 M1_1_9_0 ( .A(\MR_int[1][9] ), .B(\MR_int[1][11] ), .S(n7), .Z(
        \MR_int[2][9] ) );
  MUX2_X1 M1_1_8_0 ( .A(\MR_int[1][8] ), .B(\MR_int[1][10] ), .S(n7), .Z(
        \MR_int[2][8] ) );
  MUX2_X1 M1_1_7_0 ( .A(\MR_int[1][7] ), .B(\MR_int[1][9] ), .S(n7), .Z(
        \MR_int[2][7] ) );
  MUX2_X1 M1_1_6_0 ( .A(\MR_int[1][6] ), .B(\MR_int[1][8] ), .S(n7), .Z(
        \MR_int[2][6] ) );
  MUX2_X1 M1_1_5_0 ( .A(\MR_int[1][5] ), .B(\MR_int[1][7] ), .S(n7), .Z(
        \MR_int[2][5] ) );
  MUX2_X1 M1_1_4_0 ( .A(\MR_int[1][4] ), .B(\MR_int[1][6] ), .S(n7), .Z(
        \MR_int[2][4] ) );
  MUX2_X1 M1_1_3_0 ( .A(\MR_int[1][3] ), .B(\MR_int[1][5] ), .S(n7), .Z(
        \MR_int[2][3] ) );
  MUX2_X1 M1_1_2_0 ( .A(\MR_int[1][2] ), .B(\MR_int[1][4] ), .S(n7), .Z(
        \MR_int[2][2] ) );
  MUX2_X1 M1_1_1 ( .A(\MR_int[1][1] ), .B(\MR_int[1][3] ), .S(n7), .Z(
        \MR_int[2][1] ) );
  MUX2_X1 M1_1_0 ( .A(\MR_int[1][0] ), .B(\MR_int[1][2] ), .S(n7), .Z(
        \MR_int[2][0] ) );
  MUX2_X1 M1_0_31_0 ( .A(A[31]), .B(A[0]), .S(n6), .Z(\MR_int[1][31] ) );
  MUX2_X1 M1_0_30_0 ( .A(A[30]), .B(A[31]), .S(n6), .Z(\MR_int[1][30] ) );
  MUX2_X1 M1_0_29_0 ( .A(A[29]), .B(A[30]), .S(n6), .Z(\MR_int[1][29] ) );
  MUX2_X1 M1_0_28_0 ( .A(A[28]), .B(A[29]), .S(n6), .Z(\MR_int[1][28] ) );
  MUX2_X1 M1_0_27_0 ( .A(A[27]), .B(A[28]), .S(n6), .Z(\MR_int[1][27] ) );
  MUX2_X1 M1_0_26_0 ( .A(A[26]), .B(A[27]), .S(n6), .Z(\MR_int[1][26] ) );
  MUX2_X1 M1_0_25_0 ( .A(A[25]), .B(A[26]), .S(n6), .Z(\MR_int[1][25] ) );
  MUX2_X1 M1_0_24_0 ( .A(A[24]), .B(A[25]), .S(n6), .Z(\MR_int[1][24] ) );
  MUX2_X1 M1_0_23_0 ( .A(A[23]), .B(A[24]), .S(n6), .Z(\MR_int[1][23] ) );
  MUX2_X1 M1_0_22_0 ( .A(A[22]), .B(A[23]), .S(n6), .Z(\MR_int[1][22] ) );
  MUX2_X1 M1_0_21_0 ( .A(A[21]), .B(A[22]), .S(n5), .Z(\MR_int[1][21] ) );
  MUX2_X1 M1_0_20_0 ( .A(A[20]), .B(A[21]), .S(n5), .Z(\MR_int[1][20] ) );
  MUX2_X1 M1_0_19_0 ( .A(A[19]), .B(A[20]), .S(n5), .Z(\MR_int[1][19] ) );
  MUX2_X1 M1_0_18_0 ( .A(A[18]), .B(A[19]), .S(n5), .Z(\MR_int[1][18] ) );
  MUX2_X1 M1_0_17_0 ( .A(A[17]), .B(A[18]), .S(n5), .Z(\MR_int[1][17] ) );
  MUX2_X1 M1_0_16_0 ( .A(A[16]), .B(A[17]), .S(n5), .Z(\MR_int[1][16] ) );
  MUX2_X1 M1_0_15_0 ( .A(A[15]), .B(A[16]), .S(n5), .Z(\MR_int[1][15] ) );
  MUX2_X1 M1_0_14_0 ( .A(A[14]), .B(A[15]), .S(n5), .Z(\MR_int[1][14] ) );
  MUX2_X1 M1_0_13_0 ( .A(A[13]), .B(A[14]), .S(n5), .Z(\MR_int[1][13] ) );
  MUX2_X1 M1_0_12_0 ( .A(A[12]), .B(A[13]), .S(n5), .Z(\MR_int[1][12] ) );
  MUX2_X1 M1_0_11_0 ( .A(A[11]), .B(A[12]), .S(n5), .Z(\MR_int[1][11] ) );
  MUX2_X1 M1_0_10_0 ( .A(A[10]), .B(A[11]), .S(n4), .Z(\MR_int[1][10] ) );
  MUX2_X1 M1_0_9_0 ( .A(A[9]), .B(A[10]), .S(n4), .Z(\MR_int[1][9] ) );
  MUX2_X1 M1_0_8_0 ( .A(A[8]), .B(A[9]), .S(n4), .Z(\MR_int[1][8] ) );
  MUX2_X1 M1_0_7_0 ( .A(A[7]), .B(A[8]), .S(n4), .Z(\MR_int[1][7] ) );
  MUX2_X1 M1_0_6_0 ( .A(A[6]), .B(A[7]), .S(n4), .Z(\MR_int[1][6] ) );
  MUX2_X1 M1_0_5_0 ( .A(A[5]), .B(A[6]), .S(n4), .Z(\MR_int[1][5] ) );
  MUX2_X1 M1_0_4_0 ( .A(A[4]), .B(A[5]), .S(n4), .Z(\MR_int[1][4] ) );
  MUX2_X1 M1_0_3_0 ( .A(A[3]), .B(A[4]), .S(n4), .Z(\MR_int[1][3] ) );
  MUX2_X1 M1_0_2_0 ( .A(A[2]), .B(A[3]), .S(n4), .Z(\MR_int[1][2] ) );
  MUX2_X1 M1_0_1_0 ( .A(A[1]), .B(A[2]), .S(n4), .Z(\MR_int[1][1] ) );
  MUX2_X1 M1_0_0 ( .A(A[0]), .B(A[1]), .S(n4), .Z(\MR_int[1][0] ) );
  BUF_X1 U2 ( .A(SH[3]), .Z(n14) );
  BUF_X1 U3 ( .A(SH[3]), .Z(n13) );
  BUF_X1 U4 ( .A(SH[4]), .Z(n16) );
  BUF_X1 U5 ( .A(SH[4]), .Z(n17) );
  BUF_X1 U6 ( .A(SH[3]), .Z(n15) );
  BUF_X1 U7 ( .A(SH[4]), .Z(n18) );
  BUF_X1 U8 ( .A(SH[0]), .Z(n5) );
  BUF_X1 U9 ( .A(SH[0]), .Z(n4) );
  BUF_X1 U10 ( .A(SH[1]), .Z(n8) );
  BUF_X1 U11 ( .A(SH[1]), .Z(n7) );
  BUF_X1 U12 ( .A(SH[2]), .Z(n11) );
  BUF_X1 U13 ( .A(SH[2]), .Z(n10) );
  BUF_X1 U14 ( .A(SH[0]), .Z(n6) );
  BUF_X1 U15 ( .A(SH[1]), .Z(n9) );
  BUF_X1 U16 ( .A(SH[2]), .Z(n12) );
endmodule


module SHIFTER_GENERIC_N32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE, 
        OUTPUT );
  input [31:0] A;
  input [4:0] B;
  output [31:0] OUTPUT;
  input LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, n10, n11, n12, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108;

  SHIFTER_GENERIC_N32_DW01_ash_0 sll_49 ( .A(A), .DATA_TC(1'b0), .SH({n105, 
        n104, B[2:0]}), .SH_TC(1'b0), .B({N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, 
        N235, N234}) );
  SHIFTER_GENERIC_N32_DW_sla_0 sla_47 ( .A(A), .SH({n105, n104, B[2:0]}), 
        .SH_TC(1'b0), .B({N233, N232, N231, N230, N229, N228, N227, N226, N225, 
        N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, 
        N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202}) );
  SHIFTER_GENERIC_N32_DW_rash_0 srl_42 ( .A(A), .DATA_TC(1'b0), .SH({n105, 
        n104, B[2:0]}), .SH_TC(1'b0), .B({N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, 
        N138, N137}) );
  SHIFTER_GENERIC_N32_DW_sra_0 sra_40 ( .A(A), .SH({n105, n104, B[2:0]}), 
        .SH_TC(1'b0), .B({N136, N135, N134, N133, N132, N131, N130, N129, N128, 
        N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, 
        N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105}) );
  SHIFTER_GENERIC_N32_DW_lbsh_0 rol_33 ( .A(A), .SH({n105, n104, B[2:0]}), 
        .SH_TC(1'b0), .B({N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, 
        N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, 
        N46, N45, N44, N43, N42, N41, N40, N39}) );
  SHIFTER_GENERIC_N32_DW_rbsh_0 ror_31 ( .A(A), .SH({n105, n104, B[2:0]}), 
        .SH_TC(1'b0), .B({N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7}) );
  BUF_X1 U1 ( .A(B[3]), .Z(n104) );
  AOI222_X1 U2 ( .A1(N232), .A2(n103), .B1(N135), .B2(n99), .C1(N167), .C2(n96), .ZN(n39) );
  AOI222_X1 U3 ( .A1(N231), .A2(n102), .B1(N134), .B2(n99), .C1(N166), .C2(n96), .ZN(n43) );
  AOI222_X1 U4 ( .A1(N230), .A2(n102), .B1(N133), .B2(n99), .C1(N165), .C2(n96), .ZN(n45) );
  AOI222_X1 U11 ( .A1(N229), .A2(n102), .B1(N132), .B2(n99), .C1(N164), .C2(
        n96), .ZN(n47) );
  AOI222_X1 U12 ( .A1(N228), .A2(n102), .B1(N131), .B2(n99), .C1(N163), .C2(
        n96), .ZN(n49) );
  AOI222_X1 U13 ( .A1(N227), .A2(n102), .B1(N130), .B2(n99), .C1(N162), .C2(
        n96), .ZN(n51) );
  AOI222_X1 U14 ( .A1(N226), .A2(n102), .B1(N129), .B2(n99), .C1(N161), .C2(
        n96), .ZN(n53) );
  AOI222_X1 U15 ( .A1(N225), .A2(n102), .B1(N128), .B2(n99), .C1(N160), .C2(
        n96), .ZN(n55) );
  AOI222_X1 U16 ( .A1(N224), .A2(n102), .B1(N127), .B2(n99), .C1(N159), .C2(
        n96), .ZN(n57) );
  AOI222_X1 U17 ( .A1(N223), .A2(n102), .B1(N126), .B2(n99), .C1(N158), .C2(
        n96), .ZN(n59) );
  AOI222_X1 U18 ( .A1(N222), .A2(n102), .B1(N125), .B2(n99), .C1(N157), .C2(
        n96), .ZN(n61) );
  AOI222_X1 U19 ( .A1(N221), .A2(n101), .B1(N124), .B2(n98), .C1(N156), .C2(
        n95), .ZN(n65) );
  AOI222_X1 U20 ( .A1(N220), .A2(n101), .B1(N123), .B2(n98), .C1(N155), .C2(
        n95), .ZN(n67) );
  AOI222_X1 U21 ( .A1(N219), .A2(n101), .B1(N122), .B2(n98), .C1(N154), .C2(
        n95), .ZN(n69) );
  AOI222_X1 U22 ( .A1(N218), .A2(n101), .B1(N121), .B2(n98), .C1(N153), .C2(
        n95), .ZN(n71) );
  AOI222_X1 U23 ( .A1(N217), .A2(n101), .B1(N120), .B2(n98), .C1(N152), .C2(
        n95), .ZN(n73) );
  AOI222_X1 U24 ( .A1(N216), .A2(n101), .B1(N119), .B2(n98), .C1(N151), .C2(
        n95), .ZN(n75) );
  AOI222_X1 U25 ( .A1(N215), .A2(n101), .B1(N118), .B2(n98), .C1(N150), .C2(
        n95), .ZN(n77) );
  AOI222_X1 U26 ( .A1(N214), .A2(n101), .B1(N117), .B2(n98), .C1(N149), .C2(
        n95), .ZN(n79) );
  AOI222_X1 U27 ( .A1(N213), .A2(n101), .B1(N116), .B2(n98), .C1(N148), .C2(
        n95), .ZN(n81) );
  AOI222_X1 U28 ( .A1(N212), .A2(n101), .B1(N115), .B2(n98), .C1(N147), .C2(
        n95), .ZN(n83) );
  AOI222_X1 U29 ( .A1(N204), .A2(n103), .B1(N107), .B2(n99), .C1(N139), .C2(
        n96), .ZN(n41) );
  AOI222_X1 U30 ( .A1(N203), .A2(n102), .B1(N106), .B2(n98), .C1(N138), .C2(
        n95), .ZN(n63) );
  AOI222_X1 U31 ( .A1(N211), .A2(n103), .B1(N114), .B2(n100), .C1(N146), .C2(
        n97), .ZN(n11) );
  AOI222_X1 U32 ( .A1(N210), .A2(n103), .B1(N113), .B2(n100), .C1(N145), .C2(
        n97), .ZN(n25) );
  AOI222_X1 U33 ( .A1(N209), .A2(n103), .B1(N112), .B2(n100), .C1(N144), .C2(
        n97), .ZN(n27) );
  AOI222_X1 U34 ( .A1(N208), .A2(n103), .B1(N111), .B2(n100), .C1(N143), .C2(
        n97), .ZN(n29) );
  AOI222_X1 U35 ( .A1(N207), .A2(n103), .B1(N110), .B2(n100), .C1(N142), .C2(
        n97), .ZN(n31) );
  AOI222_X1 U36 ( .A1(N206), .A2(n103), .B1(N109), .B2(n100), .C1(N141), .C2(
        n97), .ZN(n33) );
  AOI222_X1 U37 ( .A1(N205), .A2(n103), .B1(N108), .B2(n100), .C1(N140), .C2(
        n97), .ZN(n35) );
  AOI222_X1 U38 ( .A1(N69), .A2(n94), .B1(N264), .B2(n90), .C1(N37), .C2(n87), 
        .ZN(n38) );
  AOI222_X1 U39 ( .A1(N68), .A2(n93), .B1(N263), .B2(n90), .C1(N36), .C2(n87), 
        .ZN(n42) );
  AOI222_X1 U40 ( .A1(N67), .A2(n93), .B1(N262), .B2(n90), .C1(N35), .C2(n87), 
        .ZN(n44) );
  AOI222_X1 U41 ( .A1(N66), .A2(n93), .B1(N261), .B2(n90), .C1(N34), .C2(n87), 
        .ZN(n46) );
  AOI222_X1 U42 ( .A1(N65), .A2(n93), .B1(N260), .B2(n90), .C1(N33), .C2(n87), 
        .ZN(n48) );
  AOI222_X1 U43 ( .A1(N64), .A2(n93), .B1(N259), .B2(n90), .C1(N32), .C2(n87), 
        .ZN(n50) );
  AOI222_X1 U44 ( .A1(N63), .A2(n93), .B1(N258), .B2(n90), .C1(N31), .C2(n87), 
        .ZN(n52) );
  AOI222_X1 U45 ( .A1(N62), .A2(n93), .B1(N257), .B2(n90), .C1(N30), .C2(n87), 
        .ZN(n54) );
  AOI222_X1 U46 ( .A1(N61), .A2(n93), .B1(N256), .B2(n90), .C1(N29), .C2(n87), 
        .ZN(n56) );
  AOI222_X1 U47 ( .A1(N60), .A2(n93), .B1(N255), .B2(n90), .C1(N28), .C2(n87), 
        .ZN(n58) );
  AOI222_X1 U48 ( .A1(N59), .A2(n93), .B1(N254), .B2(n90), .C1(N27), .C2(n87), 
        .ZN(n60) );
  AOI222_X1 U49 ( .A1(N58), .A2(n92), .B1(N253), .B2(n89), .C1(N26), .C2(n86), 
        .ZN(n64) );
  AOI222_X1 U50 ( .A1(N57), .A2(n92), .B1(N252), .B2(n89), .C1(N25), .C2(n86), 
        .ZN(n66) );
  AOI222_X1 U51 ( .A1(N56), .A2(n92), .B1(N251), .B2(n89), .C1(N24), .C2(n86), 
        .ZN(n68) );
  AOI222_X1 U52 ( .A1(N55), .A2(n92), .B1(N250), .B2(n89), .C1(N23), .C2(n86), 
        .ZN(n70) );
  AOI222_X1 U53 ( .A1(N54), .A2(n92), .B1(N249), .B2(n89), .C1(N22), .C2(n86), 
        .ZN(n72) );
  AOI222_X1 U54 ( .A1(N53), .A2(n92), .B1(N248), .B2(n89), .C1(N21), .C2(n86), 
        .ZN(n74) );
  AOI222_X1 U55 ( .A1(N52), .A2(n92), .B1(N247), .B2(n89), .C1(N20), .C2(n86), 
        .ZN(n76) );
  AOI222_X1 U56 ( .A1(N51), .A2(n92), .B1(N246), .B2(n89), .C1(N19), .C2(n86), 
        .ZN(n78) );
  AOI222_X1 U57 ( .A1(N50), .A2(n92), .B1(N245), .B2(n89), .C1(N18), .C2(n86), 
        .ZN(n80) );
  AOI222_X1 U58 ( .A1(N49), .A2(n92), .B1(N244), .B2(n89), .C1(N17), .C2(n86), 
        .ZN(n82) );
  AOI222_X1 U59 ( .A1(N41), .A2(n94), .B1(N236), .B2(n90), .C1(N9), .C2(n87), 
        .ZN(n40) );
  AOI222_X1 U60 ( .A1(N40), .A2(n93), .B1(N235), .B2(n89), .C1(N8), .C2(n86), 
        .ZN(n62) );
  AOI222_X1 U61 ( .A1(N39), .A2(n92), .B1(N234), .B2(n89), .C1(N7), .C2(n86), 
        .ZN(n84) );
  AOI222_X1 U62 ( .A1(N70), .A2(n94), .B1(N265), .B2(n91), .C1(N38), .C2(n88), 
        .ZN(n36) );
  AOI222_X1 U63 ( .A1(N48), .A2(n94), .B1(N243), .B2(n91), .C1(N16), .C2(n88), 
        .ZN(n10) );
  AOI222_X1 U64 ( .A1(N47), .A2(n94), .B1(N242), .B2(n91), .C1(N15), .C2(n88), 
        .ZN(n24) );
  AOI222_X1 U65 ( .A1(N46), .A2(n94), .B1(N241), .B2(n91), .C1(N14), .C2(n88), 
        .ZN(n26) );
  AOI222_X1 U66 ( .A1(N45), .A2(n94), .B1(N240), .B2(n91), .C1(N13), .C2(n88), 
        .ZN(n28) );
  AOI222_X1 U67 ( .A1(N44), .A2(n94), .B1(N239), .B2(n91), .C1(N12), .C2(n88), 
        .ZN(n30) );
  AOI222_X1 U68 ( .A1(N43), .A2(n94), .B1(N238), .B2(n91), .C1(N11), .C2(n88), 
        .ZN(n32) );
  AOI222_X1 U69 ( .A1(N42), .A2(n94), .B1(N237), .B2(n91), .C1(N10), .C2(n88), 
        .ZN(n34) );
  BUF_X1 U70 ( .A(n22), .Z(n90) );
  BUF_X1 U71 ( .A(n22), .Z(n89) );
  BUF_X1 U72 ( .A(n22), .Z(n91) );
  BUF_X1 U73 ( .A(B[4]), .Z(n105) );
  NAND2_X1 U74 ( .A1(n36), .A2(n37), .ZN(OUTPUT[31]) );
  NAND2_X1 U75 ( .A1(n38), .A2(n39), .ZN(OUTPUT[30]) );
  NAND2_X1 U76 ( .A1(n42), .A2(n43), .ZN(OUTPUT[29]) );
  NAND2_X1 U77 ( .A1(n44), .A2(n45), .ZN(OUTPUT[28]) );
  NAND2_X1 U78 ( .A1(n46), .A2(n47), .ZN(OUTPUT[27]) );
  NAND2_X1 U79 ( .A1(n48), .A2(n49), .ZN(OUTPUT[26]) );
  NAND2_X1 U80 ( .A1(n50), .A2(n51), .ZN(OUTPUT[25]) );
  NAND2_X1 U81 ( .A1(n52), .A2(n53), .ZN(OUTPUT[24]) );
  NAND2_X1 U82 ( .A1(n54), .A2(n55), .ZN(OUTPUT[23]) );
  NAND2_X1 U83 ( .A1(n56), .A2(n57), .ZN(OUTPUT[22]) );
  NAND2_X1 U84 ( .A1(n58), .A2(n59), .ZN(OUTPUT[21]) );
  NAND2_X1 U85 ( .A1(n60), .A2(n61), .ZN(OUTPUT[20]) );
  NAND2_X1 U86 ( .A1(n64), .A2(n65), .ZN(OUTPUT[19]) );
  NAND2_X1 U87 ( .A1(n66), .A2(n67), .ZN(OUTPUT[18]) );
  NAND2_X1 U88 ( .A1(n68), .A2(n69), .ZN(OUTPUT[17]) );
  NAND2_X1 U89 ( .A1(n70), .A2(n71), .ZN(OUTPUT[16]) );
  NAND2_X1 U90 ( .A1(n72), .A2(n73), .ZN(OUTPUT[15]) );
  NAND2_X1 U91 ( .A1(n74), .A2(n75), .ZN(OUTPUT[14]) );
  NAND2_X1 U92 ( .A1(n76), .A2(n77), .ZN(OUTPUT[13]) );
  NAND2_X1 U93 ( .A1(n78), .A2(n79), .ZN(OUTPUT[12]) );
  NAND2_X1 U94 ( .A1(n80), .A2(n81), .ZN(OUTPUT[11]) );
  NAND2_X1 U95 ( .A1(n82), .A2(n83), .ZN(OUTPUT[10]) );
  NAND2_X1 U96 ( .A1(n10), .A2(n11), .ZN(OUTPUT[9]) );
  NAND2_X1 U97 ( .A1(n24), .A2(n25), .ZN(OUTPUT[8]) );
  NAND2_X1 U98 ( .A1(n26), .A2(n27), .ZN(OUTPUT[7]) );
  NAND2_X1 U99 ( .A1(n28), .A2(n29), .ZN(OUTPUT[6]) );
  NAND2_X1 U100 ( .A1(n30), .A2(n31), .ZN(OUTPUT[5]) );
  NAND2_X1 U101 ( .A1(n32), .A2(n33), .ZN(OUTPUT[4]) );
  AOI222_X1 U102 ( .A1(N202), .A2(n101), .B1(N105), .B2(n98), .C1(N137), .C2(
        n95), .ZN(n85) );
  AOI222_X1 U103 ( .A1(N233), .A2(n103), .B1(N136), .B2(n100), .C1(N168), .C2(
        n97), .ZN(n37) );
  BUF_X1 U104 ( .A(n19), .Z(n99) );
  BUF_X1 U105 ( .A(n19), .Z(n98) );
  BUF_X1 U106 ( .A(n20), .Z(n96) );
  BUF_X1 U107 ( .A(n20), .Z(n95) );
  BUF_X1 U108 ( .A(n23), .Z(n87) );
  BUF_X1 U109 ( .A(n23), .Z(n86) );
  BUF_X1 U110 ( .A(n12), .Z(n102) );
  BUF_X1 U111 ( .A(n12), .Z(n101) );
  BUF_X1 U112 ( .A(n21), .Z(n93) );
  BUF_X1 U113 ( .A(n21), .Z(n92) );
  NOR3_X1 U114 ( .A1(n106), .A2(n108), .A3(n107), .ZN(n22) );
  BUF_X1 U115 ( .A(n12), .Z(n103) );
  BUF_X1 U116 ( .A(n21), .Z(n94) );
  BUF_X1 U117 ( .A(n19), .Z(n100) );
  BUF_X1 U118 ( .A(n20), .Z(n97) );
  BUF_X1 U119 ( .A(n23), .Z(n88) );
  NAND2_X1 U120 ( .A1(n34), .A2(n35), .ZN(OUTPUT[3]) );
  NAND2_X1 U121 ( .A1(n40), .A2(n41), .ZN(OUTPUT[2]) );
  NAND2_X1 U122 ( .A1(n62), .A2(n63), .ZN(OUTPUT[1]) );
  NOR3_X1 U123 ( .A1(n108), .A2(LEFT_RIGHT), .A3(n106), .ZN(n20) );
  NOR3_X1 U124 ( .A1(LEFT_RIGHT), .A2(LOGIC_ARITH), .A3(n108), .ZN(n19) );
  NOR3_X1 U125 ( .A1(n108), .A2(LOGIC_ARITH), .A3(n107), .ZN(n12) );
  NOR2_X1 U126 ( .A1(LEFT_RIGHT), .A2(SHIFT_ROTATE), .ZN(n23) );
  NOR2_X1 U127 ( .A1(n107), .A2(SHIFT_ROTATE), .ZN(n21) );
  INV_X1 U128 ( .A(LEFT_RIGHT), .ZN(n107) );
  INV_X1 U129 ( .A(LOGIC_ARITH), .ZN(n106) );
  NAND2_X1 U130 ( .A1(n84), .A2(n85), .ZN(OUTPUT[0]) );
  INV_X1 U131 ( .A(SHIFT_ROTATE), .ZN(n108) );
endmodule


module G_0 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_43 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_0 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_0 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_43 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_0 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_52 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module G_42 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_42 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_42 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_42 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_42 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_41 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_41 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_41 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_41 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_41 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_40 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_40 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_40 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_40 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_40 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_39 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_39 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_39 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_39 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_39 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_38 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_38 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_38 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_38 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_38 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_37 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_37 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_37 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_37 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_37 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_36 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_36 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_36 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_36 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_36 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_35 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_35 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_35 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_35 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_35 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_34 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_34 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_34 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_34 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_34 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_33 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_33 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_33 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_33 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_33 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_32 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_32 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_32 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_32 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_32 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_31 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_31 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_31 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_31 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_31 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_30 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_30 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_30 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_30 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_30 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_29 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_29 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_29 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_29 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_29 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_28 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_28 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_28 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_28 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_28 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_27 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_27 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_27 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_27 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_27 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_26 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_26 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_26 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_26 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_26 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_25 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_25 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_25 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_25 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_25 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_24 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_24 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_24 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_24 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_24 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_23 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_23 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_23 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_23 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_23 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_22 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_22 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_22 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_22 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_22 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_21 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_21 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_21 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_21 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_21 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_20 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_20 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_20 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_20 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_20 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_19 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_19 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_19 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_19 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_19 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_18 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_18 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_18 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_18 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_18 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_17 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_17 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_17 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_17 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_17 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_16 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_16 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_16 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_16 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_16 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_15 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_15 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_15 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_15 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_15 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_14 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_14 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_14 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_14 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_14 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_13 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_13 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_13 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_13 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_13 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_51 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module G_12 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_12 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_12 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_12 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_12 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_11 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_11 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_11 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_11 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_11 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_10 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_10 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_10 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_10 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_10 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_9 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_9 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_9 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_9 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_9 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_8 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_8 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_8 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_8 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_8 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_7 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_7 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_7 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_7 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_7 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_6 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_6 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_6 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_6 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_6 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_50 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module G_5 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_5 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_5 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_5 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_5 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_4 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_4 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_4 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_4 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_4 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_3 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_3 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_3 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_3 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_3 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_49 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module G_48 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module G_2 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_2 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_2 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_2 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_2 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_1 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module P_1 ( p1, P2, Co );
  input p1, P2;
  output Co;


  AND2_X1 U1 ( .A1(p1), .A2(P2), .ZN(Co) );
endmodule


module PG_1 ( G1, P1, G2, P2, gout, pout );
  input G1, P1, G2, P2;
  output gout, pout;


  G_1 g_comp ( .G1(G1), .P(P1), .G2(G2), .Co(gout) );
  P_1 p_comp ( .p1(P1), .P2(P2), .Co(pout) );
endmodule


module G_47 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module G_46 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module G_45 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module G_44 ( G1, P, G2, Co );
  input G1, P, G2;
  output Co;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI21_X1 U2 ( .B1(P), .B2(G2), .A(G1), .ZN(n4) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   \gi[32][4] , \gi[32][3] , \gi[32][2] , \gi[32][1] , \gi[32][0] ,
         \gi[31][0] , \gi[30][0] , \gi[29][0] , \gi[28][4] , \gi[28][2] ,
         \gi[28][1] , \gi[28][0] , \gi[27][0] , \gi[26][0] , \gi[25][0] ,
         \gi[24][3] , \gi[24][2] , \gi[24][1] , \gi[24][0] , \gi[23][0] ,
         \gi[22][0] , \gi[21][0] , \gi[20][2] , \gi[20][1] , \gi[20][0] ,
         \gi[19][0] , \gi[18][0] , \gi[17][0] , \gi[16][3] , \gi[16][2] ,
         \gi[16][1] , \gi[16][0] , \gi[15][0] , \gi[14][0] , \gi[13][0] ,
         \gi[12][2] , \gi[12][1] , \gi[12][0] , \gi[11][0] , \gi[10][0] ,
         \gi[9][0] , \gi[8][2] , \gi[8][1] , \gi[8][0] , \gi[7][0] ,
         \gi[6][0] , \gi[5][0] , \gi[4][1] , \gi[4][0] , \gi[3][0] ,
         \gi[2][1] , \gi[2][0] , \gi[1][0] , \gi[0][0] , \pi[32][4] ,
         \pi[32][3] , \pi[32][2] , \pi[32][1] , \pi[32][0] , \pi[31][0] ,
         \pi[30][0] , \pi[29][0] , \pi[28][4] , \pi[28][2] , \pi[28][1] ,
         \pi[28][0] , \pi[27][0] , \pi[26][0] , \pi[25][0] , \pi[24][3] ,
         \pi[24][2] , \pi[24][1] , \pi[24][0] , \pi[23][0] , \pi[22][0] ,
         \pi[21][0] , \pi[20][2] , \pi[20][1] , \pi[20][0] , \pi[19][0] ,
         \pi[18][0] , \pi[17][0] , \pi[16][3] , \pi[16][2] , \pi[16][1] ,
         \pi[16][0] , \pi[15][0] , \pi[14][0] , \pi[13][0] , \pi[12][2] ,
         \pi[12][1] , \pi[12][0] , \pi[11][0] , \pi[10][0] , \pi[9][0] ,
         \pi[8][2] , \pi[8][1] , \pi[8][0] , \pi[7][0] , \pi[6][0] ,
         \pi[5][0] , \pi[4][1] , \pi[4][0] , \pi[3][0] , \pi[2][0] ,
         \pi[0][0] ;

  XOR2_X1 U34 ( .A(B[8]), .B(A[8]), .Z(\pi[9][0] ) );
  XOR2_X1 U35 ( .A(B[7]), .B(A[7]), .Z(\pi[8][0] ) );
  XOR2_X1 U36 ( .A(B[6]), .B(A[6]), .Z(\pi[7][0] ) );
  XOR2_X1 U37 ( .A(B[5]), .B(A[5]), .Z(\pi[6][0] ) );
  XOR2_X1 U38 ( .A(B[4]), .B(A[4]), .Z(\pi[5][0] ) );
  XOR2_X1 U39 ( .A(B[3]), .B(A[3]), .Z(\pi[4][0] ) );
  XOR2_X1 U40 ( .A(B[2]), .B(A[2]), .Z(\pi[3][0] ) );
  XOR2_X1 U41 ( .A(B[31]), .B(A[31]), .Z(\pi[32][0] ) );
  XOR2_X1 U42 ( .A(B[30]), .B(A[30]), .Z(\pi[31][0] ) );
  XOR2_X1 U43 ( .A(B[29]), .B(A[29]), .Z(\pi[30][0] ) );
  XOR2_X1 U44 ( .A(B[1]), .B(A[1]), .Z(\pi[2][0] ) );
  XOR2_X1 U45 ( .A(B[28]), .B(A[28]), .Z(\pi[29][0] ) );
  XOR2_X1 U46 ( .A(B[27]), .B(A[27]), .Z(\pi[28][0] ) );
  XOR2_X1 U47 ( .A(B[26]), .B(A[26]), .Z(\pi[27][0] ) );
  XOR2_X1 U48 ( .A(B[25]), .B(A[25]), .Z(\pi[26][0] ) );
  XOR2_X1 U49 ( .A(B[24]), .B(A[24]), .Z(\pi[25][0] ) );
  XOR2_X1 U50 ( .A(B[23]), .B(A[23]), .Z(\pi[24][0] ) );
  XOR2_X1 U51 ( .A(B[22]), .B(A[22]), .Z(\pi[23][0] ) );
  XOR2_X1 U52 ( .A(B[21]), .B(A[21]), .Z(\pi[22][0] ) );
  XOR2_X1 U53 ( .A(B[20]), .B(A[20]), .Z(\pi[21][0] ) );
  XOR2_X1 U54 ( .A(B[19]), .B(A[19]), .Z(\pi[20][0] ) );
  XOR2_X1 U55 ( .A(B[18]), .B(A[18]), .Z(\pi[19][0] ) );
  XOR2_X1 U56 ( .A(B[17]), .B(A[17]), .Z(\pi[18][0] ) );
  XOR2_X1 U57 ( .A(B[16]), .B(A[16]), .Z(\pi[17][0] ) );
  XOR2_X1 U58 ( .A(B[15]), .B(A[15]), .Z(\pi[16][0] ) );
  XOR2_X1 U59 ( .A(B[14]), .B(A[14]), .Z(\pi[15][0] ) );
  XOR2_X1 U60 ( .A(B[13]), .B(A[13]), .Z(\pi[14][0] ) );
  XOR2_X1 U61 ( .A(B[12]), .B(A[12]), .Z(\pi[13][0] ) );
  XOR2_X1 U62 ( .A(B[11]), .B(A[11]), .Z(\pi[12][0] ) );
  XOR2_X1 U63 ( .A(B[10]), .B(A[10]), .Z(\pi[11][0] ) );
  XOR2_X1 U64 ( .A(B[9]), .B(A[9]), .Z(\pi[10][0] ) );
  XOR2_X1 U65 ( .A(B[0]), .B(A[0]), .Z(\pi[0][0] ) );
  G_0 g_port0_0_1 ( .G1(\gi[0][0] ), .P(\pi[0][0] ), .G2(Cin), .Co(\gi[1][0] )
         );
  PG_0 pg_port2_1_1 ( .G1(\gi[1][0] ), .P1(1'b0), .G2(\gi[0][0] ), .P2(
        \pi[0][0] ) );
  G_52 g_port1_1_2 ( .G1(\gi[2][0] ), .P(\pi[2][0] ), .G2(\gi[1][0] ), .Co(
        \gi[2][1] ) );
  PG_42 pg_port2_1_3 ( .G1(\gi[3][0] ), .P1(\pi[3][0] ), .G2(\gi[2][0] ), .P2(
        \pi[2][0] ) );
  PG_41 pg_port2_1_4 ( .G1(\gi[4][0] ), .P1(\pi[4][0] ), .G2(\gi[3][0] ), .P2(
        \pi[3][0] ), .gout(\gi[4][1] ), .pout(\pi[4][1] ) );
  PG_40 pg_port2_1_5 ( .G1(\gi[5][0] ), .P1(\pi[5][0] ), .G2(\gi[4][0] ), .P2(
        \pi[4][0] ) );
  PG_39 pg_port2_1_6 ( .G1(\gi[6][0] ), .P1(\pi[6][0] ), .G2(\gi[5][0] ), .P2(
        \pi[5][0] ) );
  PG_38 pg_port2_1_7 ( .G1(\gi[7][0] ), .P1(\pi[7][0] ), .G2(\gi[6][0] ), .P2(
        \pi[6][0] ) );
  PG_37 pg_port2_1_8 ( .G1(\gi[8][0] ), .P1(\pi[8][0] ), .G2(\gi[7][0] ), .P2(
        \pi[7][0] ), .gout(\gi[8][1] ), .pout(\pi[8][1] ) );
  PG_36 pg_port2_1_9 ( .G1(\gi[9][0] ), .P1(\pi[9][0] ), .G2(\gi[8][0] ), .P2(
        \pi[8][0] ) );
  PG_35 pg_port2_1_10 ( .G1(\gi[10][0] ), .P1(\pi[10][0] ), .G2(\gi[9][0] ), 
        .P2(\pi[9][0] ) );
  PG_34 pg_port2_1_11 ( .G1(\gi[11][0] ), .P1(\pi[11][0] ), .G2(\gi[10][0] ), 
        .P2(\pi[10][0] ) );
  PG_33 pg_port2_1_12 ( .G1(\gi[12][0] ), .P1(\pi[12][0] ), .G2(\gi[11][0] ), 
        .P2(\pi[11][0] ), .gout(\gi[12][1] ), .pout(\pi[12][1] ) );
  PG_32 pg_port2_1_13 ( .G1(\gi[13][0] ), .P1(\pi[13][0] ), .G2(\gi[12][0] ), 
        .P2(\pi[12][0] ) );
  PG_31 pg_port2_1_14 ( .G1(\gi[14][0] ), .P1(\pi[14][0] ), .G2(\gi[13][0] ), 
        .P2(\pi[13][0] ) );
  PG_30 pg_port2_1_15 ( .G1(\gi[15][0] ), .P1(\pi[15][0] ), .G2(\gi[14][0] ), 
        .P2(\pi[14][0] ) );
  PG_29 pg_port2_1_16 ( .G1(\gi[16][0] ), .P1(\pi[16][0] ), .G2(\gi[15][0] ), 
        .P2(\pi[15][0] ), .gout(\gi[16][1] ), .pout(\pi[16][1] ) );
  PG_28 pg_port2_1_17 ( .G1(\gi[17][0] ), .P1(\pi[17][0] ), .G2(\gi[16][0] ), 
        .P2(\pi[16][0] ) );
  PG_27 pg_port2_1_18 ( .G1(\gi[18][0] ), .P1(\pi[18][0] ), .G2(\gi[17][0] ), 
        .P2(\pi[17][0] ) );
  PG_26 pg_port2_1_19 ( .G1(\gi[19][0] ), .P1(\pi[19][0] ), .G2(\gi[18][0] ), 
        .P2(\pi[18][0] ) );
  PG_25 pg_port2_1_20 ( .G1(\gi[20][0] ), .P1(\pi[20][0] ), .G2(\gi[19][0] ), 
        .P2(\pi[19][0] ), .gout(\gi[20][1] ), .pout(\pi[20][1] ) );
  PG_24 pg_port2_1_21 ( .G1(\gi[21][0] ), .P1(\pi[21][0] ), .G2(\gi[20][0] ), 
        .P2(\pi[20][0] ) );
  PG_23 pg_port2_1_22 ( .G1(\gi[22][0] ), .P1(\pi[22][0] ), .G2(\gi[21][0] ), 
        .P2(\pi[21][0] ) );
  PG_22 pg_port2_1_23 ( .G1(\gi[23][0] ), .P1(\pi[23][0] ), .G2(\gi[22][0] ), 
        .P2(\pi[22][0] ) );
  PG_21 pg_port2_1_24 ( .G1(\gi[24][0] ), .P1(\pi[24][0] ), .G2(\gi[23][0] ), 
        .P2(\pi[23][0] ), .gout(\gi[24][1] ), .pout(\pi[24][1] ) );
  PG_20 pg_port2_1_25 ( .G1(\gi[25][0] ), .P1(\pi[25][0] ), .G2(\gi[24][0] ), 
        .P2(\pi[24][0] ) );
  PG_19 pg_port2_1_26 ( .G1(\gi[26][0] ), .P1(\pi[26][0] ), .G2(\gi[25][0] ), 
        .P2(\pi[25][0] ) );
  PG_18 pg_port2_1_27 ( .G1(\gi[27][0] ), .P1(\pi[27][0] ), .G2(\gi[26][0] ), 
        .P2(\pi[26][0] ) );
  PG_17 pg_port2_1_28 ( .G1(\gi[28][0] ), .P1(\pi[28][0] ), .G2(\gi[27][0] ), 
        .P2(\pi[27][0] ), .gout(\gi[28][1] ), .pout(\pi[28][1] ) );
  PG_16 pg_port2_1_29 ( .G1(\gi[29][0] ), .P1(\pi[29][0] ), .G2(\gi[28][0] ), 
        .P2(\pi[28][0] ) );
  PG_15 pg_port2_1_30 ( .G1(\gi[30][0] ), .P1(\pi[30][0] ), .G2(\gi[29][0] ), 
        .P2(\pi[29][0] ) );
  PG_14 pg_port2_1_31 ( .G1(\gi[31][0] ), .P1(\pi[31][0] ), .G2(\gi[30][0] ), 
        .P2(\pi[30][0] ) );
  PG_13 pg_port2_1_32 ( .G1(\gi[32][0] ), .P1(\pi[32][0] ), .G2(\gi[31][0] ), 
        .P2(\pi[31][0] ), .gout(\gi[32][1] ), .pout(\pi[32][1] ) );
  G_51 g_port_0 ( .G1(\gi[4][1] ), .P(\pi[4][1] ), .G2(\gi[2][1] ), .Co(Co[0])
         );
  PG_12 pg_port2_0_1_2 ( .G1(\gi[8][1] ), .P1(\pi[8][1] ), .G2(\gi[4][1] ), 
        .P2(\pi[4][1] ), .gout(\gi[8][2] ), .pout(\pi[8][2] ) );
  PG_11 pg_port2_0_2_3 ( .G1(\gi[12][1] ), .P1(\pi[12][1] ), .G2(\gi[8][1] ), 
        .P2(\pi[8][1] ), .gout(\gi[12][2] ), .pout(\pi[12][2] ) );
  PG_10 pg_port2_0_3_4 ( .G1(\gi[16][1] ), .P1(\pi[16][1] ), .G2(\gi[12][1] ), 
        .P2(\pi[12][1] ), .gout(\gi[16][2] ), .pout(\pi[16][2] ) );
  PG_9 pg_port2_0_4_5 ( .G1(\gi[20][1] ), .P1(\pi[20][1] ), .G2(\gi[16][1] ), 
        .P2(\pi[16][1] ), .gout(\gi[20][2] ), .pout(\pi[20][2] ) );
  PG_8 pg_port2_0_5_6 ( .G1(\gi[24][1] ), .P1(\pi[24][1] ), .G2(\gi[20][1] ), 
        .P2(\pi[20][1] ), .gout(\gi[24][2] ), .pout(\pi[24][2] ) );
  PG_7 pg_port2_0_6_7 ( .G1(\gi[28][1] ), .P1(\pi[28][1] ), .G2(\gi[24][1] ), 
        .P2(\pi[24][1] ), .gout(\gi[28][2] ), .pout(\pi[28][2] ) );
  PG_6 pg_port2_0_7_8 ( .G1(\gi[32][1] ), .P1(\pi[32][1] ), .G2(\gi[28][1] ), 
        .P2(\pi[28][1] ), .gout(\gi[32][2] ), .pout(\pi[32][2] ) );
  G_50 g_port_1_2 ( .G1(\gi[8][2] ), .P(\pi[8][2] ), .G2(Co[0]), .Co(Co[1]) );
  PG_5 pg_port2_1_1_4 ( .G1(\gi[16][2] ), .P1(\pi[16][2] ), .G2(\gi[12][2] ), 
        .P2(\pi[12][2] ), .gout(\gi[16][3] ), .pout(\pi[16][3] ) );
  PG_4 pg_port2_1_2_6 ( .G1(\gi[24][2] ), .P1(\pi[24][2] ), .G2(\gi[20][2] ), 
        .P2(\pi[20][2] ), .gout(\gi[24][3] ), .pout(\pi[24][3] ) );
  PG_3 pg_port2_1_3_8 ( .G1(\gi[32][2] ), .P1(\pi[32][2] ), .G2(\gi[28][2] ), 
        .P2(\pi[28][2] ), .gout(\gi[32][3] ), .pout(\pi[32][3] ) );
  G_49 g_port_2_3 ( .G1(\gi[12][2] ), .P(\pi[12][2] ), .G2(Co[1]), .Co(Co[2])
         );
  G_48 g_port_2_4 ( .G1(\gi[16][3] ), .P(\pi[16][3] ), .G2(Co[1]), .Co(Co[3])
         );
  PG_2 pg_port2_2_1_7 ( .G1(\gi[28][2] ), .P1(\pi[28][2] ), .G2(\gi[24][3] ), 
        .P2(\pi[24][3] ), .gout(\gi[28][4] ), .pout(\pi[28][4] ) );
  PG_1 pg_port2_2_1_8 ( .G1(\gi[32][3] ), .P1(\pi[32][3] ), .G2(\gi[24][3] ), 
        .P2(\pi[24][3] ), .gout(\gi[32][4] ), .pout(\pi[32][4] ) );
  G_47 g_port_3_5 ( .G1(\gi[20][2] ), .P(\pi[20][2] ), .G2(Co[3]), .Co(Co[4])
         );
  G_46 g_port_3_6 ( .G1(\gi[24][3] ), .P(\pi[24][3] ), .G2(Co[3]), .Co(Co[5])
         );
  G_45 g_port_3_7 ( .G1(\gi[28][4] ), .P(\pi[28][4] ), .G2(Co[3]), .Co(Co[6])
         );
  G_44 g_port_3_8 ( .G1(\gi[32][4] ), .P(\pi[32][4] ), .G2(Co[3]), .Co(Co[7])
         );
  AND2_X1 U2 ( .A1(B[31]), .A2(A[31]), .ZN(\gi[32][0] ) );
  AND2_X1 U3 ( .A1(B[15]), .A2(A[15]), .ZN(\gi[16][0] ) );
  AND2_X1 U4 ( .A1(B[14]), .A2(A[14]), .ZN(\gi[15][0] ) );
  AND2_X1 U5 ( .A1(B[23]), .A2(A[23]), .ZN(\gi[24][0] ) );
  AND2_X1 U6 ( .A1(B[22]), .A2(A[22]), .ZN(\gi[23][0] ) );
  AND2_X1 U7 ( .A1(B[19]), .A2(A[19]), .ZN(\gi[20][0] ) );
  AND2_X1 U8 ( .A1(B[18]), .A2(A[18]), .ZN(\gi[19][0] ) );
  AND2_X1 U9 ( .A1(B[0]), .A2(A[0]), .ZN(\gi[0][0] ) );
  AND2_X1 U10 ( .A1(B[3]), .A2(A[3]), .ZN(\gi[4][0] ) );
  AND2_X1 U11 ( .A1(B[2]), .A2(A[2]), .ZN(\gi[3][0] ) );
  AND2_X1 U12 ( .A1(B[7]), .A2(A[7]), .ZN(\gi[8][0] ) );
  AND2_X1 U13 ( .A1(B[6]), .A2(A[6]), .ZN(\gi[7][0] ) );
  AND2_X1 U14 ( .A1(B[11]), .A2(A[11]), .ZN(\gi[12][0] ) );
  AND2_X1 U15 ( .A1(B[10]), .A2(A[10]), .ZN(\gi[11][0] ) );
  AND2_X1 U16 ( .A1(B[27]), .A2(A[27]), .ZN(\gi[28][0] ) );
  AND2_X1 U17 ( .A1(B[26]), .A2(A[26]), .ZN(\gi[27][0] ) );
  AND2_X1 U18 ( .A1(B[30]), .A2(A[30]), .ZN(\gi[31][0] ) );
  AND2_X1 U19 ( .A1(B[1]), .A2(A[1]), .ZN(\gi[2][0] ) );
  AND2_X1 U20 ( .A1(B[4]), .A2(A[4]), .ZN(\gi[5][0] ) );
  AND2_X1 U21 ( .A1(B[5]), .A2(A[5]), .ZN(\gi[6][0] ) );
  AND2_X1 U22 ( .A1(B[8]), .A2(A[8]), .ZN(\gi[9][0] ) );
  AND2_X1 U23 ( .A1(B[9]), .A2(A[9]), .ZN(\gi[10][0] ) );
  AND2_X1 U24 ( .A1(B[12]), .A2(A[12]), .ZN(\gi[13][0] ) );
  AND2_X1 U25 ( .A1(B[13]), .A2(A[13]), .ZN(\gi[14][0] ) );
  AND2_X1 U26 ( .A1(B[16]), .A2(A[16]), .ZN(\gi[17][0] ) );
  AND2_X1 U27 ( .A1(B[17]), .A2(A[17]), .ZN(\gi[18][0] ) );
  AND2_X1 U28 ( .A1(B[20]), .A2(A[20]), .ZN(\gi[21][0] ) );
  AND2_X1 U29 ( .A1(B[21]), .A2(A[21]), .ZN(\gi[22][0] ) );
  AND2_X1 U30 ( .A1(B[24]), .A2(A[24]), .ZN(\gi[25][0] ) );
  AND2_X1 U31 ( .A1(B[25]), .A2(A[25]), .ZN(\gi[26][0] ) );
  AND2_X1 U32 ( .A1(B[28]), .A2(A[28]), .ZN(\gi[29][0] ) );
  AND2_X1 U33 ( .A1(B[29]), .A2(A[29]), .ZN(\gi[30][0] ) );
endmodule


module RCA_NBIT4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_32 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_32 UIV ( .A(S), .Y(SB) );
  ND2_96 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_95 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_94 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31 UIV ( .A(S), .Y(SB) );
  ND2_93 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_92 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_91 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30 UIV ( .A(S), .Y(SB) );
  ND2_90 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_89 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_88 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_29 UIV ( .A(S), .Y(SB) );
  ND2_87 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_86 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_85 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_32 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_29 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_0 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_28 UIV ( .A(S), .Y(SB) );
  ND2_84 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_83 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_82 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_27 UIV ( .A(S), .Y(SB) );
  ND2_81 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_80 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_79 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_26 UIV ( .A(S), .Y(SB) );
  ND2_78 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_77 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_76 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_25 UIV ( .A(S), .Y(SB) );
  ND2_75 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_74 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_73 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_28 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_27 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_26 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_25 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_7 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_24 UIV ( .A(S), .Y(SB) );
  ND2_72 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_71 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_70 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_23 UIV ( .A(S), .Y(SB) );
  ND2_69 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_68 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_67 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_22 UIV ( .A(S), .Y(SB) );
  ND2_66 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_65 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_64 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_21 UIV ( .A(S), .Y(SB) );
  ND2_63 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_62 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_61 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_24 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_23 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_22 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_21 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_6 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_20 UIV ( .A(S), .Y(SB) );
  ND2_60 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_59 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_58 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_19 UIV ( .A(S), .Y(SB) );
  ND2_57 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_56 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_55 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_18 UIV ( .A(S), .Y(SB) );
  ND2_54 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_53 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_52 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_17 UIV ( .A(S), .Y(SB) );
  ND2_51 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_50 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_49 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_20 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_19 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_18 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_17 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_5 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_16 UIV ( .A(S), .Y(SB) );
  ND2_48 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_47 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_46 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_15 UIV ( .A(S), .Y(SB) );
  ND2_45 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_44 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_43 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_14 UIV ( .A(S), .Y(SB) );
  ND2_42 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_41 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_40 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_13 UIV ( .A(S), .Y(SB) );
  ND2_39 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_38 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_37 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_16 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_15 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_14 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_13 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_4 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_12 UIV ( .A(S), .Y(SB) );
  ND2_36 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_35 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_34 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_11 UIV ( .A(S), .Y(SB) );
  ND2_33 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_32 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_31 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_10 UIV ( .A(S), .Y(SB) );
  ND2_30 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_29 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_28 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_9 UIV ( .A(S), .Y(SB) );
  ND2_27 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_26 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_25 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_12 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_11 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_10 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_9 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_3 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_8 UIV ( .A(S), .Y(SB) );
  ND2_24 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_23 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_22 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_7 UIV ( .A(S), .Y(SB) );
  ND2_21 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_20 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_19 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_6 UIV ( .A(S), .Y(SB) );
  ND2_18 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_17 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_16 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_5 UIV ( .A(S), .Y(SB) );
  ND2_15 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_14 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_13 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_8 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_7 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_6 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_5 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_2 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module RCA_NBIT4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module RCA_NBIT4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \add_1_root_add_52_2/carry[3] , \add_1_root_add_52_2/carry[2] ,
         \add_1_root_add_52_2/carry[1] ;

  FA_X1 \add_1_root_add_52_2/U1_0  ( .A(A[0]), .B(B[0]), .CI(Ci), .CO(
        \add_1_root_add_52_2/carry[1] ), .S(S[0]) );
  FA_X1 \add_1_root_add_52_2/U1_1  ( .A(A[1]), .B(B[1]), .CI(
        \add_1_root_add_52_2/carry[1] ), .CO(\add_1_root_add_52_2/carry[2] ), 
        .S(S[1]) );
  FA_X1 \add_1_root_add_52_2/U1_2  ( .A(A[2]), .B(B[2]), .CI(
        \add_1_root_add_52_2/carry[2] ), .CO(\add_1_root_add_52_2/carry[3] ), 
        .S(S[2]) );
  FA_X1 \add_1_root_add_52_2/U1_3  ( .A(A[3]), .B(B[3]), .CI(
        \add_1_root_add_52_2/carry[3] ), .CO(Co), .S(S[3]) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_4 UIV ( .A(S), .Y(SB) );
  ND2_12 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_11 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_10 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_3 UIV ( .A(S), .Y(SB) );
  ND2_9 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_8 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_7 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_2 UIV ( .A(S), .Y(SB) );
  ND2_6 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_5 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_4 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_1 UIV ( .A(S), .Y(SB) );
  ND2_3 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_2 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_1 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_4 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_3 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_2 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_1 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module CSB_NBIT4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] out_rca0;
  wire   [3:0] out_rca1;

  RCA_NBIT4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out_rca0) );
  RCA_NBIT4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out_rca1) );
  MUX21_GENERIC_NBIT4_1 MUXCin ( .A(out_rca1), .B(out_rca0), .SEL(Ci), .Y(S)
         );
endmodule


module SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSB_NBIT4_0 CSBI_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSB_NBIT4_7 CSBI_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSB_NBIT4_6 CSBI_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8]) );
  CSB_NBIT4_5 CSBI_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(S[15:12]) );
  CSB_NBIT4_4 CSBI_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(S[19:16]) );
  CSB_NBIT4_3 CSBI_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(S[23:20]) );
  CSB_NBIT4_2 CSBI_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(S[27:24]) );
  CSB_NBIT4_1 CSBI_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28]) );
endmodule


module P4_ADDER_NBIT32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [6:0] Cout_gen;

  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 carry_logic ( .A(A), .B(B), .Cin(Cin), 
        .Co({Cout, Cout_gen}) );
  SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 sum_logic ( .A(A), .B(B), .Ci({
        Cout_gen, Cin}), .S(S) );
endmodule


module ALU_N32 ( CLK, .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , 
        \FUNC[1] , \FUNC[0] }), DATA1, DATA2, OUT_ALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUT_ALU;
  input CLK, \FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   Cout_i, \OUTPUT3[0] , LOGIC_ARITH_i, LEFT_RIGHT_i, Cin_i, N139, N141,
         N142, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, n87, n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242;
  wire   [5:0] FUNC;
  wire   [31:0] OUTPUT_alu_i;
  wire   [31:0] OUTPUT4;
  wire   [31:0] OUTPUT2;
  wire   [31:0] OUTPUT1;
  wire   [31:0] data1i;
  wire   [31:0] data2i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  DLH_X1 Cin_i_reg ( .G(n164), .D(n87), .Q(Cin_i) );
  DLH_X1 \data2i_reg[31]  ( .G(n164), .D(N205), .Q(data2i[31]) );
  DLH_X1 \data2i_reg[30]  ( .G(n162), .D(N204), .Q(data2i[30]) );
  DLH_X1 \data2i_reg[29]  ( .G(n162), .D(N203), .Q(data2i[29]) );
  DLH_X1 \data2i_reg[28]  ( .G(n164), .D(N202), .Q(data2i[28]) );
  DLH_X1 \data2i_reg[27]  ( .G(n162), .D(N201), .Q(data2i[27]) );
  DLH_X1 \data2i_reg[26]  ( .G(n162), .D(N200), .Q(data2i[26]) );
  DLH_X1 \data2i_reg[25]  ( .G(n162), .D(N199), .Q(data2i[25]) );
  DLH_X1 \data2i_reg[24]  ( .G(n162), .D(N198), .Q(data2i[24]) );
  DLH_X1 \data2i_reg[23]  ( .G(n164), .D(N197), .Q(data2i[23]) );
  DLH_X1 \data2i_reg[22]  ( .G(n162), .D(N196), .Q(data2i[22]) );
  DLH_X1 \data2i_reg[21]  ( .G(n163), .D(N195), .Q(data2i[21]) );
  DLH_X1 \data2i_reg[20]  ( .G(n162), .D(N194), .Q(data2i[20]) );
  DLH_X1 \data2i_reg[19]  ( .G(n163), .D(N193), .Q(data2i[19]) );
  DLH_X1 \data2i_reg[18]  ( .G(n163), .D(N192), .Q(data2i[18]) );
  DLH_X1 \data2i_reg[17]  ( .G(n163), .D(N191), .Q(data2i[17]) );
  DLH_X1 \data2i_reg[16]  ( .G(n163), .D(N190), .Q(data2i[16]) );
  DLH_X1 \data2i_reg[15]  ( .G(n164), .D(N189), .Q(data2i[15]) );
  DLH_X1 \data2i_reg[14]  ( .G(n163), .D(N188), .Q(data2i[14]) );
  DLH_X1 \data2i_reg[13]  ( .G(n163), .D(N187), .Q(data2i[13]) );
  DLH_X1 \data2i_reg[12]  ( .G(n163), .D(N186), .Q(data2i[12]) );
  DLH_X1 \data2i_reg[11]  ( .G(n162), .D(N185), .Q(data2i[11]) );
  DLH_X1 \data2i_reg[10]  ( .G(n162), .D(N184), .Q(data2i[10]) );
  DLH_X1 \data2i_reg[9]  ( .G(n163), .D(N183), .Q(data2i[9]) );
  DLH_X1 \data2i_reg[8]  ( .G(n162), .D(N182), .Q(data2i[8]) );
  DLH_X1 \data2i_reg[7]  ( .G(n164), .D(N181), .Q(data2i[7]) );
  DLH_X1 \data2i_reg[6]  ( .G(n164), .D(N180), .Q(data2i[6]) );
  DLH_X1 \data2i_reg[5]  ( .G(n163), .D(N179), .Q(data2i[5]) );
  DLH_X1 \data2i_reg[4]  ( .G(n163), .D(N178), .Q(data2i[4]) );
  DLH_X1 \data2i_reg[3]  ( .G(n163), .D(N177), .Q(data2i[3]) );
  DLH_X1 \data2i_reg[2]  ( .G(n162), .D(N176), .Q(data2i[2]) );
  DLH_X1 \data2i_reg[1]  ( .G(n163), .D(N175), .Q(data2i[1]) );
  DLH_X1 \data2i_reg[0]  ( .G(n164), .D(N174), .Q(data2i[0]) );
  DLH_X1 \data1i_reg[31]  ( .G(n164), .D(DATA1[31]), .Q(data1i[31]) );
  DLH_X1 \data1i_reg[30]  ( .G(n162), .D(DATA1[30]), .Q(data1i[30]) );
  DLH_X1 \data1i_reg[29]  ( .G(n162), .D(DATA1[29]), .Q(data1i[29]) );
  DLH_X1 \data1i_reg[28]  ( .G(n164), .D(DATA1[28]), .Q(data1i[28]) );
  DLH_X1 \data1i_reg[27]  ( .G(n162), .D(DATA1[27]), .Q(data1i[27]) );
  DLH_X1 \data1i_reg[26]  ( .G(n162), .D(DATA1[26]), .Q(data1i[26]) );
  DLH_X1 \data1i_reg[25]  ( .G(n162), .D(DATA1[25]), .Q(data1i[25]) );
  DLH_X1 \data1i_reg[24]  ( .G(n162), .D(DATA1[24]), .Q(data1i[24]) );
  DLH_X1 \data1i_reg[23]  ( .G(n164), .D(DATA1[23]), .Q(data1i[23]) );
  DLH_X1 \data1i_reg[22]  ( .G(n162), .D(DATA1[22]), .Q(data1i[22]) );
  DLH_X1 \data1i_reg[21]  ( .G(n163), .D(DATA1[21]), .Q(data1i[21]) );
  DLH_X1 \data1i_reg[20]  ( .G(n162), .D(DATA1[20]), .Q(data1i[20]) );
  DLH_X1 \data1i_reg[19]  ( .G(n164), .D(DATA1[19]), .Q(data1i[19]) );
  DLH_X1 \data1i_reg[18]  ( .G(n163), .D(DATA1[18]), .Q(data1i[18]) );
  DLH_X1 \data1i_reg[17]  ( .G(n163), .D(DATA1[17]), .Q(data1i[17]) );
  DLH_X1 \data1i_reg[16]  ( .G(n163), .D(DATA1[16]), .Q(data1i[16]) );
  DLH_X1 \data1i_reg[15]  ( .G(n164), .D(DATA1[15]), .Q(data1i[15]) );
  DLH_X1 \data1i_reg[14]  ( .G(n163), .D(DATA1[14]), .Q(data1i[14]) );
  DLH_X1 \data1i_reg[13]  ( .G(n163), .D(DATA1[13]), .Q(data1i[13]) );
  DLH_X1 \data1i_reg[12]  ( .G(n163), .D(DATA1[12]), .Q(data1i[12]) );
  DLH_X1 \data1i_reg[11]  ( .G(n162), .D(DATA1[11]), .Q(data1i[11]) );
  DLH_X1 \data1i_reg[10]  ( .G(n162), .D(DATA1[10]), .Q(data1i[10]) );
  DLH_X1 \data1i_reg[9]  ( .G(n163), .D(DATA1[9]), .Q(data1i[9]) );
  DLH_X1 \data1i_reg[8]  ( .G(n162), .D(DATA1[8]), .Q(data1i[8]) );
  DLH_X1 \data1i_reg[7]  ( .G(n164), .D(DATA1[7]), .Q(data1i[7]) );
  DLH_X1 \data1i_reg[6]  ( .G(n164), .D(DATA1[6]), .Q(data1i[6]) );
  DLH_X1 \data1i_reg[5]  ( .G(n163), .D(DATA1[5]), .Q(data1i[5]) );
  DLH_X1 \data1i_reg[4]  ( .G(n163), .D(DATA1[4]), .Q(data1i[4]) );
  DLH_X1 \data1i_reg[3]  ( .G(n163), .D(DATA1[3]), .Q(data1i[3]) );
  DLH_X1 \data1i_reg[2]  ( .G(n163), .D(DATA1[2]), .Q(data1i[2]) );
  DLH_X1 \data1i_reg[1]  ( .G(n163), .D(DATA1[1]), .Q(data1i[1]) );
  DLH_X1 \data1i_reg[0]  ( .G(n164), .D(DATA1[0]), .Q(data1i[0]) );
  DLH_X1 LOGIC_ARITH_i_reg ( .G(n157), .D(n142), .Q(LOGIC_ARITH_i) );
  DLH_X1 LEFT_RIGHT_i_reg ( .G(n157), .D(n142), .Q(LEFT_RIGHT_i) );
  DLH_X1 \OUTPUT_alu_i_reg[0]  ( .G(n158), .D(N142), .Q(OUTPUT_alu_i[0]) );
  DFF_X1 \OUT_ALU_reg[0]  ( .D(OUTPUT_alu_i[0]), .CK(CLK), .Q(OUT_ALU[0]) );
  DLH_X1 \OUTPUT_alu_i_reg[1]  ( .G(n161), .D(n197), .Q(OUTPUT_alu_i[1]) );
  DFF_X1 \OUT_ALU_reg[1]  ( .D(OUTPUT_alu_i[1]), .CK(CLK), .Q(OUT_ALU[1]) );
  DLH_X1 \OUTPUT_alu_i_reg[2]  ( .G(n160), .D(n195), .Q(OUTPUT_alu_i[2]) );
  DFF_X1 \OUT_ALU_reg[2]  ( .D(OUTPUT_alu_i[2]), .CK(CLK), .Q(OUT_ALU[2]) );
  DLH_X1 \OUTPUT_alu_i_reg[3]  ( .G(n159), .D(n199), .Q(OUTPUT_alu_i[3]) );
  DFF_X1 \OUT_ALU_reg[3]  ( .D(OUTPUT_alu_i[3]), .CK(CLK), .Q(OUT_ALU[3]) );
  DLH_X1 \OUTPUT_alu_i_reg[4]  ( .G(n160), .D(n194), .Q(OUTPUT_alu_i[4]) );
  DFF_X1 \OUT_ALU_reg[4]  ( .D(OUTPUT_alu_i[4]), .CK(CLK), .Q(OUT_ALU[4]) );
  DLH_X1 \OUTPUT_alu_i_reg[5]  ( .G(n160), .D(n198), .Q(OUTPUT_alu_i[5]) );
  DFF_X1 \OUT_ALU_reg[5]  ( .D(OUTPUT_alu_i[5]), .CK(CLK), .Q(OUT_ALU[5]) );
  DLH_X1 \OUTPUT_alu_i_reg[6]  ( .G(n158), .D(n196), .Q(OUTPUT_alu_i[6]) );
  DFF_X1 \OUT_ALU_reg[6]  ( .D(OUTPUT_alu_i[6]), .CK(CLK), .Q(OUT_ALU[6]) );
  DLH_X1 \OUTPUT_alu_i_reg[7]  ( .G(n158), .D(n200), .Q(OUTPUT_alu_i[7]) );
  DFF_X1 \OUT_ALU_reg[7]  ( .D(OUTPUT_alu_i[7]), .CK(CLK), .Q(OUT_ALU[7]) );
  DLH_X1 \OUTPUT_alu_i_reg[8]  ( .G(n159), .D(n173), .Q(OUTPUT_alu_i[8]) );
  DFF_X1 \OUT_ALU_reg[8]  ( .D(OUTPUT_alu_i[8]), .CK(CLK), .Q(OUT_ALU[8]) );
  DLH_X1 \OUTPUT_alu_i_reg[9]  ( .G(n159), .D(n172), .Q(OUTPUT_alu_i[9]) );
  DFF_X1 \OUT_ALU_reg[9]  ( .D(OUTPUT_alu_i[9]), .CK(CLK), .Q(OUT_ALU[9]) );
  DLH_X1 \OUTPUT_alu_i_reg[10]  ( .G(n159), .D(n171), .Q(OUTPUT_alu_i[10]) );
  DFF_X1 \OUT_ALU_reg[10]  ( .D(OUTPUT_alu_i[10]), .CK(CLK), .Q(OUT_ALU[10])
         );
  DLH_X1 \OUTPUT_alu_i_reg[11]  ( .G(n159), .D(n170), .Q(OUTPUT_alu_i[11]) );
  DFF_X1 \OUT_ALU_reg[11]  ( .D(OUTPUT_alu_i[11]), .CK(CLK), .Q(OUT_ALU[11])
         );
  DLH_X1 \OUTPUT_alu_i_reg[12]  ( .G(n160), .D(n177), .Q(OUTPUT_alu_i[12]) );
  DFF_X1 \OUT_ALU_reg[12]  ( .D(OUTPUT_alu_i[12]), .CK(CLK), .Q(OUT_ALU[12])
         );
  DLH_X1 \OUTPUT_alu_i_reg[13]  ( .G(n160), .D(n176), .Q(OUTPUT_alu_i[13]) );
  DFF_X1 \OUT_ALU_reg[13]  ( .D(OUTPUT_alu_i[13]), .CK(CLK), .Q(OUT_ALU[13])
         );
  DLH_X1 \OUTPUT_alu_i_reg[14]  ( .G(n160), .D(n175), .Q(OUTPUT_alu_i[14]) );
  DFF_X1 \OUT_ALU_reg[14]  ( .D(OUTPUT_alu_i[14]), .CK(CLK), .Q(OUT_ALU[14])
         );
  DLH_X1 \OUTPUT_alu_i_reg[15]  ( .G(n158), .D(n174), .Q(OUTPUT_alu_i[15]) );
  DFF_X1 \OUT_ALU_reg[15]  ( .D(OUTPUT_alu_i[15]), .CK(CLK), .Q(OUT_ALU[15])
         );
  DLH_X1 \OUTPUT_alu_i_reg[16]  ( .G(n160), .D(n181), .Q(OUTPUT_alu_i[16]) );
  DFF_X1 \OUT_ALU_reg[16]  ( .D(OUTPUT_alu_i[16]), .CK(CLK), .Q(OUT_ALU[16])
         );
  DLH_X1 \OUTPUT_alu_i_reg[17]  ( .G(n160), .D(n180), .Q(OUTPUT_alu_i[17]) );
  DFF_X1 \OUT_ALU_reg[17]  ( .D(OUTPUT_alu_i[17]), .CK(CLK), .Q(OUT_ALU[17])
         );
  DLH_X1 \OUTPUT_alu_i_reg[18]  ( .G(n161), .D(n179), .Q(OUTPUT_alu_i[18]) );
  DFF_X1 \OUT_ALU_reg[18]  ( .D(OUTPUT_alu_i[18]), .CK(CLK), .Q(OUT_ALU[18])
         );
  DLH_X1 \OUTPUT_alu_i_reg[19]  ( .G(n158), .D(n178), .Q(OUTPUT_alu_i[19]) );
  DFF_X1 \OUT_ALU_reg[19]  ( .D(OUTPUT_alu_i[19]), .CK(CLK), .Q(OUT_ALU[19])
         );
  DLH_X1 \OUTPUT_alu_i_reg[20]  ( .G(n160), .D(n185), .Q(OUTPUT_alu_i[20]) );
  DFF_X1 \OUT_ALU_reg[20]  ( .D(OUTPUT_alu_i[20]), .CK(CLK), .Q(OUT_ALU[20])
         );
  DLH_X1 \OUTPUT_alu_i_reg[21]  ( .G(n159), .D(n184), .Q(OUTPUT_alu_i[21]) );
  DFF_X1 \OUT_ALU_reg[21]  ( .D(OUTPUT_alu_i[21]), .CK(CLK), .Q(OUT_ALU[21])
         );
  DLH_X1 \OUTPUT_alu_i_reg[22]  ( .G(n159), .D(n183), .Q(OUTPUT_alu_i[22]) );
  DFF_X1 \OUT_ALU_reg[22]  ( .D(OUTPUT_alu_i[22]), .CK(CLK), .Q(OUT_ALU[22])
         );
  DLH_X1 \OUTPUT_alu_i_reg[23]  ( .G(n158), .D(n182), .Q(OUTPUT_alu_i[23]) );
  DFF_X1 \OUT_ALU_reg[23]  ( .D(OUTPUT_alu_i[23]), .CK(CLK), .Q(OUT_ALU[23])
         );
  DLH_X1 \OUTPUT_alu_i_reg[24]  ( .G(n160), .D(n189), .Q(OUTPUT_alu_i[24]) );
  DFF_X1 \OUT_ALU_reg[24]  ( .D(OUTPUT_alu_i[24]), .CK(CLK), .Q(OUT_ALU[24])
         );
  DLH_X1 \OUTPUT_alu_i_reg[25]  ( .G(n159), .D(n188), .Q(OUTPUT_alu_i[25]) );
  DFF_X1 \OUT_ALU_reg[25]  ( .D(OUTPUT_alu_i[25]), .CK(CLK), .Q(OUT_ALU[25])
         );
  DLH_X1 \OUTPUT_alu_i_reg[26]  ( .G(n159), .D(n187), .Q(OUTPUT_alu_i[26]) );
  DFF_X1 \OUT_ALU_reg[26]  ( .D(OUTPUT_alu_i[26]), .CK(CLK), .Q(OUT_ALU[26])
         );
  DLH_X1 \OUTPUT_alu_i_reg[27]  ( .G(n159), .D(n186), .Q(OUTPUT_alu_i[27]) );
  DFF_X1 \OUT_ALU_reg[27]  ( .D(OUTPUT_alu_i[27]), .CK(CLK), .Q(OUT_ALU[27])
         );
  DLH_X1 \OUTPUT_alu_i_reg[28]  ( .G(n158), .D(n193), .Q(OUTPUT_alu_i[28]) );
  DFF_X1 \OUT_ALU_reg[28]  ( .D(OUTPUT_alu_i[28]), .CK(CLK), .Q(OUT_ALU[28])
         );
  DLH_X1 \OUTPUT_alu_i_reg[29]  ( .G(n158), .D(n192), .Q(OUTPUT_alu_i[29]) );
  DFF_X1 \OUT_ALU_reg[29]  ( .D(OUTPUT_alu_i[29]), .CK(CLK), .Q(OUT_ALU[29])
         );
  DLH_X1 \OUTPUT_alu_i_reg[30]  ( .G(n158), .D(n191), .Q(OUTPUT_alu_i[30]) );
  DFF_X1 \OUT_ALU_reg[30]  ( .D(OUTPUT_alu_i[30]), .CK(CLK), .Q(OUT_ALU[30])
         );
  DLH_X1 \OUTPUT_alu_i_reg[31]  ( .G(n158), .D(n190), .Q(OUTPUT_alu_i[31]) );
  DFF_X1 \OUT_ALU_reg[31]  ( .D(OUTPUT_alu_i[31]), .CK(CLK), .Q(OUT_ALU[31])
         );
  NAND3_X1 U177 ( .A1(n112), .A2(n113), .A3(n229), .ZN(n87) );
  OAI33_X1 U178 ( .A1(n131), .A2(n239), .A3(n240), .B1(n132), .B2(FUNC[3]), 
        .B3(FUNC[2]), .ZN(n130) );
  NAND3_X1 U179 ( .A1(n112), .A2(n113), .A3(n151), .ZN(n80) );
  NAND3_X1 U180 ( .A1(FUNC[3]), .A2(n237), .A3(FUNC[5]), .ZN(n131) );
  NAND3_X1 U181 ( .A1(n140), .A2(n126), .A3(n235), .ZN(n139) );
  logic_N32 log ( .FUNC({\FUNC[5] , \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , 
        \FUNC[0] }), .DATA1(DATA1), .DATA2(DATA2), .OUT_ALU(OUTPUT4) );
  comparator comp ( .DATA1(OUTPUT2), .DATA2i(Cout_i), .tipo({\FUNC[5] , 
        \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }), .OUTALU({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, \OUTPUT3[0] }) );
  SHIFTER_GENERIC_N32 shifter ( .A(DATA1), .B(DATA2[4:0]), .LOGIC_ARITH(
        LOGIC_ARITH_i), .LEFT_RIGHT(LEFT_RIGHT_i), .SHIFT_ROTATE(1'b1), 
        .OUTPUT(OUTPUT1) );
  P4_ADDER_NBIT32 adder ( .A(data1i), .B(data2i), .Cin(Cin_i), .S(OUTPUT2), 
        .Cout(Cout_i) );
  BUF_X1 U4 ( .A(N139), .Z(n163) );
  BUF_X1 U5 ( .A(n228), .Z(n143) );
  BUF_X1 U6 ( .A(n228), .Z(n144) );
  BUF_X1 U7 ( .A(N139), .Z(n162) );
  BUF_X1 U8 ( .A(n228), .Z(n145) );
  BUF_X1 U9 ( .A(N139), .Z(n164) );
  BUF_X1 U10 ( .A(n80), .Z(n152) );
  BUF_X1 U11 ( .A(n80), .Z(n153) );
  BUF_X1 U12 ( .A(n80), .Z(n154) );
  INV_X1 U13 ( .A(n140), .ZN(n234) );
  INV_X1 U14 ( .A(n87), .ZN(n228) );
  INV_X1 U15 ( .A(n118), .ZN(n240) );
  OR2_X1 U16 ( .A1(n154), .A2(n114), .ZN(N139) );
  OR3_X1 U17 ( .A1(n162), .A2(n155), .A3(n148), .ZN(N141) );
  INV_X1 U18 ( .A(n111), .ZN(n190) );
  AOI222_X1 U19 ( .A1(OUTPUT1[31]), .A2(n155), .B1(OUTPUT4[31]), .B2(n148), 
        .C1(OUTPUT2[31]), .C2(n154), .ZN(n111) );
  INV_X1 U20 ( .A(n110), .ZN(n191) );
  AOI222_X1 U21 ( .A1(OUTPUT1[30]), .A2(n157), .B1(OUTPUT4[30]), .B2(n148), 
        .C1(OUTPUT2[30]), .C2(n154), .ZN(n110) );
  INV_X1 U22 ( .A(n109), .ZN(n192) );
  AOI222_X1 U23 ( .A1(OUTPUT1[29]), .A2(n157), .B1(OUTPUT4[29]), .B2(n148), 
        .C1(OUTPUT2[29]), .C2(n154), .ZN(n109) );
  INV_X1 U24 ( .A(n108), .ZN(n193) );
  AOI222_X1 U25 ( .A1(OUTPUT1[28]), .A2(n157), .B1(OUTPUT4[28]), .B2(n148), 
        .C1(OUTPUT2[28]), .C2(n154), .ZN(n108) );
  INV_X1 U26 ( .A(n107), .ZN(n186) );
  AOI222_X1 U27 ( .A1(OUTPUT1[27]), .A2(n157), .B1(OUTPUT4[27]), .B2(n148), 
        .C1(OUTPUT2[27]), .C2(n154), .ZN(n107) );
  INV_X1 U28 ( .A(n106), .ZN(n187) );
  AOI222_X1 U29 ( .A1(OUTPUT1[26]), .A2(n157), .B1(OUTPUT4[26]), .B2(n148), 
        .C1(OUTPUT2[26]), .C2(n154), .ZN(n106) );
  INV_X1 U30 ( .A(n105), .ZN(n188) );
  AOI222_X1 U31 ( .A1(OUTPUT1[25]), .A2(n157), .B1(OUTPUT4[25]), .B2(n148), 
        .C1(OUTPUT2[25]), .C2(n154), .ZN(n105) );
  INV_X1 U32 ( .A(n104), .ZN(n189) );
  AOI222_X1 U33 ( .A1(OUTPUT1[24]), .A2(n157), .B1(OUTPUT4[24]), .B2(n148), 
        .C1(OUTPUT2[24]), .C2(n154), .ZN(n104) );
  INV_X1 U34 ( .A(n103), .ZN(n182) );
  AOI222_X1 U35 ( .A1(OUTPUT1[23]), .A2(n157), .B1(OUTPUT4[23]), .B2(n147), 
        .C1(OUTPUT2[23]), .C2(n153), .ZN(n103) );
  INV_X1 U36 ( .A(n102), .ZN(n183) );
  AOI222_X1 U37 ( .A1(OUTPUT1[22]), .A2(n157), .B1(OUTPUT4[22]), .B2(n147), 
        .C1(OUTPUT2[22]), .C2(n153), .ZN(n102) );
  INV_X1 U38 ( .A(n101), .ZN(n184) );
  AOI222_X1 U39 ( .A1(OUTPUT1[21]), .A2(n156), .B1(OUTPUT4[21]), .B2(n147), 
        .C1(OUTPUT2[21]), .C2(n153), .ZN(n101) );
  INV_X1 U40 ( .A(n100), .ZN(n185) );
  AOI222_X1 U41 ( .A1(OUTPUT1[20]), .A2(n156), .B1(OUTPUT4[20]), .B2(n147), 
        .C1(OUTPUT2[20]), .C2(n153), .ZN(n100) );
  INV_X1 U42 ( .A(n99), .ZN(n178) );
  AOI222_X1 U43 ( .A1(OUTPUT1[19]), .A2(n156), .B1(OUTPUT4[19]), .B2(n147), 
        .C1(OUTPUT2[19]), .C2(n153), .ZN(n99) );
  INV_X1 U44 ( .A(n98), .ZN(n179) );
  AOI222_X1 U45 ( .A1(OUTPUT1[18]), .A2(n156), .B1(OUTPUT4[18]), .B2(n147), 
        .C1(OUTPUT2[18]), .C2(n153), .ZN(n98) );
  INV_X1 U46 ( .A(n97), .ZN(n180) );
  AOI222_X1 U47 ( .A1(OUTPUT1[17]), .A2(n156), .B1(OUTPUT4[17]), .B2(n147), 
        .C1(OUTPUT2[17]), .C2(n153), .ZN(n97) );
  INV_X1 U48 ( .A(n96), .ZN(n181) );
  AOI222_X1 U49 ( .A1(OUTPUT1[16]), .A2(n156), .B1(OUTPUT4[16]), .B2(n147), 
        .C1(OUTPUT2[16]), .C2(n153), .ZN(n96) );
  INV_X1 U50 ( .A(n95), .ZN(n174) );
  AOI222_X1 U51 ( .A1(OUTPUT1[15]), .A2(n156), .B1(OUTPUT4[15]), .B2(n147), 
        .C1(OUTPUT2[15]), .C2(n153), .ZN(n95) );
  INV_X1 U52 ( .A(n94), .ZN(n175) );
  AOI222_X1 U53 ( .A1(OUTPUT1[14]), .A2(n156), .B1(OUTPUT4[14]), .B2(n147), 
        .C1(OUTPUT2[14]), .C2(n153), .ZN(n94) );
  INV_X1 U54 ( .A(n93), .ZN(n176) );
  AOI222_X1 U55 ( .A1(OUTPUT1[13]), .A2(n156), .B1(OUTPUT4[13]), .B2(n147), 
        .C1(OUTPUT2[13]), .C2(n153), .ZN(n93) );
  INV_X1 U56 ( .A(n92), .ZN(n177) );
  AOI222_X1 U57 ( .A1(OUTPUT1[12]), .A2(n156), .B1(OUTPUT4[12]), .B2(n146), 
        .C1(OUTPUT2[12]), .C2(n152), .ZN(n92) );
  INV_X1 U58 ( .A(n91), .ZN(n170) );
  AOI222_X1 U59 ( .A1(OUTPUT1[11]), .A2(n156), .B1(OUTPUT4[11]), .B2(n146), 
        .C1(OUTPUT2[11]), .C2(n152), .ZN(n91) );
  INV_X1 U60 ( .A(n90), .ZN(n171) );
  AOI222_X1 U61 ( .A1(OUTPUT1[10]), .A2(n155), .B1(OUTPUT4[10]), .B2(n146), 
        .C1(OUTPUT2[10]), .C2(n152), .ZN(n90) );
  INV_X1 U62 ( .A(n89), .ZN(n172) );
  AOI222_X1 U63 ( .A1(OUTPUT1[9]), .A2(n155), .B1(OUTPUT4[9]), .B2(n146), .C1(
        OUTPUT2[9]), .C2(n152), .ZN(n89) );
  INV_X1 U64 ( .A(n88), .ZN(n173) );
  AOI222_X1 U65 ( .A1(OUTPUT1[8]), .A2(n155), .B1(OUTPUT4[8]), .B2(n146), .C1(
        OUTPUT2[8]), .C2(n152), .ZN(n88) );
  INV_X1 U66 ( .A(n86), .ZN(n200) );
  AOI222_X1 U67 ( .A1(OUTPUT1[7]), .A2(n156), .B1(OUTPUT4[7]), .B2(n146), .C1(
        OUTPUT2[7]), .C2(n152), .ZN(n86) );
  INV_X1 U68 ( .A(n85), .ZN(n196) );
  AOI222_X1 U69 ( .A1(OUTPUT1[6]), .A2(n155), .B1(OUTPUT4[6]), .B2(n146), .C1(
        OUTPUT2[6]), .C2(n152), .ZN(n85) );
  INV_X1 U70 ( .A(n84), .ZN(n198) );
  AOI222_X1 U71 ( .A1(OUTPUT1[5]), .A2(n155), .B1(OUTPUT4[5]), .B2(n146), .C1(
        OUTPUT2[5]), .C2(n152), .ZN(n84) );
  INV_X1 U72 ( .A(n83), .ZN(n194) );
  AOI222_X1 U73 ( .A1(OUTPUT1[4]), .A2(n155), .B1(OUTPUT4[4]), .B2(n146), .C1(
        OUTPUT2[4]), .C2(n152), .ZN(n83) );
  OAI221_X1 U74 ( .B1(n241), .B2(n126), .C1(n118), .C2(n231), .A(n128), .ZN(
        n114) );
  INV_X1 U75 ( .A(n133), .ZN(n231) );
  NOR2_X1 U76 ( .A1(n129), .A2(n130), .ZN(n128) );
  AOI21_X1 U77 ( .B1(n242), .B2(n241), .A(n122), .ZN(n129) );
  NOR2_X1 U78 ( .A1(n241), .A2(n242), .ZN(n118) );
  AOI221_X1 U79 ( .B1(n127), .B2(n237), .C1(n139), .C2(n242), .A(n119), .ZN(
        n135) );
  INV_X1 U80 ( .A(n121), .ZN(n235) );
  BUF_X1 U81 ( .A(n232), .Z(n149) );
  BUF_X1 U82 ( .A(n232), .Z(n150) );
  BUF_X1 U83 ( .A(n232), .Z(n151) );
  BUF_X1 U84 ( .A(N206), .Z(n157) );
  BUF_X1 U85 ( .A(n230), .Z(n148) );
  BUF_X1 U86 ( .A(n230), .Z(n146) );
  BUF_X1 U87 ( .A(n230), .Z(n147) );
  BUF_X1 U88 ( .A(N206), .Z(n155) );
  BUF_X1 U89 ( .A(N206), .Z(n156) );
  OAI22_X1 U90 ( .A1(DATA2[0]), .A2(n143), .B1(n149), .B2(n165), .ZN(N174) );
  OAI22_X1 U91 ( .A1(DATA2[1]), .A2(n143), .B1(n149), .B2(n166), .ZN(N175) );
  OAI22_X1 U92 ( .A1(DATA2[2]), .A2(n143), .B1(n149), .B2(n167), .ZN(N176) );
  OAI22_X1 U93 ( .A1(DATA2[3]), .A2(n143), .B1(n149), .B2(n168), .ZN(N177) );
  OAI22_X1 U94 ( .A1(DATA2[4]), .A2(n143), .B1(n149), .B2(n169), .ZN(N178) );
  OAI22_X1 U95 ( .A1(DATA2[5]), .A2(n143), .B1(n149), .B2(n227), .ZN(N179) );
  INV_X1 U96 ( .A(DATA2[5]), .ZN(n227) );
  OAI22_X1 U97 ( .A1(DATA2[6]), .A2(n143), .B1(n149), .B2(n226), .ZN(N180) );
  INV_X1 U98 ( .A(DATA2[6]), .ZN(n226) );
  OAI22_X1 U99 ( .A1(DATA2[7]), .A2(n143), .B1(n149), .B2(n225), .ZN(N181) );
  INV_X1 U100 ( .A(DATA2[7]), .ZN(n225) );
  OAI22_X1 U101 ( .A1(DATA2[8]), .A2(n143), .B1(n149), .B2(n224), .ZN(N182) );
  INV_X1 U102 ( .A(DATA2[8]), .ZN(n224) );
  OAI22_X1 U103 ( .A1(DATA2[9]), .A2(n143), .B1(n149), .B2(n223), .ZN(N183) );
  INV_X1 U104 ( .A(DATA2[9]), .ZN(n223) );
  OAI22_X1 U105 ( .A1(DATA2[10]), .A2(n143), .B1(n149), .B2(n222), .ZN(N184)
         );
  INV_X1 U106 ( .A(DATA2[10]), .ZN(n222) );
  OAI22_X1 U107 ( .A1(DATA2[11]), .A2(n143), .B1(n150), .B2(n221), .ZN(N185)
         );
  INV_X1 U108 ( .A(DATA2[11]), .ZN(n221) );
  OAI22_X1 U109 ( .A1(DATA2[12]), .A2(n144), .B1(n150), .B2(n220), .ZN(N186)
         );
  INV_X1 U110 ( .A(DATA2[12]), .ZN(n220) );
  OAI22_X1 U111 ( .A1(DATA2[13]), .A2(n144), .B1(n150), .B2(n219), .ZN(N187)
         );
  INV_X1 U112 ( .A(DATA2[13]), .ZN(n219) );
  OAI22_X1 U113 ( .A1(DATA2[14]), .A2(n144), .B1(n150), .B2(n218), .ZN(N188)
         );
  INV_X1 U114 ( .A(DATA2[14]), .ZN(n218) );
  OAI22_X1 U115 ( .A1(DATA2[15]), .A2(n144), .B1(n150), .B2(n217), .ZN(N189)
         );
  INV_X1 U116 ( .A(DATA2[15]), .ZN(n217) );
  OAI22_X1 U117 ( .A1(DATA2[16]), .A2(n144), .B1(n150), .B2(n216), .ZN(N190)
         );
  INV_X1 U118 ( .A(DATA2[16]), .ZN(n216) );
  OAI22_X1 U119 ( .A1(DATA2[17]), .A2(n144), .B1(n150), .B2(n215), .ZN(N191)
         );
  INV_X1 U120 ( .A(DATA2[17]), .ZN(n215) );
  OAI22_X1 U121 ( .A1(DATA2[18]), .A2(n144), .B1(n150), .B2(n214), .ZN(N192)
         );
  INV_X1 U122 ( .A(DATA2[18]), .ZN(n214) );
  OAI22_X1 U123 ( .A1(DATA2[19]), .A2(n144), .B1(n150), .B2(n213), .ZN(N193)
         );
  INV_X1 U124 ( .A(DATA2[19]), .ZN(n213) );
  OAI22_X1 U125 ( .A1(DATA2[20]), .A2(n144), .B1(n150), .B2(n212), .ZN(N194)
         );
  INV_X1 U126 ( .A(DATA2[20]), .ZN(n212) );
  OAI22_X1 U127 ( .A1(DATA2[21]), .A2(n144), .B1(n150), .B2(n211), .ZN(N195)
         );
  INV_X1 U128 ( .A(DATA2[21]), .ZN(n211) );
  OAI22_X1 U129 ( .A1(DATA2[22]), .A2(n144), .B1(n151), .B2(n210), .ZN(N196)
         );
  INV_X1 U130 ( .A(DATA2[22]), .ZN(n210) );
  OAI22_X1 U131 ( .A1(DATA2[23]), .A2(n144), .B1(n151), .B2(n209), .ZN(N197)
         );
  INV_X1 U132 ( .A(DATA2[23]), .ZN(n209) );
  OAI22_X1 U133 ( .A1(DATA2[24]), .A2(n145), .B1(n151), .B2(n208), .ZN(N198)
         );
  INV_X1 U134 ( .A(DATA2[24]), .ZN(n208) );
  OAI22_X1 U135 ( .A1(DATA2[25]), .A2(n145), .B1(n151), .B2(n207), .ZN(N199)
         );
  INV_X1 U136 ( .A(DATA2[25]), .ZN(n207) );
  OAI22_X1 U137 ( .A1(DATA2[26]), .A2(n145), .B1(n151), .B2(n206), .ZN(N200)
         );
  INV_X1 U138 ( .A(DATA2[26]), .ZN(n206) );
  OAI22_X1 U139 ( .A1(DATA2[27]), .A2(n145), .B1(n151), .B2(n205), .ZN(N201)
         );
  INV_X1 U140 ( .A(DATA2[27]), .ZN(n205) );
  OAI22_X1 U141 ( .A1(DATA2[28]), .A2(n145), .B1(n151), .B2(n204), .ZN(N202)
         );
  INV_X1 U142 ( .A(DATA2[28]), .ZN(n204) );
  OAI22_X1 U143 ( .A1(DATA2[29]), .A2(n145), .B1(n151), .B2(n203), .ZN(N203)
         );
  INV_X1 U144 ( .A(DATA2[29]), .ZN(n203) );
  OAI22_X1 U145 ( .A1(DATA2[30]), .A2(n145), .B1(n151), .B2(n202), .ZN(N204)
         );
  INV_X1 U146 ( .A(DATA2[30]), .ZN(n202) );
  OAI22_X1 U147 ( .A1(DATA2[31]), .A2(n145), .B1(n151), .B2(n201), .ZN(N205)
         );
  INV_X1 U148 ( .A(DATA2[31]), .ZN(n201) );
  INV_X1 U149 ( .A(n127), .ZN(n236) );
  INV_X1 U150 ( .A(n114), .ZN(n229) );
  NAND2_X1 U151 ( .A1(n141), .A2(n239), .ZN(n140) );
  INV_X1 U152 ( .A(n82), .ZN(n199) );
  AOI222_X1 U153 ( .A1(OUTPUT1[3]), .A2(n155), .B1(OUTPUT4[3]), .B2(n146), 
        .C1(OUTPUT2[3]), .C2(n152), .ZN(n82) );
  INV_X1 U154 ( .A(n81), .ZN(n195) );
  AOI222_X1 U155 ( .A1(OUTPUT1[2]), .A2(n155), .B1(OUTPUT4[2]), .B2(n146), 
        .C1(OUTPUT2[2]), .C2(n152), .ZN(n81) );
  INV_X1 U156 ( .A(n79), .ZN(n197) );
  AOI222_X1 U157 ( .A1(OUTPUT1[1]), .A2(n155), .B1(OUTPUT4[1]), .B2(n147), 
        .C1(OUTPUT2[1]), .C2(n153), .ZN(n79) );
  NOR4_X1 U158 ( .A1(n239), .A2(FUNC[3]), .A3(FUNC[4]), .A4(FUNC[5]), .ZN(n121) );
  NOR4_X1 U159 ( .A1(n239), .A2(n238), .A3(FUNC[4]), .A4(FUNC[5]), .ZN(n119)
         );
  OAI21_X1 U160 ( .B1(n237), .B2(n241), .A(FUNC[5]), .ZN(n132) );
  NAND4_X1 U161 ( .A1(FUNC[3]), .A2(n239), .A3(n237), .A4(n233), .ZN(n122) );
  INV_X1 U162 ( .A(FUNC[1]), .ZN(n241) );
  NOR3_X1 U163 ( .A1(FUNC[3]), .A2(FUNC[5]), .A3(FUNC[2]), .ZN(n127) );
  INV_X1 U164 ( .A(FUNC[2]), .ZN(n239) );
  NOR3_X1 U165 ( .A1(n237), .A2(FUNC[5]), .A3(n238), .ZN(n141) );
  INV_X1 U166 ( .A(FUNC[4]), .ZN(n237) );
  OAI21_X1 U167 ( .B1(FUNC[2]), .B2(n131), .A(n138), .ZN(n133) );
  NAND4_X1 U168 ( .A1(FUNC[2]), .A2(FUNC[4]), .A3(n238), .A4(n233), .ZN(n138)
         );
  INV_X1 U169 ( .A(FUNC[3]), .ZN(n238) );
  OAI211_X1 U170 ( .C1(n241), .C2(n236), .A(n123), .B(n124), .ZN(N206) );
  OR3_X1 U171 ( .A1(n242), .A2(FUNC[1]), .A3(n126), .ZN(n123) );
  NAND4_X1 U172 ( .A1(n238), .A2(n237), .A3(FUNC[2]), .A4(n125), .ZN(n124) );
  NOR2_X1 U173 ( .A1(n240), .A2(n233), .ZN(n125) );
  INV_X1 U174 ( .A(FUNC[5]), .ZN(n233) );
  NAND2_X1 U175 ( .A1(n141), .A2(FUNC[2]), .ZN(n126) );
  INV_X1 U176 ( .A(FUNC[0]), .ZN(n242) );
  OAI211_X1 U182 ( .C1(n119), .C2(n234), .A(n242), .B(FUNC[1]), .ZN(n113) );
  NOR3_X1 U183 ( .A1(n241), .A2(FUNC[0]), .A3(n236), .ZN(n142) );
  OAI211_X1 U184 ( .C1(n234), .C2(n121), .A(n241), .B(FUNC[0]), .ZN(n112) );
  INV_X1 U185 ( .A(n117), .ZN(n230) );
  AOI222_X1 U186 ( .A1(n118), .A2(n119), .B1(n241), .B2(n120), .C1(FUNC[1]), 
        .C2(n121), .ZN(n117) );
  OAI22_X1 U187 ( .A1(n236), .A2(n237), .B1(n122), .B2(FUNC[0]), .ZN(n120) );
  INV_X1 U188 ( .A(n134), .ZN(n232) );
  OAI211_X1 U189 ( .C1(FUNC[1]), .C2(n135), .A(n136), .B(n137), .ZN(n134) );
  OR3_X1 U190 ( .A1(n239), .A2(n118), .A3(n131), .ZN(n137) );
  OAI21_X1 U191 ( .B1(n234), .B2(n133), .A(n118), .ZN(n136) );
  INV_X1 U192 ( .A(DATA2[2]), .ZN(n167) );
  INV_X1 U193 ( .A(DATA2[1]), .ZN(n166) );
  NAND2_X1 U194 ( .A1(n115), .A2(n116), .ZN(N142) );
  AOI22_X1 U195 ( .A1(OUTPUT2[0]), .A2(n152), .B1(OUTPUT1[0]), .B2(n155), .ZN(
        n115) );
  AOI22_X1 U196 ( .A1(OUTPUT4[0]), .A2(n146), .B1(\OUTPUT3[0] ), .B2(n114), 
        .ZN(n116) );
  CLKBUF_X1 U197 ( .A(N141), .Z(n158) );
  CLKBUF_X1 U198 ( .A(N141), .Z(n159) );
  CLKBUF_X1 U199 ( .A(N141), .Z(n160) );
  CLKBUF_X1 U200 ( .A(N141), .Z(n161) );
  INV_X1 U201 ( .A(DATA2[0]), .ZN(n165) );
  INV_X1 U202 ( .A(DATA2[3]), .ZN(n168) );
  INV_X1 U203 ( .A(DATA2[4]), .ZN(n169) );
endmodule


module zero_eval_NBIT32 ( \input , res );
  input [31:0] \input ;
  output res;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(\input [23]), .A2(\input [22]), .A3(\input [21]), .A4(
        \input [20]), .ZN(n6) );
  NOR4_X1 U2 ( .A1(\input [9]), .A2(\input [8]), .A3(\input [7]), .A4(
        \input [6]), .ZN(n10) );
  NOR4_X1 U3 ( .A1(\input [5]), .A2(\input [4]), .A3(\input [3]), .A4(
        \input [31]), .ZN(n9) );
  NOR4_X1 U4 ( .A1(\input [30]), .A2(\input [2]), .A3(\input [29]), .A4(
        \input [28]), .ZN(n8) );
  NOR4_X1 U5 ( .A1(\input [27]), .A2(\input [26]), .A3(\input [25]), .A4(
        \input [24]), .ZN(n7) );
  NAND4_X1 U6 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NOR4_X1 U7 ( .A1(\input [12]), .A2(\input [11]), .A3(\input [10]), .A4(
        \input [0]), .ZN(n3) );
  NOR4_X1 U8 ( .A1(\input [16]), .A2(\input [15]), .A3(\input [14]), .A4(
        \input [13]), .ZN(n4) );
  NOR4_X1 U9 ( .A1(\input [1]), .A2(\input [19]), .A3(\input [18]), .A4(
        \input [17]), .ZN(n5) );
  NOR2_X1 U10 ( .A1(n1), .A2(n2), .ZN(res) );
  NAND4_X1 U11 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
endmodule


module COND_BT_NBIT32 ( ZERO_BIT, OPCODE_0, branch_op, con_sign );
  input ZERO_BIT, OPCODE_0, branch_op;
  output con_sign;
  wire   n1;

  XOR2_X1 U3 ( .A(ZERO_BIT), .B(OPCODE_0), .Z(n1) );
  AND2_X1 U2 ( .A1(branch_op), .A2(n1), .ZN(con_sign) );
endmodule


module IV_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_160 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_160 UIV ( .A(S), .Y(SB) );
  ND2_480 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_479 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_478 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_159 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_159 UIV ( .A(S), .Y(SB) );
  ND2_477 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_476 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_475 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_158 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_158 UIV ( .A(S), .Y(SB) );
  ND2_474 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_473 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_472 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_157 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_157 UIV ( .A(S), .Y(SB) );
  ND2_471 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_470 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_469 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_156 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_156 UIV ( .A(S), .Y(SB) );
  ND2_468 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_467 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_466 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_155 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_155 UIV ( .A(S), .Y(SB) );
  ND2_465 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_464 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_463 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_154 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_154 UIV ( .A(S), .Y(SB) );
  ND2_462 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_461 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_460 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_153 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_153 UIV ( .A(S), .Y(SB) );
  ND2_459 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_458 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_457 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_152 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_152 UIV ( .A(S), .Y(SB) );
  ND2_456 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_455 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_454 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_151 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_151 UIV ( .A(S), .Y(SB) );
  ND2_453 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_452 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_451 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_150 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_150 UIV ( .A(S), .Y(SB) );
  ND2_450 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_449 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_448 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_149 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_149 UIV ( .A(S), .Y(SB) );
  ND2_447 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_446 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_445 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_148 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_148 UIV ( .A(S), .Y(SB) );
  ND2_444 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_443 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_442 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_147 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_147 UIV ( .A(S), .Y(SB) );
  ND2_441 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_440 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_439 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_146 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_146 UIV ( .A(S), .Y(SB) );
  ND2_438 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_437 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_436 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_145 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_145 UIV ( .A(S), .Y(SB) );
  ND2_435 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_434 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_433 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_144 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_144 UIV ( .A(S), .Y(SB) );
  ND2_432 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_431 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_430 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_143 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_143 UIV ( .A(S), .Y(SB) );
  ND2_429 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_428 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_427 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_142 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_142 UIV ( .A(S), .Y(SB) );
  ND2_426 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_425 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_424 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_141 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_141 UIV ( .A(S), .Y(SB) );
  ND2_423 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_422 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_421 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_140 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_140 UIV ( .A(S), .Y(SB) );
  ND2_420 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_419 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_418 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_139 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_139 UIV ( .A(S), .Y(SB) );
  ND2_417 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_416 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_415 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_138 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_138 UIV ( .A(S), .Y(SB) );
  ND2_414 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_413 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_412 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_137 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_137 UIV ( .A(S), .Y(SB) );
  ND2_411 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_410 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_409 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_136 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_136 UIV ( .A(S), .Y(SB) );
  ND2_408 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_407 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_406 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_135 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_135 UIV ( .A(S), .Y(SB) );
  ND2_405 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_404 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_403 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_134 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_134 UIV ( .A(S), .Y(SB) );
  ND2_402 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_401 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_400 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_133 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_133 UIV ( .A(S), .Y(SB) );
  ND2_399 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_398 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_397 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_132 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_132 UIV ( .A(S), .Y(SB) );
  ND2_396 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_395 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_394 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_131 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_131 UIV ( .A(S), .Y(SB) );
  ND2_393 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_392 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_391 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_130 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_130 UIV ( .A(S), .Y(SB) );
  ND2_390 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_389 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_388 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_129 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_129 UIV ( .A(S), .Y(SB) );
  ND2_387 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_386 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_385 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_160 gen1_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_159 gen1_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_158 gen1_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_157 gen1_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_156 gen1_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_155 gen1_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_154 gen1_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_153 gen1_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_152 gen1_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_151 gen1_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_150 gen1_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_149 gen1_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_148 gen1_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_147 gen1_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_146 gen1_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_145 gen1_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_144 gen1_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_143 gen1_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_142 gen1_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_141 gen1_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_140 gen1_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_139 gen1_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_138 gen1_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_137 gen1_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_136 gen1_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_135 gen1_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_134 gen1_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_133 gen1_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_132 gen1_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_131 gen1_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_130 gen1_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_129 gen1_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module FF_6 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n2, n3, n5, n6;

  DFF_X1 Q_reg ( .D(n2), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n3), .ZN(n2) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n5), .B2(Q), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n5) );
  INV_X1 U6 ( .A(RESET), .ZN(n3) );
endmodule


module regFFD_NBIT32_5 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U52 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U53 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U54 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U55 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U56 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U57 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U58 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U59 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U60 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U61 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U62 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U63 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U64 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U65 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U66 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
  OAI21_X1 U67 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U68 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
endmodule


module FF_5 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n2, n3, n5, n6;

  DFF_X1 Q_reg ( .D(n2), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n3), .ZN(n2) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n5), .B2(Q), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n5) );
  INV_X1 U6 ( .A(RESET), .ZN(n3) );
endmodule


module regFFD_NBIT32_4 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n65) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n66) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n67) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n68) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n69) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n98), .Q(Q[26]), .QN(n70) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n98), .Q(Q[25]), .QN(n71) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n98), .Q(Q[24]), .QN(n72) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n73) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n74) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n75) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n99), .Q(Q[20]), .QN(n76) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n97), .Q(Q[19]), .QN(n77) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n99), .Q(Q[18]), .QN(n78) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n99), .Q(Q[17]), .QN(n79) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n99), .Q(Q[16]), .QN(n80) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n97), .Q(Q[15]), .QN(n81) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n99), .Q(Q[14]), .QN(n82) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n99), .Q(Q[13]), .QN(n83) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n99), .Q(Q[12]), .QN(n84) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n85) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n86) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n98), .Q(Q[9]), .QN(n87) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n98), .Q(Q[8]), .QN(n88) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n97), .Q(Q[7]), .QN(n89) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n97), .Q(Q[6]), .QN(n90) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n91) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n92) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n98), .Q(Q[3]), .QN(n93) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n98), .Q(Q[2]), .QN(n94) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n95) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n97), .Q(Q[0]), .QN(n96) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n96), .B2(ENABLE), .A(n39), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n39) );
  OAI21_X1 U7 ( .B1(n95), .B2(ENABLE), .A(n40), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n40) );
  OAI21_X1 U9 ( .B1(n94), .B2(ENABLE), .A(n41), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n41) );
  OAI21_X1 U11 ( .B1(n93), .B2(ENABLE), .A(n43), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n43) );
  OAI21_X1 U13 ( .B1(n92), .B2(ENABLE), .A(n44), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n44) );
  OAI21_X1 U15 ( .B1(n91), .B2(ENABLE), .A(n45), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n45) );
  OAI21_X1 U17 ( .B1(n90), .B2(ENABLE), .A(n46), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n46) );
  OAI21_X1 U19 ( .B1(n89), .B2(ENABLE), .A(n47), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n47) );
  OAI21_X1 U21 ( .B1(n88), .B2(ENABLE), .A(n48), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n48) );
  OAI21_X1 U23 ( .B1(n87), .B2(ENABLE), .A(n49), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n49) );
  OAI21_X1 U25 ( .B1(n86), .B2(ENABLE), .A(n50), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n50) );
  OAI21_X1 U27 ( .B1(n85), .B2(ENABLE), .A(n51), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n51) );
  OAI21_X1 U29 ( .B1(n84), .B2(ENABLE), .A(n52), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n52) );
  OAI21_X1 U31 ( .B1(n83), .B2(ENABLE), .A(n54), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n54) );
  OAI21_X1 U33 ( .B1(n82), .B2(ENABLE), .A(n55), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n55) );
  OAI21_X1 U35 ( .B1(n81), .B2(ENABLE), .A(n56), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n56) );
  OAI21_X1 U37 ( .B1(n80), .B2(ENABLE), .A(n57), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n57) );
  OAI21_X1 U39 ( .B1(n79), .B2(ENABLE), .A(n58), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n58) );
  OAI21_X1 U41 ( .B1(n78), .B2(ENABLE), .A(n59), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n59) );
  OAI21_X1 U43 ( .B1(n77), .B2(ENABLE), .A(n60), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n60) );
  OAI21_X1 U45 ( .B1(n76), .B2(ENABLE), .A(n61), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n61) );
  OAI21_X1 U47 ( .B1(n75), .B2(ENABLE), .A(n62), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n62) );
  OAI21_X1 U49 ( .B1(n74), .B2(ENABLE), .A(n63), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n63) );
  OAI21_X1 U51 ( .B1(n72), .B2(ENABLE), .A(n34), .ZN(n8) );
  NAND2_X1 U52 ( .A1(D[24]), .A2(ENABLE), .ZN(n34) );
  OAI21_X1 U53 ( .B1(n71), .B2(ENABLE), .A(n35), .ZN(n7) );
  NAND2_X1 U54 ( .A1(D[25]), .A2(ENABLE), .ZN(n35) );
  OAI21_X1 U55 ( .B1(n70), .B2(ENABLE), .A(n36), .ZN(n6) );
  NAND2_X1 U56 ( .A1(D[26]), .A2(ENABLE), .ZN(n36) );
  OAI21_X1 U57 ( .B1(n69), .B2(ENABLE), .A(n37), .ZN(n5) );
  NAND2_X1 U58 ( .A1(D[27]), .A2(ENABLE), .ZN(n37) );
  OAI21_X1 U59 ( .B1(n68), .B2(ENABLE), .A(n38), .ZN(n4) );
  NAND2_X1 U60 ( .A1(D[28]), .A2(ENABLE), .ZN(n38) );
  OAI21_X1 U61 ( .B1(n67), .B2(ENABLE), .A(n42), .ZN(n3) );
  NAND2_X1 U62 ( .A1(D[29]), .A2(ENABLE), .ZN(n42) );
  OAI21_X1 U63 ( .B1(n66), .B2(ENABLE), .A(n53), .ZN(n2) );
  NAND2_X1 U64 ( .A1(D[30]), .A2(ENABLE), .ZN(n53) );
  OAI21_X1 U65 ( .B1(n65), .B2(ENABLE), .A(n64), .ZN(n1) );
  NAND2_X1 U66 ( .A1(D[31]), .A2(ENABLE), .ZN(n64) );
  OAI21_X1 U67 ( .B1(n73), .B2(ENABLE), .A(n33), .ZN(n9) );
  NAND2_X1 U68 ( .A1(ENABLE), .A2(D[23]), .ZN(n33) );
endmodule


module regFFD_NBIT5_2 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n20) );
  DFFR_X1 \Q_reg[3]  ( .D(n2), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n19) );
  DFFR_X1 \Q_reg[2]  ( .D(n3), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n18) );
  DFFR_X1 \Q_reg[1]  ( .D(n4), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n17) );
  DFFR_X1 \Q_reg[0]  ( .D(n5), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n16) );
  OAI21_X1 U2 ( .B1(n16), .B2(ENABLE), .A(n25), .ZN(n5) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n25) );
  OAI21_X1 U4 ( .B1(n17), .B2(ENABLE), .A(n24), .ZN(n4) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n24) );
  OAI21_X1 U6 ( .B1(n18), .B2(ENABLE), .A(n23), .ZN(n3) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n23) );
  OAI21_X1 U8 ( .B1(n19), .B2(ENABLE), .A(n22), .ZN(n2) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n22) );
  OAI21_X1 U10 ( .B1(n20), .B2(ENABLE), .A(n21), .ZN(n1) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n21) );
endmodule


module FF_4 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n5, n6;

  SDFF_X1 Q_reg ( .D(RESET), .SI(1'b0), .SE(n6), .CK(CLK), .Q(Q) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n5), .B2(Q), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n5) );
endmodule


module regFFD_NBIT6_1 ( CK, RESET, ENABLE, D, Q );
  input [5:0] D;
  output [5:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30;

  DFFR_X1 \Q_reg[5]  ( .D(n1), .CK(CK), .RN(RESET), .Q(Q[5]), .QN(n24) );
  DFFR_X1 \Q_reg[4]  ( .D(n2), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n23) );
  DFFR_X1 \Q_reg[3]  ( .D(n3), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n22) );
  DFFR_X1 \Q_reg[2]  ( .D(n4), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n21) );
  DFFR_X1 \Q_reg[1]  ( .D(n5), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n20) );
  DFFR_X1 \Q_reg[0]  ( .D(n6), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n19) );
  OAI21_X1 U2 ( .B1(n19), .B2(ENABLE), .A(n30), .ZN(n6) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n30) );
  OAI21_X1 U4 ( .B1(n20), .B2(ENABLE), .A(n29), .ZN(n5) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n29) );
  OAI21_X1 U6 ( .B1(n21), .B2(ENABLE), .A(n28), .ZN(n4) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n28) );
  OAI21_X1 U8 ( .B1(n22), .B2(ENABLE), .A(n27), .ZN(n3) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n27) );
  OAI21_X1 U10 ( .B1(n23), .B2(ENABLE), .A(n26), .ZN(n2) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n26) );
  OAI21_X1 U12 ( .B1(n24), .B2(ENABLE), .A(n25), .ZN(n1) );
  NAND2_X1 U13 ( .A1(D[5]), .A2(ENABLE), .ZN(n25) );
endmodule


module IV_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_128 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_128 UIV ( .A(S), .Y(SB) );
  ND2_384 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_383 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_382 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_127 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_127 UIV ( .A(S), .Y(SB) );
  ND2_381 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_380 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_379 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_126 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_126 UIV ( .A(S), .Y(SB) );
  ND2_378 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_377 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_376 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_125 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_125 UIV ( .A(S), .Y(SB) );
  ND2_375 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_374 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_373 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_124 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_124 UIV ( .A(S), .Y(SB) );
  ND2_372 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_371 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_370 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_123 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_123 UIV ( .A(S), .Y(SB) );
  ND2_369 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_368 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_367 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_122 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_122 UIV ( .A(S), .Y(SB) );
  ND2_366 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_365 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_364 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_121 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_121 UIV ( .A(S), .Y(SB) );
  ND2_363 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_362 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_361 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_120 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_120 UIV ( .A(S), .Y(SB) );
  ND2_360 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_359 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_358 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_119 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_119 UIV ( .A(S), .Y(SB) );
  ND2_357 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_356 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_355 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_118 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_118 UIV ( .A(S), .Y(SB) );
  ND2_354 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_353 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_352 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_117 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_117 UIV ( .A(S), .Y(SB) );
  ND2_351 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_350 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_349 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_116 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_116 UIV ( .A(S), .Y(SB) );
  ND2_348 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_347 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_346 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_115 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_115 UIV ( .A(S), .Y(SB) );
  ND2_345 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_344 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_343 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_114 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_114 UIV ( .A(S), .Y(SB) );
  ND2_342 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_341 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_340 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_113 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_113 UIV ( .A(S), .Y(SB) );
  ND2_339 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_338 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_337 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_112 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_112 UIV ( .A(S), .Y(SB) );
  ND2_336 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_335 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_334 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_111 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_111 UIV ( .A(S), .Y(SB) );
  ND2_333 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_332 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_331 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_110 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_110 UIV ( .A(S), .Y(SB) );
  ND2_330 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_329 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_328 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_109 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_109 UIV ( .A(S), .Y(SB) );
  ND2_327 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_326 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_325 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_108 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_108 UIV ( .A(S), .Y(SB) );
  ND2_324 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_323 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_322 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_107 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_107 UIV ( .A(S), .Y(SB) );
  ND2_321 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_320 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_319 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_106 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_106 UIV ( .A(S), .Y(SB) );
  ND2_318 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_317 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_316 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_105 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_105 UIV ( .A(S), .Y(SB) );
  ND2_315 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_314 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_313 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_104 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_104 UIV ( .A(S), .Y(SB) );
  ND2_312 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_311 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_310 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_103 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_103 UIV ( .A(S), .Y(SB) );
  ND2_309 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_308 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_307 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_102 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_102 UIV ( .A(S), .Y(SB) );
  ND2_306 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_305 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_304 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_101 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_101 UIV ( .A(S), .Y(SB) );
  ND2_303 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_302 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_301 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_100 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_100 UIV ( .A(S), .Y(SB) );
  ND2_300 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_299 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_298 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_99 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_99 UIV ( .A(S), .Y(SB) );
  ND2_297 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_296 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_295 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_98 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_98 UIV ( .A(S), .Y(SB) );
  ND2_294 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_293 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_292 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_97 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_97 UIV ( .A(S), .Y(SB) );
  ND2_291 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_290 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_289 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n4, n5, n6;

  MUX21_128 gen1_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_127 gen1_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_126 gen1_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_125 gen1_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_124 gen1_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_123 gen1_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_122 gen1_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_121 gen1_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_120 gen1_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_119 gen1_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_118 gen1_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_117 gen1_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_116 gen1_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_115 gen1_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_114 gen1_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_113 gen1_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_112 gen1_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_111 gen1_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_110 gen1_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_109 gen1_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_108 gen1_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_107 gen1_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_106 gen1_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_105 gen1_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_104 gen1_24 ( .A(A[24]), .B(B[24]), .S(n6), .Y(Y[24]) );
  MUX21_103 gen1_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_102 gen1_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_101 gen1_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_100 gen1_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_99 gen1_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_98 gen1_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_97 gen1_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n4) );
  BUF_X1 U2 ( .A(SEL), .Z(n5) );
  BUF_X1 U3 ( .A(SEL), .Z(n6) );
endmodule


module load_data ( data_in, signed_val, load_op, load_type, data_out );
  input [31:0] data_in;
  input [1:0] load_type;
  output [31:0] data_out;
  input signed_val, load_op;
  wire   N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34;

  DLH_X1 \data_out_reg[31]  ( .G(load_op), .D(N67), .Q(data_out[31]) );
  DLH_X1 \data_out_reg[30]  ( .G(load_op), .D(N66), .Q(data_out[30]) );
  DLH_X1 \data_out_reg[29]  ( .G(load_op), .D(N65), .Q(data_out[29]) );
  DLH_X1 \data_out_reg[28]  ( .G(load_op), .D(N64), .Q(data_out[28]) );
  DLH_X1 \data_out_reg[27]  ( .G(load_op), .D(N63), .Q(data_out[27]) );
  DLH_X1 \data_out_reg[26]  ( .G(load_op), .D(N62), .Q(data_out[26]) );
  DLH_X1 \data_out_reg[25]  ( .G(load_op), .D(N61), .Q(data_out[25]) );
  DLH_X1 \data_out_reg[24]  ( .G(load_op), .D(N60), .Q(data_out[24]) );
  DLH_X1 \data_out_reg[23]  ( .G(load_op), .D(N59), .Q(data_out[23]) );
  DLH_X1 \data_out_reg[22]  ( .G(load_op), .D(N58), .Q(data_out[22]) );
  DLH_X1 \data_out_reg[21]  ( .G(load_op), .D(N57), .Q(data_out[21]) );
  DLH_X1 \data_out_reg[20]  ( .G(load_op), .D(N56), .Q(data_out[20]) );
  DLH_X1 \data_out_reg[19]  ( .G(load_op), .D(N55), .Q(data_out[19]) );
  DLH_X1 \data_out_reg[18]  ( .G(load_op), .D(N54), .Q(data_out[18]) );
  DLH_X1 \data_out_reg[17]  ( .G(load_op), .D(N53), .Q(data_out[17]) );
  DLH_X1 \data_out_reg[16]  ( .G(load_op), .D(N52), .Q(data_out[16]) );
  DLH_X1 \data_out_reg[15]  ( .G(load_op), .D(N51), .Q(data_out[15]) );
  DLH_X1 \data_out_reg[14]  ( .G(load_op), .D(N50), .Q(data_out[14]) );
  DLH_X1 \data_out_reg[13]  ( .G(load_op), .D(N49), .Q(data_out[13]) );
  DLH_X1 \data_out_reg[12]  ( .G(load_op), .D(N48), .Q(data_out[12]) );
  DLH_X1 \data_out_reg[11]  ( .G(load_op), .D(N47), .Q(data_out[11]) );
  DLH_X1 \data_out_reg[10]  ( .G(load_op), .D(N46), .Q(data_out[10]) );
  DLH_X1 \data_out_reg[9]  ( .G(load_op), .D(N45), .Q(data_out[9]) );
  DLH_X1 \data_out_reg[8]  ( .G(load_op), .D(N44), .Q(data_out[8]) );
  DLH_X1 \data_out_reg[7]  ( .G(load_op), .D(N43), .Q(data_out[7]) );
  DLH_X1 \data_out_reg[6]  ( .G(load_op), .D(N42), .Q(data_out[6]) );
  DLH_X1 \data_out_reg[5]  ( .G(load_op), .D(N41), .Q(data_out[5]) );
  DLH_X1 \data_out_reg[4]  ( .G(load_op), .D(N40), .Q(data_out[4]) );
  DLH_X1 \data_out_reg[3]  ( .G(load_op), .D(N39), .Q(data_out[3]) );
  DLH_X1 \data_out_reg[2]  ( .G(load_op), .D(N38), .Q(data_out[2]) );
  DLH_X1 \data_out_reg[1]  ( .G(load_op), .D(N37), .Q(data_out[1]) );
  DLH_X1 \data_out_reg[0]  ( .G(load_op), .D(N36), .Q(data_out[0]) );
  INV_X1 U2 ( .A(n4), .ZN(n32) );
  BUF_X1 U3 ( .A(n5), .Z(n30) );
  BUF_X1 U4 ( .A(n5), .Z(n31) );
  OAI21_X1 U5 ( .B1(n4), .B2(n34), .A(n30), .ZN(N67) );
  NAND2_X1 U6 ( .A1(load_type[1]), .A2(n33), .ZN(n29) );
  INV_X1 U7 ( .A(load_type[0]), .ZN(n33) );
  NAND2_X1 U8 ( .A1(load_type[1]), .A2(load_type[0]), .ZN(n4) );
  OR4_X1 U9 ( .A1(load_type[0]), .A2(n34), .A3(signed_val), .A4(load_type[1]), 
        .ZN(n5) );
  INV_X1 U10 ( .A(data_in[31]), .ZN(n34) );
  NAND2_X1 U11 ( .A1(n31), .A2(n28), .ZN(N44) );
  NAND2_X1 U12 ( .A1(data_in[8]), .A2(load_type[0]), .ZN(n28) );
  NAND2_X1 U13 ( .A1(n31), .A2(n27), .ZN(N45) );
  NAND2_X1 U14 ( .A1(data_in[9]), .A2(load_type[0]), .ZN(n27) );
  NAND2_X1 U15 ( .A1(n31), .A2(n26), .ZN(N46) );
  NAND2_X1 U16 ( .A1(data_in[10]), .A2(load_type[0]), .ZN(n26) );
  NAND2_X1 U17 ( .A1(n31), .A2(n25), .ZN(N47) );
  NAND2_X1 U18 ( .A1(data_in[11]), .A2(load_type[0]), .ZN(n25) );
  NAND2_X1 U19 ( .A1(n31), .A2(n24), .ZN(N48) );
  NAND2_X1 U20 ( .A1(data_in[12]), .A2(load_type[0]), .ZN(n24) );
  NAND2_X1 U21 ( .A1(n31), .A2(n23), .ZN(N49) );
  NAND2_X1 U22 ( .A1(data_in[13]), .A2(load_type[0]), .ZN(n23) );
  NAND2_X1 U23 ( .A1(n31), .A2(n22), .ZN(N50) );
  NAND2_X1 U24 ( .A1(data_in[14]), .A2(load_type[0]), .ZN(n22) );
  NAND2_X1 U25 ( .A1(n31), .A2(n21), .ZN(N51) );
  NAND2_X1 U26 ( .A1(data_in[15]), .A2(load_type[0]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(n30), .A2(n16), .ZN(N56) );
  NAND2_X1 U28 ( .A1(data_in[20]), .A2(n32), .ZN(n16) );
  NAND2_X1 U29 ( .A1(n30), .A2(n15), .ZN(N57) );
  NAND2_X1 U30 ( .A1(data_in[21]), .A2(n32), .ZN(n15) );
  NAND2_X1 U31 ( .A1(n30), .A2(n14), .ZN(N58) );
  NAND2_X1 U32 ( .A1(data_in[22]), .A2(n32), .ZN(n14) );
  NAND2_X1 U33 ( .A1(n30), .A2(n13), .ZN(N59) );
  NAND2_X1 U34 ( .A1(data_in[23]), .A2(n32), .ZN(n13) );
  NAND2_X1 U35 ( .A1(n30), .A2(n12), .ZN(N60) );
  NAND2_X1 U36 ( .A1(data_in[24]), .A2(n32), .ZN(n12) );
  NAND2_X1 U37 ( .A1(n30), .A2(n11), .ZN(N61) );
  NAND2_X1 U38 ( .A1(data_in[25]), .A2(n32), .ZN(n11) );
  NAND2_X1 U39 ( .A1(n30), .A2(n10), .ZN(N62) );
  NAND2_X1 U40 ( .A1(data_in[26]), .A2(n32), .ZN(n10) );
  NAND2_X1 U41 ( .A1(n30), .A2(n9), .ZN(N63) );
  NAND2_X1 U42 ( .A1(data_in[27]), .A2(n32), .ZN(n9) );
  NAND2_X1 U43 ( .A1(n30), .A2(n8), .ZN(N64) );
  NAND2_X1 U44 ( .A1(data_in[28]), .A2(n32), .ZN(n8) );
  NAND2_X1 U45 ( .A1(n30), .A2(n7), .ZN(N65) );
  NAND2_X1 U46 ( .A1(data_in[29]), .A2(n32), .ZN(n7) );
  NAND2_X1 U47 ( .A1(n30), .A2(n6), .ZN(N66) );
  NAND2_X1 U48 ( .A1(data_in[30]), .A2(n32), .ZN(n6) );
  NAND2_X1 U49 ( .A1(n31), .A2(n20), .ZN(N52) );
  NAND2_X1 U50 ( .A1(data_in[16]), .A2(n32), .ZN(n20) );
  NAND2_X1 U51 ( .A1(n31), .A2(n19), .ZN(N53) );
  NAND2_X1 U52 ( .A1(data_in[17]), .A2(n32), .ZN(n19) );
  NAND2_X1 U53 ( .A1(n31), .A2(n18), .ZN(N54) );
  NAND2_X1 U54 ( .A1(data_in[18]), .A2(n32), .ZN(n18) );
  NAND2_X1 U55 ( .A1(n31), .A2(n17), .ZN(N55) );
  NAND2_X1 U56 ( .A1(data_in[19]), .A2(n32), .ZN(n17) );
  AND2_X1 U57 ( .A1(data_in[0]), .A2(n29), .ZN(N36) );
  AND2_X1 U58 ( .A1(data_in[1]), .A2(n29), .ZN(N37) );
  AND2_X1 U59 ( .A1(data_in[2]), .A2(n29), .ZN(N38) );
  AND2_X1 U60 ( .A1(data_in[3]), .A2(n29), .ZN(N39) );
  AND2_X1 U61 ( .A1(data_in[4]), .A2(n29), .ZN(N40) );
  AND2_X1 U62 ( .A1(data_in[5]), .A2(n29), .ZN(N41) );
  AND2_X1 U63 ( .A1(data_in[6]), .A2(n29), .ZN(N42) );
  AND2_X1 U64 ( .A1(data_in[7]), .A2(n29), .ZN(N43) );
endmodule


module regFFD_NBIT32_3 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n99), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n99), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n99), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n99), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n98), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n98), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n98), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n98), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n99), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n98), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n98), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n97), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n99), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n97), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n97), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n97), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n99), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n97), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n97), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n97), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n98), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n98), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n97), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n97), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n98), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n97), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n97), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n97) );
  BUF_X1 U3 ( .A(RESET), .Z(n98) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U6 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U7 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U8 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U9 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U10 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U11 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U12 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U13 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U14 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U15 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U16 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U17 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U18 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U19 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U20 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U21 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U22 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
  OAI21_X1 U23 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U24 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U25 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U26 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U27 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U28 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U29 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U30 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U31 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U32 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U33 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U34 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U35 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U36 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U37 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U38 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U39 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U40 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U41 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U42 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U43 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U44 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U45 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U46 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U47 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U48 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U49 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U50 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U51 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U52 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U53 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U54 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U55 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U56 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U57 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U58 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U59 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U60 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U61 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U62 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U63 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U64 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U65 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U66 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U67 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U68 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
endmodule


module regFFD_NBIT32_2 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U52 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
  OAI21_X1 U53 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U54 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U55 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U56 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U57 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U58 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U59 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U60 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U61 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U62 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U63 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U64 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U65 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U66 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U67 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U68 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
endmodule


module regFFD_NBIT5_1 ( CK, RESET, ENABLE, D, Q );
  input [4:0] D;
  output [4:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(CK), .RN(RESET), .Q(Q[4]), .QN(n20) );
  DFFR_X1 \Q_reg[3]  ( .D(n2), .CK(CK), .RN(RESET), .Q(Q[3]), .QN(n19) );
  DFFR_X1 \Q_reg[2]  ( .D(n3), .CK(CK), .RN(RESET), .Q(Q[2]), .QN(n18) );
  DFFR_X1 \Q_reg[1]  ( .D(n4), .CK(CK), .RN(RESET), .Q(Q[1]), .QN(n17) );
  DFFR_X1 \Q_reg[0]  ( .D(n5), .CK(CK), .RN(RESET), .Q(Q[0]), .QN(n16) );
  OAI21_X1 U2 ( .B1(n16), .B2(ENABLE), .A(n25), .ZN(n5) );
  NAND2_X1 U3 ( .A1(ENABLE), .A2(D[0]), .ZN(n25) );
  OAI21_X1 U4 ( .B1(n17), .B2(ENABLE), .A(n24), .ZN(n4) );
  NAND2_X1 U5 ( .A1(D[1]), .A2(ENABLE), .ZN(n24) );
  OAI21_X1 U6 ( .B1(n18), .B2(ENABLE), .A(n23), .ZN(n3) );
  NAND2_X1 U7 ( .A1(D[2]), .A2(ENABLE), .ZN(n23) );
  OAI21_X1 U8 ( .B1(n19), .B2(ENABLE), .A(n22), .ZN(n2) );
  NAND2_X1 U9 ( .A1(D[3]), .A2(ENABLE), .ZN(n22) );
  OAI21_X1 U10 ( .B1(n20), .B2(ENABLE), .A(n21), .ZN(n1) );
  NAND2_X1 U11 ( .A1(D[4]), .A2(ENABLE), .ZN(n21) );
endmodule


module FF_3 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n2, n3, n5, n6;

  DFF_X1 Q_reg ( .D(n2), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n3), .ZN(n2) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n5), .B2(Q), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n5) );
  INV_X1 U6 ( .A(RESET), .ZN(n3) );
endmodule


module FF_2 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n2, n3, n5, n6;

  DFF_X1 Q_reg ( .D(n2), .CK(CLK), .Q(Q) );
  NOR2_X1 U3 ( .A1(n6), .A2(n3), .ZN(n2) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n5), .B2(Q), .ZN(n6) );
  INV_X1 U5 ( .A(EN), .ZN(n5) );
  INV_X1 U6 ( .A(RESET), .ZN(n3) );
endmodule


module FF_1 ( CLK, RESET, EN, D, Q );
  input CLK, RESET, EN, D;
  output Q;
  wire   n6, n5, n3, n7, n8;
  assign Q = n6;

  DFF_X1 Q_reg ( .D(n5), .CK(CLK), .Q(n6) );
  NOR2_X1 U3 ( .A1(n3), .A2(n7), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n6), .B2(n8), .ZN(n3) );
  INV_X1 U5 ( .A(EN), .ZN(n8) );
  INV_X1 U6 ( .A(RESET), .ZN(n7) );
endmodule


module regFFD_NBIT32_1 ( CK, RESET, ENABLE, D, Q );
  input [31:0] D;
  output [31:0] Q;
  input CK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CK), .RN(n97), .Q(Q[31]), .QN(n131) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CK), .RN(n97), .Q(Q[30]), .QN(n130) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CK), .RN(n97), .Q(Q[29]), .QN(n129) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CK), .RN(n97), .Q(Q[28]), .QN(n128) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CK), .RN(n97), .Q(Q[27]), .QN(n127) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CK), .RN(n97), .Q(Q[26]), .QN(n126) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CK), .RN(n97), .Q(Q[25]), .QN(n125) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CK), .RN(n97), .Q(Q[24]), .QN(n124) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CK), .RN(n97), .Q(Q[23]), .QN(n123) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CK), .RN(n97), .Q(Q[22]), .QN(n122) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CK), .RN(n97), .Q(Q[21]), .QN(n121) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CK), .RN(n98), .Q(Q[20]), .QN(n120) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CK), .RN(n98), .Q(Q[19]), .QN(n119) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CK), .RN(n98), .Q(Q[18]), .QN(n118) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CK), .RN(n98), .Q(Q[17]), .QN(n117) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CK), .RN(n98), .Q(Q[16]), .QN(n116) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CK), .RN(n98), .Q(Q[15]), .QN(n115) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CK), .RN(n98), .Q(Q[14]), .QN(n114) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CK), .RN(n98), .Q(Q[13]), .QN(n113) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CK), .RN(n98), .Q(Q[12]), .QN(n112) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CK), .RN(n98), .Q(Q[11]), .QN(n111) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CK), .RN(n98), .Q(Q[10]), .QN(n110) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CK), .RN(n99), .Q(Q[9]), .QN(n109) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CK), .RN(n99), .Q(Q[8]), .QN(n108) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CK), .RN(n99), .Q(Q[7]), .QN(n107) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CK), .RN(n99), .Q(Q[6]), .QN(n106) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CK), .RN(n99), .Q(Q[5]), .QN(n105) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CK), .RN(n99), .Q(Q[4]), .QN(n104) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CK), .RN(n99), .Q(Q[3]), .QN(n103) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CK), .RN(n99), .Q(Q[2]), .QN(n102) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CK), .RN(n99), .Q(Q[1]), .QN(n101) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CK), .RN(n99), .Q(Q[0]), .QN(n100) );
  BUF_X1 U2 ( .A(RESET), .Z(n98) );
  BUF_X1 U3 ( .A(RESET), .Z(n97) );
  BUF_X1 U4 ( .A(RESET), .Z(n99) );
  OAI21_X1 U5 ( .B1(n100), .B2(ENABLE), .A(n157), .ZN(n32) );
  NAND2_X1 U6 ( .A1(D[0]), .A2(ENABLE), .ZN(n157) );
  OAI21_X1 U7 ( .B1(n101), .B2(ENABLE), .A(n156), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(ENABLE), .ZN(n156) );
  OAI21_X1 U9 ( .B1(n102), .B2(ENABLE), .A(n155), .ZN(n30) );
  NAND2_X1 U10 ( .A1(D[2]), .A2(ENABLE), .ZN(n155) );
  OAI21_X1 U11 ( .B1(n103), .B2(ENABLE), .A(n153), .ZN(n29) );
  NAND2_X1 U12 ( .A1(D[3]), .A2(ENABLE), .ZN(n153) );
  OAI21_X1 U13 ( .B1(n104), .B2(ENABLE), .A(n152), .ZN(n28) );
  NAND2_X1 U14 ( .A1(D[4]), .A2(ENABLE), .ZN(n152) );
  OAI21_X1 U15 ( .B1(n105), .B2(ENABLE), .A(n151), .ZN(n27) );
  NAND2_X1 U16 ( .A1(D[5]), .A2(ENABLE), .ZN(n151) );
  OAI21_X1 U17 ( .B1(n106), .B2(ENABLE), .A(n150), .ZN(n26) );
  NAND2_X1 U18 ( .A1(D[6]), .A2(ENABLE), .ZN(n150) );
  OAI21_X1 U19 ( .B1(n107), .B2(ENABLE), .A(n149), .ZN(n25) );
  NAND2_X1 U20 ( .A1(D[7]), .A2(ENABLE), .ZN(n149) );
  OAI21_X1 U21 ( .B1(n108), .B2(ENABLE), .A(n148), .ZN(n24) );
  NAND2_X1 U22 ( .A1(D[8]), .A2(ENABLE), .ZN(n148) );
  OAI21_X1 U23 ( .B1(n109), .B2(ENABLE), .A(n147), .ZN(n23) );
  NAND2_X1 U24 ( .A1(D[9]), .A2(ENABLE), .ZN(n147) );
  OAI21_X1 U25 ( .B1(n110), .B2(ENABLE), .A(n146), .ZN(n22) );
  NAND2_X1 U26 ( .A1(D[10]), .A2(ENABLE), .ZN(n146) );
  OAI21_X1 U27 ( .B1(n111), .B2(ENABLE), .A(n145), .ZN(n21) );
  NAND2_X1 U28 ( .A1(D[11]), .A2(ENABLE), .ZN(n145) );
  OAI21_X1 U29 ( .B1(n112), .B2(ENABLE), .A(n144), .ZN(n20) );
  NAND2_X1 U30 ( .A1(D[12]), .A2(ENABLE), .ZN(n144) );
  OAI21_X1 U31 ( .B1(n113), .B2(ENABLE), .A(n142), .ZN(n19) );
  NAND2_X1 U32 ( .A1(D[13]), .A2(ENABLE), .ZN(n142) );
  OAI21_X1 U33 ( .B1(n114), .B2(ENABLE), .A(n141), .ZN(n18) );
  NAND2_X1 U34 ( .A1(D[14]), .A2(ENABLE), .ZN(n141) );
  OAI21_X1 U35 ( .B1(n115), .B2(ENABLE), .A(n140), .ZN(n17) );
  NAND2_X1 U36 ( .A1(D[15]), .A2(ENABLE), .ZN(n140) );
  OAI21_X1 U37 ( .B1(n116), .B2(ENABLE), .A(n139), .ZN(n16) );
  NAND2_X1 U38 ( .A1(D[16]), .A2(ENABLE), .ZN(n139) );
  OAI21_X1 U39 ( .B1(n117), .B2(ENABLE), .A(n138), .ZN(n15) );
  NAND2_X1 U40 ( .A1(D[17]), .A2(ENABLE), .ZN(n138) );
  OAI21_X1 U41 ( .B1(n118), .B2(ENABLE), .A(n137), .ZN(n14) );
  NAND2_X1 U42 ( .A1(D[18]), .A2(ENABLE), .ZN(n137) );
  OAI21_X1 U43 ( .B1(n119), .B2(ENABLE), .A(n136), .ZN(n13) );
  NAND2_X1 U44 ( .A1(D[19]), .A2(ENABLE), .ZN(n136) );
  OAI21_X1 U45 ( .B1(n120), .B2(ENABLE), .A(n135), .ZN(n12) );
  NAND2_X1 U46 ( .A1(D[20]), .A2(ENABLE), .ZN(n135) );
  OAI21_X1 U47 ( .B1(n121), .B2(ENABLE), .A(n134), .ZN(n11) );
  NAND2_X1 U48 ( .A1(D[21]), .A2(ENABLE), .ZN(n134) );
  OAI21_X1 U49 ( .B1(n122), .B2(ENABLE), .A(n133), .ZN(n10) );
  NAND2_X1 U50 ( .A1(D[22]), .A2(ENABLE), .ZN(n133) );
  OAI21_X1 U51 ( .B1(n124), .B2(ENABLE), .A(n162), .ZN(n8) );
  NAND2_X1 U52 ( .A1(D[24]), .A2(ENABLE), .ZN(n162) );
  OAI21_X1 U53 ( .B1(n125), .B2(ENABLE), .A(n161), .ZN(n7) );
  NAND2_X1 U54 ( .A1(D[25]), .A2(ENABLE), .ZN(n161) );
  OAI21_X1 U55 ( .B1(n126), .B2(ENABLE), .A(n160), .ZN(n6) );
  NAND2_X1 U56 ( .A1(D[26]), .A2(ENABLE), .ZN(n160) );
  OAI21_X1 U57 ( .B1(n127), .B2(ENABLE), .A(n159), .ZN(n5) );
  NAND2_X1 U58 ( .A1(D[27]), .A2(ENABLE), .ZN(n159) );
  OAI21_X1 U59 ( .B1(n128), .B2(ENABLE), .A(n158), .ZN(n4) );
  NAND2_X1 U60 ( .A1(D[28]), .A2(ENABLE), .ZN(n158) );
  OAI21_X1 U61 ( .B1(n129), .B2(ENABLE), .A(n154), .ZN(n3) );
  NAND2_X1 U62 ( .A1(D[29]), .A2(ENABLE), .ZN(n154) );
  OAI21_X1 U63 ( .B1(n130), .B2(ENABLE), .A(n143), .ZN(n2) );
  NAND2_X1 U64 ( .A1(D[30]), .A2(ENABLE), .ZN(n143) );
  OAI21_X1 U65 ( .B1(n131), .B2(ENABLE), .A(n132), .ZN(n1) );
  NAND2_X1 U66 ( .A1(D[31]), .A2(ENABLE), .ZN(n132) );
  OAI21_X1 U67 ( .B1(n123), .B2(ENABLE), .A(n163), .ZN(n9) );
  NAND2_X1 U68 ( .A1(ENABLE), .A2(D[23]), .ZN(n163) );
endmodule


module IV_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_96 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_96 UIV ( .A(S), .Y(SB) );
  ND2_288 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_287 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_286 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_95 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_95 UIV ( .A(S), .Y(SB) );
  ND2_285 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_284 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_283 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_94 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_94 UIV ( .A(S), .Y(SB) );
  ND2_282 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_281 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_280 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_93 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_93 UIV ( .A(S), .Y(SB) );
  ND2_279 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_278 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_277 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_92 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_92 UIV ( .A(S), .Y(SB) );
  ND2_276 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_275 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_274 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_91 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_91 UIV ( .A(S), .Y(SB) );
  ND2_273 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_272 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_271 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_90 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_90 UIV ( .A(S), .Y(SB) );
  ND2_270 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_269 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_268 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_89 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_89 UIV ( .A(S), .Y(SB) );
  ND2_267 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_266 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_265 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_88 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_88 UIV ( .A(S), .Y(SB) );
  ND2_264 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_263 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_262 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_87 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_87 UIV ( .A(S), .Y(SB) );
  ND2_261 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_260 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_259 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_86 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_86 UIV ( .A(S), .Y(SB) );
  ND2_258 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_257 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_256 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_85 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_85 UIV ( .A(S), .Y(SB) );
  ND2_255 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_254 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_253 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_84 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_84 UIV ( .A(S), .Y(SB) );
  ND2_252 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_251 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_250 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_83 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_83 UIV ( .A(S), .Y(SB) );
  ND2_249 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_248 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_247 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_82 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_82 UIV ( .A(S), .Y(SB) );
  ND2_246 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_245 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_244 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_81 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_81 UIV ( .A(S), .Y(SB) );
  ND2_243 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_242 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_241 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_80 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_80 UIV ( .A(S), .Y(SB) );
  ND2_240 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_239 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_238 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_79 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_79 UIV ( .A(S), .Y(SB) );
  ND2_237 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_236 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_235 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_78 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_78 UIV ( .A(S), .Y(SB) );
  ND2_234 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_233 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_232 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_77 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_77 UIV ( .A(S), .Y(SB) );
  ND2_231 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_230 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_229 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_76 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_76 UIV ( .A(S), .Y(SB) );
  ND2_228 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_227 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_226 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_75 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_75 UIV ( .A(S), .Y(SB) );
  ND2_225 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_224 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_223 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_74 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_74 UIV ( .A(S), .Y(SB) );
  ND2_222 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_221 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_220 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_73 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_73 UIV ( .A(S), .Y(SB) );
  ND2_219 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_218 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_217 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_72 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_72 UIV ( .A(S), .Y(SB) );
  ND2_216 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_215 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_214 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_71 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_71 UIV ( .A(S), .Y(SB) );
  ND2_213 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_212 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_211 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_70 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_70 UIV ( .A(S), .Y(SB) );
  ND2_210 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_209 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_208 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_69 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_69 UIV ( .A(S), .Y(SB) );
  ND2_207 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_206 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_205 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_68 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_68 UIV ( .A(S), .Y(SB) );
  ND2_204 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_203 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_202 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_67 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_67 UIV ( .A(S), .Y(SB) );
  ND2_201 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_200 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_199 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_66 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_66 UIV ( .A(S), .Y(SB) );
  ND2_198 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_197 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_196 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_65 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_65 UIV ( .A(S), .Y(SB) );
  ND2_195 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_194 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_193 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;


  MUX21_96 gen1_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_95 gen1_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_94 gen1_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_93 gen1_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_92 gen1_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_91 gen1_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_90 gen1_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_89 gen1_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
  MUX21_88 gen1_8 ( .A(A[8]), .B(B[8]), .S(SEL), .Y(Y[8]) );
  MUX21_87 gen1_9 ( .A(A[9]), .B(B[9]), .S(SEL), .Y(Y[9]) );
  MUX21_86 gen1_10 ( .A(A[10]), .B(B[10]), .S(SEL), .Y(Y[10]) );
  MUX21_85 gen1_11 ( .A(A[11]), .B(B[11]), .S(SEL), .Y(Y[11]) );
  MUX21_84 gen1_12 ( .A(A[12]), .B(B[12]), .S(SEL), .Y(Y[12]) );
  MUX21_83 gen1_13 ( .A(A[13]), .B(B[13]), .S(SEL), .Y(Y[13]) );
  MUX21_82 gen1_14 ( .A(A[14]), .B(B[14]), .S(SEL), .Y(Y[14]) );
  MUX21_81 gen1_15 ( .A(A[15]), .B(B[15]), .S(SEL), .Y(Y[15]) );
  MUX21_80 gen1_16 ( .A(A[16]), .B(B[16]), .S(SEL), .Y(Y[16]) );
  MUX21_79 gen1_17 ( .A(A[17]), .B(B[17]), .S(SEL), .Y(Y[17]) );
  MUX21_78 gen1_18 ( .A(A[18]), .B(B[18]), .S(SEL), .Y(Y[18]) );
  MUX21_77 gen1_19 ( .A(A[19]), .B(B[19]), .S(SEL), .Y(Y[19]) );
  MUX21_76 gen1_20 ( .A(A[20]), .B(B[20]), .S(SEL), .Y(Y[20]) );
  MUX21_75 gen1_21 ( .A(A[21]), .B(B[21]), .S(SEL), .Y(Y[21]) );
  MUX21_74 gen1_22 ( .A(A[22]), .B(B[22]), .S(SEL), .Y(Y[22]) );
  MUX21_73 gen1_23 ( .A(A[23]), .B(B[23]), .S(SEL), .Y(Y[23]) );
  MUX21_72 gen1_24 ( .A(A[24]), .B(B[24]), .S(SEL), .Y(Y[24]) );
  MUX21_71 gen1_25 ( .A(A[25]), .B(B[25]), .S(SEL), .Y(Y[25]) );
  MUX21_70 gen1_26 ( .A(A[26]), .B(B[26]), .S(SEL), .Y(Y[26]) );
  MUX21_69 gen1_27 ( .A(A[27]), .B(B[27]), .S(SEL), .Y(Y[27]) );
  MUX21_68 gen1_28 ( .A(A[28]), .B(B[28]), .S(SEL), .Y(Y[28]) );
  MUX21_67 gen1_29 ( .A(A[29]), .B(B[29]), .S(SEL), .Y(Y[29]) );
  MUX21_66 gen1_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_65 gen1_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
endmodule


module IV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_64 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_64 UIV ( .A(S), .Y(SB) );
  ND2_192 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_191 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_190 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_63 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_63 UIV ( .A(S), .Y(SB) );
  ND2_189 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_188 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_187 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_62 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_62 UIV ( .A(S), .Y(SB) );
  ND2_186 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_185 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_184 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_61 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_61 UIV ( .A(S), .Y(SB) );
  ND2_183 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_182 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_181 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_60 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_60 UIV ( .A(S), .Y(SB) );
  ND2_180 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_179 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_178 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_59 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_59 UIV ( .A(S), .Y(SB) );
  ND2_177 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_176 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_175 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_58 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_58 UIV ( .A(S), .Y(SB) );
  ND2_174 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_173 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_172 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_57 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_57 UIV ( .A(S), .Y(SB) );
  ND2_171 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_170 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_169 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_56 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_56 UIV ( .A(S), .Y(SB) );
  ND2_168 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_167 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_166 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_55 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_55 UIV ( .A(S), .Y(SB) );
  ND2_165 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_164 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_163 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_54 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_54 UIV ( .A(S), .Y(SB) );
  ND2_162 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_161 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_160 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_53 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_53 UIV ( .A(S), .Y(SB) );
  ND2_159 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_158 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_157 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_52 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_52 UIV ( .A(S), .Y(SB) );
  ND2_156 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_155 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_154 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_51 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_51 UIV ( .A(S), .Y(SB) );
  ND2_153 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_152 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_151 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_50 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_50 UIV ( .A(S), .Y(SB) );
  ND2_150 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_149 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_148 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_49 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_49 UIV ( .A(S), .Y(SB) );
  ND2_147 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_146 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_145 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_48 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_48 UIV ( .A(S), .Y(SB) );
  ND2_144 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_143 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_142 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_47 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_47 UIV ( .A(S), .Y(SB) );
  ND2_141 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_140 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_139 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_46 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_46 UIV ( .A(S), .Y(SB) );
  ND2_138 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_137 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_136 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_45 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_45 UIV ( .A(S), .Y(SB) );
  ND2_135 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_134 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_133 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_44 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_44 UIV ( .A(S), .Y(SB) );
  ND2_132 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_131 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_130 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_43 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_43 UIV ( .A(S), .Y(SB) );
  ND2_129 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_128 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_127 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_42 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_42 UIV ( .A(S), .Y(SB) );
  ND2_126 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_125 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_124 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_41 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_41 UIV ( .A(S), .Y(SB) );
  ND2_123 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_122 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_121 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_40 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_40 UIV ( .A(S), .Y(SB) );
  ND2_120 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_119 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_118 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_39 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_39 UIV ( .A(S), .Y(SB) );
  ND2_117 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_116 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_115 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_38 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_38 UIV ( .A(S), .Y(SB) );
  ND2_114 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_113 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_112 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_37 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_37 UIV ( .A(S), .Y(SB) );
  ND2_111 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_110 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_109 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_36 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_36 UIV ( .A(S), .Y(SB) );
  ND2_108 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_107 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_106 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_35 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_35 UIV ( .A(S), .Y(SB) );
  ND2_105 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_104 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_103 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_34 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_34 UIV ( .A(S), .Y(SB) );
  ND2_102 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_101 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_100 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_33 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_33 UIV ( .A(S), .Y(SB) );
  ND2_99 UND1 ( .A(A), .B(S), .Y(Y1) );
  ND2_98 UND2 ( .A(B), .B(SB), .Y(Y2) );
  ND2_97 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_64 gen1_0 ( .A(A[0]), .B(B[0]), .S(n3), .Y(Y[0]) );
  MUX21_63 gen1_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_62 gen1_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_61 gen1_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_60 gen1_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_59 gen1_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_58 gen1_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_57 gen1_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_56 gen1_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_55 gen1_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_54 gen1_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_53 gen1_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_52 gen1_12 ( .A(A[12]), .B(B[12]), .S(n1), .Y(Y[12]) );
  MUX21_51 gen1_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_50 gen1_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_49 gen1_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_48 gen1_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_47 gen1_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_46 gen1_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_45 gen1_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_44 gen1_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_43 gen1_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_42 gen1_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_41 gen1_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_40 gen1_24 ( .A(A[24]), .B(B[24]), .S(n2), .Y(Y[24]) );
  MUX21_39 gen1_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_38 gen1_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_37 gen1_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_36 gen1_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_35 gen1_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_34 gen1_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_33 gen1_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U2 ( .A(carry[31]), .B(A[31]), .Z(SUM[31]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module DATAPTH_NBIT32_REG_BIT5 ( CLK, RST, PC, IR, PC_OUT, NPC_LATCH_EN, 
        ir_LATCH_EN, signed_op, trap_cs, ret_cs, RF1, RF2, WF1, 
        regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond, sb_op, RM, 
        WM, EN3, S3, .instruction_alu({\instruction_alu[5] , 
        \instruction_alu[4] , \instruction_alu[3] , \instruction_alu[2] , 
        \instruction_alu[1] , \instruction_alu[0] }), DATA_MEM_ADDR, 
        DATA_MEM_IN, DATA_MEM_OUT, DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM
 );
  input [31:0] PC;
  input [31:0] IR;
  output [31:0] PC_OUT;
  output [31:0] DATA_MEM_ADDR;
  output [31:0] DATA_MEM_IN;
  input [31:0] DATA_MEM_OUT;
  input CLK, RST, NPC_LATCH_EN, ir_LATCH_EN, signed_op, trap_cs, ret_cs, RF1,
         RF2, WF1, regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond,
         sb_op, RM, WM, EN3, S3, \instruction_alu[5] , \instruction_alu[4] ,
         \instruction_alu[3] , \instruction_alu[2] , \instruction_alu[1] ,
         \instruction_alu[0] ;
  output DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM;
  wire   RM, WM, sel_npc, wr_signal_wb, signed_op_ex, wr_signal_exe, is_zero,
         cond, signed_op_mem, cond_mem, wr_signal_mem, sel_saved_reg, N13,
         wr_signal_mem1, sel_saved_reg_wb, n34, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55;
  wire   [5:0] instruction_alu;
  wire   [31:0] PC_fetch0;
  wire   [31:0] NPC;
  wire   [31:0] NPC_fetch1;
  wire   [31:0] PC_fetch1;
  wire   [31:0] PC_OUT_i;
  wire   [31:0] NPC_fetch;
  wire   [31:0] PC_fetch;
  wire   [31:0] ir_fetch;
  wire   [31:0] NPC_Dec;
  wire   [31:0] IR_Dec;
  wire   [4:0] RS1;
  wire   [4:0] RS2;
  wire   [4:0] RD;
  wire   [31:0] Imm;
  wire   [4:0] RD_wb;
  wire   [31:0] OUT_wb;
  wire   [31:0] regA;
  wire   [31:0] regB;
  wire   [31:0] NPC_ex;
  wire   [31:0] regA_ex;
  wire   [31:0] regB_ex;
  wire   [31:0] Imm_ex;
  wire   [4:0] RD_ex;
  wire   [5:0] IR_26_ex;
  wire   [31:0] LHI_ex1;
  wire   [31:0] LHI_ex;
  wire   [31:0] input1_ALU;
  wire   [31:0] input2_ALU;
  wire   [31:0] ALU_out;
  wire   [31:0] ALU_ex;
  wire   [31:0] NPC_mem;
  wire   [31:8] regB_mem;
  wire   [4:0] RD_mem;
  wire   [5:0] IR_26_mem;
  wire   [31:0] LMD_out;
  wire   [31:0] ALU_wb;
  wire   [31:0] LMD_wb;
  wire   [31:0] NPC_wb;
  wire   [31:0] OUT_data;
  assign DATA_MEM_RM = RM;
  assign DATA_MEM_WM = WM;

  DLH_X1 \DATA_MEM_ADDR_reg[31]  ( .G(n43), .D(ALU_ex[31]), .Q(
        DATA_MEM_ADDR[31]) );
  DLH_X1 \DATA_MEM_ADDR_reg[30]  ( .G(n42), .D(ALU_ex[30]), .Q(
        DATA_MEM_ADDR[30]) );
  DLH_X1 \DATA_MEM_ADDR_reg[29]  ( .G(n42), .D(ALU_ex[29]), .Q(
        DATA_MEM_ADDR[29]) );
  DLH_X1 \DATA_MEM_ADDR_reg[28]  ( .G(n42), .D(ALU_ex[28]), .Q(
        DATA_MEM_ADDR[28]) );
  DLH_X1 \DATA_MEM_ADDR_reg[27]  ( .G(n42), .D(ALU_ex[27]), .Q(
        DATA_MEM_ADDR[27]) );
  DLH_X1 \DATA_MEM_ADDR_reg[26]  ( .G(n41), .D(ALU_ex[26]), .Q(
        DATA_MEM_ADDR[26]) );
  DLH_X1 \DATA_MEM_ADDR_reg[25]  ( .G(n41), .D(ALU_ex[25]), .Q(
        DATA_MEM_ADDR[25]) );
  DLH_X1 \DATA_MEM_ADDR_reg[24]  ( .G(n41), .D(ALU_ex[24]), .Q(
        DATA_MEM_ADDR[24]) );
  DLH_X1 \DATA_MEM_ADDR_reg[23]  ( .G(n42), .D(ALU_ex[23]), .Q(
        DATA_MEM_ADDR[23]) );
  DLH_X1 \DATA_MEM_ADDR_reg[22]  ( .G(n41), .D(ALU_ex[22]), .Q(
        DATA_MEM_ADDR[22]) );
  DLH_X1 \DATA_MEM_ADDR_reg[21]  ( .G(n41), .D(ALU_ex[21]), .Q(
        DATA_MEM_ADDR[21]) );
  DLH_X1 \DATA_MEM_ADDR_reg[20]  ( .G(n40), .D(ALU_ex[20]), .Q(
        DATA_MEM_ADDR[20]) );
  DLH_X1 \DATA_MEM_ADDR_reg[19]  ( .G(n42), .D(ALU_ex[19]), .Q(
        DATA_MEM_ADDR[19]) );
  DLH_X1 \DATA_MEM_ADDR_reg[18]  ( .G(n40), .D(ALU_ex[18]), .Q(
        DATA_MEM_ADDR[18]) );
  DLH_X1 \DATA_MEM_ADDR_reg[17]  ( .G(n40), .D(ALU_ex[17]), .Q(
        DATA_MEM_ADDR[17]) );
  DLH_X1 \DATA_MEM_ADDR_reg[16]  ( .G(n40), .D(ALU_ex[16]), .Q(
        DATA_MEM_ADDR[16]) );
  DLH_X1 \DATA_MEM_ADDR_reg[15]  ( .G(n42), .D(ALU_ex[15]), .Q(
        DATA_MEM_ADDR[15]) );
  DLH_X1 \DATA_MEM_ADDR_reg[14]  ( .G(n40), .D(ALU_ex[14]), .Q(
        DATA_MEM_ADDR[14]) );
  DLH_X1 \DATA_MEM_ADDR_reg[13]  ( .G(n40), .D(ALU_ex[13]), .Q(
        DATA_MEM_ADDR[13]) );
  DLH_X1 \DATA_MEM_ADDR_reg[12]  ( .G(n40), .D(ALU_ex[12]), .Q(
        DATA_MEM_ADDR[12]) );
  DLH_X1 \DATA_MEM_ADDR_reg[11]  ( .G(n41), .D(ALU_ex[11]), .Q(
        DATA_MEM_ADDR[11]) );
  DLH_X1 \DATA_MEM_ADDR_reg[10]  ( .G(n41), .D(ALU_ex[10]), .Q(
        DATA_MEM_ADDR[10]) );
  DLH_X1 \DATA_MEM_ADDR_reg[9]  ( .G(n41), .D(ALU_ex[9]), .Q(DATA_MEM_ADDR[9])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[8]  ( .G(n41), .D(ALU_ex[8]), .Q(DATA_MEM_ADDR[8])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[7]  ( .G(n42), .D(ALU_ex[7]), .Q(DATA_MEM_ADDR[7])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[6]  ( .G(n42), .D(ALU_ex[6]), .Q(DATA_MEM_ADDR[6])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[5]  ( .G(n40), .D(ALU_ex[5]), .Q(DATA_MEM_ADDR[5])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[4]  ( .G(n40), .D(ALU_ex[4]), .Q(DATA_MEM_ADDR[4])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[3]  ( .G(n42), .D(ALU_ex[3]), .Q(DATA_MEM_ADDR[3])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[2]  ( .G(n41), .D(ALU_ex[2]), .Q(DATA_MEM_ADDR[2])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[1]  ( .G(n40), .D(ALU_ex[1]), .Q(DATA_MEM_ADDR[1])
         );
  DLH_X1 \DATA_MEM_ADDR_reg[0]  ( .G(n43), .D(ALU_ex[0]), .Q(DATA_MEM_ADDR[0])
         );
  XOR2_X1 U62 ( .A(IR_Dec[27]), .B(IR_Dec[26]), .Z(n15) );
  NAND3_X1 U63 ( .A1(instruction_alu[2]), .A2(instruction_alu[1]), .A3(
        instruction_alu[4]), .ZN(n31) );
  regFFD_NBIT32_0 pipeline_PCING ( .CK(CLK), .RESET(n45), .ENABLE(1'b1), .D(PC), .Q(PC_fetch0) );
  regFFD_NBIT32_19 pipeline_fetch1_NPC ( .CK(CLK), .RESET(n45), .ENABLE(
        NPC_LATCH_EN), .D(NPC), .Q(NPC_fetch1) );
  regFFD_NBIT32_18 pipeline_fetch1_PC ( .CK(CLK), .RESET(n45), .ENABLE(
        ir_LATCH_EN), .D(PC_fetch0), .Q(PC_fetch1) );
  MUX21_GENERIC_NBIT32_0 MUX_PC1 ( .A(PC_OUT_i), .B(NPC_fetch1), .SEL(sel_npc), 
        .Y(PC_OUT) );
  regFFD_NBIT32_17 pipeline_fetch_NPC ( .CK(CLK), .RESET(n45), .ENABLE(
        NPC_LATCH_EN), .D(NPC_fetch1), .Q(NPC_fetch) );
  regFFD_NBIT32_16 pipeline_fetch_PC ( .CK(CLK), .RESET(n45), .ENABLE(
        ir_LATCH_EN), .D(PC_fetch1), .Q(PC_fetch) );
  regFFD_NBIT32_15 pipeline_fetch_ir ( .CK(CLK), .RESET(n45), .ENABLE(
        ir_LATCH_EN), .D(IR), .Q(ir_fetch) );
  regFFD_NBIT32_14 pipeline_newpc1 ( .CK(CLK), .RESET(n45), .ENABLE(
        NPC_LATCH_EN), .D(NPC_fetch), .Q(NPC_Dec) );
  regFFD_NBIT32_13 pipeline_pc1 ( .CK(CLK), .RESET(n45), .ENABLE(ir_LATCH_EN), 
        .D(PC_fetch) );
  regFFD_NBIT32_12 pipeline_IR1 ( .CK(CLK), .RESET(n45), .ENABLE(ir_LATCH_EN), 
        .D(ir_fetch), .Q(IR_Dec) );
  IR_DECODE_NBIT32_opBIT6_regBIT5 IR_OP ( .CLK(CLK), .IR_26(IR_Dec[25:0]), 
        .OPCODE(IR_Dec[31:26]), .is_signed(signed_op), .RS1(RS1), .RS2(RS2), 
        .RD(RD), .IMMEDIATE(Imm) );
  windRF_M8_N8_F5_NBIT32 RF ( .CLK(CLK), .RESET(n44), .ENABLE(1'b1), .CALL(
        trap_cs), .RETRN(ret_cs), .BUSin({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .RD1(RF1), .RD2(RF2), .WR(WF1), .ADD_WR(RD_wb), 
        .ADD_RD1(RS1), .ADD_RD2(RS2), .DATAIN(OUT_wb), .OUT1(regA), .OUT2(regB), .wr_signal(wr_signal_wb) );
  FF_0 pipeline_sign2 ( .CLK(CLK), .RESET(n45), .EN(1'b1), .D(signed_op), .Q(
        signed_op_ex) );
  regFFD_NBIT32_11 pipeline_newpc2 ( .CK(CLK), .RESET(n45), .ENABLE(1'b1), .D(
        NPC_Dec), .Q(NPC_ex) );
  regFFD_NBIT32_10 pipeline_A2 ( .CK(CLK), .RESET(n44), .ENABLE(RF1), .D(regA), 
        .Q(regA_ex) );
  regFFD_NBIT32_9 pipeline_B2 ( .CK(CLK), .RESET(n44), .ENABLE(RF2), .D(regB), 
        .Q(regB_ex) );
  regFFD_NBIT32_8 pipeline_IMM2 ( .CK(CLK), .RESET(n44), .ENABLE(
        regImm_LATCH_EN), .D(Imm), .Q(Imm_ex) );
  regFFD_NBIT5_0 pipeline_RD2 ( .CK(CLK), .RESET(n44), .ENABLE(1'b1), .D(RD), 
        .Q(RD_ex) );
  FF_7 pipeline_wr_signal ( .CLK(CLK), .RESET(n45), .EN(1'b1), .D(n34), .Q(
        wr_signal_exe) );
  regFFD_NBIT6_0 pipeline_IR2 ( .CK(CLK), .RESET(n44), .ENABLE(1'b1), .D({n36, 
        IR_Dec[30], n35, IR_Dec[28:26]}), .Q(IR_26_ex) );
  regFFD_NBIT32_7 pipeline_LHI2 ( .CK(CLK), .RESET(n45), .ENABLE(1'b1), .D({
        Imm[15:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Q(LHI_ex1) );
  regFFD_NBIT32_6 pipeline_LHI3 ( .CK(CLK), .RESET(n45), .ENABLE(1'b1), .D(
        LHI_ex1), .Q(LHI_ex) );
  MUX21_GENERIC_NBIT32_6 MUX_ALU_A ( .A(NPC_ex), .B(regA_ex), .SEL(S1), .Y(
        input1_ALU) );
  MUX21_GENERIC_NBIT32_5 MUX_ALU_B ( .A(Imm_ex), .B(regB_ex), .SEL(S2), .Y(
        input2_ALU) );
  ALU_N32 ALU_OP ( .CLK(CLK), .FUNC({\instruction_alu[5] , 
        \instruction_alu[4] , \instruction_alu[3] , \instruction_alu[2] , 
        \instruction_alu[1] , \instruction_alu[0] }), .DATA1(input1_ALU), 
        .DATA2(input2_ALU), .OUT_ALU(ALU_out) );
  zero_eval_NBIT32 ZERO_OP ( .\input (regA_ex), .res(is_zero) );
  COND_BT_NBIT32 COND_OP ( .ZERO_BIT(is_zero), .OPCODE_0(IR_26_ex[0]), 
        .branch_op(branch_cond), .con_sign(cond) );
  MUX21_GENERIC_NBIT32_4 MUX_alu_out ( .A(LHI_ex), .B(ALU_out), .SEL(lhi_sel), 
        .Y(ALU_ex) );
  FF_6 pipeline_sign3 ( .CLK(CLK), .RESET(n45), .EN(1'b1), .D(signed_op_ex), 
        .Q(signed_op_mem) );
  regFFD_NBIT32_5 pipeline_newpc3 ( .CK(CLK), .RESET(n45), .ENABLE(1'b1), .D(
        NPC_ex), .Q(NPC_mem) );
  FF_5 pipeline_cond3 ( .CLK(CLK), .RESET(n45), .EN(1'b1), .D(cond), .Q(
        cond_mem) );
  regFFD_NBIT32_4 pipeline_B3 ( .CK(CLK), .RESET(n44), .ENABLE(1'b1), .D(
        regB_ex), .Q({regB_mem, DATA_MEM_IN[7:0]}) );
  regFFD_NBIT5_2 pipeline_RD3 ( .CK(CLK), .RESET(n44), .ENABLE(1'b1), .D(RD_ex), .Q(RD_mem) );
  FF_4 pipeline_wr_signal2 ( .CLK(CLK), .RESET(n45), .EN(1'b1), .D(
        wr_signal_exe), .Q(wr_signal_mem) );
  regFFD_NBIT6_1 pipeline_IR3 ( .CK(CLK), .RESET(n44), .ENABLE(1'b1), .D(
        IR_26_ex), .Q(IR_26_mem) );
  MUX21_GENERIC_NBIT32_3 MUX_PC ( .A(ALU_ex), .B(NPC_mem), .SEL(sel_npc), .Y(
        PC_OUT_i) );
  load_data LOAD_DATA_OUT ( .data_in(DATA_MEM_OUT), .signed_val(signed_op_mem), 
        .load_op(RM), .load_type(IR_26_mem[1:0]), .data_out(LMD_out) );
  regFFD_NBIT32_3 pipeline_alu4 ( .CK(CLK), .RESET(n45), .ENABLE(1'b1), .D(
        ALU_ex), .Q(ALU_wb) );
  regFFD_NBIT32_2 pipeline_LMD4 ( .CK(CLK), .RESET(n45), .ENABLE(RM), .D(
        LMD_out), .Q(LMD_wb) );
  regFFD_NBIT5_1 pipeline_RD4 ( .CK(CLK), .RESET(n44), .ENABLE(1'b1), .D(
        RD_mem), .Q(RD_wb) );
  FF_3 pipeline_wr_signal3 ( .CLK(CLK), .RESET(n45), .EN(1'b1), .D(
        wr_signal_mem1), .Q(wr_signal_wb) );
  FF_2 pipeline_WM ( .CLK(CLK), .RESET(n45), .EN(1'b1), .D(WM) );
  FF_1 pipeline_JAL ( .CLK(CLK), .RESET(n45), .EN(1'b1), .D(sel_saved_reg), 
        .Q(sel_saved_reg_wb) );
  regFFD_NBIT32_1 pipeline_NPC_wb ( .CK(CLK), .RESET(n45), .ENABLE(1'b1), .D(
        NPC_mem), .Q(NPC_wb) );
  MUX21_GENERIC_NBIT32_2 MUX_WB ( .A(ALU_wb), .B(LMD_wb), .SEL(S3), .Y(
        OUT_data) );
  MUX21_GENERIC_NBIT32_1 MUX_jal ( .A(NPC_wb), .B(OUT_data), .SEL(
        sel_saved_reg_wb), .Y(OUT_wb) );
  DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 add_240 ( .A(PC_fetch0), .SUM(NPC) );
  INV_X1 U3 ( .A(n49), .ZN(n35) );
  INV_X1 U4 ( .A(n48), .ZN(n36) );
  BUF_X2 U5 ( .A(RST), .Z(n45) );
  BUF_X1 U6 ( .A(n55), .Z(n38) );
  BUF_X1 U7 ( .A(n55), .Z(n37) );
  BUF_X1 U8 ( .A(n55), .Z(n39) );
  NOR4_X1 U9 ( .A1(n23), .A2(IR_Dec[22]), .A3(IR_Dec[24]), .A4(IR_Dec[23]), 
        .ZN(n20) );
  OR4_X1 U10 ( .A1(IR_Dec[26]), .A2(IR_Dec[25]), .A3(IR_Dec[2]), .A4(
        IR_Dec[28]), .ZN(n23) );
  OAI22_X1 U11 ( .A1(IR_Dec[31]), .A2(n13), .B1(n14), .B2(n48), .ZN(n34) );
  INV_X1 U12 ( .A(IR_Dec[31]), .ZN(n48) );
  NOR4_X1 U13 ( .A1(IR_Dec[30]), .A2(IR_Dec[28]), .A3(n49), .A4(n15), .ZN(n14)
         );
  AOI211_X1 U14 ( .C1(n16), .C2(n17), .A(n35), .B(IR_Dec[27]), .ZN(n13) );
  NAND4_X1 U15 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .ZN(n17) );
  NOR4_X1 U16 ( .A1(n22), .A2(IR_Dec[3]), .A3(IR_Dec[5]), .A4(IR_Dec[4]), .ZN(
        n21) );
  NOR4_X1 U17 ( .A1(n24), .A2(IR_Dec[16]), .A3(IR_Dec[18]), .A4(IR_Dec[17]), 
        .ZN(n19) );
  NOR4_X1 U18 ( .A1(n25), .A2(IR_Dec[0]), .A3(IR_Dec[11]), .A4(IR_Dec[10]), 
        .ZN(n18) );
  AOI21_X1 U19 ( .B1(jump_en), .B2(n11), .A(n47), .ZN(wr_signal_mem1) );
  NAND4_X1 U20 ( .A1(IR_26_mem[1]), .A2(IR_26_mem[0]), .A3(n12), .A4(n46), 
        .ZN(n11) );
  INV_X1 U21 ( .A(wr_signal_mem), .ZN(n47) );
  INV_X1 U22 ( .A(IR_26_mem[2]), .ZN(n46) );
  OR4_X1 U23 ( .A1(IR_Dec[13]), .A2(IR_Dec[12]), .A3(IR_Dec[15]), .A4(
        IR_Dec[14]), .ZN(n25) );
  OR4_X1 U24 ( .A1(IR_Dec[1]), .A2(IR_Dec[19]), .A3(IR_Dec[21]), .A4(
        IR_Dec[20]), .ZN(n24) );
  OR4_X1 U25 ( .A1(IR_Dec[7]), .A2(IR_Dec[6]), .A3(IR_Dec[9]), .A4(IR_Dec[8]), 
        .ZN(n22) );
  OAI21_X1 U26 ( .B1(IR_Dec[26]), .B2(n50), .A(IR_Dec[30]), .ZN(n16) );
  INV_X1 U27 ( .A(IR_Dec[28]), .ZN(n50) );
  INV_X1 U28 ( .A(IR_Dec[29]), .ZN(n49) );
  AOI22_X1 U29 ( .A1(n30), .A2(instruction_alu[1]), .B1(instruction_alu[2]), 
        .B2(n53), .ZN(n29) );
  INV_X1 U30 ( .A(instruction_alu[1]), .ZN(n53) );
  NOR2_X1 U31 ( .A1(instruction_alu[2]), .A2(n54), .ZN(n30) );
  NAND4_X1 U32 ( .A1(IR_26_mem[2]), .A2(IR_26_mem[0]), .A3(IR_26_mem[4]), .A4(
        n26), .ZN(N13) );
  NOR3_X1 U33 ( .A1(IR_26_mem[1]), .A2(IR_26_mem[5]), .A3(IR_26_mem[3]), .ZN(
        n26) );
  BUF_X2 U34 ( .A(RST), .Z(n44) );
  INV_X1 U35 ( .A(instruction_alu[3]), .ZN(n52) );
  INV_X1 U36 ( .A(instruction_alu[5]), .ZN(n51) );
  OR2_X1 U37 ( .A1(cond_mem), .A2(jump_en), .ZN(sel_npc) );
  INV_X1 U38 ( .A(instruction_alu[0]), .ZN(n54) );
  NOR2_X1 U39 ( .A1(IR_26_mem[5]), .A2(IR_26_mem[3]), .ZN(n12) );
  OR4_X1 U40 ( .A1(n27), .A2(n28), .A3(WM), .A4(RM), .ZN(DATA_MEM_ENABLE) );
  NOR4_X1 U41 ( .A1(n31), .A2(n54), .A3(instruction_alu[5]), .A4(
        instruction_alu[3]), .ZN(n27) );
  NOR4_X1 U42 ( .A1(instruction_alu[4]), .A2(n29), .A3(n52), .A4(n51), .ZN(n28) );
  AND2_X1 U43 ( .A1(IR_26_mem[0]), .A2(jump_en), .ZN(sel_saved_reg) );
  INV_X1 U44 ( .A(sb_op), .ZN(n55) );
  AND2_X1 U45 ( .A1(regB_mem[31]), .A2(n37), .ZN(DATA_MEM_IN[31]) );
  AND2_X1 U46 ( .A1(regB_mem[30]), .A2(n37), .ZN(DATA_MEM_IN[30]) );
  AND2_X1 U47 ( .A1(regB_mem[29]), .A2(n37), .ZN(DATA_MEM_IN[29]) );
  AND2_X1 U48 ( .A1(regB_mem[28]), .A2(n37), .ZN(DATA_MEM_IN[28]) );
  AND2_X1 U49 ( .A1(regB_mem[27]), .A2(n37), .ZN(DATA_MEM_IN[27]) );
  AND2_X1 U50 ( .A1(regB_mem[26]), .A2(n37), .ZN(DATA_MEM_IN[26]) );
  AND2_X1 U51 ( .A1(regB_mem[25]), .A2(n37), .ZN(DATA_MEM_IN[25]) );
  AND2_X1 U52 ( .A1(regB_mem[24]), .A2(n37), .ZN(DATA_MEM_IN[24]) );
  AND2_X1 U53 ( .A1(regB_mem[23]), .A2(n37), .ZN(DATA_MEM_IN[23]) );
  AND2_X1 U54 ( .A1(regB_mem[22]), .A2(n38), .ZN(DATA_MEM_IN[22]) );
  AND2_X1 U55 ( .A1(regB_mem[21]), .A2(n38), .ZN(DATA_MEM_IN[21]) );
  AND2_X1 U56 ( .A1(regB_mem[20]), .A2(n38), .ZN(DATA_MEM_IN[20]) );
  AND2_X1 U57 ( .A1(regB_mem[19]), .A2(n38), .ZN(DATA_MEM_IN[19]) );
  AND2_X1 U58 ( .A1(regB_mem[18]), .A2(n38), .ZN(DATA_MEM_IN[18]) );
  AND2_X1 U59 ( .A1(regB_mem[17]), .A2(n38), .ZN(DATA_MEM_IN[17]) );
  AND2_X1 U60 ( .A1(regB_mem[16]), .A2(n38), .ZN(DATA_MEM_IN[16]) );
  AND2_X1 U61 ( .A1(regB_mem[15]), .A2(n38), .ZN(DATA_MEM_IN[15]) );
  AND2_X1 U64 ( .A1(regB_mem[14]), .A2(n38), .ZN(DATA_MEM_IN[14]) );
  AND2_X1 U65 ( .A1(regB_mem[13]), .A2(n38), .ZN(DATA_MEM_IN[13]) );
  AND2_X1 U66 ( .A1(regB_mem[12]), .A2(n38), .ZN(DATA_MEM_IN[12]) );
  AND2_X1 U67 ( .A1(regB_mem[9]), .A2(n37), .ZN(DATA_MEM_IN[9]) );
  AND2_X1 U68 ( .A1(regB_mem[8]), .A2(n37), .ZN(DATA_MEM_IN[8]) );
  AND2_X1 U69 ( .A1(regB_mem[11]), .A2(n39), .ZN(DATA_MEM_IN[11]) );
  AND2_X1 U70 ( .A1(regB_mem[10]), .A2(n39), .ZN(DATA_MEM_IN[10]) );
  CLKBUF_X1 U71 ( .A(N13), .Z(n40) );
  CLKBUF_X1 U72 ( .A(N13), .Z(n41) );
  CLKBUF_X1 U73 ( .A(N13), .Z(n42) );
  CLKBUF_X1 U74 ( .A(N13), .Z(n43) );
endmodule


module DLX_IR_SIZE32_PC_SIZE32 ( CLK, RST, IRAM_ADDRESS, IRAM_ISSUE, 
        IRAM_READY, IRAM_DATA, DRAM_ADDRESS, DRAM_ISSUE, DRAM_READNOTWRITE, 
        DRAM_READY, DRAM_DATA );
  output [31:0] IRAM_ADDRESS;
  input [63:0] IRAM_DATA;
  output [31:0] DRAM_ADDRESS;
  inout [63:0] DRAM_DATA;
  input CLK, RST, IRAM_READY, DRAM_READY;
  output IRAM_ISSUE, DRAM_ISSUE, DRAM_READNOTWRITE;
  wire   signed_unsigned_i, lhi_sel_i, sb_op_i, trap_cs_i, ret_cs_i,
         DATA_MEM_WM_i, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272;
  wire   [31:0] IR;
  wire   [31:0] PC;
  wire   [5:0] ALU_OPCODE_i;
  wire   [31:0] DATA_MEM_IN_i;
  wire   [31:0] dram_data_i;
  tri   [63:0] DRAM_DATA;
  assign IRAM_ADDRESS[31] = 1'b0;
  assign IRAM_ADDRESS[30] = 1'b0;
  assign IRAM_ADDRESS[29] = 1'b0;
  assign IRAM_ADDRESS[28] = 1'b0;
  assign IRAM_ADDRESS[27] = 1'b0;
  assign IRAM_ADDRESS[26] = 1'b0;
  assign IRAM_ADDRESS[25] = 1'b0;
  assign IRAM_ADDRESS[24] = 1'b0;
  assign IRAM_ADDRESS[23] = 1'b0;
  assign IRAM_ADDRESS[22] = 1'b0;
  assign IRAM_ADDRESS[21] = 1'b0;
  assign IRAM_ADDRESS[20] = 1'b0;
  assign IRAM_ADDRESS[19] = 1'b0;
  assign IRAM_ADDRESS[18] = 1'b0;
  assign IRAM_ADDRESS[17] = 1'b0;
  assign IRAM_ADDRESS[16] = 1'b0;
  assign IRAM_ADDRESS[15] = 1'b0;
  assign IRAM_ADDRESS[14] = 1'b0;
  assign IRAM_ADDRESS[13] = 1'b0;
  assign IRAM_ADDRESS[12] = 1'b0;
  assign IRAM_ADDRESS[11] = 1'b0;
  assign IRAM_ADDRESS[10] = 1'b0;
  assign IRAM_ADDRESS[9] = 1'b0;
  assign IRAM_ADDRESS[8] = 1'b0;
  assign IRAM_ADDRESS[7] = 1'b0;
  assign IRAM_ADDRESS[6] = 1'b0;
  assign IRAM_ADDRESS[5] = 1'b0;
  assign IRAM_ADDRESS[4] = 1'b0;
  assign IRAM_ADDRESS[3] = 1'b0;
  assign IRAM_ADDRESS[2] = 1'b0;
  assign IRAM_ADDRESS[1] = 1'b0;
  assign IRAM_ADDRESS[0] = 1'b0;

  DFF_X1 DRAM_READNOTWRITE_reg ( .D(n271), .CK(CLK), .Q(DRAM_READNOTWRITE) );
  dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 CU_I ( 
        .Clk(CLK), .Rst(RST), .IR_IN({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .ALU_OPCODE(ALU_OPCODE_i), .signed_unsigned(signed_unsigned_i), 
        .lhi_sel(lhi_sel_i), .sb_op(sb_op_i), .s_trap(trap_cs_i), .s_ret(
        ret_cs_i) );
  DATAPTH_NBIT32_REG_BIT5 DTPTH_I ( .CLK(CLK), .RST(RST), .PC({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IR({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .NPC_LATCH_EN(1'b0), .ir_LATCH_EN(1'b0), 
        .signed_op(signed_unsigned_i), .trap_cs(trap_cs_i), .ret_cs(ret_cs_i), 
        .RF1(1'b0), .RF2(1'b0), .WF1(1'b0), .regImm_LATCH_EN(1'b0), .S1(1'b0), 
        .S2(1'b0), .EN2(1'b0), .lhi_sel(lhi_sel_i), .jump_en(1'b0), 
        .branch_cond(1'b0), .sb_op(sb_op_i), .RM(1'b0), .WM(1'b0), .EN3(1'b0), 
        .S3(1'b0), .instruction_alu(ALU_OPCODE_i), .DATA_MEM_ADDR(DRAM_ADDRESS), .DATA_MEM_IN(DATA_MEM_IN_i), .DATA_MEM_OUT(dram_data_i), .DATA_MEM_ENABLE(
        DRAM_ISSUE), .DATA_MEM_WM(DATA_MEM_WM_i) );
  TBUF_X1 \DRAM_DATA_tri[32]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[32]) );
  TBUF_X1 \DRAM_DATA_tri[33]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[33]) );
  TBUF_X1 \DRAM_DATA_tri[34]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[34]) );
  TBUF_X1 \DRAM_DATA_tri[35]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[35]) );
  TBUF_X1 \DRAM_DATA_tri[36]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[36]) );
  TBUF_X1 \DRAM_DATA_tri[37]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[37]) );
  TBUF_X1 \DRAM_DATA_tri[38]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[38]) );
  TBUF_X1 \DRAM_DATA_tri[39]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[39]) );
  TBUF_X1 \DRAM_DATA_tri[40]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[40]) );
  TBUF_X1 \DRAM_DATA_tri[41]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[41]) );
  TBUF_X1 \DRAM_DATA_tri[42]  ( .A(1'b0), .EN(n264), .Z(DRAM_DATA[42]) );
  TBUF_X1 \DRAM_DATA_tri[43]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[43]) );
  TBUF_X1 \DRAM_DATA_tri[44]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[44]) );
  TBUF_X1 \DRAM_DATA_tri[45]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[45]) );
  TBUF_X1 \DRAM_DATA_tri[46]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[46]) );
  TBUF_X1 \DRAM_DATA_tri[47]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[47]) );
  TBUF_X1 \DRAM_DATA_tri[48]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[48]) );
  TBUF_X1 \DRAM_DATA_tri[49]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[49]) );
  TBUF_X1 \DRAM_DATA_tri[50]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[50]) );
  TBUF_X1 \DRAM_DATA_tri[51]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[51]) );
  TBUF_X1 \DRAM_DATA_tri[52]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[52]) );
  TBUF_X1 \DRAM_DATA_tri[53]  ( .A(1'b0), .EN(n265), .Z(DRAM_DATA[53]) );
  TBUF_X1 \DRAM_DATA_tri[54]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[54]) );
  TBUF_X1 \DRAM_DATA_tri[55]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[55]) );
  TBUF_X1 \DRAM_DATA_tri[56]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[56]) );
  TBUF_X1 \DRAM_DATA_tri[57]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[57]) );
  TBUF_X1 \DRAM_DATA_tri[58]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[58]) );
  TBUF_X1 \DRAM_DATA_tri[59]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[59]) );
  TBUF_X1 \DRAM_DATA_tri[60]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[60]) );
  TBUF_X1 \DRAM_DATA_tri[61]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[61]) );
  TBUF_X1 \DRAM_DATA_tri[62]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[62]) );
  TBUF_X1 \DRAM_DATA_tri[63]  ( .A(1'b0), .EN(n266), .Z(DRAM_DATA[63]) );
  TBUF_X1 \DRAM_DATA_tri[8]  ( .A(DATA_MEM_IN_i[8]), .EN(n267), .Z(
        DRAM_DATA[8]) );
  TBUF_X1 \DRAM_DATA_tri[9]  ( .A(DATA_MEM_IN_i[9]), .EN(n267), .Z(
        DRAM_DATA[9]) );
  TBUF_X1 \DRAM_DATA_tri[10]  ( .A(DATA_MEM_IN_i[10]), .EN(n267), .Z(
        DRAM_DATA[10]) );
  TBUF_X1 \DRAM_DATA_tri[11]  ( .A(DATA_MEM_IN_i[11]), .EN(n267), .Z(
        DRAM_DATA[11]) );
  TBUF_X1 \DRAM_DATA_tri[12]  ( .A(DATA_MEM_IN_i[12]), .EN(n268), .Z(
        DRAM_DATA[12]) );
  TBUF_X1 \DRAM_DATA_tri[13]  ( .A(DATA_MEM_IN_i[13]), .EN(n268), .Z(
        DRAM_DATA[13]) );
  TBUF_X1 \DRAM_DATA_tri[14]  ( .A(DATA_MEM_IN_i[14]), .EN(n268), .Z(
        DRAM_DATA[14]) );
  TBUF_X1 \DRAM_DATA_tri[15]  ( .A(DATA_MEM_IN_i[15]), .EN(n268), .Z(
        DRAM_DATA[15]) );
  TBUF_X1 \DRAM_DATA_tri[16]  ( .A(DATA_MEM_IN_i[16]), .EN(n268), .Z(
        DRAM_DATA[16]) );
  TBUF_X1 \DRAM_DATA_tri[17]  ( .A(DATA_MEM_IN_i[17]), .EN(n268), .Z(
        DRAM_DATA[17]) );
  TBUF_X1 \DRAM_DATA_tri[18]  ( .A(DATA_MEM_IN_i[18]), .EN(n268), .Z(
        DRAM_DATA[18]) );
  TBUF_X1 \DRAM_DATA_tri[19]  ( .A(DATA_MEM_IN_i[19]), .EN(n268), .Z(
        DRAM_DATA[19]) );
  TBUF_X1 \DRAM_DATA_tri[20]  ( .A(DATA_MEM_IN_i[20]), .EN(n268), .Z(
        DRAM_DATA[20]) );
  TBUF_X1 \DRAM_DATA_tri[21]  ( .A(DATA_MEM_IN_i[21]), .EN(n268), .Z(
        DRAM_DATA[21]) );
  TBUF_X1 \DRAM_DATA_tri[22]  ( .A(DATA_MEM_IN_i[22]), .EN(n268), .Z(
        DRAM_DATA[22]) );
  TBUF_X1 \DRAM_DATA_tri[23]  ( .A(DATA_MEM_IN_i[23]), .EN(n269), .Z(
        DRAM_DATA[23]) );
  TBUF_X1 \DRAM_DATA_tri[24]  ( .A(DATA_MEM_IN_i[24]), .EN(n269), .Z(
        DRAM_DATA[24]) );
  TBUF_X1 \DRAM_DATA_tri[25]  ( .A(DATA_MEM_IN_i[25]), .EN(n269), .Z(
        DRAM_DATA[25]) );
  TBUF_X1 \DRAM_DATA_tri[26]  ( .A(DATA_MEM_IN_i[26]), .EN(n269), .Z(
        DRAM_DATA[26]) );
  TBUF_X1 \DRAM_DATA_tri[27]  ( .A(DATA_MEM_IN_i[27]), .EN(n269), .Z(
        DRAM_DATA[27]) );
  TBUF_X1 \DRAM_DATA_tri[28]  ( .A(DATA_MEM_IN_i[28]), .EN(n269), .Z(
        DRAM_DATA[28]) );
  TBUF_X1 \DRAM_DATA_tri[29]  ( .A(DATA_MEM_IN_i[29]), .EN(n269), .Z(
        DRAM_DATA[29]) );
  TBUF_X1 \DRAM_DATA_tri[30]  ( .A(DATA_MEM_IN_i[30]), .EN(n269), .Z(
        DRAM_DATA[30]) );
  TBUF_X1 \DRAM_DATA_tri[31]  ( .A(DATA_MEM_IN_i[31]), .EN(n269), .Z(
        DRAM_DATA[31]) );
  TBUF_X1 \DRAM_DATA_tri[0]  ( .A(DATA_MEM_IN_i[0]), .EN(n266), .Z(
        DRAM_DATA[0]) );
  TBUF_X1 \DRAM_DATA_tri[1]  ( .A(DATA_MEM_IN_i[1]), .EN(n267), .Z(
        DRAM_DATA[1]) );
  TBUF_X1 \DRAM_DATA_tri[2]  ( .A(DATA_MEM_IN_i[2]), .EN(n267), .Z(
        DRAM_DATA[2]) );
  TBUF_X1 \DRAM_DATA_tri[3]  ( .A(DATA_MEM_IN_i[3]), .EN(n267), .Z(
        DRAM_DATA[3]) );
  TBUF_X1 \DRAM_DATA_tri[4]  ( .A(DATA_MEM_IN_i[4]), .EN(n267), .Z(
        DRAM_DATA[4]) );
  TBUF_X1 \DRAM_DATA_tri[5]  ( .A(DATA_MEM_IN_i[5]), .EN(n267), .Z(
        DRAM_DATA[5]) );
  TBUF_X1 \DRAM_DATA_tri[6]  ( .A(DATA_MEM_IN_i[6]), .EN(n267), .Z(
        DRAM_DATA[6]) );
  TBUF_X1 \DRAM_DATA_tri[7]  ( .A(DATA_MEM_IN_i[7]), .EN(n267), .Z(
        DRAM_DATA[7]) );
  BUF_X1 U342 ( .A(n263), .Z(n270) );
  BUF_X1 U343 ( .A(n263), .Z(n269) );
  BUF_X1 U344 ( .A(n263), .Z(n268) );
  BUF_X1 U345 ( .A(n262), .Z(n267) );
  BUF_X1 U346 ( .A(n262), .Z(n266) );
  BUF_X1 U347 ( .A(n262), .Z(n265) );
  BUF_X1 U348 ( .A(n262), .Z(n264) );
  BUF_X1 U349 ( .A(n263), .Z(n271) );
  BUF_X1 U350 ( .A(n272), .Z(n262) );
  BUF_X1 U351 ( .A(n272), .Z(n263) );
  AND2_X1 U352 ( .A1(DRAM_DATA[63]), .A2(n271), .ZN(dram_data_i[31]) );
  AND2_X1 U353 ( .A1(DRAM_DATA[40]), .A2(n271), .ZN(dram_data_i[8]) );
  AND2_X1 U354 ( .A1(DRAM_DATA[41]), .A2(n271), .ZN(dram_data_i[9]) );
  AND2_X1 U355 ( .A1(DRAM_DATA[42]), .A2(n269), .ZN(dram_data_i[10]) );
  AND2_X1 U356 ( .A1(DRAM_DATA[43]), .A2(n269), .ZN(dram_data_i[11]) );
  AND2_X1 U357 ( .A1(DRAM_DATA[44]), .A2(n270), .ZN(dram_data_i[12]) );
  AND2_X1 U358 ( .A1(DRAM_DATA[45]), .A2(n270), .ZN(dram_data_i[13]) );
  AND2_X1 U359 ( .A1(DRAM_DATA[46]), .A2(n270), .ZN(dram_data_i[14]) );
  AND2_X1 U360 ( .A1(DRAM_DATA[47]), .A2(n270), .ZN(dram_data_i[15]) );
  AND2_X1 U361 ( .A1(DRAM_DATA[52]), .A2(n270), .ZN(dram_data_i[20]) );
  AND2_X1 U362 ( .A1(DRAM_DATA[53]), .A2(n270), .ZN(dram_data_i[21]) );
  AND2_X1 U363 ( .A1(DRAM_DATA[54]), .A2(n270), .ZN(dram_data_i[22]) );
  AND2_X1 U364 ( .A1(DRAM_DATA[55]), .A2(n270), .ZN(dram_data_i[23]) );
  AND2_X1 U365 ( .A1(DRAM_DATA[56]), .A2(n270), .ZN(dram_data_i[24]) );
  AND2_X1 U366 ( .A1(DRAM_DATA[57]), .A2(n270), .ZN(dram_data_i[25]) );
  AND2_X1 U367 ( .A1(DRAM_DATA[58]), .A2(n270), .ZN(dram_data_i[26]) );
  AND2_X1 U368 ( .A1(DRAM_DATA[59]), .A2(n271), .ZN(dram_data_i[27]) );
  AND2_X1 U369 ( .A1(DRAM_DATA[60]), .A2(n271), .ZN(dram_data_i[28]) );
  AND2_X1 U370 ( .A1(DRAM_DATA[61]), .A2(n271), .ZN(dram_data_i[29]) );
  AND2_X1 U371 ( .A1(DRAM_DATA[62]), .A2(n271), .ZN(dram_data_i[30]) );
  AND2_X1 U372 ( .A1(DRAM_DATA[48]), .A2(n270), .ZN(dram_data_i[16]) );
  AND2_X1 U373 ( .A1(DRAM_DATA[49]), .A2(n270), .ZN(dram_data_i[17]) );
  AND2_X1 U374 ( .A1(DRAM_DATA[50]), .A2(n270), .ZN(dram_data_i[18]) );
  AND2_X1 U375 ( .A1(DRAM_DATA[51]), .A2(n270), .ZN(dram_data_i[19]) );
  AND2_X1 U376 ( .A1(DRAM_DATA[32]), .A2(n269), .ZN(dram_data_i[0]) );
  AND2_X1 U377 ( .A1(DRAM_DATA[33]), .A2(n270), .ZN(dram_data_i[1]) );
  AND2_X1 U378 ( .A1(DRAM_DATA[34]), .A2(n271), .ZN(dram_data_i[2]) );
  AND2_X1 U379 ( .A1(DRAM_DATA[35]), .A2(n271), .ZN(dram_data_i[3]) );
  AND2_X1 U380 ( .A1(DRAM_DATA[36]), .A2(n271), .ZN(dram_data_i[4]) );
  AND2_X1 U381 ( .A1(DRAM_DATA[37]), .A2(n271), .ZN(dram_data_i[5]) );
  AND2_X1 U382 ( .A1(DRAM_DATA[38]), .A2(n271), .ZN(dram_data_i[6]) );
  AND2_X1 U383 ( .A1(DRAM_DATA[39]), .A2(n271), .ZN(dram_data_i[7]) );
  INV_X1 U384 ( .A(DATA_MEM_WM_i), .ZN(n272) );
endmodule

